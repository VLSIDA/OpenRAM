**************************************************
* OpenRAM generated memory.
* Words: 1024
* Data bits: 32
* Banks: 1
* Column mux: 4:1
**************************************************

* ptx M{0} {1} nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p

* ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p

.SUBCKT pnand2_1 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand2_1

.SUBCKT pnand3_1 A B C Z vdd gnd
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand3_1

* ptx M{0} {1} nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p

* ptx M{0} {1} pmos_vtg m=1 w=0.405u l=0.05u pd=0.91u ps=0.91u as=0.050625p ad=0.050625p

.SUBCKT pnor2_1 A B Z vdd gnd
Mpnor2_pmos1 vdd A net1 vdd pmos_vtg m=1 w=0.405u l=0.05u pd=0.91u ps=0.91u as=0.050625p ad=0.050625p
Mpnor2_pmos2 net1 B Z vdd pmos_vtg m=1 w=0.405u l=0.05u pd=0.91u ps=0.91u as=0.050625p ad=0.050625p
Mpnor2_nmos1 Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
Mpnor2_nmos2 Z B gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pnor2_1

.SUBCKT pinv_1 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_1

* ptx M{0} {1} nmos_vtg m=2 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p

* ptx M{0} {1} pmos_vtg m=2 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p

.SUBCKT pinv_2 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=2 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=2 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_2

* ptx M{0} {1} nmos_vtg m=3 w=0.12u l=0.05u pd=0.34u ps=0.34u as=0.015p ad=0.015p

* ptx M{0} {1} pmos_vtg m=3 w=0.36u l=0.05u pd=0.82u ps=0.82u as=0.045p ad=0.045p

.SUBCKT pinv_3 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=3 w=0.36u l=0.05u pd=0.82u ps=0.82u as=0.045p ad=0.045p
Mpinv_nmos Z A gnd gnd nmos_vtg m=3 w=0.12u l=0.05u pd=0.34u ps=0.34u as=0.015p ad=0.015p
.ENDS pinv_3

* ptx M{0} {1} nmos_vtg m=6 w=0.12u l=0.05u pd=0.34u ps=0.34u as=0.015p ad=0.015p

* ptx M{0} {1} pmos_vtg m=6 w=0.36u l=0.05u pd=0.82u ps=0.82u as=0.045p ad=0.045p

.SUBCKT pinv_4 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=6 w=0.36u l=0.05u pd=0.82u ps=0.82u as=0.045p ad=0.045p
Mpinv_nmos Z A gnd gnd nmos_vtg m=6 w=0.12u l=0.05u pd=0.34u ps=0.34u as=0.015p ad=0.015p
.ENDS pinv_4

* ptx M{0} {1} nmos_vtg m=12 w=0.12u l=0.05u pd=0.34u ps=0.34u as=0.015p ad=0.015p

* ptx M{0} {1} pmos_vtg m=12 w=0.36u l=0.05u pd=0.82u ps=0.82u as=0.045p ad=0.045p

.SUBCKT pinv_5 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=12 w=0.36u l=0.05u pd=0.82u ps=0.82u as=0.045p ad=0.045p
Mpinv_nmos Z A gnd gnd nmos_vtg m=12 w=0.12u l=0.05u pd=0.34u ps=0.34u as=0.015p ad=0.015p
.ENDS pinv_5
*master-slave flip-flop with both output and inverted ouput

.SUBCKT ms_flop din dout dout_bar clk vdd gnd
xmaster din mout mout_bar clk clk_bar vdd gnd dlatch
xslave mout_bar dout_bar dout clk_bar clk_nn vdd gnd dlatch
.ENDS flop

.SUBCKT dlatch din dout dout_bar clk clk_bar vdd gnd
*clk inverter
mPff1 clk_bar clk vdd vdd PMOS_VTG W=180.0n L=50n m=1
mNff1 clk_bar clk gnd gnd NMOS_VTG W=90n L=50n m=1

*transmission gate 1
mtmP1 din clk int1 vdd PMOS_VTG W=180.0n L=50n m=1
mtmN1 din clk_bar int1 gnd NMOS_VTG W=90n L=50n m=1

*foward inverter
mPff3 dout_bar int1 vdd vdd PMOS_VTG W=180.0n L=50n m=1
mNff3 dout_bar int1 gnd gnd NMOS_VTG W=90n L=50n m=1

*backward inverter
mPff4 dout dout_bar vdd vdd PMOS_VTG W=180.0n L=50n m=1
mNf4 dout dout_bar gnd gnd NMOS_VTG W=90n L=50n m=1

*transmission gate 2
mtmP2 int1 clk_bar dout vdd PMOS_VTG W=180.0n L=50n m=1
mtmN2 int1 clk dout gnd NMOS_VTG W=90n L=50n m=1
.ENDS dlatch


.SUBCKT msf_control din[0] din[1] din[2] dout[0] dout_bar[0] dout[1] dout_bar[1] dout[2] dout_bar[2] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
XXdff1 din[1] dout[1] dout_bar[1] clk vdd gnd ms_flop
XXdff2 din[2] dout[2] dout_bar[2] clk vdd gnd ms_flop
.ENDS msf_control

.SUBCKT replica_cell_6t bl br wl vdd gnd
MM3 bl wl gnd gnd NMOS_VTG W=135.00n L=50n
MM2 br wl net4 gnd NMOS_VTG W=135.00n L=50n
MM1 gnd net4 gnd gnd NMOS_VTG W=205.00n L=50n
MM0 net4 gnd gnd gnd NMOS_VTG W=205.00n L=50n
MM5 gnd net4 vdd vdd PMOS_VTG W=90n L=50n
MM4 net4 gnd vdd vdd PMOS_VTG W=90n L=50n
.ENDS replica_cell_6t


.SUBCKT cell_6t bl br wl vdd gnd
MM3 bl wl net10 gnd NMOS_VTG W=135.00n L=50n
MM2 br wl net4 gnd NMOS_VTG W=135.00n L=50n
MM1 net10 net4 gnd gnd NMOS_VTG W=205.00n L=50n
MM0 net4 net10 gnd gnd NMOS_VTG W=205.00n L=50n
MM5 net10 net4 vdd vdd PMOS_VTG W=90n L=50n
MM4 net4 net10 vdd vdd PMOS_VTG W=90n L=50n
.ENDS cell_6t


.SUBCKT bitline_load bl[0] br[0] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] vdd gnd
Xbit_r0_c0 bl[0] br[0] wl[0] vdd gnd cell_6t
Xbit_r1_c0 bl[0] br[0] wl[1] vdd gnd cell_6t
Xbit_r2_c0 bl[0] br[0] wl[2] vdd gnd cell_6t
Xbit_r3_c0 bl[0] br[0] wl[3] vdd gnd cell_6t
Xbit_r4_c0 bl[0] br[0] wl[4] vdd gnd cell_6t
Xbit_r5_c0 bl[0] br[0] wl[5] vdd gnd cell_6t
Xbit_r6_c0 bl[0] br[0] wl[6] vdd gnd cell_6t
Xbit_r7_c0 bl[0] br[0] wl[7] vdd gnd cell_6t
Xbit_r8_c0 bl[0] br[0] wl[8] vdd gnd cell_6t
Xbit_r9_c0 bl[0] br[0] wl[9] vdd gnd cell_6t
Xbit_r10_c0 bl[0] br[0] wl[10] vdd gnd cell_6t
Xbit_r11_c0 bl[0] br[0] wl[11] vdd gnd cell_6t
Xbit_r12_c0 bl[0] br[0] wl[12] vdd gnd cell_6t
Xbit_r13_c0 bl[0] br[0] wl[13] vdd gnd cell_6t
Xbit_r14_c0 bl[0] br[0] wl[14] vdd gnd cell_6t
Xbit_r15_c0 bl[0] br[0] wl[15] vdd gnd cell_6t
Xbit_r16_c0 bl[0] br[0] wl[16] vdd gnd cell_6t
Xbit_r17_c0 bl[0] br[0] wl[17] vdd gnd cell_6t
Xbit_r18_c0 bl[0] br[0] wl[18] vdd gnd cell_6t
Xbit_r19_c0 bl[0] br[0] wl[19] vdd gnd cell_6t
Xbit_r20_c0 bl[0] br[0] wl[20] vdd gnd cell_6t
Xbit_r21_c0 bl[0] br[0] wl[21] vdd gnd cell_6t
Xbit_r22_c0 bl[0] br[0] wl[22] vdd gnd cell_6t
Xbit_r23_c0 bl[0] br[0] wl[23] vdd gnd cell_6t
Xbit_r24_c0 bl[0] br[0] wl[24] vdd gnd cell_6t
Xbit_r25_c0 bl[0] br[0] wl[25] vdd gnd cell_6t
Xbit_r26_c0 bl[0] br[0] wl[26] vdd gnd cell_6t
Xbit_r27_c0 bl[0] br[0] wl[27] vdd gnd cell_6t
Xbit_r28_c0 bl[0] br[0] wl[28] vdd gnd cell_6t
Xbit_r29_c0 bl[0] br[0] wl[29] vdd gnd cell_6t
Xbit_r30_c0 bl[0] br[0] wl[30] vdd gnd cell_6t
Xbit_r31_c0 bl[0] br[0] wl[31] vdd gnd cell_6t
Xbit_r32_c0 bl[0] br[0] wl[32] vdd gnd cell_6t
Xbit_r33_c0 bl[0] br[0] wl[33] vdd gnd cell_6t
Xbit_r34_c0 bl[0] br[0] wl[34] vdd gnd cell_6t
Xbit_r35_c0 bl[0] br[0] wl[35] vdd gnd cell_6t
Xbit_r36_c0 bl[0] br[0] wl[36] vdd gnd cell_6t
Xbit_r37_c0 bl[0] br[0] wl[37] vdd gnd cell_6t
Xbit_r38_c0 bl[0] br[0] wl[38] vdd gnd cell_6t
Xbit_r39_c0 bl[0] br[0] wl[39] vdd gnd cell_6t
Xbit_r40_c0 bl[0] br[0] wl[40] vdd gnd cell_6t
Xbit_r41_c0 bl[0] br[0] wl[41] vdd gnd cell_6t
Xbit_r42_c0 bl[0] br[0] wl[42] vdd gnd cell_6t
Xbit_r43_c0 bl[0] br[0] wl[43] vdd gnd cell_6t
Xbit_r44_c0 bl[0] br[0] wl[44] vdd gnd cell_6t
Xbit_r45_c0 bl[0] br[0] wl[45] vdd gnd cell_6t
Xbit_r46_c0 bl[0] br[0] wl[46] vdd gnd cell_6t
Xbit_r47_c0 bl[0] br[0] wl[47] vdd gnd cell_6t
Xbit_r48_c0 bl[0] br[0] wl[48] vdd gnd cell_6t
Xbit_r49_c0 bl[0] br[0] wl[49] vdd gnd cell_6t
Xbit_r50_c0 bl[0] br[0] wl[50] vdd gnd cell_6t
Xbit_r51_c0 bl[0] br[0] wl[51] vdd gnd cell_6t
.ENDS bitline_load

.SUBCKT pinv_6 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_6

.SUBCKT delay_chain in out vdd gnd
Xdinv0 in s1 vdd gnd pinv_6
Xdinv1 s1 s2n1 vdd gnd pinv_6
Xdinv2 s1 s2n2 vdd gnd pinv_6
Xdinv3 s1 s2 vdd gnd pinv_6
Xdinv4 s2 s3n1 vdd gnd pinv_6
Xdinv5 s2 s3n2 vdd gnd pinv_6
Xdinv6 s2 s3 vdd gnd pinv_6
Xdinv7 s3 s4n1 vdd gnd pinv_6
Xdinv8 s3 s4n2 vdd gnd pinv_6
Xdinv9 s3 s4 vdd gnd pinv_6
Xdinv10 s4 s5n1 vdd gnd pinv_6
Xdinv11 s4 s5n2 vdd gnd pinv_6
Xdinv12 s4 out vdd gnd pinv_6
.ENDS delay_chain

.SUBCKT pinv_7 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_7

* ptx M{0} {1} pmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p

.SUBCKT replica_bitline en out vdd gnd
Xrbl_inv bl[0] out vdd gnd pinv_7
Mrbl_access_tx vdd delayed_en bl[0] vdd pmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
Xdelay_chain en delayed_en vdd gnd delay_chain
Xbitcell bl[0] br[0] delayed_en vdd gnd replica_cell_6t
Xload bl[0] br[0] gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd vdd gnd bitline_load
.ENDS replica_bitline

.SUBCKT control_logic csb web oeb clk s_en w_en tri_en tri_en_bar clk_bar clk_buf vdd gnd
Xmsf_control oeb csb web oe_bar oe cs_bar cs we_bar we clk_buf vdd gnd msf_control
Xinv_clk1_bar clk clk1_bar vdd gnd pinv_2
Xinv_clk2 clk1_bar clk2 vdd gnd pinv_3
Xinv_clk_bar clk2 clk_bar vdd gnd pinv_4
Xinv_clk_buf clk_bar clk_buf vdd gnd pinv_5
Xnand3_rblk_bar clk_bar oe cs rblk_bar vdd gnd pnand3_1
Xinv_rblk rblk_bar rblk vdd gnd pinv_1
Xnor2_tri_en clk_buf oe_bar tri_en vdd gnd pnor2_1
Xnand2_tri_en clk_bar oe tri_en_bar vdd gnd pnand2_1
Xinv_s_en pre_s_en_bar s_en vdd gnd pinv_1
Xinv_pre_s_en_bar pre_s_en pre_s_en_bar vdd gnd pinv_1
Xnand3_w_en_bar clk_bar cs we w_en_bar vdd gnd pnand3_1
Xinv_pre_w_en w_en_bar pre_w_en vdd gnd pinv_1
Xinv_pre_w_en_bar pre_w_en pre_w_en_bar vdd gnd pinv_1
Xinv_w_en2 pre_w_en_bar w_en vdd gnd pinv_1
Xreplica_bitline rblk pre_s_en vdd gnd replica_bitline
.ENDS control_logic

.SUBCKT bitcell_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] vdd gnd
Xbit_r0_c0 bl[0] br[0] wl[0] vdd gnd cell_6t
Xbit_r1_c0 bl[0] br[0] wl[1] vdd gnd cell_6t
Xbit_r2_c0 bl[0] br[0] wl[2] vdd gnd cell_6t
Xbit_r3_c0 bl[0] br[0] wl[3] vdd gnd cell_6t
Xbit_r4_c0 bl[0] br[0] wl[4] vdd gnd cell_6t
Xbit_r5_c0 bl[0] br[0] wl[5] vdd gnd cell_6t
Xbit_r6_c0 bl[0] br[0] wl[6] vdd gnd cell_6t
Xbit_r7_c0 bl[0] br[0] wl[7] vdd gnd cell_6t
Xbit_r8_c0 bl[0] br[0] wl[8] vdd gnd cell_6t
Xbit_r9_c0 bl[0] br[0] wl[9] vdd gnd cell_6t
Xbit_r10_c0 bl[0] br[0] wl[10] vdd gnd cell_6t
Xbit_r11_c0 bl[0] br[0] wl[11] vdd gnd cell_6t
Xbit_r12_c0 bl[0] br[0] wl[12] vdd gnd cell_6t
Xbit_r13_c0 bl[0] br[0] wl[13] vdd gnd cell_6t
Xbit_r14_c0 bl[0] br[0] wl[14] vdd gnd cell_6t
Xbit_r15_c0 bl[0] br[0] wl[15] vdd gnd cell_6t
Xbit_r16_c0 bl[0] br[0] wl[16] vdd gnd cell_6t
Xbit_r17_c0 bl[0] br[0] wl[17] vdd gnd cell_6t
Xbit_r18_c0 bl[0] br[0] wl[18] vdd gnd cell_6t
Xbit_r19_c0 bl[0] br[0] wl[19] vdd gnd cell_6t
Xbit_r20_c0 bl[0] br[0] wl[20] vdd gnd cell_6t
Xbit_r21_c0 bl[0] br[0] wl[21] vdd gnd cell_6t
Xbit_r22_c0 bl[0] br[0] wl[22] vdd gnd cell_6t
Xbit_r23_c0 bl[0] br[0] wl[23] vdd gnd cell_6t
Xbit_r24_c0 bl[0] br[0] wl[24] vdd gnd cell_6t
Xbit_r25_c0 bl[0] br[0] wl[25] vdd gnd cell_6t
Xbit_r26_c0 bl[0] br[0] wl[26] vdd gnd cell_6t
Xbit_r27_c0 bl[0] br[0] wl[27] vdd gnd cell_6t
Xbit_r28_c0 bl[0] br[0] wl[28] vdd gnd cell_6t
Xbit_r29_c0 bl[0] br[0] wl[29] vdd gnd cell_6t
Xbit_r30_c0 bl[0] br[0] wl[30] vdd gnd cell_6t
Xbit_r31_c0 bl[0] br[0] wl[31] vdd gnd cell_6t
Xbit_r32_c0 bl[0] br[0] wl[32] vdd gnd cell_6t
Xbit_r33_c0 bl[0] br[0] wl[33] vdd gnd cell_6t
Xbit_r34_c0 bl[0] br[0] wl[34] vdd gnd cell_6t
Xbit_r35_c0 bl[0] br[0] wl[35] vdd gnd cell_6t
Xbit_r36_c0 bl[0] br[0] wl[36] vdd gnd cell_6t
Xbit_r37_c0 bl[0] br[0] wl[37] vdd gnd cell_6t
Xbit_r38_c0 bl[0] br[0] wl[38] vdd gnd cell_6t
Xbit_r39_c0 bl[0] br[0] wl[39] vdd gnd cell_6t
Xbit_r40_c0 bl[0] br[0] wl[40] vdd gnd cell_6t
Xbit_r41_c0 bl[0] br[0] wl[41] vdd gnd cell_6t
Xbit_r42_c0 bl[0] br[0] wl[42] vdd gnd cell_6t
Xbit_r43_c0 bl[0] br[0] wl[43] vdd gnd cell_6t
Xbit_r44_c0 bl[0] br[0] wl[44] vdd gnd cell_6t
Xbit_r45_c0 bl[0] br[0] wl[45] vdd gnd cell_6t
Xbit_r46_c0 bl[0] br[0] wl[46] vdd gnd cell_6t
Xbit_r47_c0 bl[0] br[0] wl[47] vdd gnd cell_6t
Xbit_r48_c0 bl[0] br[0] wl[48] vdd gnd cell_6t
Xbit_r49_c0 bl[0] br[0] wl[49] vdd gnd cell_6t
Xbit_r50_c0 bl[0] br[0] wl[50] vdd gnd cell_6t
Xbit_r51_c0 bl[0] br[0] wl[51] vdd gnd cell_6t
Xbit_r52_c0 bl[0] br[0] wl[52] vdd gnd cell_6t
Xbit_r53_c0 bl[0] br[0] wl[53] vdd gnd cell_6t
Xbit_r54_c0 bl[0] br[0] wl[54] vdd gnd cell_6t
Xbit_r55_c0 bl[0] br[0] wl[55] vdd gnd cell_6t
Xbit_r56_c0 bl[0] br[0] wl[56] vdd gnd cell_6t
Xbit_r57_c0 bl[0] br[0] wl[57] vdd gnd cell_6t
Xbit_r58_c0 bl[0] br[0] wl[58] vdd gnd cell_6t
Xbit_r59_c0 bl[0] br[0] wl[59] vdd gnd cell_6t
Xbit_r60_c0 bl[0] br[0] wl[60] vdd gnd cell_6t
Xbit_r61_c0 bl[0] br[0] wl[61] vdd gnd cell_6t
Xbit_r62_c0 bl[0] br[0] wl[62] vdd gnd cell_6t
Xbit_r63_c0 bl[0] br[0] wl[63] vdd gnd cell_6t
Xbit_r64_c0 bl[0] br[0] wl[64] vdd gnd cell_6t
Xbit_r65_c0 bl[0] br[0] wl[65] vdd gnd cell_6t
Xbit_r66_c0 bl[0] br[0] wl[66] vdd gnd cell_6t
Xbit_r67_c0 bl[0] br[0] wl[67] vdd gnd cell_6t
Xbit_r68_c0 bl[0] br[0] wl[68] vdd gnd cell_6t
Xbit_r69_c0 bl[0] br[0] wl[69] vdd gnd cell_6t
Xbit_r70_c0 bl[0] br[0] wl[70] vdd gnd cell_6t
Xbit_r71_c0 bl[0] br[0] wl[71] vdd gnd cell_6t
Xbit_r72_c0 bl[0] br[0] wl[72] vdd gnd cell_6t
Xbit_r73_c0 bl[0] br[0] wl[73] vdd gnd cell_6t
Xbit_r74_c0 bl[0] br[0] wl[74] vdd gnd cell_6t
Xbit_r75_c0 bl[0] br[0] wl[75] vdd gnd cell_6t
Xbit_r76_c0 bl[0] br[0] wl[76] vdd gnd cell_6t
Xbit_r77_c0 bl[0] br[0] wl[77] vdd gnd cell_6t
Xbit_r78_c0 bl[0] br[0] wl[78] vdd gnd cell_6t
Xbit_r79_c0 bl[0] br[0] wl[79] vdd gnd cell_6t
Xbit_r80_c0 bl[0] br[0] wl[80] vdd gnd cell_6t
Xbit_r81_c0 bl[0] br[0] wl[81] vdd gnd cell_6t
Xbit_r82_c0 bl[0] br[0] wl[82] vdd gnd cell_6t
Xbit_r83_c0 bl[0] br[0] wl[83] vdd gnd cell_6t
Xbit_r84_c0 bl[0] br[0] wl[84] vdd gnd cell_6t
Xbit_r85_c0 bl[0] br[0] wl[85] vdd gnd cell_6t
Xbit_r86_c0 bl[0] br[0] wl[86] vdd gnd cell_6t
Xbit_r87_c0 bl[0] br[0] wl[87] vdd gnd cell_6t
Xbit_r88_c0 bl[0] br[0] wl[88] vdd gnd cell_6t
Xbit_r89_c0 bl[0] br[0] wl[89] vdd gnd cell_6t
Xbit_r90_c0 bl[0] br[0] wl[90] vdd gnd cell_6t
Xbit_r91_c0 bl[0] br[0] wl[91] vdd gnd cell_6t
Xbit_r92_c0 bl[0] br[0] wl[92] vdd gnd cell_6t
Xbit_r93_c0 bl[0] br[0] wl[93] vdd gnd cell_6t
Xbit_r94_c0 bl[0] br[0] wl[94] vdd gnd cell_6t
Xbit_r95_c0 bl[0] br[0] wl[95] vdd gnd cell_6t
Xbit_r96_c0 bl[0] br[0] wl[96] vdd gnd cell_6t
Xbit_r97_c0 bl[0] br[0] wl[97] vdd gnd cell_6t
Xbit_r98_c0 bl[0] br[0] wl[98] vdd gnd cell_6t
Xbit_r99_c0 bl[0] br[0] wl[99] vdd gnd cell_6t
Xbit_r100_c0 bl[0] br[0] wl[100] vdd gnd cell_6t
Xbit_r101_c0 bl[0] br[0] wl[101] vdd gnd cell_6t
Xbit_r102_c0 bl[0] br[0] wl[102] vdd gnd cell_6t
Xbit_r103_c0 bl[0] br[0] wl[103] vdd gnd cell_6t
Xbit_r104_c0 bl[0] br[0] wl[104] vdd gnd cell_6t
Xbit_r105_c0 bl[0] br[0] wl[105] vdd gnd cell_6t
Xbit_r106_c0 bl[0] br[0] wl[106] vdd gnd cell_6t
Xbit_r107_c0 bl[0] br[0] wl[107] vdd gnd cell_6t
Xbit_r108_c0 bl[0] br[0] wl[108] vdd gnd cell_6t
Xbit_r109_c0 bl[0] br[0] wl[109] vdd gnd cell_6t
Xbit_r110_c0 bl[0] br[0] wl[110] vdd gnd cell_6t
Xbit_r111_c0 bl[0] br[0] wl[111] vdd gnd cell_6t
Xbit_r112_c0 bl[0] br[0] wl[112] vdd gnd cell_6t
Xbit_r113_c0 bl[0] br[0] wl[113] vdd gnd cell_6t
Xbit_r114_c0 bl[0] br[0] wl[114] vdd gnd cell_6t
Xbit_r115_c0 bl[0] br[0] wl[115] vdd gnd cell_6t
Xbit_r116_c0 bl[0] br[0] wl[116] vdd gnd cell_6t
Xbit_r117_c0 bl[0] br[0] wl[117] vdd gnd cell_6t
Xbit_r118_c0 bl[0] br[0] wl[118] vdd gnd cell_6t
Xbit_r119_c0 bl[0] br[0] wl[119] vdd gnd cell_6t
Xbit_r120_c0 bl[0] br[0] wl[120] vdd gnd cell_6t
Xbit_r121_c0 bl[0] br[0] wl[121] vdd gnd cell_6t
Xbit_r122_c0 bl[0] br[0] wl[122] vdd gnd cell_6t
Xbit_r123_c0 bl[0] br[0] wl[123] vdd gnd cell_6t
Xbit_r124_c0 bl[0] br[0] wl[124] vdd gnd cell_6t
Xbit_r125_c0 bl[0] br[0] wl[125] vdd gnd cell_6t
Xbit_r126_c0 bl[0] br[0] wl[126] vdd gnd cell_6t
Xbit_r127_c0 bl[0] br[0] wl[127] vdd gnd cell_6t
Xbit_r128_c0 bl[0] br[0] wl[128] vdd gnd cell_6t
Xbit_r129_c0 bl[0] br[0] wl[129] vdd gnd cell_6t
Xbit_r130_c0 bl[0] br[0] wl[130] vdd gnd cell_6t
Xbit_r131_c0 bl[0] br[0] wl[131] vdd gnd cell_6t
Xbit_r132_c0 bl[0] br[0] wl[132] vdd gnd cell_6t
Xbit_r133_c0 bl[0] br[0] wl[133] vdd gnd cell_6t
Xbit_r134_c0 bl[0] br[0] wl[134] vdd gnd cell_6t
Xbit_r135_c0 bl[0] br[0] wl[135] vdd gnd cell_6t
Xbit_r136_c0 bl[0] br[0] wl[136] vdd gnd cell_6t
Xbit_r137_c0 bl[0] br[0] wl[137] vdd gnd cell_6t
Xbit_r138_c0 bl[0] br[0] wl[138] vdd gnd cell_6t
Xbit_r139_c0 bl[0] br[0] wl[139] vdd gnd cell_6t
Xbit_r140_c0 bl[0] br[0] wl[140] vdd gnd cell_6t
Xbit_r141_c0 bl[0] br[0] wl[141] vdd gnd cell_6t
Xbit_r142_c0 bl[0] br[0] wl[142] vdd gnd cell_6t
Xbit_r143_c0 bl[0] br[0] wl[143] vdd gnd cell_6t
Xbit_r144_c0 bl[0] br[0] wl[144] vdd gnd cell_6t
Xbit_r145_c0 bl[0] br[0] wl[145] vdd gnd cell_6t
Xbit_r146_c0 bl[0] br[0] wl[146] vdd gnd cell_6t
Xbit_r147_c0 bl[0] br[0] wl[147] vdd gnd cell_6t
Xbit_r148_c0 bl[0] br[0] wl[148] vdd gnd cell_6t
Xbit_r149_c0 bl[0] br[0] wl[149] vdd gnd cell_6t
Xbit_r150_c0 bl[0] br[0] wl[150] vdd gnd cell_6t
Xbit_r151_c0 bl[0] br[0] wl[151] vdd gnd cell_6t
Xbit_r152_c0 bl[0] br[0] wl[152] vdd gnd cell_6t
Xbit_r153_c0 bl[0] br[0] wl[153] vdd gnd cell_6t
Xbit_r154_c0 bl[0] br[0] wl[154] vdd gnd cell_6t
Xbit_r155_c0 bl[0] br[0] wl[155] vdd gnd cell_6t
Xbit_r156_c0 bl[0] br[0] wl[156] vdd gnd cell_6t
Xbit_r157_c0 bl[0] br[0] wl[157] vdd gnd cell_6t
Xbit_r158_c0 bl[0] br[0] wl[158] vdd gnd cell_6t
Xbit_r159_c0 bl[0] br[0] wl[159] vdd gnd cell_6t
Xbit_r160_c0 bl[0] br[0] wl[160] vdd gnd cell_6t
Xbit_r161_c0 bl[0] br[0] wl[161] vdd gnd cell_6t
Xbit_r162_c0 bl[0] br[0] wl[162] vdd gnd cell_6t
Xbit_r163_c0 bl[0] br[0] wl[163] vdd gnd cell_6t
Xbit_r164_c0 bl[0] br[0] wl[164] vdd gnd cell_6t
Xbit_r165_c0 bl[0] br[0] wl[165] vdd gnd cell_6t
Xbit_r166_c0 bl[0] br[0] wl[166] vdd gnd cell_6t
Xbit_r167_c0 bl[0] br[0] wl[167] vdd gnd cell_6t
Xbit_r168_c0 bl[0] br[0] wl[168] vdd gnd cell_6t
Xbit_r169_c0 bl[0] br[0] wl[169] vdd gnd cell_6t
Xbit_r170_c0 bl[0] br[0] wl[170] vdd gnd cell_6t
Xbit_r171_c0 bl[0] br[0] wl[171] vdd gnd cell_6t
Xbit_r172_c0 bl[0] br[0] wl[172] vdd gnd cell_6t
Xbit_r173_c0 bl[0] br[0] wl[173] vdd gnd cell_6t
Xbit_r174_c0 bl[0] br[0] wl[174] vdd gnd cell_6t
Xbit_r175_c0 bl[0] br[0] wl[175] vdd gnd cell_6t
Xbit_r176_c0 bl[0] br[0] wl[176] vdd gnd cell_6t
Xbit_r177_c0 bl[0] br[0] wl[177] vdd gnd cell_6t
Xbit_r178_c0 bl[0] br[0] wl[178] vdd gnd cell_6t
Xbit_r179_c0 bl[0] br[0] wl[179] vdd gnd cell_6t
Xbit_r180_c0 bl[0] br[0] wl[180] vdd gnd cell_6t
Xbit_r181_c0 bl[0] br[0] wl[181] vdd gnd cell_6t
Xbit_r182_c0 bl[0] br[0] wl[182] vdd gnd cell_6t
Xbit_r183_c0 bl[0] br[0] wl[183] vdd gnd cell_6t
Xbit_r184_c0 bl[0] br[0] wl[184] vdd gnd cell_6t
Xbit_r185_c0 bl[0] br[0] wl[185] vdd gnd cell_6t
Xbit_r186_c0 bl[0] br[0] wl[186] vdd gnd cell_6t
Xbit_r187_c0 bl[0] br[0] wl[187] vdd gnd cell_6t
Xbit_r188_c0 bl[0] br[0] wl[188] vdd gnd cell_6t
Xbit_r189_c0 bl[0] br[0] wl[189] vdd gnd cell_6t
Xbit_r190_c0 bl[0] br[0] wl[190] vdd gnd cell_6t
Xbit_r191_c0 bl[0] br[0] wl[191] vdd gnd cell_6t
Xbit_r192_c0 bl[0] br[0] wl[192] vdd gnd cell_6t
Xbit_r193_c0 bl[0] br[0] wl[193] vdd gnd cell_6t
Xbit_r194_c0 bl[0] br[0] wl[194] vdd gnd cell_6t
Xbit_r195_c0 bl[0] br[0] wl[195] vdd gnd cell_6t
Xbit_r196_c0 bl[0] br[0] wl[196] vdd gnd cell_6t
Xbit_r197_c0 bl[0] br[0] wl[197] vdd gnd cell_6t
Xbit_r198_c0 bl[0] br[0] wl[198] vdd gnd cell_6t
Xbit_r199_c0 bl[0] br[0] wl[199] vdd gnd cell_6t
Xbit_r200_c0 bl[0] br[0] wl[200] vdd gnd cell_6t
Xbit_r201_c0 bl[0] br[0] wl[201] vdd gnd cell_6t
Xbit_r202_c0 bl[0] br[0] wl[202] vdd gnd cell_6t
Xbit_r203_c0 bl[0] br[0] wl[203] vdd gnd cell_6t
Xbit_r204_c0 bl[0] br[0] wl[204] vdd gnd cell_6t
Xbit_r205_c0 bl[0] br[0] wl[205] vdd gnd cell_6t
Xbit_r206_c0 bl[0] br[0] wl[206] vdd gnd cell_6t
Xbit_r207_c0 bl[0] br[0] wl[207] vdd gnd cell_6t
Xbit_r208_c0 bl[0] br[0] wl[208] vdd gnd cell_6t
Xbit_r209_c0 bl[0] br[0] wl[209] vdd gnd cell_6t
Xbit_r210_c0 bl[0] br[0] wl[210] vdd gnd cell_6t
Xbit_r211_c0 bl[0] br[0] wl[211] vdd gnd cell_6t
Xbit_r212_c0 bl[0] br[0] wl[212] vdd gnd cell_6t
Xbit_r213_c0 bl[0] br[0] wl[213] vdd gnd cell_6t
Xbit_r214_c0 bl[0] br[0] wl[214] vdd gnd cell_6t
Xbit_r215_c0 bl[0] br[0] wl[215] vdd gnd cell_6t
Xbit_r216_c0 bl[0] br[0] wl[216] vdd gnd cell_6t
Xbit_r217_c0 bl[0] br[0] wl[217] vdd gnd cell_6t
Xbit_r218_c0 bl[0] br[0] wl[218] vdd gnd cell_6t
Xbit_r219_c0 bl[0] br[0] wl[219] vdd gnd cell_6t
Xbit_r220_c0 bl[0] br[0] wl[220] vdd gnd cell_6t
Xbit_r221_c0 bl[0] br[0] wl[221] vdd gnd cell_6t
Xbit_r222_c0 bl[0] br[0] wl[222] vdd gnd cell_6t
Xbit_r223_c0 bl[0] br[0] wl[223] vdd gnd cell_6t
Xbit_r224_c0 bl[0] br[0] wl[224] vdd gnd cell_6t
Xbit_r225_c0 bl[0] br[0] wl[225] vdd gnd cell_6t
Xbit_r226_c0 bl[0] br[0] wl[226] vdd gnd cell_6t
Xbit_r227_c0 bl[0] br[0] wl[227] vdd gnd cell_6t
Xbit_r228_c0 bl[0] br[0] wl[228] vdd gnd cell_6t
Xbit_r229_c0 bl[0] br[0] wl[229] vdd gnd cell_6t
Xbit_r230_c0 bl[0] br[0] wl[230] vdd gnd cell_6t
Xbit_r231_c0 bl[0] br[0] wl[231] vdd gnd cell_6t
Xbit_r232_c0 bl[0] br[0] wl[232] vdd gnd cell_6t
Xbit_r233_c0 bl[0] br[0] wl[233] vdd gnd cell_6t
Xbit_r234_c0 bl[0] br[0] wl[234] vdd gnd cell_6t
Xbit_r235_c0 bl[0] br[0] wl[235] vdd gnd cell_6t
Xbit_r236_c0 bl[0] br[0] wl[236] vdd gnd cell_6t
Xbit_r237_c0 bl[0] br[0] wl[237] vdd gnd cell_6t
Xbit_r238_c0 bl[0] br[0] wl[238] vdd gnd cell_6t
Xbit_r239_c0 bl[0] br[0] wl[239] vdd gnd cell_6t
Xbit_r240_c0 bl[0] br[0] wl[240] vdd gnd cell_6t
Xbit_r241_c0 bl[0] br[0] wl[241] vdd gnd cell_6t
Xbit_r242_c0 bl[0] br[0] wl[242] vdd gnd cell_6t
Xbit_r243_c0 bl[0] br[0] wl[243] vdd gnd cell_6t
Xbit_r244_c0 bl[0] br[0] wl[244] vdd gnd cell_6t
Xbit_r245_c0 bl[0] br[0] wl[245] vdd gnd cell_6t
Xbit_r246_c0 bl[0] br[0] wl[246] vdd gnd cell_6t
Xbit_r247_c0 bl[0] br[0] wl[247] vdd gnd cell_6t
Xbit_r248_c0 bl[0] br[0] wl[248] vdd gnd cell_6t
Xbit_r249_c0 bl[0] br[0] wl[249] vdd gnd cell_6t
Xbit_r250_c0 bl[0] br[0] wl[250] vdd gnd cell_6t
Xbit_r251_c0 bl[0] br[0] wl[251] vdd gnd cell_6t
Xbit_r252_c0 bl[0] br[0] wl[252] vdd gnd cell_6t
Xbit_r253_c0 bl[0] br[0] wl[253] vdd gnd cell_6t
Xbit_r254_c0 bl[0] br[0] wl[254] vdd gnd cell_6t
Xbit_r255_c0 bl[0] br[0] wl[255] vdd gnd cell_6t
Xbit_r0_c1 bl[1] br[1] wl[0] vdd gnd cell_6t
Xbit_r1_c1 bl[1] br[1] wl[1] vdd gnd cell_6t
Xbit_r2_c1 bl[1] br[1] wl[2] vdd gnd cell_6t
Xbit_r3_c1 bl[1] br[1] wl[3] vdd gnd cell_6t
Xbit_r4_c1 bl[1] br[1] wl[4] vdd gnd cell_6t
Xbit_r5_c1 bl[1] br[1] wl[5] vdd gnd cell_6t
Xbit_r6_c1 bl[1] br[1] wl[6] vdd gnd cell_6t
Xbit_r7_c1 bl[1] br[1] wl[7] vdd gnd cell_6t
Xbit_r8_c1 bl[1] br[1] wl[8] vdd gnd cell_6t
Xbit_r9_c1 bl[1] br[1] wl[9] vdd gnd cell_6t
Xbit_r10_c1 bl[1] br[1] wl[10] vdd gnd cell_6t
Xbit_r11_c1 bl[1] br[1] wl[11] vdd gnd cell_6t
Xbit_r12_c1 bl[1] br[1] wl[12] vdd gnd cell_6t
Xbit_r13_c1 bl[1] br[1] wl[13] vdd gnd cell_6t
Xbit_r14_c1 bl[1] br[1] wl[14] vdd gnd cell_6t
Xbit_r15_c1 bl[1] br[1] wl[15] vdd gnd cell_6t
Xbit_r16_c1 bl[1] br[1] wl[16] vdd gnd cell_6t
Xbit_r17_c1 bl[1] br[1] wl[17] vdd gnd cell_6t
Xbit_r18_c1 bl[1] br[1] wl[18] vdd gnd cell_6t
Xbit_r19_c1 bl[1] br[1] wl[19] vdd gnd cell_6t
Xbit_r20_c1 bl[1] br[1] wl[20] vdd gnd cell_6t
Xbit_r21_c1 bl[1] br[1] wl[21] vdd gnd cell_6t
Xbit_r22_c1 bl[1] br[1] wl[22] vdd gnd cell_6t
Xbit_r23_c1 bl[1] br[1] wl[23] vdd gnd cell_6t
Xbit_r24_c1 bl[1] br[1] wl[24] vdd gnd cell_6t
Xbit_r25_c1 bl[1] br[1] wl[25] vdd gnd cell_6t
Xbit_r26_c1 bl[1] br[1] wl[26] vdd gnd cell_6t
Xbit_r27_c1 bl[1] br[1] wl[27] vdd gnd cell_6t
Xbit_r28_c1 bl[1] br[1] wl[28] vdd gnd cell_6t
Xbit_r29_c1 bl[1] br[1] wl[29] vdd gnd cell_6t
Xbit_r30_c1 bl[1] br[1] wl[30] vdd gnd cell_6t
Xbit_r31_c1 bl[1] br[1] wl[31] vdd gnd cell_6t
Xbit_r32_c1 bl[1] br[1] wl[32] vdd gnd cell_6t
Xbit_r33_c1 bl[1] br[1] wl[33] vdd gnd cell_6t
Xbit_r34_c1 bl[1] br[1] wl[34] vdd gnd cell_6t
Xbit_r35_c1 bl[1] br[1] wl[35] vdd gnd cell_6t
Xbit_r36_c1 bl[1] br[1] wl[36] vdd gnd cell_6t
Xbit_r37_c1 bl[1] br[1] wl[37] vdd gnd cell_6t
Xbit_r38_c1 bl[1] br[1] wl[38] vdd gnd cell_6t
Xbit_r39_c1 bl[1] br[1] wl[39] vdd gnd cell_6t
Xbit_r40_c1 bl[1] br[1] wl[40] vdd gnd cell_6t
Xbit_r41_c1 bl[1] br[1] wl[41] vdd gnd cell_6t
Xbit_r42_c1 bl[1] br[1] wl[42] vdd gnd cell_6t
Xbit_r43_c1 bl[1] br[1] wl[43] vdd gnd cell_6t
Xbit_r44_c1 bl[1] br[1] wl[44] vdd gnd cell_6t
Xbit_r45_c1 bl[1] br[1] wl[45] vdd gnd cell_6t
Xbit_r46_c1 bl[1] br[1] wl[46] vdd gnd cell_6t
Xbit_r47_c1 bl[1] br[1] wl[47] vdd gnd cell_6t
Xbit_r48_c1 bl[1] br[1] wl[48] vdd gnd cell_6t
Xbit_r49_c1 bl[1] br[1] wl[49] vdd gnd cell_6t
Xbit_r50_c1 bl[1] br[1] wl[50] vdd gnd cell_6t
Xbit_r51_c1 bl[1] br[1] wl[51] vdd gnd cell_6t
Xbit_r52_c1 bl[1] br[1] wl[52] vdd gnd cell_6t
Xbit_r53_c1 bl[1] br[1] wl[53] vdd gnd cell_6t
Xbit_r54_c1 bl[1] br[1] wl[54] vdd gnd cell_6t
Xbit_r55_c1 bl[1] br[1] wl[55] vdd gnd cell_6t
Xbit_r56_c1 bl[1] br[1] wl[56] vdd gnd cell_6t
Xbit_r57_c1 bl[1] br[1] wl[57] vdd gnd cell_6t
Xbit_r58_c1 bl[1] br[1] wl[58] vdd gnd cell_6t
Xbit_r59_c1 bl[1] br[1] wl[59] vdd gnd cell_6t
Xbit_r60_c1 bl[1] br[1] wl[60] vdd gnd cell_6t
Xbit_r61_c1 bl[1] br[1] wl[61] vdd gnd cell_6t
Xbit_r62_c1 bl[1] br[1] wl[62] vdd gnd cell_6t
Xbit_r63_c1 bl[1] br[1] wl[63] vdd gnd cell_6t
Xbit_r64_c1 bl[1] br[1] wl[64] vdd gnd cell_6t
Xbit_r65_c1 bl[1] br[1] wl[65] vdd gnd cell_6t
Xbit_r66_c1 bl[1] br[1] wl[66] vdd gnd cell_6t
Xbit_r67_c1 bl[1] br[1] wl[67] vdd gnd cell_6t
Xbit_r68_c1 bl[1] br[1] wl[68] vdd gnd cell_6t
Xbit_r69_c1 bl[1] br[1] wl[69] vdd gnd cell_6t
Xbit_r70_c1 bl[1] br[1] wl[70] vdd gnd cell_6t
Xbit_r71_c1 bl[1] br[1] wl[71] vdd gnd cell_6t
Xbit_r72_c1 bl[1] br[1] wl[72] vdd gnd cell_6t
Xbit_r73_c1 bl[1] br[1] wl[73] vdd gnd cell_6t
Xbit_r74_c1 bl[1] br[1] wl[74] vdd gnd cell_6t
Xbit_r75_c1 bl[1] br[1] wl[75] vdd gnd cell_6t
Xbit_r76_c1 bl[1] br[1] wl[76] vdd gnd cell_6t
Xbit_r77_c1 bl[1] br[1] wl[77] vdd gnd cell_6t
Xbit_r78_c1 bl[1] br[1] wl[78] vdd gnd cell_6t
Xbit_r79_c1 bl[1] br[1] wl[79] vdd gnd cell_6t
Xbit_r80_c1 bl[1] br[1] wl[80] vdd gnd cell_6t
Xbit_r81_c1 bl[1] br[1] wl[81] vdd gnd cell_6t
Xbit_r82_c1 bl[1] br[1] wl[82] vdd gnd cell_6t
Xbit_r83_c1 bl[1] br[1] wl[83] vdd gnd cell_6t
Xbit_r84_c1 bl[1] br[1] wl[84] vdd gnd cell_6t
Xbit_r85_c1 bl[1] br[1] wl[85] vdd gnd cell_6t
Xbit_r86_c1 bl[1] br[1] wl[86] vdd gnd cell_6t
Xbit_r87_c1 bl[1] br[1] wl[87] vdd gnd cell_6t
Xbit_r88_c1 bl[1] br[1] wl[88] vdd gnd cell_6t
Xbit_r89_c1 bl[1] br[1] wl[89] vdd gnd cell_6t
Xbit_r90_c1 bl[1] br[1] wl[90] vdd gnd cell_6t
Xbit_r91_c1 bl[1] br[1] wl[91] vdd gnd cell_6t
Xbit_r92_c1 bl[1] br[1] wl[92] vdd gnd cell_6t
Xbit_r93_c1 bl[1] br[1] wl[93] vdd gnd cell_6t
Xbit_r94_c1 bl[1] br[1] wl[94] vdd gnd cell_6t
Xbit_r95_c1 bl[1] br[1] wl[95] vdd gnd cell_6t
Xbit_r96_c1 bl[1] br[1] wl[96] vdd gnd cell_6t
Xbit_r97_c1 bl[1] br[1] wl[97] vdd gnd cell_6t
Xbit_r98_c1 bl[1] br[1] wl[98] vdd gnd cell_6t
Xbit_r99_c1 bl[1] br[1] wl[99] vdd gnd cell_6t
Xbit_r100_c1 bl[1] br[1] wl[100] vdd gnd cell_6t
Xbit_r101_c1 bl[1] br[1] wl[101] vdd gnd cell_6t
Xbit_r102_c1 bl[1] br[1] wl[102] vdd gnd cell_6t
Xbit_r103_c1 bl[1] br[1] wl[103] vdd gnd cell_6t
Xbit_r104_c1 bl[1] br[1] wl[104] vdd gnd cell_6t
Xbit_r105_c1 bl[1] br[1] wl[105] vdd gnd cell_6t
Xbit_r106_c1 bl[1] br[1] wl[106] vdd gnd cell_6t
Xbit_r107_c1 bl[1] br[1] wl[107] vdd gnd cell_6t
Xbit_r108_c1 bl[1] br[1] wl[108] vdd gnd cell_6t
Xbit_r109_c1 bl[1] br[1] wl[109] vdd gnd cell_6t
Xbit_r110_c1 bl[1] br[1] wl[110] vdd gnd cell_6t
Xbit_r111_c1 bl[1] br[1] wl[111] vdd gnd cell_6t
Xbit_r112_c1 bl[1] br[1] wl[112] vdd gnd cell_6t
Xbit_r113_c1 bl[1] br[1] wl[113] vdd gnd cell_6t
Xbit_r114_c1 bl[1] br[1] wl[114] vdd gnd cell_6t
Xbit_r115_c1 bl[1] br[1] wl[115] vdd gnd cell_6t
Xbit_r116_c1 bl[1] br[1] wl[116] vdd gnd cell_6t
Xbit_r117_c1 bl[1] br[1] wl[117] vdd gnd cell_6t
Xbit_r118_c1 bl[1] br[1] wl[118] vdd gnd cell_6t
Xbit_r119_c1 bl[1] br[1] wl[119] vdd gnd cell_6t
Xbit_r120_c1 bl[1] br[1] wl[120] vdd gnd cell_6t
Xbit_r121_c1 bl[1] br[1] wl[121] vdd gnd cell_6t
Xbit_r122_c1 bl[1] br[1] wl[122] vdd gnd cell_6t
Xbit_r123_c1 bl[1] br[1] wl[123] vdd gnd cell_6t
Xbit_r124_c1 bl[1] br[1] wl[124] vdd gnd cell_6t
Xbit_r125_c1 bl[1] br[1] wl[125] vdd gnd cell_6t
Xbit_r126_c1 bl[1] br[1] wl[126] vdd gnd cell_6t
Xbit_r127_c1 bl[1] br[1] wl[127] vdd gnd cell_6t
Xbit_r128_c1 bl[1] br[1] wl[128] vdd gnd cell_6t
Xbit_r129_c1 bl[1] br[1] wl[129] vdd gnd cell_6t
Xbit_r130_c1 bl[1] br[1] wl[130] vdd gnd cell_6t
Xbit_r131_c1 bl[1] br[1] wl[131] vdd gnd cell_6t
Xbit_r132_c1 bl[1] br[1] wl[132] vdd gnd cell_6t
Xbit_r133_c1 bl[1] br[1] wl[133] vdd gnd cell_6t
Xbit_r134_c1 bl[1] br[1] wl[134] vdd gnd cell_6t
Xbit_r135_c1 bl[1] br[1] wl[135] vdd gnd cell_6t
Xbit_r136_c1 bl[1] br[1] wl[136] vdd gnd cell_6t
Xbit_r137_c1 bl[1] br[1] wl[137] vdd gnd cell_6t
Xbit_r138_c1 bl[1] br[1] wl[138] vdd gnd cell_6t
Xbit_r139_c1 bl[1] br[1] wl[139] vdd gnd cell_6t
Xbit_r140_c1 bl[1] br[1] wl[140] vdd gnd cell_6t
Xbit_r141_c1 bl[1] br[1] wl[141] vdd gnd cell_6t
Xbit_r142_c1 bl[1] br[1] wl[142] vdd gnd cell_6t
Xbit_r143_c1 bl[1] br[1] wl[143] vdd gnd cell_6t
Xbit_r144_c1 bl[1] br[1] wl[144] vdd gnd cell_6t
Xbit_r145_c1 bl[1] br[1] wl[145] vdd gnd cell_6t
Xbit_r146_c1 bl[1] br[1] wl[146] vdd gnd cell_6t
Xbit_r147_c1 bl[1] br[1] wl[147] vdd gnd cell_6t
Xbit_r148_c1 bl[1] br[1] wl[148] vdd gnd cell_6t
Xbit_r149_c1 bl[1] br[1] wl[149] vdd gnd cell_6t
Xbit_r150_c1 bl[1] br[1] wl[150] vdd gnd cell_6t
Xbit_r151_c1 bl[1] br[1] wl[151] vdd gnd cell_6t
Xbit_r152_c1 bl[1] br[1] wl[152] vdd gnd cell_6t
Xbit_r153_c1 bl[1] br[1] wl[153] vdd gnd cell_6t
Xbit_r154_c1 bl[1] br[1] wl[154] vdd gnd cell_6t
Xbit_r155_c1 bl[1] br[1] wl[155] vdd gnd cell_6t
Xbit_r156_c1 bl[1] br[1] wl[156] vdd gnd cell_6t
Xbit_r157_c1 bl[1] br[1] wl[157] vdd gnd cell_6t
Xbit_r158_c1 bl[1] br[1] wl[158] vdd gnd cell_6t
Xbit_r159_c1 bl[1] br[1] wl[159] vdd gnd cell_6t
Xbit_r160_c1 bl[1] br[1] wl[160] vdd gnd cell_6t
Xbit_r161_c1 bl[1] br[1] wl[161] vdd gnd cell_6t
Xbit_r162_c1 bl[1] br[1] wl[162] vdd gnd cell_6t
Xbit_r163_c1 bl[1] br[1] wl[163] vdd gnd cell_6t
Xbit_r164_c1 bl[1] br[1] wl[164] vdd gnd cell_6t
Xbit_r165_c1 bl[1] br[1] wl[165] vdd gnd cell_6t
Xbit_r166_c1 bl[1] br[1] wl[166] vdd gnd cell_6t
Xbit_r167_c1 bl[1] br[1] wl[167] vdd gnd cell_6t
Xbit_r168_c1 bl[1] br[1] wl[168] vdd gnd cell_6t
Xbit_r169_c1 bl[1] br[1] wl[169] vdd gnd cell_6t
Xbit_r170_c1 bl[1] br[1] wl[170] vdd gnd cell_6t
Xbit_r171_c1 bl[1] br[1] wl[171] vdd gnd cell_6t
Xbit_r172_c1 bl[1] br[1] wl[172] vdd gnd cell_6t
Xbit_r173_c1 bl[1] br[1] wl[173] vdd gnd cell_6t
Xbit_r174_c1 bl[1] br[1] wl[174] vdd gnd cell_6t
Xbit_r175_c1 bl[1] br[1] wl[175] vdd gnd cell_6t
Xbit_r176_c1 bl[1] br[1] wl[176] vdd gnd cell_6t
Xbit_r177_c1 bl[1] br[1] wl[177] vdd gnd cell_6t
Xbit_r178_c1 bl[1] br[1] wl[178] vdd gnd cell_6t
Xbit_r179_c1 bl[1] br[1] wl[179] vdd gnd cell_6t
Xbit_r180_c1 bl[1] br[1] wl[180] vdd gnd cell_6t
Xbit_r181_c1 bl[1] br[1] wl[181] vdd gnd cell_6t
Xbit_r182_c1 bl[1] br[1] wl[182] vdd gnd cell_6t
Xbit_r183_c1 bl[1] br[1] wl[183] vdd gnd cell_6t
Xbit_r184_c1 bl[1] br[1] wl[184] vdd gnd cell_6t
Xbit_r185_c1 bl[1] br[1] wl[185] vdd gnd cell_6t
Xbit_r186_c1 bl[1] br[1] wl[186] vdd gnd cell_6t
Xbit_r187_c1 bl[1] br[1] wl[187] vdd gnd cell_6t
Xbit_r188_c1 bl[1] br[1] wl[188] vdd gnd cell_6t
Xbit_r189_c1 bl[1] br[1] wl[189] vdd gnd cell_6t
Xbit_r190_c1 bl[1] br[1] wl[190] vdd gnd cell_6t
Xbit_r191_c1 bl[1] br[1] wl[191] vdd gnd cell_6t
Xbit_r192_c1 bl[1] br[1] wl[192] vdd gnd cell_6t
Xbit_r193_c1 bl[1] br[1] wl[193] vdd gnd cell_6t
Xbit_r194_c1 bl[1] br[1] wl[194] vdd gnd cell_6t
Xbit_r195_c1 bl[1] br[1] wl[195] vdd gnd cell_6t
Xbit_r196_c1 bl[1] br[1] wl[196] vdd gnd cell_6t
Xbit_r197_c1 bl[1] br[1] wl[197] vdd gnd cell_6t
Xbit_r198_c1 bl[1] br[1] wl[198] vdd gnd cell_6t
Xbit_r199_c1 bl[1] br[1] wl[199] vdd gnd cell_6t
Xbit_r200_c1 bl[1] br[1] wl[200] vdd gnd cell_6t
Xbit_r201_c1 bl[1] br[1] wl[201] vdd gnd cell_6t
Xbit_r202_c1 bl[1] br[1] wl[202] vdd gnd cell_6t
Xbit_r203_c1 bl[1] br[1] wl[203] vdd gnd cell_6t
Xbit_r204_c1 bl[1] br[1] wl[204] vdd gnd cell_6t
Xbit_r205_c1 bl[1] br[1] wl[205] vdd gnd cell_6t
Xbit_r206_c1 bl[1] br[1] wl[206] vdd gnd cell_6t
Xbit_r207_c1 bl[1] br[1] wl[207] vdd gnd cell_6t
Xbit_r208_c1 bl[1] br[1] wl[208] vdd gnd cell_6t
Xbit_r209_c1 bl[1] br[1] wl[209] vdd gnd cell_6t
Xbit_r210_c1 bl[1] br[1] wl[210] vdd gnd cell_6t
Xbit_r211_c1 bl[1] br[1] wl[211] vdd gnd cell_6t
Xbit_r212_c1 bl[1] br[1] wl[212] vdd gnd cell_6t
Xbit_r213_c1 bl[1] br[1] wl[213] vdd gnd cell_6t
Xbit_r214_c1 bl[1] br[1] wl[214] vdd gnd cell_6t
Xbit_r215_c1 bl[1] br[1] wl[215] vdd gnd cell_6t
Xbit_r216_c1 bl[1] br[1] wl[216] vdd gnd cell_6t
Xbit_r217_c1 bl[1] br[1] wl[217] vdd gnd cell_6t
Xbit_r218_c1 bl[1] br[1] wl[218] vdd gnd cell_6t
Xbit_r219_c1 bl[1] br[1] wl[219] vdd gnd cell_6t
Xbit_r220_c1 bl[1] br[1] wl[220] vdd gnd cell_6t
Xbit_r221_c1 bl[1] br[1] wl[221] vdd gnd cell_6t
Xbit_r222_c1 bl[1] br[1] wl[222] vdd gnd cell_6t
Xbit_r223_c1 bl[1] br[1] wl[223] vdd gnd cell_6t
Xbit_r224_c1 bl[1] br[1] wl[224] vdd gnd cell_6t
Xbit_r225_c1 bl[1] br[1] wl[225] vdd gnd cell_6t
Xbit_r226_c1 bl[1] br[1] wl[226] vdd gnd cell_6t
Xbit_r227_c1 bl[1] br[1] wl[227] vdd gnd cell_6t
Xbit_r228_c1 bl[1] br[1] wl[228] vdd gnd cell_6t
Xbit_r229_c1 bl[1] br[1] wl[229] vdd gnd cell_6t
Xbit_r230_c1 bl[1] br[1] wl[230] vdd gnd cell_6t
Xbit_r231_c1 bl[1] br[1] wl[231] vdd gnd cell_6t
Xbit_r232_c1 bl[1] br[1] wl[232] vdd gnd cell_6t
Xbit_r233_c1 bl[1] br[1] wl[233] vdd gnd cell_6t
Xbit_r234_c1 bl[1] br[1] wl[234] vdd gnd cell_6t
Xbit_r235_c1 bl[1] br[1] wl[235] vdd gnd cell_6t
Xbit_r236_c1 bl[1] br[1] wl[236] vdd gnd cell_6t
Xbit_r237_c1 bl[1] br[1] wl[237] vdd gnd cell_6t
Xbit_r238_c1 bl[1] br[1] wl[238] vdd gnd cell_6t
Xbit_r239_c1 bl[1] br[1] wl[239] vdd gnd cell_6t
Xbit_r240_c1 bl[1] br[1] wl[240] vdd gnd cell_6t
Xbit_r241_c1 bl[1] br[1] wl[241] vdd gnd cell_6t
Xbit_r242_c1 bl[1] br[1] wl[242] vdd gnd cell_6t
Xbit_r243_c1 bl[1] br[1] wl[243] vdd gnd cell_6t
Xbit_r244_c1 bl[1] br[1] wl[244] vdd gnd cell_6t
Xbit_r245_c1 bl[1] br[1] wl[245] vdd gnd cell_6t
Xbit_r246_c1 bl[1] br[1] wl[246] vdd gnd cell_6t
Xbit_r247_c1 bl[1] br[1] wl[247] vdd gnd cell_6t
Xbit_r248_c1 bl[1] br[1] wl[248] vdd gnd cell_6t
Xbit_r249_c1 bl[1] br[1] wl[249] vdd gnd cell_6t
Xbit_r250_c1 bl[1] br[1] wl[250] vdd gnd cell_6t
Xbit_r251_c1 bl[1] br[1] wl[251] vdd gnd cell_6t
Xbit_r252_c1 bl[1] br[1] wl[252] vdd gnd cell_6t
Xbit_r253_c1 bl[1] br[1] wl[253] vdd gnd cell_6t
Xbit_r254_c1 bl[1] br[1] wl[254] vdd gnd cell_6t
Xbit_r255_c1 bl[1] br[1] wl[255] vdd gnd cell_6t
Xbit_r0_c2 bl[2] br[2] wl[0] vdd gnd cell_6t
Xbit_r1_c2 bl[2] br[2] wl[1] vdd gnd cell_6t
Xbit_r2_c2 bl[2] br[2] wl[2] vdd gnd cell_6t
Xbit_r3_c2 bl[2] br[2] wl[3] vdd gnd cell_6t
Xbit_r4_c2 bl[2] br[2] wl[4] vdd gnd cell_6t
Xbit_r5_c2 bl[2] br[2] wl[5] vdd gnd cell_6t
Xbit_r6_c2 bl[2] br[2] wl[6] vdd gnd cell_6t
Xbit_r7_c2 bl[2] br[2] wl[7] vdd gnd cell_6t
Xbit_r8_c2 bl[2] br[2] wl[8] vdd gnd cell_6t
Xbit_r9_c2 bl[2] br[2] wl[9] vdd gnd cell_6t
Xbit_r10_c2 bl[2] br[2] wl[10] vdd gnd cell_6t
Xbit_r11_c2 bl[2] br[2] wl[11] vdd gnd cell_6t
Xbit_r12_c2 bl[2] br[2] wl[12] vdd gnd cell_6t
Xbit_r13_c2 bl[2] br[2] wl[13] vdd gnd cell_6t
Xbit_r14_c2 bl[2] br[2] wl[14] vdd gnd cell_6t
Xbit_r15_c2 bl[2] br[2] wl[15] vdd gnd cell_6t
Xbit_r16_c2 bl[2] br[2] wl[16] vdd gnd cell_6t
Xbit_r17_c2 bl[2] br[2] wl[17] vdd gnd cell_6t
Xbit_r18_c2 bl[2] br[2] wl[18] vdd gnd cell_6t
Xbit_r19_c2 bl[2] br[2] wl[19] vdd gnd cell_6t
Xbit_r20_c2 bl[2] br[2] wl[20] vdd gnd cell_6t
Xbit_r21_c2 bl[2] br[2] wl[21] vdd gnd cell_6t
Xbit_r22_c2 bl[2] br[2] wl[22] vdd gnd cell_6t
Xbit_r23_c2 bl[2] br[2] wl[23] vdd gnd cell_6t
Xbit_r24_c2 bl[2] br[2] wl[24] vdd gnd cell_6t
Xbit_r25_c2 bl[2] br[2] wl[25] vdd gnd cell_6t
Xbit_r26_c2 bl[2] br[2] wl[26] vdd gnd cell_6t
Xbit_r27_c2 bl[2] br[2] wl[27] vdd gnd cell_6t
Xbit_r28_c2 bl[2] br[2] wl[28] vdd gnd cell_6t
Xbit_r29_c2 bl[2] br[2] wl[29] vdd gnd cell_6t
Xbit_r30_c2 bl[2] br[2] wl[30] vdd gnd cell_6t
Xbit_r31_c2 bl[2] br[2] wl[31] vdd gnd cell_6t
Xbit_r32_c2 bl[2] br[2] wl[32] vdd gnd cell_6t
Xbit_r33_c2 bl[2] br[2] wl[33] vdd gnd cell_6t
Xbit_r34_c2 bl[2] br[2] wl[34] vdd gnd cell_6t
Xbit_r35_c2 bl[2] br[2] wl[35] vdd gnd cell_6t
Xbit_r36_c2 bl[2] br[2] wl[36] vdd gnd cell_6t
Xbit_r37_c2 bl[2] br[2] wl[37] vdd gnd cell_6t
Xbit_r38_c2 bl[2] br[2] wl[38] vdd gnd cell_6t
Xbit_r39_c2 bl[2] br[2] wl[39] vdd gnd cell_6t
Xbit_r40_c2 bl[2] br[2] wl[40] vdd gnd cell_6t
Xbit_r41_c2 bl[2] br[2] wl[41] vdd gnd cell_6t
Xbit_r42_c2 bl[2] br[2] wl[42] vdd gnd cell_6t
Xbit_r43_c2 bl[2] br[2] wl[43] vdd gnd cell_6t
Xbit_r44_c2 bl[2] br[2] wl[44] vdd gnd cell_6t
Xbit_r45_c2 bl[2] br[2] wl[45] vdd gnd cell_6t
Xbit_r46_c2 bl[2] br[2] wl[46] vdd gnd cell_6t
Xbit_r47_c2 bl[2] br[2] wl[47] vdd gnd cell_6t
Xbit_r48_c2 bl[2] br[2] wl[48] vdd gnd cell_6t
Xbit_r49_c2 bl[2] br[2] wl[49] vdd gnd cell_6t
Xbit_r50_c2 bl[2] br[2] wl[50] vdd gnd cell_6t
Xbit_r51_c2 bl[2] br[2] wl[51] vdd gnd cell_6t
Xbit_r52_c2 bl[2] br[2] wl[52] vdd gnd cell_6t
Xbit_r53_c2 bl[2] br[2] wl[53] vdd gnd cell_6t
Xbit_r54_c2 bl[2] br[2] wl[54] vdd gnd cell_6t
Xbit_r55_c2 bl[2] br[2] wl[55] vdd gnd cell_6t
Xbit_r56_c2 bl[2] br[2] wl[56] vdd gnd cell_6t
Xbit_r57_c2 bl[2] br[2] wl[57] vdd gnd cell_6t
Xbit_r58_c2 bl[2] br[2] wl[58] vdd gnd cell_6t
Xbit_r59_c2 bl[2] br[2] wl[59] vdd gnd cell_6t
Xbit_r60_c2 bl[2] br[2] wl[60] vdd gnd cell_6t
Xbit_r61_c2 bl[2] br[2] wl[61] vdd gnd cell_6t
Xbit_r62_c2 bl[2] br[2] wl[62] vdd gnd cell_6t
Xbit_r63_c2 bl[2] br[2] wl[63] vdd gnd cell_6t
Xbit_r64_c2 bl[2] br[2] wl[64] vdd gnd cell_6t
Xbit_r65_c2 bl[2] br[2] wl[65] vdd gnd cell_6t
Xbit_r66_c2 bl[2] br[2] wl[66] vdd gnd cell_6t
Xbit_r67_c2 bl[2] br[2] wl[67] vdd gnd cell_6t
Xbit_r68_c2 bl[2] br[2] wl[68] vdd gnd cell_6t
Xbit_r69_c2 bl[2] br[2] wl[69] vdd gnd cell_6t
Xbit_r70_c2 bl[2] br[2] wl[70] vdd gnd cell_6t
Xbit_r71_c2 bl[2] br[2] wl[71] vdd gnd cell_6t
Xbit_r72_c2 bl[2] br[2] wl[72] vdd gnd cell_6t
Xbit_r73_c2 bl[2] br[2] wl[73] vdd gnd cell_6t
Xbit_r74_c2 bl[2] br[2] wl[74] vdd gnd cell_6t
Xbit_r75_c2 bl[2] br[2] wl[75] vdd gnd cell_6t
Xbit_r76_c2 bl[2] br[2] wl[76] vdd gnd cell_6t
Xbit_r77_c2 bl[2] br[2] wl[77] vdd gnd cell_6t
Xbit_r78_c2 bl[2] br[2] wl[78] vdd gnd cell_6t
Xbit_r79_c2 bl[2] br[2] wl[79] vdd gnd cell_6t
Xbit_r80_c2 bl[2] br[2] wl[80] vdd gnd cell_6t
Xbit_r81_c2 bl[2] br[2] wl[81] vdd gnd cell_6t
Xbit_r82_c2 bl[2] br[2] wl[82] vdd gnd cell_6t
Xbit_r83_c2 bl[2] br[2] wl[83] vdd gnd cell_6t
Xbit_r84_c2 bl[2] br[2] wl[84] vdd gnd cell_6t
Xbit_r85_c2 bl[2] br[2] wl[85] vdd gnd cell_6t
Xbit_r86_c2 bl[2] br[2] wl[86] vdd gnd cell_6t
Xbit_r87_c2 bl[2] br[2] wl[87] vdd gnd cell_6t
Xbit_r88_c2 bl[2] br[2] wl[88] vdd gnd cell_6t
Xbit_r89_c2 bl[2] br[2] wl[89] vdd gnd cell_6t
Xbit_r90_c2 bl[2] br[2] wl[90] vdd gnd cell_6t
Xbit_r91_c2 bl[2] br[2] wl[91] vdd gnd cell_6t
Xbit_r92_c2 bl[2] br[2] wl[92] vdd gnd cell_6t
Xbit_r93_c2 bl[2] br[2] wl[93] vdd gnd cell_6t
Xbit_r94_c2 bl[2] br[2] wl[94] vdd gnd cell_6t
Xbit_r95_c2 bl[2] br[2] wl[95] vdd gnd cell_6t
Xbit_r96_c2 bl[2] br[2] wl[96] vdd gnd cell_6t
Xbit_r97_c2 bl[2] br[2] wl[97] vdd gnd cell_6t
Xbit_r98_c2 bl[2] br[2] wl[98] vdd gnd cell_6t
Xbit_r99_c2 bl[2] br[2] wl[99] vdd gnd cell_6t
Xbit_r100_c2 bl[2] br[2] wl[100] vdd gnd cell_6t
Xbit_r101_c2 bl[2] br[2] wl[101] vdd gnd cell_6t
Xbit_r102_c2 bl[2] br[2] wl[102] vdd gnd cell_6t
Xbit_r103_c2 bl[2] br[2] wl[103] vdd gnd cell_6t
Xbit_r104_c2 bl[2] br[2] wl[104] vdd gnd cell_6t
Xbit_r105_c2 bl[2] br[2] wl[105] vdd gnd cell_6t
Xbit_r106_c2 bl[2] br[2] wl[106] vdd gnd cell_6t
Xbit_r107_c2 bl[2] br[2] wl[107] vdd gnd cell_6t
Xbit_r108_c2 bl[2] br[2] wl[108] vdd gnd cell_6t
Xbit_r109_c2 bl[2] br[2] wl[109] vdd gnd cell_6t
Xbit_r110_c2 bl[2] br[2] wl[110] vdd gnd cell_6t
Xbit_r111_c2 bl[2] br[2] wl[111] vdd gnd cell_6t
Xbit_r112_c2 bl[2] br[2] wl[112] vdd gnd cell_6t
Xbit_r113_c2 bl[2] br[2] wl[113] vdd gnd cell_6t
Xbit_r114_c2 bl[2] br[2] wl[114] vdd gnd cell_6t
Xbit_r115_c2 bl[2] br[2] wl[115] vdd gnd cell_6t
Xbit_r116_c2 bl[2] br[2] wl[116] vdd gnd cell_6t
Xbit_r117_c2 bl[2] br[2] wl[117] vdd gnd cell_6t
Xbit_r118_c2 bl[2] br[2] wl[118] vdd gnd cell_6t
Xbit_r119_c2 bl[2] br[2] wl[119] vdd gnd cell_6t
Xbit_r120_c2 bl[2] br[2] wl[120] vdd gnd cell_6t
Xbit_r121_c2 bl[2] br[2] wl[121] vdd gnd cell_6t
Xbit_r122_c2 bl[2] br[2] wl[122] vdd gnd cell_6t
Xbit_r123_c2 bl[2] br[2] wl[123] vdd gnd cell_6t
Xbit_r124_c2 bl[2] br[2] wl[124] vdd gnd cell_6t
Xbit_r125_c2 bl[2] br[2] wl[125] vdd gnd cell_6t
Xbit_r126_c2 bl[2] br[2] wl[126] vdd gnd cell_6t
Xbit_r127_c2 bl[2] br[2] wl[127] vdd gnd cell_6t
Xbit_r128_c2 bl[2] br[2] wl[128] vdd gnd cell_6t
Xbit_r129_c2 bl[2] br[2] wl[129] vdd gnd cell_6t
Xbit_r130_c2 bl[2] br[2] wl[130] vdd gnd cell_6t
Xbit_r131_c2 bl[2] br[2] wl[131] vdd gnd cell_6t
Xbit_r132_c2 bl[2] br[2] wl[132] vdd gnd cell_6t
Xbit_r133_c2 bl[2] br[2] wl[133] vdd gnd cell_6t
Xbit_r134_c2 bl[2] br[2] wl[134] vdd gnd cell_6t
Xbit_r135_c2 bl[2] br[2] wl[135] vdd gnd cell_6t
Xbit_r136_c2 bl[2] br[2] wl[136] vdd gnd cell_6t
Xbit_r137_c2 bl[2] br[2] wl[137] vdd gnd cell_6t
Xbit_r138_c2 bl[2] br[2] wl[138] vdd gnd cell_6t
Xbit_r139_c2 bl[2] br[2] wl[139] vdd gnd cell_6t
Xbit_r140_c2 bl[2] br[2] wl[140] vdd gnd cell_6t
Xbit_r141_c2 bl[2] br[2] wl[141] vdd gnd cell_6t
Xbit_r142_c2 bl[2] br[2] wl[142] vdd gnd cell_6t
Xbit_r143_c2 bl[2] br[2] wl[143] vdd gnd cell_6t
Xbit_r144_c2 bl[2] br[2] wl[144] vdd gnd cell_6t
Xbit_r145_c2 bl[2] br[2] wl[145] vdd gnd cell_6t
Xbit_r146_c2 bl[2] br[2] wl[146] vdd gnd cell_6t
Xbit_r147_c2 bl[2] br[2] wl[147] vdd gnd cell_6t
Xbit_r148_c2 bl[2] br[2] wl[148] vdd gnd cell_6t
Xbit_r149_c2 bl[2] br[2] wl[149] vdd gnd cell_6t
Xbit_r150_c2 bl[2] br[2] wl[150] vdd gnd cell_6t
Xbit_r151_c2 bl[2] br[2] wl[151] vdd gnd cell_6t
Xbit_r152_c2 bl[2] br[2] wl[152] vdd gnd cell_6t
Xbit_r153_c2 bl[2] br[2] wl[153] vdd gnd cell_6t
Xbit_r154_c2 bl[2] br[2] wl[154] vdd gnd cell_6t
Xbit_r155_c2 bl[2] br[2] wl[155] vdd gnd cell_6t
Xbit_r156_c2 bl[2] br[2] wl[156] vdd gnd cell_6t
Xbit_r157_c2 bl[2] br[2] wl[157] vdd gnd cell_6t
Xbit_r158_c2 bl[2] br[2] wl[158] vdd gnd cell_6t
Xbit_r159_c2 bl[2] br[2] wl[159] vdd gnd cell_6t
Xbit_r160_c2 bl[2] br[2] wl[160] vdd gnd cell_6t
Xbit_r161_c2 bl[2] br[2] wl[161] vdd gnd cell_6t
Xbit_r162_c2 bl[2] br[2] wl[162] vdd gnd cell_6t
Xbit_r163_c2 bl[2] br[2] wl[163] vdd gnd cell_6t
Xbit_r164_c2 bl[2] br[2] wl[164] vdd gnd cell_6t
Xbit_r165_c2 bl[2] br[2] wl[165] vdd gnd cell_6t
Xbit_r166_c2 bl[2] br[2] wl[166] vdd gnd cell_6t
Xbit_r167_c2 bl[2] br[2] wl[167] vdd gnd cell_6t
Xbit_r168_c2 bl[2] br[2] wl[168] vdd gnd cell_6t
Xbit_r169_c2 bl[2] br[2] wl[169] vdd gnd cell_6t
Xbit_r170_c2 bl[2] br[2] wl[170] vdd gnd cell_6t
Xbit_r171_c2 bl[2] br[2] wl[171] vdd gnd cell_6t
Xbit_r172_c2 bl[2] br[2] wl[172] vdd gnd cell_6t
Xbit_r173_c2 bl[2] br[2] wl[173] vdd gnd cell_6t
Xbit_r174_c2 bl[2] br[2] wl[174] vdd gnd cell_6t
Xbit_r175_c2 bl[2] br[2] wl[175] vdd gnd cell_6t
Xbit_r176_c2 bl[2] br[2] wl[176] vdd gnd cell_6t
Xbit_r177_c2 bl[2] br[2] wl[177] vdd gnd cell_6t
Xbit_r178_c2 bl[2] br[2] wl[178] vdd gnd cell_6t
Xbit_r179_c2 bl[2] br[2] wl[179] vdd gnd cell_6t
Xbit_r180_c2 bl[2] br[2] wl[180] vdd gnd cell_6t
Xbit_r181_c2 bl[2] br[2] wl[181] vdd gnd cell_6t
Xbit_r182_c2 bl[2] br[2] wl[182] vdd gnd cell_6t
Xbit_r183_c2 bl[2] br[2] wl[183] vdd gnd cell_6t
Xbit_r184_c2 bl[2] br[2] wl[184] vdd gnd cell_6t
Xbit_r185_c2 bl[2] br[2] wl[185] vdd gnd cell_6t
Xbit_r186_c2 bl[2] br[2] wl[186] vdd gnd cell_6t
Xbit_r187_c2 bl[2] br[2] wl[187] vdd gnd cell_6t
Xbit_r188_c2 bl[2] br[2] wl[188] vdd gnd cell_6t
Xbit_r189_c2 bl[2] br[2] wl[189] vdd gnd cell_6t
Xbit_r190_c2 bl[2] br[2] wl[190] vdd gnd cell_6t
Xbit_r191_c2 bl[2] br[2] wl[191] vdd gnd cell_6t
Xbit_r192_c2 bl[2] br[2] wl[192] vdd gnd cell_6t
Xbit_r193_c2 bl[2] br[2] wl[193] vdd gnd cell_6t
Xbit_r194_c2 bl[2] br[2] wl[194] vdd gnd cell_6t
Xbit_r195_c2 bl[2] br[2] wl[195] vdd gnd cell_6t
Xbit_r196_c2 bl[2] br[2] wl[196] vdd gnd cell_6t
Xbit_r197_c2 bl[2] br[2] wl[197] vdd gnd cell_6t
Xbit_r198_c2 bl[2] br[2] wl[198] vdd gnd cell_6t
Xbit_r199_c2 bl[2] br[2] wl[199] vdd gnd cell_6t
Xbit_r200_c2 bl[2] br[2] wl[200] vdd gnd cell_6t
Xbit_r201_c2 bl[2] br[2] wl[201] vdd gnd cell_6t
Xbit_r202_c2 bl[2] br[2] wl[202] vdd gnd cell_6t
Xbit_r203_c2 bl[2] br[2] wl[203] vdd gnd cell_6t
Xbit_r204_c2 bl[2] br[2] wl[204] vdd gnd cell_6t
Xbit_r205_c2 bl[2] br[2] wl[205] vdd gnd cell_6t
Xbit_r206_c2 bl[2] br[2] wl[206] vdd gnd cell_6t
Xbit_r207_c2 bl[2] br[2] wl[207] vdd gnd cell_6t
Xbit_r208_c2 bl[2] br[2] wl[208] vdd gnd cell_6t
Xbit_r209_c2 bl[2] br[2] wl[209] vdd gnd cell_6t
Xbit_r210_c2 bl[2] br[2] wl[210] vdd gnd cell_6t
Xbit_r211_c2 bl[2] br[2] wl[211] vdd gnd cell_6t
Xbit_r212_c2 bl[2] br[2] wl[212] vdd gnd cell_6t
Xbit_r213_c2 bl[2] br[2] wl[213] vdd gnd cell_6t
Xbit_r214_c2 bl[2] br[2] wl[214] vdd gnd cell_6t
Xbit_r215_c2 bl[2] br[2] wl[215] vdd gnd cell_6t
Xbit_r216_c2 bl[2] br[2] wl[216] vdd gnd cell_6t
Xbit_r217_c2 bl[2] br[2] wl[217] vdd gnd cell_6t
Xbit_r218_c2 bl[2] br[2] wl[218] vdd gnd cell_6t
Xbit_r219_c2 bl[2] br[2] wl[219] vdd gnd cell_6t
Xbit_r220_c2 bl[2] br[2] wl[220] vdd gnd cell_6t
Xbit_r221_c2 bl[2] br[2] wl[221] vdd gnd cell_6t
Xbit_r222_c2 bl[2] br[2] wl[222] vdd gnd cell_6t
Xbit_r223_c2 bl[2] br[2] wl[223] vdd gnd cell_6t
Xbit_r224_c2 bl[2] br[2] wl[224] vdd gnd cell_6t
Xbit_r225_c2 bl[2] br[2] wl[225] vdd gnd cell_6t
Xbit_r226_c2 bl[2] br[2] wl[226] vdd gnd cell_6t
Xbit_r227_c2 bl[2] br[2] wl[227] vdd gnd cell_6t
Xbit_r228_c2 bl[2] br[2] wl[228] vdd gnd cell_6t
Xbit_r229_c2 bl[2] br[2] wl[229] vdd gnd cell_6t
Xbit_r230_c2 bl[2] br[2] wl[230] vdd gnd cell_6t
Xbit_r231_c2 bl[2] br[2] wl[231] vdd gnd cell_6t
Xbit_r232_c2 bl[2] br[2] wl[232] vdd gnd cell_6t
Xbit_r233_c2 bl[2] br[2] wl[233] vdd gnd cell_6t
Xbit_r234_c2 bl[2] br[2] wl[234] vdd gnd cell_6t
Xbit_r235_c2 bl[2] br[2] wl[235] vdd gnd cell_6t
Xbit_r236_c2 bl[2] br[2] wl[236] vdd gnd cell_6t
Xbit_r237_c2 bl[2] br[2] wl[237] vdd gnd cell_6t
Xbit_r238_c2 bl[2] br[2] wl[238] vdd gnd cell_6t
Xbit_r239_c2 bl[2] br[2] wl[239] vdd gnd cell_6t
Xbit_r240_c2 bl[2] br[2] wl[240] vdd gnd cell_6t
Xbit_r241_c2 bl[2] br[2] wl[241] vdd gnd cell_6t
Xbit_r242_c2 bl[2] br[2] wl[242] vdd gnd cell_6t
Xbit_r243_c2 bl[2] br[2] wl[243] vdd gnd cell_6t
Xbit_r244_c2 bl[2] br[2] wl[244] vdd gnd cell_6t
Xbit_r245_c2 bl[2] br[2] wl[245] vdd gnd cell_6t
Xbit_r246_c2 bl[2] br[2] wl[246] vdd gnd cell_6t
Xbit_r247_c2 bl[2] br[2] wl[247] vdd gnd cell_6t
Xbit_r248_c2 bl[2] br[2] wl[248] vdd gnd cell_6t
Xbit_r249_c2 bl[2] br[2] wl[249] vdd gnd cell_6t
Xbit_r250_c2 bl[2] br[2] wl[250] vdd gnd cell_6t
Xbit_r251_c2 bl[2] br[2] wl[251] vdd gnd cell_6t
Xbit_r252_c2 bl[2] br[2] wl[252] vdd gnd cell_6t
Xbit_r253_c2 bl[2] br[2] wl[253] vdd gnd cell_6t
Xbit_r254_c2 bl[2] br[2] wl[254] vdd gnd cell_6t
Xbit_r255_c2 bl[2] br[2] wl[255] vdd gnd cell_6t
Xbit_r0_c3 bl[3] br[3] wl[0] vdd gnd cell_6t
Xbit_r1_c3 bl[3] br[3] wl[1] vdd gnd cell_6t
Xbit_r2_c3 bl[3] br[3] wl[2] vdd gnd cell_6t
Xbit_r3_c3 bl[3] br[3] wl[3] vdd gnd cell_6t
Xbit_r4_c3 bl[3] br[3] wl[4] vdd gnd cell_6t
Xbit_r5_c3 bl[3] br[3] wl[5] vdd gnd cell_6t
Xbit_r6_c3 bl[3] br[3] wl[6] vdd gnd cell_6t
Xbit_r7_c3 bl[3] br[3] wl[7] vdd gnd cell_6t
Xbit_r8_c3 bl[3] br[3] wl[8] vdd gnd cell_6t
Xbit_r9_c3 bl[3] br[3] wl[9] vdd gnd cell_6t
Xbit_r10_c3 bl[3] br[3] wl[10] vdd gnd cell_6t
Xbit_r11_c3 bl[3] br[3] wl[11] vdd gnd cell_6t
Xbit_r12_c3 bl[3] br[3] wl[12] vdd gnd cell_6t
Xbit_r13_c3 bl[3] br[3] wl[13] vdd gnd cell_6t
Xbit_r14_c3 bl[3] br[3] wl[14] vdd gnd cell_6t
Xbit_r15_c3 bl[3] br[3] wl[15] vdd gnd cell_6t
Xbit_r16_c3 bl[3] br[3] wl[16] vdd gnd cell_6t
Xbit_r17_c3 bl[3] br[3] wl[17] vdd gnd cell_6t
Xbit_r18_c3 bl[3] br[3] wl[18] vdd gnd cell_6t
Xbit_r19_c3 bl[3] br[3] wl[19] vdd gnd cell_6t
Xbit_r20_c3 bl[3] br[3] wl[20] vdd gnd cell_6t
Xbit_r21_c3 bl[3] br[3] wl[21] vdd gnd cell_6t
Xbit_r22_c3 bl[3] br[3] wl[22] vdd gnd cell_6t
Xbit_r23_c3 bl[3] br[3] wl[23] vdd gnd cell_6t
Xbit_r24_c3 bl[3] br[3] wl[24] vdd gnd cell_6t
Xbit_r25_c3 bl[3] br[3] wl[25] vdd gnd cell_6t
Xbit_r26_c3 bl[3] br[3] wl[26] vdd gnd cell_6t
Xbit_r27_c3 bl[3] br[3] wl[27] vdd gnd cell_6t
Xbit_r28_c3 bl[3] br[3] wl[28] vdd gnd cell_6t
Xbit_r29_c3 bl[3] br[3] wl[29] vdd gnd cell_6t
Xbit_r30_c3 bl[3] br[3] wl[30] vdd gnd cell_6t
Xbit_r31_c3 bl[3] br[3] wl[31] vdd gnd cell_6t
Xbit_r32_c3 bl[3] br[3] wl[32] vdd gnd cell_6t
Xbit_r33_c3 bl[3] br[3] wl[33] vdd gnd cell_6t
Xbit_r34_c3 bl[3] br[3] wl[34] vdd gnd cell_6t
Xbit_r35_c3 bl[3] br[3] wl[35] vdd gnd cell_6t
Xbit_r36_c3 bl[3] br[3] wl[36] vdd gnd cell_6t
Xbit_r37_c3 bl[3] br[3] wl[37] vdd gnd cell_6t
Xbit_r38_c3 bl[3] br[3] wl[38] vdd gnd cell_6t
Xbit_r39_c3 bl[3] br[3] wl[39] vdd gnd cell_6t
Xbit_r40_c3 bl[3] br[3] wl[40] vdd gnd cell_6t
Xbit_r41_c3 bl[3] br[3] wl[41] vdd gnd cell_6t
Xbit_r42_c3 bl[3] br[3] wl[42] vdd gnd cell_6t
Xbit_r43_c3 bl[3] br[3] wl[43] vdd gnd cell_6t
Xbit_r44_c3 bl[3] br[3] wl[44] vdd gnd cell_6t
Xbit_r45_c3 bl[3] br[3] wl[45] vdd gnd cell_6t
Xbit_r46_c3 bl[3] br[3] wl[46] vdd gnd cell_6t
Xbit_r47_c3 bl[3] br[3] wl[47] vdd gnd cell_6t
Xbit_r48_c3 bl[3] br[3] wl[48] vdd gnd cell_6t
Xbit_r49_c3 bl[3] br[3] wl[49] vdd gnd cell_6t
Xbit_r50_c3 bl[3] br[3] wl[50] vdd gnd cell_6t
Xbit_r51_c3 bl[3] br[3] wl[51] vdd gnd cell_6t
Xbit_r52_c3 bl[3] br[3] wl[52] vdd gnd cell_6t
Xbit_r53_c3 bl[3] br[3] wl[53] vdd gnd cell_6t
Xbit_r54_c3 bl[3] br[3] wl[54] vdd gnd cell_6t
Xbit_r55_c3 bl[3] br[3] wl[55] vdd gnd cell_6t
Xbit_r56_c3 bl[3] br[3] wl[56] vdd gnd cell_6t
Xbit_r57_c3 bl[3] br[3] wl[57] vdd gnd cell_6t
Xbit_r58_c3 bl[3] br[3] wl[58] vdd gnd cell_6t
Xbit_r59_c3 bl[3] br[3] wl[59] vdd gnd cell_6t
Xbit_r60_c3 bl[3] br[3] wl[60] vdd gnd cell_6t
Xbit_r61_c3 bl[3] br[3] wl[61] vdd gnd cell_6t
Xbit_r62_c3 bl[3] br[3] wl[62] vdd gnd cell_6t
Xbit_r63_c3 bl[3] br[3] wl[63] vdd gnd cell_6t
Xbit_r64_c3 bl[3] br[3] wl[64] vdd gnd cell_6t
Xbit_r65_c3 bl[3] br[3] wl[65] vdd gnd cell_6t
Xbit_r66_c3 bl[3] br[3] wl[66] vdd gnd cell_6t
Xbit_r67_c3 bl[3] br[3] wl[67] vdd gnd cell_6t
Xbit_r68_c3 bl[3] br[3] wl[68] vdd gnd cell_6t
Xbit_r69_c3 bl[3] br[3] wl[69] vdd gnd cell_6t
Xbit_r70_c3 bl[3] br[3] wl[70] vdd gnd cell_6t
Xbit_r71_c3 bl[3] br[3] wl[71] vdd gnd cell_6t
Xbit_r72_c3 bl[3] br[3] wl[72] vdd gnd cell_6t
Xbit_r73_c3 bl[3] br[3] wl[73] vdd gnd cell_6t
Xbit_r74_c3 bl[3] br[3] wl[74] vdd gnd cell_6t
Xbit_r75_c3 bl[3] br[3] wl[75] vdd gnd cell_6t
Xbit_r76_c3 bl[3] br[3] wl[76] vdd gnd cell_6t
Xbit_r77_c3 bl[3] br[3] wl[77] vdd gnd cell_6t
Xbit_r78_c3 bl[3] br[3] wl[78] vdd gnd cell_6t
Xbit_r79_c3 bl[3] br[3] wl[79] vdd gnd cell_6t
Xbit_r80_c3 bl[3] br[3] wl[80] vdd gnd cell_6t
Xbit_r81_c3 bl[3] br[3] wl[81] vdd gnd cell_6t
Xbit_r82_c3 bl[3] br[3] wl[82] vdd gnd cell_6t
Xbit_r83_c3 bl[3] br[3] wl[83] vdd gnd cell_6t
Xbit_r84_c3 bl[3] br[3] wl[84] vdd gnd cell_6t
Xbit_r85_c3 bl[3] br[3] wl[85] vdd gnd cell_6t
Xbit_r86_c3 bl[3] br[3] wl[86] vdd gnd cell_6t
Xbit_r87_c3 bl[3] br[3] wl[87] vdd gnd cell_6t
Xbit_r88_c3 bl[3] br[3] wl[88] vdd gnd cell_6t
Xbit_r89_c3 bl[3] br[3] wl[89] vdd gnd cell_6t
Xbit_r90_c3 bl[3] br[3] wl[90] vdd gnd cell_6t
Xbit_r91_c3 bl[3] br[3] wl[91] vdd gnd cell_6t
Xbit_r92_c3 bl[3] br[3] wl[92] vdd gnd cell_6t
Xbit_r93_c3 bl[3] br[3] wl[93] vdd gnd cell_6t
Xbit_r94_c3 bl[3] br[3] wl[94] vdd gnd cell_6t
Xbit_r95_c3 bl[3] br[3] wl[95] vdd gnd cell_6t
Xbit_r96_c3 bl[3] br[3] wl[96] vdd gnd cell_6t
Xbit_r97_c3 bl[3] br[3] wl[97] vdd gnd cell_6t
Xbit_r98_c3 bl[3] br[3] wl[98] vdd gnd cell_6t
Xbit_r99_c3 bl[3] br[3] wl[99] vdd gnd cell_6t
Xbit_r100_c3 bl[3] br[3] wl[100] vdd gnd cell_6t
Xbit_r101_c3 bl[3] br[3] wl[101] vdd gnd cell_6t
Xbit_r102_c3 bl[3] br[3] wl[102] vdd gnd cell_6t
Xbit_r103_c3 bl[3] br[3] wl[103] vdd gnd cell_6t
Xbit_r104_c3 bl[3] br[3] wl[104] vdd gnd cell_6t
Xbit_r105_c3 bl[3] br[3] wl[105] vdd gnd cell_6t
Xbit_r106_c3 bl[3] br[3] wl[106] vdd gnd cell_6t
Xbit_r107_c3 bl[3] br[3] wl[107] vdd gnd cell_6t
Xbit_r108_c3 bl[3] br[3] wl[108] vdd gnd cell_6t
Xbit_r109_c3 bl[3] br[3] wl[109] vdd gnd cell_6t
Xbit_r110_c3 bl[3] br[3] wl[110] vdd gnd cell_6t
Xbit_r111_c3 bl[3] br[3] wl[111] vdd gnd cell_6t
Xbit_r112_c3 bl[3] br[3] wl[112] vdd gnd cell_6t
Xbit_r113_c3 bl[3] br[3] wl[113] vdd gnd cell_6t
Xbit_r114_c3 bl[3] br[3] wl[114] vdd gnd cell_6t
Xbit_r115_c3 bl[3] br[3] wl[115] vdd gnd cell_6t
Xbit_r116_c3 bl[3] br[3] wl[116] vdd gnd cell_6t
Xbit_r117_c3 bl[3] br[3] wl[117] vdd gnd cell_6t
Xbit_r118_c3 bl[3] br[3] wl[118] vdd gnd cell_6t
Xbit_r119_c3 bl[3] br[3] wl[119] vdd gnd cell_6t
Xbit_r120_c3 bl[3] br[3] wl[120] vdd gnd cell_6t
Xbit_r121_c3 bl[3] br[3] wl[121] vdd gnd cell_6t
Xbit_r122_c3 bl[3] br[3] wl[122] vdd gnd cell_6t
Xbit_r123_c3 bl[3] br[3] wl[123] vdd gnd cell_6t
Xbit_r124_c3 bl[3] br[3] wl[124] vdd gnd cell_6t
Xbit_r125_c3 bl[3] br[3] wl[125] vdd gnd cell_6t
Xbit_r126_c3 bl[3] br[3] wl[126] vdd gnd cell_6t
Xbit_r127_c3 bl[3] br[3] wl[127] vdd gnd cell_6t
Xbit_r128_c3 bl[3] br[3] wl[128] vdd gnd cell_6t
Xbit_r129_c3 bl[3] br[3] wl[129] vdd gnd cell_6t
Xbit_r130_c3 bl[3] br[3] wl[130] vdd gnd cell_6t
Xbit_r131_c3 bl[3] br[3] wl[131] vdd gnd cell_6t
Xbit_r132_c3 bl[3] br[3] wl[132] vdd gnd cell_6t
Xbit_r133_c3 bl[3] br[3] wl[133] vdd gnd cell_6t
Xbit_r134_c3 bl[3] br[3] wl[134] vdd gnd cell_6t
Xbit_r135_c3 bl[3] br[3] wl[135] vdd gnd cell_6t
Xbit_r136_c3 bl[3] br[3] wl[136] vdd gnd cell_6t
Xbit_r137_c3 bl[3] br[3] wl[137] vdd gnd cell_6t
Xbit_r138_c3 bl[3] br[3] wl[138] vdd gnd cell_6t
Xbit_r139_c3 bl[3] br[3] wl[139] vdd gnd cell_6t
Xbit_r140_c3 bl[3] br[3] wl[140] vdd gnd cell_6t
Xbit_r141_c3 bl[3] br[3] wl[141] vdd gnd cell_6t
Xbit_r142_c3 bl[3] br[3] wl[142] vdd gnd cell_6t
Xbit_r143_c3 bl[3] br[3] wl[143] vdd gnd cell_6t
Xbit_r144_c3 bl[3] br[3] wl[144] vdd gnd cell_6t
Xbit_r145_c3 bl[3] br[3] wl[145] vdd gnd cell_6t
Xbit_r146_c3 bl[3] br[3] wl[146] vdd gnd cell_6t
Xbit_r147_c3 bl[3] br[3] wl[147] vdd gnd cell_6t
Xbit_r148_c3 bl[3] br[3] wl[148] vdd gnd cell_6t
Xbit_r149_c3 bl[3] br[3] wl[149] vdd gnd cell_6t
Xbit_r150_c3 bl[3] br[3] wl[150] vdd gnd cell_6t
Xbit_r151_c3 bl[3] br[3] wl[151] vdd gnd cell_6t
Xbit_r152_c3 bl[3] br[3] wl[152] vdd gnd cell_6t
Xbit_r153_c3 bl[3] br[3] wl[153] vdd gnd cell_6t
Xbit_r154_c3 bl[3] br[3] wl[154] vdd gnd cell_6t
Xbit_r155_c3 bl[3] br[3] wl[155] vdd gnd cell_6t
Xbit_r156_c3 bl[3] br[3] wl[156] vdd gnd cell_6t
Xbit_r157_c3 bl[3] br[3] wl[157] vdd gnd cell_6t
Xbit_r158_c3 bl[3] br[3] wl[158] vdd gnd cell_6t
Xbit_r159_c3 bl[3] br[3] wl[159] vdd gnd cell_6t
Xbit_r160_c3 bl[3] br[3] wl[160] vdd gnd cell_6t
Xbit_r161_c3 bl[3] br[3] wl[161] vdd gnd cell_6t
Xbit_r162_c3 bl[3] br[3] wl[162] vdd gnd cell_6t
Xbit_r163_c3 bl[3] br[3] wl[163] vdd gnd cell_6t
Xbit_r164_c3 bl[3] br[3] wl[164] vdd gnd cell_6t
Xbit_r165_c3 bl[3] br[3] wl[165] vdd gnd cell_6t
Xbit_r166_c3 bl[3] br[3] wl[166] vdd gnd cell_6t
Xbit_r167_c3 bl[3] br[3] wl[167] vdd gnd cell_6t
Xbit_r168_c3 bl[3] br[3] wl[168] vdd gnd cell_6t
Xbit_r169_c3 bl[3] br[3] wl[169] vdd gnd cell_6t
Xbit_r170_c3 bl[3] br[3] wl[170] vdd gnd cell_6t
Xbit_r171_c3 bl[3] br[3] wl[171] vdd gnd cell_6t
Xbit_r172_c3 bl[3] br[3] wl[172] vdd gnd cell_6t
Xbit_r173_c3 bl[3] br[3] wl[173] vdd gnd cell_6t
Xbit_r174_c3 bl[3] br[3] wl[174] vdd gnd cell_6t
Xbit_r175_c3 bl[3] br[3] wl[175] vdd gnd cell_6t
Xbit_r176_c3 bl[3] br[3] wl[176] vdd gnd cell_6t
Xbit_r177_c3 bl[3] br[3] wl[177] vdd gnd cell_6t
Xbit_r178_c3 bl[3] br[3] wl[178] vdd gnd cell_6t
Xbit_r179_c3 bl[3] br[3] wl[179] vdd gnd cell_6t
Xbit_r180_c3 bl[3] br[3] wl[180] vdd gnd cell_6t
Xbit_r181_c3 bl[3] br[3] wl[181] vdd gnd cell_6t
Xbit_r182_c3 bl[3] br[3] wl[182] vdd gnd cell_6t
Xbit_r183_c3 bl[3] br[3] wl[183] vdd gnd cell_6t
Xbit_r184_c3 bl[3] br[3] wl[184] vdd gnd cell_6t
Xbit_r185_c3 bl[3] br[3] wl[185] vdd gnd cell_6t
Xbit_r186_c3 bl[3] br[3] wl[186] vdd gnd cell_6t
Xbit_r187_c3 bl[3] br[3] wl[187] vdd gnd cell_6t
Xbit_r188_c3 bl[3] br[3] wl[188] vdd gnd cell_6t
Xbit_r189_c3 bl[3] br[3] wl[189] vdd gnd cell_6t
Xbit_r190_c3 bl[3] br[3] wl[190] vdd gnd cell_6t
Xbit_r191_c3 bl[3] br[3] wl[191] vdd gnd cell_6t
Xbit_r192_c3 bl[3] br[3] wl[192] vdd gnd cell_6t
Xbit_r193_c3 bl[3] br[3] wl[193] vdd gnd cell_6t
Xbit_r194_c3 bl[3] br[3] wl[194] vdd gnd cell_6t
Xbit_r195_c3 bl[3] br[3] wl[195] vdd gnd cell_6t
Xbit_r196_c3 bl[3] br[3] wl[196] vdd gnd cell_6t
Xbit_r197_c3 bl[3] br[3] wl[197] vdd gnd cell_6t
Xbit_r198_c3 bl[3] br[3] wl[198] vdd gnd cell_6t
Xbit_r199_c3 bl[3] br[3] wl[199] vdd gnd cell_6t
Xbit_r200_c3 bl[3] br[3] wl[200] vdd gnd cell_6t
Xbit_r201_c3 bl[3] br[3] wl[201] vdd gnd cell_6t
Xbit_r202_c3 bl[3] br[3] wl[202] vdd gnd cell_6t
Xbit_r203_c3 bl[3] br[3] wl[203] vdd gnd cell_6t
Xbit_r204_c3 bl[3] br[3] wl[204] vdd gnd cell_6t
Xbit_r205_c3 bl[3] br[3] wl[205] vdd gnd cell_6t
Xbit_r206_c3 bl[3] br[3] wl[206] vdd gnd cell_6t
Xbit_r207_c3 bl[3] br[3] wl[207] vdd gnd cell_6t
Xbit_r208_c3 bl[3] br[3] wl[208] vdd gnd cell_6t
Xbit_r209_c3 bl[3] br[3] wl[209] vdd gnd cell_6t
Xbit_r210_c3 bl[3] br[3] wl[210] vdd gnd cell_6t
Xbit_r211_c3 bl[3] br[3] wl[211] vdd gnd cell_6t
Xbit_r212_c3 bl[3] br[3] wl[212] vdd gnd cell_6t
Xbit_r213_c3 bl[3] br[3] wl[213] vdd gnd cell_6t
Xbit_r214_c3 bl[3] br[3] wl[214] vdd gnd cell_6t
Xbit_r215_c3 bl[3] br[3] wl[215] vdd gnd cell_6t
Xbit_r216_c3 bl[3] br[3] wl[216] vdd gnd cell_6t
Xbit_r217_c3 bl[3] br[3] wl[217] vdd gnd cell_6t
Xbit_r218_c3 bl[3] br[3] wl[218] vdd gnd cell_6t
Xbit_r219_c3 bl[3] br[3] wl[219] vdd gnd cell_6t
Xbit_r220_c3 bl[3] br[3] wl[220] vdd gnd cell_6t
Xbit_r221_c3 bl[3] br[3] wl[221] vdd gnd cell_6t
Xbit_r222_c3 bl[3] br[3] wl[222] vdd gnd cell_6t
Xbit_r223_c3 bl[3] br[3] wl[223] vdd gnd cell_6t
Xbit_r224_c3 bl[3] br[3] wl[224] vdd gnd cell_6t
Xbit_r225_c3 bl[3] br[3] wl[225] vdd gnd cell_6t
Xbit_r226_c3 bl[3] br[3] wl[226] vdd gnd cell_6t
Xbit_r227_c3 bl[3] br[3] wl[227] vdd gnd cell_6t
Xbit_r228_c3 bl[3] br[3] wl[228] vdd gnd cell_6t
Xbit_r229_c3 bl[3] br[3] wl[229] vdd gnd cell_6t
Xbit_r230_c3 bl[3] br[3] wl[230] vdd gnd cell_6t
Xbit_r231_c3 bl[3] br[3] wl[231] vdd gnd cell_6t
Xbit_r232_c3 bl[3] br[3] wl[232] vdd gnd cell_6t
Xbit_r233_c3 bl[3] br[3] wl[233] vdd gnd cell_6t
Xbit_r234_c3 bl[3] br[3] wl[234] vdd gnd cell_6t
Xbit_r235_c3 bl[3] br[3] wl[235] vdd gnd cell_6t
Xbit_r236_c3 bl[3] br[3] wl[236] vdd gnd cell_6t
Xbit_r237_c3 bl[3] br[3] wl[237] vdd gnd cell_6t
Xbit_r238_c3 bl[3] br[3] wl[238] vdd gnd cell_6t
Xbit_r239_c3 bl[3] br[3] wl[239] vdd gnd cell_6t
Xbit_r240_c3 bl[3] br[3] wl[240] vdd gnd cell_6t
Xbit_r241_c3 bl[3] br[3] wl[241] vdd gnd cell_6t
Xbit_r242_c3 bl[3] br[3] wl[242] vdd gnd cell_6t
Xbit_r243_c3 bl[3] br[3] wl[243] vdd gnd cell_6t
Xbit_r244_c3 bl[3] br[3] wl[244] vdd gnd cell_6t
Xbit_r245_c3 bl[3] br[3] wl[245] vdd gnd cell_6t
Xbit_r246_c3 bl[3] br[3] wl[246] vdd gnd cell_6t
Xbit_r247_c3 bl[3] br[3] wl[247] vdd gnd cell_6t
Xbit_r248_c3 bl[3] br[3] wl[248] vdd gnd cell_6t
Xbit_r249_c3 bl[3] br[3] wl[249] vdd gnd cell_6t
Xbit_r250_c3 bl[3] br[3] wl[250] vdd gnd cell_6t
Xbit_r251_c3 bl[3] br[3] wl[251] vdd gnd cell_6t
Xbit_r252_c3 bl[3] br[3] wl[252] vdd gnd cell_6t
Xbit_r253_c3 bl[3] br[3] wl[253] vdd gnd cell_6t
Xbit_r254_c3 bl[3] br[3] wl[254] vdd gnd cell_6t
Xbit_r255_c3 bl[3] br[3] wl[255] vdd gnd cell_6t
Xbit_r0_c4 bl[4] br[4] wl[0] vdd gnd cell_6t
Xbit_r1_c4 bl[4] br[4] wl[1] vdd gnd cell_6t
Xbit_r2_c4 bl[4] br[4] wl[2] vdd gnd cell_6t
Xbit_r3_c4 bl[4] br[4] wl[3] vdd gnd cell_6t
Xbit_r4_c4 bl[4] br[4] wl[4] vdd gnd cell_6t
Xbit_r5_c4 bl[4] br[4] wl[5] vdd gnd cell_6t
Xbit_r6_c4 bl[4] br[4] wl[6] vdd gnd cell_6t
Xbit_r7_c4 bl[4] br[4] wl[7] vdd gnd cell_6t
Xbit_r8_c4 bl[4] br[4] wl[8] vdd gnd cell_6t
Xbit_r9_c4 bl[4] br[4] wl[9] vdd gnd cell_6t
Xbit_r10_c4 bl[4] br[4] wl[10] vdd gnd cell_6t
Xbit_r11_c4 bl[4] br[4] wl[11] vdd gnd cell_6t
Xbit_r12_c4 bl[4] br[4] wl[12] vdd gnd cell_6t
Xbit_r13_c4 bl[4] br[4] wl[13] vdd gnd cell_6t
Xbit_r14_c4 bl[4] br[4] wl[14] vdd gnd cell_6t
Xbit_r15_c4 bl[4] br[4] wl[15] vdd gnd cell_6t
Xbit_r16_c4 bl[4] br[4] wl[16] vdd gnd cell_6t
Xbit_r17_c4 bl[4] br[4] wl[17] vdd gnd cell_6t
Xbit_r18_c4 bl[4] br[4] wl[18] vdd gnd cell_6t
Xbit_r19_c4 bl[4] br[4] wl[19] vdd gnd cell_6t
Xbit_r20_c4 bl[4] br[4] wl[20] vdd gnd cell_6t
Xbit_r21_c4 bl[4] br[4] wl[21] vdd gnd cell_6t
Xbit_r22_c4 bl[4] br[4] wl[22] vdd gnd cell_6t
Xbit_r23_c4 bl[4] br[4] wl[23] vdd gnd cell_6t
Xbit_r24_c4 bl[4] br[4] wl[24] vdd gnd cell_6t
Xbit_r25_c4 bl[4] br[4] wl[25] vdd gnd cell_6t
Xbit_r26_c4 bl[4] br[4] wl[26] vdd gnd cell_6t
Xbit_r27_c4 bl[4] br[4] wl[27] vdd gnd cell_6t
Xbit_r28_c4 bl[4] br[4] wl[28] vdd gnd cell_6t
Xbit_r29_c4 bl[4] br[4] wl[29] vdd gnd cell_6t
Xbit_r30_c4 bl[4] br[4] wl[30] vdd gnd cell_6t
Xbit_r31_c4 bl[4] br[4] wl[31] vdd gnd cell_6t
Xbit_r32_c4 bl[4] br[4] wl[32] vdd gnd cell_6t
Xbit_r33_c4 bl[4] br[4] wl[33] vdd gnd cell_6t
Xbit_r34_c4 bl[4] br[4] wl[34] vdd gnd cell_6t
Xbit_r35_c4 bl[4] br[4] wl[35] vdd gnd cell_6t
Xbit_r36_c4 bl[4] br[4] wl[36] vdd gnd cell_6t
Xbit_r37_c4 bl[4] br[4] wl[37] vdd gnd cell_6t
Xbit_r38_c4 bl[4] br[4] wl[38] vdd gnd cell_6t
Xbit_r39_c4 bl[4] br[4] wl[39] vdd gnd cell_6t
Xbit_r40_c4 bl[4] br[4] wl[40] vdd gnd cell_6t
Xbit_r41_c4 bl[4] br[4] wl[41] vdd gnd cell_6t
Xbit_r42_c4 bl[4] br[4] wl[42] vdd gnd cell_6t
Xbit_r43_c4 bl[4] br[4] wl[43] vdd gnd cell_6t
Xbit_r44_c4 bl[4] br[4] wl[44] vdd gnd cell_6t
Xbit_r45_c4 bl[4] br[4] wl[45] vdd gnd cell_6t
Xbit_r46_c4 bl[4] br[4] wl[46] vdd gnd cell_6t
Xbit_r47_c4 bl[4] br[4] wl[47] vdd gnd cell_6t
Xbit_r48_c4 bl[4] br[4] wl[48] vdd gnd cell_6t
Xbit_r49_c4 bl[4] br[4] wl[49] vdd gnd cell_6t
Xbit_r50_c4 bl[4] br[4] wl[50] vdd gnd cell_6t
Xbit_r51_c4 bl[4] br[4] wl[51] vdd gnd cell_6t
Xbit_r52_c4 bl[4] br[4] wl[52] vdd gnd cell_6t
Xbit_r53_c4 bl[4] br[4] wl[53] vdd gnd cell_6t
Xbit_r54_c4 bl[4] br[4] wl[54] vdd gnd cell_6t
Xbit_r55_c4 bl[4] br[4] wl[55] vdd gnd cell_6t
Xbit_r56_c4 bl[4] br[4] wl[56] vdd gnd cell_6t
Xbit_r57_c4 bl[4] br[4] wl[57] vdd gnd cell_6t
Xbit_r58_c4 bl[4] br[4] wl[58] vdd gnd cell_6t
Xbit_r59_c4 bl[4] br[4] wl[59] vdd gnd cell_6t
Xbit_r60_c4 bl[4] br[4] wl[60] vdd gnd cell_6t
Xbit_r61_c4 bl[4] br[4] wl[61] vdd gnd cell_6t
Xbit_r62_c4 bl[4] br[4] wl[62] vdd gnd cell_6t
Xbit_r63_c4 bl[4] br[4] wl[63] vdd gnd cell_6t
Xbit_r64_c4 bl[4] br[4] wl[64] vdd gnd cell_6t
Xbit_r65_c4 bl[4] br[4] wl[65] vdd gnd cell_6t
Xbit_r66_c4 bl[4] br[4] wl[66] vdd gnd cell_6t
Xbit_r67_c4 bl[4] br[4] wl[67] vdd gnd cell_6t
Xbit_r68_c4 bl[4] br[4] wl[68] vdd gnd cell_6t
Xbit_r69_c4 bl[4] br[4] wl[69] vdd gnd cell_6t
Xbit_r70_c4 bl[4] br[4] wl[70] vdd gnd cell_6t
Xbit_r71_c4 bl[4] br[4] wl[71] vdd gnd cell_6t
Xbit_r72_c4 bl[4] br[4] wl[72] vdd gnd cell_6t
Xbit_r73_c4 bl[4] br[4] wl[73] vdd gnd cell_6t
Xbit_r74_c4 bl[4] br[4] wl[74] vdd gnd cell_6t
Xbit_r75_c4 bl[4] br[4] wl[75] vdd gnd cell_6t
Xbit_r76_c4 bl[4] br[4] wl[76] vdd gnd cell_6t
Xbit_r77_c4 bl[4] br[4] wl[77] vdd gnd cell_6t
Xbit_r78_c4 bl[4] br[4] wl[78] vdd gnd cell_6t
Xbit_r79_c4 bl[4] br[4] wl[79] vdd gnd cell_6t
Xbit_r80_c4 bl[4] br[4] wl[80] vdd gnd cell_6t
Xbit_r81_c4 bl[4] br[4] wl[81] vdd gnd cell_6t
Xbit_r82_c4 bl[4] br[4] wl[82] vdd gnd cell_6t
Xbit_r83_c4 bl[4] br[4] wl[83] vdd gnd cell_6t
Xbit_r84_c4 bl[4] br[4] wl[84] vdd gnd cell_6t
Xbit_r85_c4 bl[4] br[4] wl[85] vdd gnd cell_6t
Xbit_r86_c4 bl[4] br[4] wl[86] vdd gnd cell_6t
Xbit_r87_c4 bl[4] br[4] wl[87] vdd gnd cell_6t
Xbit_r88_c4 bl[4] br[4] wl[88] vdd gnd cell_6t
Xbit_r89_c4 bl[4] br[4] wl[89] vdd gnd cell_6t
Xbit_r90_c4 bl[4] br[4] wl[90] vdd gnd cell_6t
Xbit_r91_c4 bl[4] br[4] wl[91] vdd gnd cell_6t
Xbit_r92_c4 bl[4] br[4] wl[92] vdd gnd cell_6t
Xbit_r93_c4 bl[4] br[4] wl[93] vdd gnd cell_6t
Xbit_r94_c4 bl[4] br[4] wl[94] vdd gnd cell_6t
Xbit_r95_c4 bl[4] br[4] wl[95] vdd gnd cell_6t
Xbit_r96_c4 bl[4] br[4] wl[96] vdd gnd cell_6t
Xbit_r97_c4 bl[4] br[4] wl[97] vdd gnd cell_6t
Xbit_r98_c4 bl[4] br[4] wl[98] vdd gnd cell_6t
Xbit_r99_c4 bl[4] br[4] wl[99] vdd gnd cell_6t
Xbit_r100_c4 bl[4] br[4] wl[100] vdd gnd cell_6t
Xbit_r101_c4 bl[4] br[4] wl[101] vdd gnd cell_6t
Xbit_r102_c4 bl[4] br[4] wl[102] vdd gnd cell_6t
Xbit_r103_c4 bl[4] br[4] wl[103] vdd gnd cell_6t
Xbit_r104_c4 bl[4] br[4] wl[104] vdd gnd cell_6t
Xbit_r105_c4 bl[4] br[4] wl[105] vdd gnd cell_6t
Xbit_r106_c4 bl[4] br[4] wl[106] vdd gnd cell_6t
Xbit_r107_c4 bl[4] br[4] wl[107] vdd gnd cell_6t
Xbit_r108_c4 bl[4] br[4] wl[108] vdd gnd cell_6t
Xbit_r109_c4 bl[4] br[4] wl[109] vdd gnd cell_6t
Xbit_r110_c4 bl[4] br[4] wl[110] vdd gnd cell_6t
Xbit_r111_c4 bl[4] br[4] wl[111] vdd gnd cell_6t
Xbit_r112_c4 bl[4] br[4] wl[112] vdd gnd cell_6t
Xbit_r113_c4 bl[4] br[4] wl[113] vdd gnd cell_6t
Xbit_r114_c4 bl[4] br[4] wl[114] vdd gnd cell_6t
Xbit_r115_c4 bl[4] br[4] wl[115] vdd gnd cell_6t
Xbit_r116_c4 bl[4] br[4] wl[116] vdd gnd cell_6t
Xbit_r117_c4 bl[4] br[4] wl[117] vdd gnd cell_6t
Xbit_r118_c4 bl[4] br[4] wl[118] vdd gnd cell_6t
Xbit_r119_c4 bl[4] br[4] wl[119] vdd gnd cell_6t
Xbit_r120_c4 bl[4] br[4] wl[120] vdd gnd cell_6t
Xbit_r121_c4 bl[4] br[4] wl[121] vdd gnd cell_6t
Xbit_r122_c4 bl[4] br[4] wl[122] vdd gnd cell_6t
Xbit_r123_c4 bl[4] br[4] wl[123] vdd gnd cell_6t
Xbit_r124_c4 bl[4] br[4] wl[124] vdd gnd cell_6t
Xbit_r125_c4 bl[4] br[4] wl[125] vdd gnd cell_6t
Xbit_r126_c4 bl[4] br[4] wl[126] vdd gnd cell_6t
Xbit_r127_c4 bl[4] br[4] wl[127] vdd gnd cell_6t
Xbit_r128_c4 bl[4] br[4] wl[128] vdd gnd cell_6t
Xbit_r129_c4 bl[4] br[4] wl[129] vdd gnd cell_6t
Xbit_r130_c4 bl[4] br[4] wl[130] vdd gnd cell_6t
Xbit_r131_c4 bl[4] br[4] wl[131] vdd gnd cell_6t
Xbit_r132_c4 bl[4] br[4] wl[132] vdd gnd cell_6t
Xbit_r133_c4 bl[4] br[4] wl[133] vdd gnd cell_6t
Xbit_r134_c4 bl[4] br[4] wl[134] vdd gnd cell_6t
Xbit_r135_c4 bl[4] br[4] wl[135] vdd gnd cell_6t
Xbit_r136_c4 bl[4] br[4] wl[136] vdd gnd cell_6t
Xbit_r137_c4 bl[4] br[4] wl[137] vdd gnd cell_6t
Xbit_r138_c4 bl[4] br[4] wl[138] vdd gnd cell_6t
Xbit_r139_c4 bl[4] br[4] wl[139] vdd gnd cell_6t
Xbit_r140_c4 bl[4] br[4] wl[140] vdd gnd cell_6t
Xbit_r141_c4 bl[4] br[4] wl[141] vdd gnd cell_6t
Xbit_r142_c4 bl[4] br[4] wl[142] vdd gnd cell_6t
Xbit_r143_c4 bl[4] br[4] wl[143] vdd gnd cell_6t
Xbit_r144_c4 bl[4] br[4] wl[144] vdd gnd cell_6t
Xbit_r145_c4 bl[4] br[4] wl[145] vdd gnd cell_6t
Xbit_r146_c4 bl[4] br[4] wl[146] vdd gnd cell_6t
Xbit_r147_c4 bl[4] br[4] wl[147] vdd gnd cell_6t
Xbit_r148_c4 bl[4] br[4] wl[148] vdd gnd cell_6t
Xbit_r149_c4 bl[4] br[4] wl[149] vdd gnd cell_6t
Xbit_r150_c4 bl[4] br[4] wl[150] vdd gnd cell_6t
Xbit_r151_c4 bl[4] br[4] wl[151] vdd gnd cell_6t
Xbit_r152_c4 bl[4] br[4] wl[152] vdd gnd cell_6t
Xbit_r153_c4 bl[4] br[4] wl[153] vdd gnd cell_6t
Xbit_r154_c4 bl[4] br[4] wl[154] vdd gnd cell_6t
Xbit_r155_c4 bl[4] br[4] wl[155] vdd gnd cell_6t
Xbit_r156_c4 bl[4] br[4] wl[156] vdd gnd cell_6t
Xbit_r157_c4 bl[4] br[4] wl[157] vdd gnd cell_6t
Xbit_r158_c4 bl[4] br[4] wl[158] vdd gnd cell_6t
Xbit_r159_c4 bl[4] br[4] wl[159] vdd gnd cell_6t
Xbit_r160_c4 bl[4] br[4] wl[160] vdd gnd cell_6t
Xbit_r161_c4 bl[4] br[4] wl[161] vdd gnd cell_6t
Xbit_r162_c4 bl[4] br[4] wl[162] vdd gnd cell_6t
Xbit_r163_c4 bl[4] br[4] wl[163] vdd gnd cell_6t
Xbit_r164_c4 bl[4] br[4] wl[164] vdd gnd cell_6t
Xbit_r165_c4 bl[4] br[4] wl[165] vdd gnd cell_6t
Xbit_r166_c4 bl[4] br[4] wl[166] vdd gnd cell_6t
Xbit_r167_c4 bl[4] br[4] wl[167] vdd gnd cell_6t
Xbit_r168_c4 bl[4] br[4] wl[168] vdd gnd cell_6t
Xbit_r169_c4 bl[4] br[4] wl[169] vdd gnd cell_6t
Xbit_r170_c4 bl[4] br[4] wl[170] vdd gnd cell_6t
Xbit_r171_c4 bl[4] br[4] wl[171] vdd gnd cell_6t
Xbit_r172_c4 bl[4] br[4] wl[172] vdd gnd cell_6t
Xbit_r173_c4 bl[4] br[4] wl[173] vdd gnd cell_6t
Xbit_r174_c4 bl[4] br[4] wl[174] vdd gnd cell_6t
Xbit_r175_c4 bl[4] br[4] wl[175] vdd gnd cell_6t
Xbit_r176_c4 bl[4] br[4] wl[176] vdd gnd cell_6t
Xbit_r177_c4 bl[4] br[4] wl[177] vdd gnd cell_6t
Xbit_r178_c4 bl[4] br[4] wl[178] vdd gnd cell_6t
Xbit_r179_c4 bl[4] br[4] wl[179] vdd gnd cell_6t
Xbit_r180_c4 bl[4] br[4] wl[180] vdd gnd cell_6t
Xbit_r181_c4 bl[4] br[4] wl[181] vdd gnd cell_6t
Xbit_r182_c4 bl[4] br[4] wl[182] vdd gnd cell_6t
Xbit_r183_c4 bl[4] br[4] wl[183] vdd gnd cell_6t
Xbit_r184_c4 bl[4] br[4] wl[184] vdd gnd cell_6t
Xbit_r185_c4 bl[4] br[4] wl[185] vdd gnd cell_6t
Xbit_r186_c4 bl[4] br[4] wl[186] vdd gnd cell_6t
Xbit_r187_c4 bl[4] br[4] wl[187] vdd gnd cell_6t
Xbit_r188_c4 bl[4] br[4] wl[188] vdd gnd cell_6t
Xbit_r189_c4 bl[4] br[4] wl[189] vdd gnd cell_6t
Xbit_r190_c4 bl[4] br[4] wl[190] vdd gnd cell_6t
Xbit_r191_c4 bl[4] br[4] wl[191] vdd gnd cell_6t
Xbit_r192_c4 bl[4] br[4] wl[192] vdd gnd cell_6t
Xbit_r193_c4 bl[4] br[4] wl[193] vdd gnd cell_6t
Xbit_r194_c4 bl[4] br[4] wl[194] vdd gnd cell_6t
Xbit_r195_c4 bl[4] br[4] wl[195] vdd gnd cell_6t
Xbit_r196_c4 bl[4] br[4] wl[196] vdd gnd cell_6t
Xbit_r197_c4 bl[4] br[4] wl[197] vdd gnd cell_6t
Xbit_r198_c4 bl[4] br[4] wl[198] vdd gnd cell_6t
Xbit_r199_c4 bl[4] br[4] wl[199] vdd gnd cell_6t
Xbit_r200_c4 bl[4] br[4] wl[200] vdd gnd cell_6t
Xbit_r201_c4 bl[4] br[4] wl[201] vdd gnd cell_6t
Xbit_r202_c4 bl[4] br[4] wl[202] vdd gnd cell_6t
Xbit_r203_c4 bl[4] br[4] wl[203] vdd gnd cell_6t
Xbit_r204_c4 bl[4] br[4] wl[204] vdd gnd cell_6t
Xbit_r205_c4 bl[4] br[4] wl[205] vdd gnd cell_6t
Xbit_r206_c4 bl[4] br[4] wl[206] vdd gnd cell_6t
Xbit_r207_c4 bl[4] br[4] wl[207] vdd gnd cell_6t
Xbit_r208_c4 bl[4] br[4] wl[208] vdd gnd cell_6t
Xbit_r209_c4 bl[4] br[4] wl[209] vdd gnd cell_6t
Xbit_r210_c4 bl[4] br[4] wl[210] vdd gnd cell_6t
Xbit_r211_c4 bl[4] br[4] wl[211] vdd gnd cell_6t
Xbit_r212_c4 bl[4] br[4] wl[212] vdd gnd cell_6t
Xbit_r213_c4 bl[4] br[4] wl[213] vdd gnd cell_6t
Xbit_r214_c4 bl[4] br[4] wl[214] vdd gnd cell_6t
Xbit_r215_c4 bl[4] br[4] wl[215] vdd gnd cell_6t
Xbit_r216_c4 bl[4] br[4] wl[216] vdd gnd cell_6t
Xbit_r217_c4 bl[4] br[4] wl[217] vdd gnd cell_6t
Xbit_r218_c4 bl[4] br[4] wl[218] vdd gnd cell_6t
Xbit_r219_c4 bl[4] br[4] wl[219] vdd gnd cell_6t
Xbit_r220_c4 bl[4] br[4] wl[220] vdd gnd cell_6t
Xbit_r221_c4 bl[4] br[4] wl[221] vdd gnd cell_6t
Xbit_r222_c4 bl[4] br[4] wl[222] vdd gnd cell_6t
Xbit_r223_c4 bl[4] br[4] wl[223] vdd gnd cell_6t
Xbit_r224_c4 bl[4] br[4] wl[224] vdd gnd cell_6t
Xbit_r225_c4 bl[4] br[4] wl[225] vdd gnd cell_6t
Xbit_r226_c4 bl[4] br[4] wl[226] vdd gnd cell_6t
Xbit_r227_c4 bl[4] br[4] wl[227] vdd gnd cell_6t
Xbit_r228_c4 bl[4] br[4] wl[228] vdd gnd cell_6t
Xbit_r229_c4 bl[4] br[4] wl[229] vdd gnd cell_6t
Xbit_r230_c4 bl[4] br[4] wl[230] vdd gnd cell_6t
Xbit_r231_c4 bl[4] br[4] wl[231] vdd gnd cell_6t
Xbit_r232_c4 bl[4] br[4] wl[232] vdd gnd cell_6t
Xbit_r233_c4 bl[4] br[4] wl[233] vdd gnd cell_6t
Xbit_r234_c4 bl[4] br[4] wl[234] vdd gnd cell_6t
Xbit_r235_c4 bl[4] br[4] wl[235] vdd gnd cell_6t
Xbit_r236_c4 bl[4] br[4] wl[236] vdd gnd cell_6t
Xbit_r237_c4 bl[4] br[4] wl[237] vdd gnd cell_6t
Xbit_r238_c4 bl[4] br[4] wl[238] vdd gnd cell_6t
Xbit_r239_c4 bl[4] br[4] wl[239] vdd gnd cell_6t
Xbit_r240_c4 bl[4] br[4] wl[240] vdd gnd cell_6t
Xbit_r241_c4 bl[4] br[4] wl[241] vdd gnd cell_6t
Xbit_r242_c4 bl[4] br[4] wl[242] vdd gnd cell_6t
Xbit_r243_c4 bl[4] br[4] wl[243] vdd gnd cell_6t
Xbit_r244_c4 bl[4] br[4] wl[244] vdd gnd cell_6t
Xbit_r245_c4 bl[4] br[4] wl[245] vdd gnd cell_6t
Xbit_r246_c4 bl[4] br[4] wl[246] vdd gnd cell_6t
Xbit_r247_c4 bl[4] br[4] wl[247] vdd gnd cell_6t
Xbit_r248_c4 bl[4] br[4] wl[248] vdd gnd cell_6t
Xbit_r249_c4 bl[4] br[4] wl[249] vdd gnd cell_6t
Xbit_r250_c4 bl[4] br[4] wl[250] vdd gnd cell_6t
Xbit_r251_c4 bl[4] br[4] wl[251] vdd gnd cell_6t
Xbit_r252_c4 bl[4] br[4] wl[252] vdd gnd cell_6t
Xbit_r253_c4 bl[4] br[4] wl[253] vdd gnd cell_6t
Xbit_r254_c4 bl[4] br[4] wl[254] vdd gnd cell_6t
Xbit_r255_c4 bl[4] br[4] wl[255] vdd gnd cell_6t
Xbit_r0_c5 bl[5] br[5] wl[0] vdd gnd cell_6t
Xbit_r1_c5 bl[5] br[5] wl[1] vdd gnd cell_6t
Xbit_r2_c5 bl[5] br[5] wl[2] vdd gnd cell_6t
Xbit_r3_c5 bl[5] br[5] wl[3] vdd gnd cell_6t
Xbit_r4_c5 bl[5] br[5] wl[4] vdd gnd cell_6t
Xbit_r5_c5 bl[5] br[5] wl[5] vdd gnd cell_6t
Xbit_r6_c5 bl[5] br[5] wl[6] vdd gnd cell_6t
Xbit_r7_c5 bl[5] br[5] wl[7] vdd gnd cell_6t
Xbit_r8_c5 bl[5] br[5] wl[8] vdd gnd cell_6t
Xbit_r9_c5 bl[5] br[5] wl[9] vdd gnd cell_6t
Xbit_r10_c5 bl[5] br[5] wl[10] vdd gnd cell_6t
Xbit_r11_c5 bl[5] br[5] wl[11] vdd gnd cell_6t
Xbit_r12_c5 bl[5] br[5] wl[12] vdd gnd cell_6t
Xbit_r13_c5 bl[5] br[5] wl[13] vdd gnd cell_6t
Xbit_r14_c5 bl[5] br[5] wl[14] vdd gnd cell_6t
Xbit_r15_c5 bl[5] br[5] wl[15] vdd gnd cell_6t
Xbit_r16_c5 bl[5] br[5] wl[16] vdd gnd cell_6t
Xbit_r17_c5 bl[5] br[5] wl[17] vdd gnd cell_6t
Xbit_r18_c5 bl[5] br[5] wl[18] vdd gnd cell_6t
Xbit_r19_c5 bl[5] br[5] wl[19] vdd gnd cell_6t
Xbit_r20_c5 bl[5] br[5] wl[20] vdd gnd cell_6t
Xbit_r21_c5 bl[5] br[5] wl[21] vdd gnd cell_6t
Xbit_r22_c5 bl[5] br[5] wl[22] vdd gnd cell_6t
Xbit_r23_c5 bl[5] br[5] wl[23] vdd gnd cell_6t
Xbit_r24_c5 bl[5] br[5] wl[24] vdd gnd cell_6t
Xbit_r25_c5 bl[5] br[5] wl[25] vdd gnd cell_6t
Xbit_r26_c5 bl[5] br[5] wl[26] vdd gnd cell_6t
Xbit_r27_c5 bl[5] br[5] wl[27] vdd gnd cell_6t
Xbit_r28_c5 bl[5] br[5] wl[28] vdd gnd cell_6t
Xbit_r29_c5 bl[5] br[5] wl[29] vdd gnd cell_6t
Xbit_r30_c5 bl[5] br[5] wl[30] vdd gnd cell_6t
Xbit_r31_c5 bl[5] br[5] wl[31] vdd gnd cell_6t
Xbit_r32_c5 bl[5] br[5] wl[32] vdd gnd cell_6t
Xbit_r33_c5 bl[5] br[5] wl[33] vdd gnd cell_6t
Xbit_r34_c5 bl[5] br[5] wl[34] vdd gnd cell_6t
Xbit_r35_c5 bl[5] br[5] wl[35] vdd gnd cell_6t
Xbit_r36_c5 bl[5] br[5] wl[36] vdd gnd cell_6t
Xbit_r37_c5 bl[5] br[5] wl[37] vdd gnd cell_6t
Xbit_r38_c5 bl[5] br[5] wl[38] vdd gnd cell_6t
Xbit_r39_c5 bl[5] br[5] wl[39] vdd gnd cell_6t
Xbit_r40_c5 bl[5] br[5] wl[40] vdd gnd cell_6t
Xbit_r41_c5 bl[5] br[5] wl[41] vdd gnd cell_6t
Xbit_r42_c5 bl[5] br[5] wl[42] vdd gnd cell_6t
Xbit_r43_c5 bl[5] br[5] wl[43] vdd gnd cell_6t
Xbit_r44_c5 bl[5] br[5] wl[44] vdd gnd cell_6t
Xbit_r45_c5 bl[5] br[5] wl[45] vdd gnd cell_6t
Xbit_r46_c5 bl[5] br[5] wl[46] vdd gnd cell_6t
Xbit_r47_c5 bl[5] br[5] wl[47] vdd gnd cell_6t
Xbit_r48_c5 bl[5] br[5] wl[48] vdd gnd cell_6t
Xbit_r49_c5 bl[5] br[5] wl[49] vdd gnd cell_6t
Xbit_r50_c5 bl[5] br[5] wl[50] vdd gnd cell_6t
Xbit_r51_c5 bl[5] br[5] wl[51] vdd gnd cell_6t
Xbit_r52_c5 bl[5] br[5] wl[52] vdd gnd cell_6t
Xbit_r53_c5 bl[5] br[5] wl[53] vdd gnd cell_6t
Xbit_r54_c5 bl[5] br[5] wl[54] vdd gnd cell_6t
Xbit_r55_c5 bl[5] br[5] wl[55] vdd gnd cell_6t
Xbit_r56_c5 bl[5] br[5] wl[56] vdd gnd cell_6t
Xbit_r57_c5 bl[5] br[5] wl[57] vdd gnd cell_6t
Xbit_r58_c5 bl[5] br[5] wl[58] vdd gnd cell_6t
Xbit_r59_c5 bl[5] br[5] wl[59] vdd gnd cell_6t
Xbit_r60_c5 bl[5] br[5] wl[60] vdd gnd cell_6t
Xbit_r61_c5 bl[5] br[5] wl[61] vdd gnd cell_6t
Xbit_r62_c5 bl[5] br[5] wl[62] vdd gnd cell_6t
Xbit_r63_c5 bl[5] br[5] wl[63] vdd gnd cell_6t
Xbit_r64_c5 bl[5] br[5] wl[64] vdd gnd cell_6t
Xbit_r65_c5 bl[5] br[5] wl[65] vdd gnd cell_6t
Xbit_r66_c5 bl[5] br[5] wl[66] vdd gnd cell_6t
Xbit_r67_c5 bl[5] br[5] wl[67] vdd gnd cell_6t
Xbit_r68_c5 bl[5] br[5] wl[68] vdd gnd cell_6t
Xbit_r69_c5 bl[5] br[5] wl[69] vdd gnd cell_6t
Xbit_r70_c5 bl[5] br[5] wl[70] vdd gnd cell_6t
Xbit_r71_c5 bl[5] br[5] wl[71] vdd gnd cell_6t
Xbit_r72_c5 bl[5] br[5] wl[72] vdd gnd cell_6t
Xbit_r73_c5 bl[5] br[5] wl[73] vdd gnd cell_6t
Xbit_r74_c5 bl[5] br[5] wl[74] vdd gnd cell_6t
Xbit_r75_c5 bl[5] br[5] wl[75] vdd gnd cell_6t
Xbit_r76_c5 bl[5] br[5] wl[76] vdd gnd cell_6t
Xbit_r77_c5 bl[5] br[5] wl[77] vdd gnd cell_6t
Xbit_r78_c5 bl[5] br[5] wl[78] vdd gnd cell_6t
Xbit_r79_c5 bl[5] br[5] wl[79] vdd gnd cell_6t
Xbit_r80_c5 bl[5] br[5] wl[80] vdd gnd cell_6t
Xbit_r81_c5 bl[5] br[5] wl[81] vdd gnd cell_6t
Xbit_r82_c5 bl[5] br[5] wl[82] vdd gnd cell_6t
Xbit_r83_c5 bl[5] br[5] wl[83] vdd gnd cell_6t
Xbit_r84_c5 bl[5] br[5] wl[84] vdd gnd cell_6t
Xbit_r85_c5 bl[5] br[5] wl[85] vdd gnd cell_6t
Xbit_r86_c5 bl[5] br[5] wl[86] vdd gnd cell_6t
Xbit_r87_c5 bl[5] br[5] wl[87] vdd gnd cell_6t
Xbit_r88_c5 bl[5] br[5] wl[88] vdd gnd cell_6t
Xbit_r89_c5 bl[5] br[5] wl[89] vdd gnd cell_6t
Xbit_r90_c5 bl[5] br[5] wl[90] vdd gnd cell_6t
Xbit_r91_c5 bl[5] br[5] wl[91] vdd gnd cell_6t
Xbit_r92_c5 bl[5] br[5] wl[92] vdd gnd cell_6t
Xbit_r93_c5 bl[5] br[5] wl[93] vdd gnd cell_6t
Xbit_r94_c5 bl[5] br[5] wl[94] vdd gnd cell_6t
Xbit_r95_c5 bl[5] br[5] wl[95] vdd gnd cell_6t
Xbit_r96_c5 bl[5] br[5] wl[96] vdd gnd cell_6t
Xbit_r97_c5 bl[5] br[5] wl[97] vdd gnd cell_6t
Xbit_r98_c5 bl[5] br[5] wl[98] vdd gnd cell_6t
Xbit_r99_c5 bl[5] br[5] wl[99] vdd gnd cell_6t
Xbit_r100_c5 bl[5] br[5] wl[100] vdd gnd cell_6t
Xbit_r101_c5 bl[5] br[5] wl[101] vdd gnd cell_6t
Xbit_r102_c5 bl[5] br[5] wl[102] vdd gnd cell_6t
Xbit_r103_c5 bl[5] br[5] wl[103] vdd gnd cell_6t
Xbit_r104_c5 bl[5] br[5] wl[104] vdd gnd cell_6t
Xbit_r105_c5 bl[5] br[5] wl[105] vdd gnd cell_6t
Xbit_r106_c5 bl[5] br[5] wl[106] vdd gnd cell_6t
Xbit_r107_c5 bl[5] br[5] wl[107] vdd gnd cell_6t
Xbit_r108_c5 bl[5] br[5] wl[108] vdd gnd cell_6t
Xbit_r109_c5 bl[5] br[5] wl[109] vdd gnd cell_6t
Xbit_r110_c5 bl[5] br[5] wl[110] vdd gnd cell_6t
Xbit_r111_c5 bl[5] br[5] wl[111] vdd gnd cell_6t
Xbit_r112_c5 bl[5] br[5] wl[112] vdd gnd cell_6t
Xbit_r113_c5 bl[5] br[5] wl[113] vdd gnd cell_6t
Xbit_r114_c5 bl[5] br[5] wl[114] vdd gnd cell_6t
Xbit_r115_c5 bl[5] br[5] wl[115] vdd gnd cell_6t
Xbit_r116_c5 bl[5] br[5] wl[116] vdd gnd cell_6t
Xbit_r117_c5 bl[5] br[5] wl[117] vdd gnd cell_6t
Xbit_r118_c5 bl[5] br[5] wl[118] vdd gnd cell_6t
Xbit_r119_c5 bl[5] br[5] wl[119] vdd gnd cell_6t
Xbit_r120_c5 bl[5] br[5] wl[120] vdd gnd cell_6t
Xbit_r121_c5 bl[5] br[5] wl[121] vdd gnd cell_6t
Xbit_r122_c5 bl[5] br[5] wl[122] vdd gnd cell_6t
Xbit_r123_c5 bl[5] br[5] wl[123] vdd gnd cell_6t
Xbit_r124_c5 bl[5] br[5] wl[124] vdd gnd cell_6t
Xbit_r125_c5 bl[5] br[5] wl[125] vdd gnd cell_6t
Xbit_r126_c5 bl[5] br[5] wl[126] vdd gnd cell_6t
Xbit_r127_c5 bl[5] br[5] wl[127] vdd gnd cell_6t
Xbit_r128_c5 bl[5] br[5] wl[128] vdd gnd cell_6t
Xbit_r129_c5 bl[5] br[5] wl[129] vdd gnd cell_6t
Xbit_r130_c5 bl[5] br[5] wl[130] vdd gnd cell_6t
Xbit_r131_c5 bl[5] br[5] wl[131] vdd gnd cell_6t
Xbit_r132_c5 bl[5] br[5] wl[132] vdd gnd cell_6t
Xbit_r133_c5 bl[5] br[5] wl[133] vdd gnd cell_6t
Xbit_r134_c5 bl[5] br[5] wl[134] vdd gnd cell_6t
Xbit_r135_c5 bl[5] br[5] wl[135] vdd gnd cell_6t
Xbit_r136_c5 bl[5] br[5] wl[136] vdd gnd cell_6t
Xbit_r137_c5 bl[5] br[5] wl[137] vdd gnd cell_6t
Xbit_r138_c5 bl[5] br[5] wl[138] vdd gnd cell_6t
Xbit_r139_c5 bl[5] br[5] wl[139] vdd gnd cell_6t
Xbit_r140_c5 bl[5] br[5] wl[140] vdd gnd cell_6t
Xbit_r141_c5 bl[5] br[5] wl[141] vdd gnd cell_6t
Xbit_r142_c5 bl[5] br[5] wl[142] vdd gnd cell_6t
Xbit_r143_c5 bl[5] br[5] wl[143] vdd gnd cell_6t
Xbit_r144_c5 bl[5] br[5] wl[144] vdd gnd cell_6t
Xbit_r145_c5 bl[5] br[5] wl[145] vdd gnd cell_6t
Xbit_r146_c5 bl[5] br[5] wl[146] vdd gnd cell_6t
Xbit_r147_c5 bl[5] br[5] wl[147] vdd gnd cell_6t
Xbit_r148_c5 bl[5] br[5] wl[148] vdd gnd cell_6t
Xbit_r149_c5 bl[5] br[5] wl[149] vdd gnd cell_6t
Xbit_r150_c5 bl[5] br[5] wl[150] vdd gnd cell_6t
Xbit_r151_c5 bl[5] br[5] wl[151] vdd gnd cell_6t
Xbit_r152_c5 bl[5] br[5] wl[152] vdd gnd cell_6t
Xbit_r153_c5 bl[5] br[5] wl[153] vdd gnd cell_6t
Xbit_r154_c5 bl[5] br[5] wl[154] vdd gnd cell_6t
Xbit_r155_c5 bl[5] br[5] wl[155] vdd gnd cell_6t
Xbit_r156_c5 bl[5] br[5] wl[156] vdd gnd cell_6t
Xbit_r157_c5 bl[5] br[5] wl[157] vdd gnd cell_6t
Xbit_r158_c5 bl[5] br[5] wl[158] vdd gnd cell_6t
Xbit_r159_c5 bl[5] br[5] wl[159] vdd gnd cell_6t
Xbit_r160_c5 bl[5] br[5] wl[160] vdd gnd cell_6t
Xbit_r161_c5 bl[5] br[5] wl[161] vdd gnd cell_6t
Xbit_r162_c5 bl[5] br[5] wl[162] vdd gnd cell_6t
Xbit_r163_c5 bl[5] br[5] wl[163] vdd gnd cell_6t
Xbit_r164_c5 bl[5] br[5] wl[164] vdd gnd cell_6t
Xbit_r165_c5 bl[5] br[5] wl[165] vdd gnd cell_6t
Xbit_r166_c5 bl[5] br[5] wl[166] vdd gnd cell_6t
Xbit_r167_c5 bl[5] br[5] wl[167] vdd gnd cell_6t
Xbit_r168_c5 bl[5] br[5] wl[168] vdd gnd cell_6t
Xbit_r169_c5 bl[5] br[5] wl[169] vdd gnd cell_6t
Xbit_r170_c5 bl[5] br[5] wl[170] vdd gnd cell_6t
Xbit_r171_c5 bl[5] br[5] wl[171] vdd gnd cell_6t
Xbit_r172_c5 bl[5] br[5] wl[172] vdd gnd cell_6t
Xbit_r173_c5 bl[5] br[5] wl[173] vdd gnd cell_6t
Xbit_r174_c5 bl[5] br[5] wl[174] vdd gnd cell_6t
Xbit_r175_c5 bl[5] br[5] wl[175] vdd gnd cell_6t
Xbit_r176_c5 bl[5] br[5] wl[176] vdd gnd cell_6t
Xbit_r177_c5 bl[5] br[5] wl[177] vdd gnd cell_6t
Xbit_r178_c5 bl[5] br[5] wl[178] vdd gnd cell_6t
Xbit_r179_c5 bl[5] br[5] wl[179] vdd gnd cell_6t
Xbit_r180_c5 bl[5] br[5] wl[180] vdd gnd cell_6t
Xbit_r181_c5 bl[5] br[5] wl[181] vdd gnd cell_6t
Xbit_r182_c5 bl[5] br[5] wl[182] vdd gnd cell_6t
Xbit_r183_c5 bl[5] br[5] wl[183] vdd gnd cell_6t
Xbit_r184_c5 bl[5] br[5] wl[184] vdd gnd cell_6t
Xbit_r185_c5 bl[5] br[5] wl[185] vdd gnd cell_6t
Xbit_r186_c5 bl[5] br[5] wl[186] vdd gnd cell_6t
Xbit_r187_c5 bl[5] br[5] wl[187] vdd gnd cell_6t
Xbit_r188_c5 bl[5] br[5] wl[188] vdd gnd cell_6t
Xbit_r189_c5 bl[5] br[5] wl[189] vdd gnd cell_6t
Xbit_r190_c5 bl[5] br[5] wl[190] vdd gnd cell_6t
Xbit_r191_c5 bl[5] br[5] wl[191] vdd gnd cell_6t
Xbit_r192_c5 bl[5] br[5] wl[192] vdd gnd cell_6t
Xbit_r193_c5 bl[5] br[5] wl[193] vdd gnd cell_6t
Xbit_r194_c5 bl[5] br[5] wl[194] vdd gnd cell_6t
Xbit_r195_c5 bl[5] br[5] wl[195] vdd gnd cell_6t
Xbit_r196_c5 bl[5] br[5] wl[196] vdd gnd cell_6t
Xbit_r197_c5 bl[5] br[5] wl[197] vdd gnd cell_6t
Xbit_r198_c5 bl[5] br[5] wl[198] vdd gnd cell_6t
Xbit_r199_c5 bl[5] br[5] wl[199] vdd gnd cell_6t
Xbit_r200_c5 bl[5] br[5] wl[200] vdd gnd cell_6t
Xbit_r201_c5 bl[5] br[5] wl[201] vdd gnd cell_6t
Xbit_r202_c5 bl[5] br[5] wl[202] vdd gnd cell_6t
Xbit_r203_c5 bl[5] br[5] wl[203] vdd gnd cell_6t
Xbit_r204_c5 bl[5] br[5] wl[204] vdd gnd cell_6t
Xbit_r205_c5 bl[5] br[5] wl[205] vdd gnd cell_6t
Xbit_r206_c5 bl[5] br[5] wl[206] vdd gnd cell_6t
Xbit_r207_c5 bl[5] br[5] wl[207] vdd gnd cell_6t
Xbit_r208_c5 bl[5] br[5] wl[208] vdd gnd cell_6t
Xbit_r209_c5 bl[5] br[5] wl[209] vdd gnd cell_6t
Xbit_r210_c5 bl[5] br[5] wl[210] vdd gnd cell_6t
Xbit_r211_c5 bl[5] br[5] wl[211] vdd gnd cell_6t
Xbit_r212_c5 bl[5] br[5] wl[212] vdd gnd cell_6t
Xbit_r213_c5 bl[5] br[5] wl[213] vdd gnd cell_6t
Xbit_r214_c5 bl[5] br[5] wl[214] vdd gnd cell_6t
Xbit_r215_c5 bl[5] br[5] wl[215] vdd gnd cell_6t
Xbit_r216_c5 bl[5] br[5] wl[216] vdd gnd cell_6t
Xbit_r217_c5 bl[5] br[5] wl[217] vdd gnd cell_6t
Xbit_r218_c5 bl[5] br[5] wl[218] vdd gnd cell_6t
Xbit_r219_c5 bl[5] br[5] wl[219] vdd gnd cell_6t
Xbit_r220_c5 bl[5] br[5] wl[220] vdd gnd cell_6t
Xbit_r221_c5 bl[5] br[5] wl[221] vdd gnd cell_6t
Xbit_r222_c5 bl[5] br[5] wl[222] vdd gnd cell_6t
Xbit_r223_c5 bl[5] br[5] wl[223] vdd gnd cell_6t
Xbit_r224_c5 bl[5] br[5] wl[224] vdd gnd cell_6t
Xbit_r225_c5 bl[5] br[5] wl[225] vdd gnd cell_6t
Xbit_r226_c5 bl[5] br[5] wl[226] vdd gnd cell_6t
Xbit_r227_c5 bl[5] br[5] wl[227] vdd gnd cell_6t
Xbit_r228_c5 bl[5] br[5] wl[228] vdd gnd cell_6t
Xbit_r229_c5 bl[5] br[5] wl[229] vdd gnd cell_6t
Xbit_r230_c5 bl[5] br[5] wl[230] vdd gnd cell_6t
Xbit_r231_c5 bl[5] br[5] wl[231] vdd gnd cell_6t
Xbit_r232_c5 bl[5] br[5] wl[232] vdd gnd cell_6t
Xbit_r233_c5 bl[5] br[5] wl[233] vdd gnd cell_6t
Xbit_r234_c5 bl[5] br[5] wl[234] vdd gnd cell_6t
Xbit_r235_c5 bl[5] br[5] wl[235] vdd gnd cell_6t
Xbit_r236_c5 bl[5] br[5] wl[236] vdd gnd cell_6t
Xbit_r237_c5 bl[5] br[5] wl[237] vdd gnd cell_6t
Xbit_r238_c5 bl[5] br[5] wl[238] vdd gnd cell_6t
Xbit_r239_c5 bl[5] br[5] wl[239] vdd gnd cell_6t
Xbit_r240_c5 bl[5] br[5] wl[240] vdd gnd cell_6t
Xbit_r241_c5 bl[5] br[5] wl[241] vdd gnd cell_6t
Xbit_r242_c5 bl[5] br[5] wl[242] vdd gnd cell_6t
Xbit_r243_c5 bl[5] br[5] wl[243] vdd gnd cell_6t
Xbit_r244_c5 bl[5] br[5] wl[244] vdd gnd cell_6t
Xbit_r245_c5 bl[5] br[5] wl[245] vdd gnd cell_6t
Xbit_r246_c5 bl[5] br[5] wl[246] vdd gnd cell_6t
Xbit_r247_c5 bl[5] br[5] wl[247] vdd gnd cell_6t
Xbit_r248_c5 bl[5] br[5] wl[248] vdd gnd cell_6t
Xbit_r249_c5 bl[5] br[5] wl[249] vdd gnd cell_6t
Xbit_r250_c5 bl[5] br[5] wl[250] vdd gnd cell_6t
Xbit_r251_c5 bl[5] br[5] wl[251] vdd gnd cell_6t
Xbit_r252_c5 bl[5] br[5] wl[252] vdd gnd cell_6t
Xbit_r253_c5 bl[5] br[5] wl[253] vdd gnd cell_6t
Xbit_r254_c5 bl[5] br[5] wl[254] vdd gnd cell_6t
Xbit_r255_c5 bl[5] br[5] wl[255] vdd gnd cell_6t
Xbit_r0_c6 bl[6] br[6] wl[0] vdd gnd cell_6t
Xbit_r1_c6 bl[6] br[6] wl[1] vdd gnd cell_6t
Xbit_r2_c6 bl[6] br[6] wl[2] vdd gnd cell_6t
Xbit_r3_c6 bl[6] br[6] wl[3] vdd gnd cell_6t
Xbit_r4_c6 bl[6] br[6] wl[4] vdd gnd cell_6t
Xbit_r5_c6 bl[6] br[6] wl[5] vdd gnd cell_6t
Xbit_r6_c6 bl[6] br[6] wl[6] vdd gnd cell_6t
Xbit_r7_c6 bl[6] br[6] wl[7] vdd gnd cell_6t
Xbit_r8_c6 bl[6] br[6] wl[8] vdd gnd cell_6t
Xbit_r9_c6 bl[6] br[6] wl[9] vdd gnd cell_6t
Xbit_r10_c6 bl[6] br[6] wl[10] vdd gnd cell_6t
Xbit_r11_c6 bl[6] br[6] wl[11] vdd gnd cell_6t
Xbit_r12_c6 bl[6] br[6] wl[12] vdd gnd cell_6t
Xbit_r13_c6 bl[6] br[6] wl[13] vdd gnd cell_6t
Xbit_r14_c6 bl[6] br[6] wl[14] vdd gnd cell_6t
Xbit_r15_c6 bl[6] br[6] wl[15] vdd gnd cell_6t
Xbit_r16_c6 bl[6] br[6] wl[16] vdd gnd cell_6t
Xbit_r17_c6 bl[6] br[6] wl[17] vdd gnd cell_6t
Xbit_r18_c6 bl[6] br[6] wl[18] vdd gnd cell_6t
Xbit_r19_c6 bl[6] br[6] wl[19] vdd gnd cell_6t
Xbit_r20_c6 bl[6] br[6] wl[20] vdd gnd cell_6t
Xbit_r21_c6 bl[6] br[6] wl[21] vdd gnd cell_6t
Xbit_r22_c6 bl[6] br[6] wl[22] vdd gnd cell_6t
Xbit_r23_c6 bl[6] br[6] wl[23] vdd gnd cell_6t
Xbit_r24_c6 bl[6] br[6] wl[24] vdd gnd cell_6t
Xbit_r25_c6 bl[6] br[6] wl[25] vdd gnd cell_6t
Xbit_r26_c6 bl[6] br[6] wl[26] vdd gnd cell_6t
Xbit_r27_c6 bl[6] br[6] wl[27] vdd gnd cell_6t
Xbit_r28_c6 bl[6] br[6] wl[28] vdd gnd cell_6t
Xbit_r29_c6 bl[6] br[6] wl[29] vdd gnd cell_6t
Xbit_r30_c6 bl[6] br[6] wl[30] vdd gnd cell_6t
Xbit_r31_c6 bl[6] br[6] wl[31] vdd gnd cell_6t
Xbit_r32_c6 bl[6] br[6] wl[32] vdd gnd cell_6t
Xbit_r33_c6 bl[6] br[6] wl[33] vdd gnd cell_6t
Xbit_r34_c6 bl[6] br[6] wl[34] vdd gnd cell_6t
Xbit_r35_c6 bl[6] br[6] wl[35] vdd gnd cell_6t
Xbit_r36_c6 bl[6] br[6] wl[36] vdd gnd cell_6t
Xbit_r37_c6 bl[6] br[6] wl[37] vdd gnd cell_6t
Xbit_r38_c6 bl[6] br[6] wl[38] vdd gnd cell_6t
Xbit_r39_c6 bl[6] br[6] wl[39] vdd gnd cell_6t
Xbit_r40_c6 bl[6] br[6] wl[40] vdd gnd cell_6t
Xbit_r41_c6 bl[6] br[6] wl[41] vdd gnd cell_6t
Xbit_r42_c6 bl[6] br[6] wl[42] vdd gnd cell_6t
Xbit_r43_c6 bl[6] br[6] wl[43] vdd gnd cell_6t
Xbit_r44_c6 bl[6] br[6] wl[44] vdd gnd cell_6t
Xbit_r45_c6 bl[6] br[6] wl[45] vdd gnd cell_6t
Xbit_r46_c6 bl[6] br[6] wl[46] vdd gnd cell_6t
Xbit_r47_c6 bl[6] br[6] wl[47] vdd gnd cell_6t
Xbit_r48_c6 bl[6] br[6] wl[48] vdd gnd cell_6t
Xbit_r49_c6 bl[6] br[6] wl[49] vdd gnd cell_6t
Xbit_r50_c6 bl[6] br[6] wl[50] vdd gnd cell_6t
Xbit_r51_c6 bl[6] br[6] wl[51] vdd gnd cell_6t
Xbit_r52_c6 bl[6] br[6] wl[52] vdd gnd cell_6t
Xbit_r53_c6 bl[6] br[6] wl[53] vdd gnd cell_6t
Xbit_r54_c6 bl[6] br[6] wl[54] vdd gnd cell_6t
Xbit_r55_c6 bl[6] br[6] wl[55] vdd gnd cell_6t
Xbit_r56_c6 bl[6] br[6] wl[56] vdd gnd cell_6t
Xbit_r57_c6 bl[6] br[6] wl[57] vdd gnd cell_6t
Xbit_r58_c6 bl[6] br[6] wl[58] vdd gnd cell_6t
Xbit_r59_c6 bl[6] br[6] wl[59] vdd gnd cell_6t
Xbit_r60_c6 bl[6] br[6] wl[60] vdd gnd cell_6t
Xbit_r61_c6 bl[6] br[6] wl[61] vdd gnd cell_6t
Xbit_r62_c6 bl[6] br[6] wl[62] vdd gnd cell_6t
Xbit_r63_c6 bl[6] br[6] wl[63] vdd gnd cell_6t
Xbit_r64_c6 bl[6] br[6] wl[64] vdd gnd cell_6t
Xbit_r65_c6 bl[6] br[6] wl[65] vdd gnd cell_6t
Xbit_r66_c6 bl[6] br[6] wl[66] vdd gnd cell_6t
Xbit_r67_c6 bl[6] br[6] wl[67] vdd gnd cell_6t
Xbit_r68_c6 bl[6] br[6] wl[68] vdd gnd cell_6t
Xbit_r69_c6 bl[6] br[6] wl[69] vdd gnd cell_6t
Xbit_r70_c6 bl[6] br[6] wl[70] vdd gnd cell_6t
Xbit_r71_c6 bl[6] br[6] wl[71] vdd gnd cell_6t
Xbit_r72_c6 bl[6] br[6] wl[72] vdd gnd cell_6t
Xbit_r73_c6 bl[6] br[6] wl[73] vdd gnd cell_6t
Xbit_r74_c6 bl[6] br[6] wl[74] vdd gnd cell_6t
Xbit_r75_c6 bl[6] br[6] wl[75] vdd gnd cell_6t
Xbit_r76_c6 bl[6] br[6] wl[76] vdd gnd cell_6t
Xbit_r77_c6 bl[6] br[6] wl[77] vdd gnd cell_6t
Xbit_r78_c6 bl[6] br[6] wl[78] vdd gnd cell_6t
Xbit_r79_c6 bl[6] br[6] wl[79] vdd gnd cell_6t
Xbit_r80_c6 bl[6] br[6] wl[80] vdd gnd cell_6t
Xbit_r81_c6 bl[6] br[6] wl[81] vdd gnd cell_6t
Xbit_r82_c6 bl[6] br[6] wl[82] vdd gnd cell_6t
Xbit_r83_c6 bl[6] br[6] wl[83] vdd gnd cell_6t
Xbit_r84_c6 bl[6] br[6] wl[84] vdd gnd cell_6t
Xbit_r85_c6 bl[6] br[6] wl[85] vdd gnd cell_6t
Xbit_r86_c6 bl[6] br[6] wl[86] vdd gnd cell_6t
Xbit_r87_c6 bl[6] br[6] wl[87] vdd gnd cell_6t
Xbit_r88_c6 bl[6] br[6] wl[88] vdd gnd cell_6t
Xbit_r89_c6 bl[6] br[6] wl[89] vdd gnd cell_6t
Xbit_r90_c6 bl[6] br[6] wl[90] vdd gnd cell_6t
Xbit_r91_c6 bl[6] br[6] wl[91] vdd gnd cell_6t
Xbit_r92_c6 bl[6] br[6] wl[92] vdd gnd cell_6t
Xbit_r93_c6 bl[6] br[6] wl[93] vdd gnd cell_6t
Xbit_r94_c6 bl[6] br[6] wl[94] vdd gnd cell_6t
Xbit_r95_c6 bl[6] br[6] wl[95] vdd gnd cell_6t
Xbit_r96_c6 bl[6] br[6] wl[96] vdd gnd cell_6t
Xbit_r97_c6 bl[6] br[6] wl[97] vdd gnd cell_6t
Xbit_r98_c6 bl[6] br[6] wl[98] vdd gnd cell_6t
Xbit_r99_c6 bl[6] br[6] wl[99] vdd gnd cell_6t
Xbit_r100_c6 bl[6] br[6] wl[100] vdd gnd cell_6t
Xbit_r101_c6 bl[6] br[6] wl[101] vdd gnd cell_6t
Xbit_r102_c6 bl[6] br[6] wl[102] vdd gnd cell_6t
Xbit_r103_c6 bl[6] br[6] wl[103] vdd gnd cell_6t
Xbit_r104_c6 bl[6] br[6] wl[104] vdd gnd cell_6t
Xbit_r105_c6 bl[6] br[6] wl[105] vdd gnd cell_6t
Xbit_r106_c6 bl[6] br[6] wl[106] vdd gnd cell_6t
Xbit_r107_c6 bl[6] br[6] wl[107] vdd gnd cell_6t
Xbit_r108_c6 bl[6] br[6] wl[108] vdd gnd cell_6t
Xbit_r109_c6 bl[6] br[6] wl[109] vdd gnd cell_6t
Xbit_r110_c6 bl[6] br[6] wl[110] vdd gnd cell_6t
Xbit_r111_c6 bl[6] br[6] wl[111] vdd gnd cell_6t
Xbit_r112_c6 bl[6] br[6] wl[112] vdd gnd cell_6t
Xbit_r113_c6 bl[6] br[6] wl[113] vdd gnd cell_6t
Xbit_r114_c6 bl[6] br[6] wl[114] vdd gnd cell_6t
Xbit_r115_c6 bl[6] br[6] wl[115] vdd gnd cell_6t
Xbit_r116_c6 bl[6] br[6] wl[116] vdd gnd cell_6t
Xbit_r117_c6 bl[6] br[6] wl[117] vdd gnd cell_6t
Xbit_r118_c6 bl[6] br[6] wl[118] vdd gnd cell_6t
Xbit_r119_c6 bl[6] br[6] wl[119] vdd gnd cell_6t
Xbit_r120_c6 bl[6] br[6] wl[120] vdd gnd cell_6t
Xbit_r121_c6 bl[6] br[6] wl[121] vdd gnd cell_6t
Xbit_r122_c6 bl[6] br[6] wl[122] vdd gnd cell_6t
Xbit_r123_c6 bl[6] br[6] wl[123] vdd gnd cell_6t
Xbit_r124_c6 bl[6] br[6] wl[124] vdd gnd cell_6t
Xbit_r125_c6 bl[6] br[6] wl[125] vdd gnd cell_6t
Xbit_r126_c6 bl[6] br[6] wl[126] vdd gnd cell_6t
Xbit_r127_c6 bl[6] br[6] wl[127] vdd gnd cell_6t
Xbit_r128_c6 bl[6] br[6] wl[128] vdd gnd cell_6t
Xbit_r129_c6 bl[6] br[6] wl[129] vdd gnd cell_6t
Xbit_r130_c6 bl[6] br[6] wl[130] vdd gnd cell_6t
Xbit_r131_c6 bl[6] br[6] wl[131] vdd gnd cell_6t
Xbit_r132_c6 bl[6] br[6] wl[132] vdd gnd cell_6t
Xbit_r133_c6 bl[6] br[6] wl[133] vdd gnd cell_6t
Xbit_r134_c6 bl[6] br[6] wl[134] vdd gnd cell_6t
Xbit_r135_c6 bl[6] br[6] wl[135] vdd gnd cell_6t
Xbit_r136_c6 bl[6] br[6] wl[136] vdd gnd cell_6t
Xbit_r137_c6 bl[6] br[6] wl[137] vdd gnd cell_6t
Xbit_r138_c6 bl[6] br[6] wl[138] vdd gnd cell_6t
Xbit_r139_c6 bl[6] br[6] wl[139] vdd gnd cell_6t
Xbit_r140_c6 bl[6] br[6] wl[140] vdd gnd cell_6t
Xbit_r141_c6 bl[6] br[6] wl[141] vdd gnd cell_6t
Xbit_r142_c6 bl[6] br[6] wl[142] vdd gnd cell_6t
Xbit_r143_c6 bl[6] br[6] wl[143] vdd gnd cell_6t
Xbit_r144_c6 bl[6] br[6] wl[144] vdd gnd cell_6t
Xbit_r145_c6 bl[6] br[6] wl[145] vdd gnd cell_6t
Xbit_r146_c6 bl[6] br[6] wl[146] vdd gnd cell_6t
Xbit_r147_c6 bl[6] br[6] wl[147] vdd gnd cell_6t
Xbit_r148_c6 bl[6] br[6] wl[148] vdd gnd cell_6t
Xbit_r149_c6 bl[6] br[6] wl[149] vdd gnd cell_6t
Xbit_r150_c6 bl[6] br[6] wl[150] vdd gnd cell_6t
Xbit_r151_c6 bl[6] br[6] wl[151] vdd gnd cell_6t
Xbit_r152_c6 bl[6] br[6] wl[152] vdd gnd cell_6t
Xbit_r153_c6 bl[6] br[6] wl[153] vdd gnd cell_6t
Xbit_r154_c6 bl[6] br[6] wl[154] vdd gnd cell_6t
Xbit_r155_c6 bl[6] br[6] wl[155] vdd gnd cell_6t
Xbit_r156_c6 bl[6] br[6] wl[156] vdd gnd cell_6t
Xbit_r157_c6 bl[6] br[6] wl[157] vdd gnd cell_6t
Xbit_r158_c6 bl[6] br[6] wl[158] vdd gnd cell_6t
Xbit_r159_c6 bl[6] br[6] wl[159] vdd gnd cell_6t
Xbit_r160_c6 bl[6] br[6] wl[160] vdd gnd cell_6t
Xbit_r161_c6 bl[6] br[6] wl[161] vdd gnd cell_6t
Xbit_r162_c6 bl[6] br[6] wl[162] vdd gnd cell_6t
Xbit_r163_c6 bl[6] br[6] wl[163] vdd gnd cell_6t
Xbit_r164_c6 bl[6] br[6] wl[164] vdd gnd cell_6t
Xbit_r165_c6 bl[6] br[6] wl[165] vdd gnd cell_6t
Xbit_r166_c6 bl[6] br[6] wl[166] vdd gnd cell_6t
Xbit_r167_c6 bl[6] br[6] wl[167] vdd gnd cell_6t
Xbit_r168_c6 bl[6] br[6] wl[168] vdd gnd cell_6t
Xbit_r169_c6 bl[6] br[6] wl[169] vdd gnd cell_6t
Xbit_r170_c6 bl[6] br[6] wl[170] vdd gnd cell_6t
Xbit_r171_c6 bl[6] br[6] wl[171] vdd gnd cell_6t
Xbit_r172_c6 bl[6] br[6] wl[172] vdd gnd cell_6t
Xbit_r173_c6 bl[6] br[6] wl[173] vdd gnd cell_6t
Xbit_r174_c6 bl[6] br[6] wl[174] vdd gnd cell_6t
Xbit_r175_c6 bl[6] br[6] wl[175] vdd gnd cell_6t
Xbit_r176_c6 bl[6] br[6] wl[176] vdd gnd cell_6t
Xbit_r177_c6 bl[6] br[6] wl[177] vdd gnd cell_6t
Xbit_r178_c6 bl[6] br[6] wl[178] vdd gnd cell_6t
Xbit_r179_c6 bl[6] br[6] wl[179] vdd gnd cell_6t
Xbit_r180_c6 bl[6] br[6] wl[180] vdd gnd cell_6t
Xbit_r181_c6 bl[6] br[6] wl[181] vdd gnd cell_6t
Xbit_r182_c6 bl[6] br[6] wl[182] vdd gnd cell_6t
Xbit_r183_c6 bl[6] br[6] wl[183] vdd gnd cell_6t
Xbit_r184_c6 bl[6] br[6] wl[184] vdd gnd cell_6t
Xbit_r185_c6 bl[6] br[6] wl[185] vdd gnd cell_6t
Xbit_r186_c6 bl[6] br[6] wl[186] vdd gnd cell_6t
Xbit_r187_c6 bl[6] br[6] wl[187] vdd gnd cell_6t
Xbit_r188_c6 bl[6] br[6] wl[188] vdd gnd cell_6t
Xbit_r189_c6 bl[6] br[6] wl[189] vdd gnd cell_6t
Xbit_r190_c6 bl[6] br[6] wl[190] vdd gnd cell_6t
Xbit_r191_c6 bl[6] br[6] wl[191] vdd gnd cell_6t
Xbit_r192_c6 bl[6] br[6] wl[192] vdd gnd cell_6t
Xbit_r193_c6 bl[6] br[6] wl[193] vdd gnd cell_6t
Xbit_r194_c6 bl[6] br[6] wl[194] vdd gnd cell_6t
Xbit_r195_c6 bl[6] br[6] wl[195] vdd gnd cell_6t
Xbit_r196_c6 bl[6] br[6] wl[196] vdd gnd cell_6t
Xbit_r197_c6 bl[6] br[6] wl[197] vdd gnd cell_6t
Xbit_r198_c6 bl[6] br[6] wl[198] vdd gnd cell_6t
Xbit_r199_c6 bl[6] br[6] wl[199] vdd gnd cell_6t
Xbit_r200_c6 bl[6] br[6] wl[200] vdd gnd cell_6t
Xbit_r201_c6 bl[6] br[6] wl[201] vdd gnd cell_6t
Xbit_r202_c6 bl[6] br[6] wl[202] vdd gnd cell_6t
Xbit_r203_c6 bl[6] br[6] wl[203] vdd gnd cell_6t
Xbit_r204_c6 bl[6] br[6] wl[204] vdd gnd cell_6t
Xbit_r205_c6 bl[6] br[6] wl[205] vdd gnd cell_6t
Xbit_r206_c6 bl[6] br[6] wl[206] vdd gnd cell_6t
Xbit_r207_c6 bl[6] br[6] wl[207] vdd gnd cell_6t
Xbit_r208_c6 bl[6] br[6] wl[208] vdd gnd cell_6t
Xbit_r209_c6 bl[6] br[6] wl[209] vdd gnd cell_6t
Xbit_r210_c6 bl[6] br[6] wl[210] vdd gnd cell_6t
Xbit_r211_c6 bl[6] br[6] wl[211] vdd gnd cell_6t
Xbit_r212_c6 bl[6] br[6] wl[212] vdd gnd cell_6t
Xbit_r213_c6 bl[6] br[6] wl[213] vdd gnd cell_6t
Xbit_r214_c6 bl[6] br[6] wl[214] vdd gnd cell_6t
Xbit_r215_c6 bl[6] br[6] wl[215] vdd gnd cell_6t
Xbit_r216_c6 bl[6] br[6] wl[216] vdd gnd cell_6t
Xbit_r217_c6 bl[6] br[6] wl[217] vdd gnd cell_6t
Xbit_r218_c6 bl[6] br[6] wl[218] vdd gnd cell_6t
Xbit_r219_c6 bl[6] br[6] wl[219] vdd gnd cell_6t
Xbit_r220_c6 bl[6] br[6] wl[220] vdd gnd cell_6t
Xbit_r221_c6 bl[6] br[6] wl[221] vdd gnd cell_6t
Xbit_r222_c6 bl[6] br[6] wl[222] vdd gnd cell_6t
Xbit_r223_c6 bl[6] br[6] wl[223] vdd gnd cell_6t
Xbit_r224_c6 bl[6] br[6] wl[224] vdd gnd cell_6t
Xbit_r225_c6 bl[6] br[6] wl[225] vdd gnd cell_6t
Xbit_r226_c6 bl[6] br[6] wl[226] vdd gnd cell_6t
Xbit_r227_c6 bl[6] br[6] wl[227] vdd gnd cell_6t
Xbit_r228_c6 bl[6] br[6] wl[228] vdd gnd cell_6t
Xbit_r229_c6 bl[6] br[6] wl[229] vdd gnd cell_6t
Xbit_r230_c6 bl[6] br[6] wl[230] vdd gnd cell_6t
Xbit_r231_c6 bl[6] br[6] wl[231] vdd gnd cell_6t
Xbit_r232_c6 bl[6] br[6] wl[232] vdd gnd cell_6t
Xbit_r233_c6 bl[6] br[6] wl[233] vdd gnd cell_6t
Xbit_r234_c6 bl[6] br[6] wl[234] vdd gnd cell_6t
Xbit_r235_c6 bl[6] br[6] wl[235] vdd gnd cell_6t
Xbit_r236_c6 bl[6] br[6] wl[236] vdd gnd cell_6t
Xbit_r237_c6 bl[6] br[6] wl[237] vdd gnd cell_6t
Xbit_r238_c6 bl[6] br[6] wl[238] vdd gnd cell_6t
Xbit_r239_c6 bl[6] br[6] wl[239] vdd gnd cell_6t
Xbit_r240_c6 bl[6] br[6] wl[240] vdd gnd cell_6t
Xbit_r241_c6 bl[6] br[6] wl[241] vdd gnd cell_6t
Xbit_r242_c6 bl[6] br[6] wl[242] vdd gnd cell_6t
Xbit_r243_c6 bl[6] br[6] wl[243] vdd gnd cell_6t
Xbit_r244_c6 bl[6] br[6] wl[244] vdd gnd cell_6t
Xbit_r245_c6 bl[6] br[6] wl[245] vdd gnd cell_6t
Xbit_r246_c6 bl[6] br[6] wl[246] vdd gnd cell_6t
Xbit_r247_c6 bl[6] br[6] wl[247] vdd gnd cell_6t
Xbit_r248_c6 bl[6] br[6] wl[248] vdd gnd cell_6t
Xbit_r249_c6 bl[6] br[6] wl[249] vdd gnd cell_6t
Xbit_r250_c6 bl[6] br[6] wl[250] vdd gnd cell_6t
Xbit_r251_c6 bl[6] br[6] wl[251] vdd gnd cell_6t
Xbit_r252_c6 bl[6] br[6] wl[252] vdd gnd cell_6t
Xbit_r253_c6 bl[6] br[6] wl[253] vdd gnd cell_6t
Xbit_r254_c6 bl[6] br[6] wl[254] vdd gnd cell_6t
Xbit_r255_c6 bl[6] br[6] wl[255] vdd gnd cell_6t
Xbit_r0_c7 bl[7] br[7] wl[0] vdd gnd cell_6t
Xbit_r1_c7 bl[7] br[7] wl[1] vdd gnd cell_6t
Xbit_r2_c7 bl[7] br[7] wl[2] vdd gnd cell_6t
Xbit_r3_c7 bl[7] br[7] wl[3] vdd gnd cell_6t
Xbit_r4_c7 bl[7] br[7] wl[4] vdd gnd cell_6t
Xbit_r5_c7 bl[7] br[7] wl[5] vdd gnd cell_6t
Xbit_r6_c7 bl[7] br[7] wl[6] vdd gnd cell_6t
Xbit_r7_c7 bl[7] br[7] wl[7] vdd gnd cell_6t
Xbit_r8_c7 bl[7] br[7] wl[8] vdd gnd cell_6t
Xbit_r9_c7 bl[7] br[7] wl[9] vdd gnd cell_6t
Xbit_r10_c7 bl[7] br[7] wl[10] vdd gnd cell_6t
Xbit_r11_c7 bl[7] br[7] wl[11] vdd gnd cell_6t
Xbit_r12_c7 bl[7] br[7] wl[12] vdd gnd cell_6t
Xbit_r13_c7 bl[7] br[7] wl[13] vdd gnd cell_6t
Xbit_r14_c7 bl[7] br[7] wl[14] vdd gnd cell_6t
Xbit_r15_c7 bl[7] br[7] wl[15] vdd gnd cell_6t
Xbit_r16_c7 bl[7] br[7] wl[16] vdd gnd cell_6t
Xbit_r17_c7 bl[7] br[7] wl[17] vdd gnd cell_6t
Xbit_r18_c7 bl[7] br[7] wl[18] vdd gnd cell_6t
Xbit_r19_c7 bl[7] br[7] wl[19] vdd gnd cell_6t
Xbit_r20_c7 bl[7] br[7] wl[20] vdd gnd cell_6t
Xbit_r21_c7 bl[7] br[7] wl[21] vdd gnd cell_6t
Xbit_r22_c7 bl[7] br[7] wl[22] vdd gnd cell_6t
Xbit_r23_c7 bl[7] br[7] wl[23] vdd gnd cell_6t
Xbit_r24_c7 bl[7] br[7] wl[24] vdd gnd cell_6t
Xbit_r25_c7 bl[7] br[7] wl[25] vdd gnd cell_6t
Xbit_r26_c7 bl[7] br[7] wl[26] vdd gnd cell_6t
Xbit_r27_c7 bl[7] br[7] wl[27] vdd gnd cell_6t
Xbit_r28_c7 bl[7] br[7] wl[28] vdd gnd cell_6t
Xbit_r29_c7 bl[7] br[7] wl[29] vdd gnd cell_6t
Xbit_r30_c7 bl[7] br[7] wl[30] vdd gnd cell_6t
Xbit_r31_c7 bl[7] br[7] wl[31] vdd gnd cell_6t
Xbit_r32_c7 bl[7] br[7] wl[32] vdd gnd cell_6t
Xbit_r33_c7 bl[7] br[7] wl[33] vdd gnd cell_6t
Xbit_r34_c7 bl[7] br[7] wl[34] vdd gnd cell_6t
Xbit_r35_c7 bl[7] br[7] wl[35] vdd gnd cell_6t
Xbit_r36_c7 bl[7] br[7] wl[36] vdd gnd cell_6t
Xbit_r37_c7 bl[7] br[7] wl[37] vdd gnd cell_6t
Xbit_r38_c7 bl[7] br[7] wl[38] vdd gnd cell_6t
Xbit_r39_c7 bl[7] br[7] wl[39] vdd gnd cell_6t
Xbit_r40_c7 bl[7] br[7] wl[40] vdd gnd cell_6t
Xbit_r41_c7 bl[7] br[7] wl[41] vdd gnd cell_6t
Xbit_r42_c7 bl[7] br[7] wl[42] vdd gnd cell_6t
Xbit_r43_c7 bl[7] br[7] wl[43] vdd gnd cell_6t
Xbit_r44_c7 bl[7] br[7] wl[44] vdd gnd cell_6t
Xbit_r45_c7 bl[7] br[7] wl[45] vdd gnd cell_6t
Xbit_r46_c7 bl[7] br[7] wl[46] vdd gnd cell_6t
Xbit_r47_c7 bl[7] br[7] wl[47] vdd gnd cell_6t
Xbit_r48_c7 bl[7] br[7] wl[48] vdd gnd cell_6t
Xbit_r49_c7 bl[7] br[7] wl[49] vdd gnd cell_6t
Xbit_r50_c7 bl[7] br[7] wl[50] vdd gnd cell_6t
Xbit_r51_c7 bl[7] br[7] wl[51] vdd gnd cell_6t
Xbit_r52_c7 bl[7] br[7] wl[52] vdd gnd cell_6t
Xbit_r53_c7 bl[7] br[7] wl[53] vdd gnd cell_6t
Xbit_r54_c7 bl[7] br[7] wl[54] vdd gnd cell_6t
Xbit_r55_c7 bl[7] br[7] wl[55] vdd gnd cell_6t
Xbit_r56_c7 bl[7] br[7] wl[56] vdd gnd cell_6t
Xbit_r57_c7 bl[7] br[7] wl[57] vdd gnd cell_6t
Xbit_r58_c7 bl[7] br[7] wl[58] vdd gnd cell_6t
Xbit_r59_c7 bl[7] br[7] wl[59] vdd gnd cell_6t
Xbit_r60_c7 bl[7] br[7] wl[60] vdd gnd cell_6t
Xbit_r61_c7 bl[7] br[7] wl[61] vdd gnd cell_6t
Xbit_r62_c7 bl[7] br[7] wl[62] vdd gnd cell_6t
Xbit_r63_c7 bl[7] br[7] wl[63] vdd gnd cell_6t
Xbit_r64_c7 bl[7] br[7] wl[64] vdd gnd cell_6t
Xbit_r65_c7 bl[7] br[7] wl[65] vdd gnd cell_6t
Xbit_r66_c7 bl[7] br[7] wl[66] vdd gnd cell_6t
Xbit_r67_c7 bl[7] br[7] wl[67] vdd gnd cell_6t
Xbit_r68_c7 bl[7] br[7] wl[68] vdd gnd cell_6t
Xbit_r69_c7 bl[7] br[7] wl[69] vdd gnd cell_6t
Xbit_r70_c7 bl[7] br[7] wl[70] vdd gnd cell_6t
Xbit_r71_c7 bl[7] br[7] wl[71] vdd gnd cell_6t
Xbit_r72_c7 bl[7] br[7] wl[72] vdd gnd cell_6t
Xbit_r73_c7 bl[7] br[7] wl[73] vdd gnd cell_6t
Xbit_r74_c7 bl[7] br[7] wl[74] vdd gnd cell_6t
Xbit_r75_c7 bl[7] br[7] wl[75] vdd gnd cell_6t
Xbit_r76_c7 bl[7] br[7] wl[76] vdd gnd cell_6t
Xbit_r77_c7 bl[7] br[7] wl[77] vdd gnd cell_6t
Xbit_r78_c7 bl[7] br[7] wl[78] vdd gnd cell_6t
Xbit_r79_c7 bl[7] br[7] wl[79] vdd gnd cell_6t
Xbit_r80_c7 bl[7] br[7] wl[80] vdd gnd cell_6t
Xbit_r81_c7 bl[7] br[7] wl[81] vdd gnd cell_6t
Xbit_r82_c7 bl[7] br[7] wl[82] vdd gnd cell_6t
Xbit_r83_c7 bl[7] br[7] wl[83] vdd gnd cell_6t
Xbit_r84_c7 bl[7] br[7] wl[84] vdd gnd cell_6t
Xbit_r85_c7 bl[7] br[7] wl[85] vdd gnd cell_6t
Xbit_r86_c7 bl[7] br[7] wl[86] vdd gnd cell_6t
Xbit_r87_c7 bl[7] br[7] wl[87] vdd gnd cell_6t
Xbit_r88_c7 bl[7] br[7] wl[88] vdd gnd cell_6t
Xbit_r89_c7 bl[7] br[7] wl[89] vdd gnd cell_6t
Xbit_r90_c7 bl[7] br[7] wl[90] vdd gnd cell_6t
Xbit_r91_c7 bl[7] br[7] wl[91] vdd gnd cell_6t
Xbit_r92_c7 bl[7] br[7] wl[92] vdd gnd cell_6t
Xbit_r93_c7 bl[7] br[7] wl[93] vdd gnd cell_6t
Xbit_r94_c7 bl[7] br[7] wl[94] vdd gnd cell_6t
Xbit_r95_c7 bl[7] br[7] wl[95] vdd gnd cell_6t
Xbit_r96_c7 bl[7] br[7] wl[96] vdd gnd cell_6t
Xbit_r97_c7 bl[7] br[7] wl[97] vdd gnd cell_6t
Xbit_r98_c7 bl[7] br[7] wl[98] vdd gnd cell_6t
Xbit_r99_c7 bl[7] br[7] wl[99] vdd gnd cell_6t
Xbit_r100_c7 bl[7] br[7] wl[100] vdd gnd cell_6t
Xbit_r101_c7 bl[7] br[7] wl[101] vdd gnd cell_6t
Xbit_r102_c7 bl[7] br[7] wl[102] vdd gnd cell_6t
Xbit_r103_c7 bl[7] br[7] wl[103] vdd gnd cell_6t
Xbit_r104_c7 bl[7] br[7] wl[104] vdd gnd cell_6t
Xbit_r105_c7 bl[7] br[7] wl[105] vdd gnd cell_6t
Xbit_r106_c7 bl[7] br[7] wl[106] vdd gnd cell_6t
Xbit_r107_c7 bl[7] br[7] wl[107] vdd gnd cell_6t
Xbit_r108_c7 bl[7] br[7] wl[108] vdd gnd cell_6t
Xbit_r109_c7 bl[7] br[7] wl[109] vdd gnd cell_6t
Xbit_r110_c7 bl[7] br[7] wl[110] vdd gnd cell_6t
Xbit_r111_c7 bl[7] br[7] wl[111] vdd gnd cell_6t
Xbit_r112_c7 bl[7] br[7] wl[112] vdd gnd cell_6t
Xbit_r113_c7 bl[7] br[7] wl[113] vdd gnd cell_6t
Xbit_r114_c7 bl[7] br[7] wl[114] vdd gnd cell_6t
Xbit_r115_c7 bl[7] br[7] wl[115] vdd gnd cell_6t
Xbit_r116_c7 bl[7] br[7] wl[116] vdd gnd cell_6t
Xbit_r117_c7 bl[7] br[7] wl[117] vdd gnd cell_6t
Xbit_r118_c7 bl[7] br[7] wl[118] vdd gnd cell_6t
Xbit_r119_c7 bl[7] br[7] wl[119] vdd gnd cell_6t
Xbit_r120_c7 bl[7] br[7] wl[120] vdd gnd cell_6t
Xbit_r121_c7 bl[7] br[7] wl[121] vdd gnd cell_6t
Xbit_r122_c7 bl[7] br[7] wl[122] vdd gnd cell_6t
Xbit_r123_c7 bl[7] br[7] wl[123] vdd gnd cell_6t
Xbit_r124_c7 bl[7] br[7] wl[124] vdd gnd cell_6t
Xbit_r125_c7 bl[7] br[7] wl[125] vdd gnd cell_6t
Xbit_r126_c7 bl[7] br[7] wl[126] vdd gnd cell_6t
Xbit_r127_c7 bl[7] br[7] wl[127] vdd gnd cell_6t
Xbit_r128_c7 bl[7] br[7] wl[128] vdd gnd cell_6t
Xbit_r129_c7 bl[7] br[7] wl[129] vdd gnd cell_6t
Xbit_r130_c7 bl[7] br[7] wl[130] vdd gnd cell_6t
Xbit_r131_c7 bl[7] br[7] wl[131] vdd gnd cell_6t
Xbit_r132_c7 bl[7] br[7] wl[132] vdd gnd cell_6t
Xbit_r133_c7 bl[7] br[7] wl[133] vdd gnd cell_6t
Xbit_r134_c7 bl[7] br[7] wl[134] vdd gnd cell_6t
Xbit_r135_c7 bl[7] br[7] wl[135] vdd gnd cell_6t
Xbit_r136_c7 bl[7] br[7] wl[136] vdd gnd cell_6t
Xbit_r137_c7 bl[7] br[7] wl[137] vdd gnd cell_6t
Xbit_r138_c7 bl[7] br[7] wl[138] vdd gnd cell_6t
Xbit_r139_c7 bl[7] br[7] wl[139] vdd gnd cell_6t
Xbit_r140_c7 bl[7] br[7] wl[140] vdd gnd cell_6t
Xbit_r141_c7 bl[7] br[7] wl[141] vdd gnd cell_6t
Xbit_r142_c7 bl[7] br[7] wl[142] vdd gnd cell_6t
Xbit_r143_c7 bl[7] br[7] wl[143] vdd gnd cell_6t
Xbit_r144_c7 bl[7] br[7] wl[144] vdd gnd cell_6t
Xbit_r145_c7 bl[7] br[7] wl[145] vdd gnd cell_6t
Xbit_r146_c7 bl[7] br[7] wl[146] vdd gnd cell_6t
Xbit_r147_c7 bl[7] br[7] wl[147] vdd gnd cell_6t
Xbit_r148_c7 bl[7] br[7] wl[148] vdd gnd cell_6t
Xbit_r149_c7 bl[7] br[7] wl[149] vdd gnd cell_6t
Xbit_r150_c7 bl[7] br[7] wl[150] vdd gnd cell_6t
Xbit_r151_c7 bl[7] br[7] wl[151] vdd gnd cell_6t
Xbit_r152_c7 bl[7] br[7] wl[152] vdd gnd cell_6t
Xbit_r153_c7 bl[7] br[7] wl[153] vdd gnd cell_6t
Xbit_r154_c7 bl[7] br[7] wl[154] vdd gnd cell_6t
Xbit_r155_c7 bl[7] br[7] wl[155] vdd gnd cell_6t
Xbit_r156_c7 bl[7] br[7] wl[156] vdd gnd cell_6t
Xbit_r157_c7 bl[7] br[7] wl[157] vdd gnd cell_6t
Xbit_r158_c7 bl[7] br[7] wl[158] vdd gnd cell_6t
Xbit_r159_c7 bl[7] br[7] wl[159] vdd gnd cell_6t
Xbit_r160_c7 bl[7] br[7] wl[160] vdd gnd cell_6t
Xbit_r161_c7 bl[7] br[7] wl[161] vdd gnd cell_6t
Xbit_r162_c7 bl[7] br[7] wl[162] vdd gnd cell_6t
Xbit_r163_c7 bl[7] br[7] wl[163] vdd gnd cell_6t
Xbit_r164_c7 bl[7] br[7] wl[164] vdd gnd cell_6t
Xbit_r165_c7 bl[7] br[7] wl[165] vdd gnd cell_6t
Xbit_r166_c7 bl[7] br[7] wl[166] vdd gnd cell_6t
Xbit_r167_c7 bl[7] br[7] wl[167] vdd gnd cell_6t
Xbit_r168_c7 bl[7] br[7] wl[168] vdd gnd cell_6t
Xbit_r169_c7 bl[7] br[7] wl[169] vdd gnd cell_6t
Xbit_r170_c7 bl[7] br[7] wl[170] vdd gnd cell_6t
Xbit_r171_c7 bl[7] br[7] wl[171] vdd gnd cell_6t
Xbit_r172_c7 bl[7] br[7] wl[172] vdd gnd cell_6t
Xbit_r173_c7 bl[7] br[7] wl[173] vdd gnd cell_6t
Xbit_r174_c7 bl[7] br[7] wl[174] vdd gnd cell_6t
Xbit_r175_c7 bl[7] br[7] wl[175] vdd gnd cell_6t
Xbit_r176_c7 bl[7] br[7] wl[176] vdd gnd cell_6t
Xbit_r177_c7 bl[7] br[7] wl[177] vdd gnd cell_6t
Xbit_r178_c7 bl[7] br[7] wl[178] vdd gnd cell_6t
Xbit_r179_c7 bl[7] br[7] wl[179] vdd gnd cell_6t
Xbit_r180_c7 bl[7] br[7] wl[180] vdd gnd cell_6t
Xbit_r181_c7 bl[7] br[7] wl[181] vdd gnd cell_6t
Xbit_r182_c7 bl[7] br[7] wl[182] vdd gnd cell_6t
Xbit_r183_c7 bl[7] br[7] wl[183] vdd gnd cell_6t
Xbit_r184_c7 bl[7] br[7] wl[184] vdd gnd cell_6t
Xbit_r185_c7 bl[7] br[7] wl[185] vdd gnd cell_6t
Xbit_r186_c7 bl[7] br[7] wl[186] vdd gnd cell_6t
Xbit_r187_c7 bl[7] br[7] wl[187] vdd gnd cell_6t
Xbit_r188_c7 bl[7] br[7] wl[188] vdd gnd cell_6t
Xbit_r189_c7 bl[7] br[7] wl[189] vdd gnd cell_6t
Xbit_r190_c7 bl[7] br[7] wl[190] vdd gnd cell_6t
Xbit_r191_c7 bl[7] br[7] wl[191] vdd gnd cell_6t
Xbit_r192_c7 bl[7] br[7] wl[192] vdd gnd cell_6t
Xbit_r193_c7 bl[7] br[7] wl[193] vdd gnd cell_6t
Xbit_r194_c7 bl[7] br[7] wl[194] vdd gnd cell_6t
Xbit_r195_c7 bl[7] br[7] wl[195] vdd gnd cell_6t
Xbit_r196_c7 bl[7] br[7] wl[196] vdd gnd cell_6t
Xbit_r197_c7 bl[7] br[7] wl[197] vdd gnd cell_6t
Xbit_r198_c7 bl[7] br[7] wl[198] vdd gnd cell_6t
Xbit_r199_c7 bl[7] br[7] wl[199] vdd gnd cell_6t
Xbit_r200_c7 bl[7] br[7] wl[200] vdd gnd cell_6t
Xbit_r201_c7 bl[7] br[7] wl[201] vdd gnd cell_6t
Xbit_r202_c7 bl[7] br[7] wl[202] vdd gnd cell_6t
Xbit_r203_c7 bl[7] br[7] wl[203] vdd gnd cell_6t
Xbit_r204_c7 bl[7] br[7] wl[204] vdd gnd cell_6t
Xbit_r205_c7 bl[7] br[7] wl[205] vdd gnd cell_6t
Xbit_r206_c7 bl[7] br[7] wl[206] vdd gnd cell_6t
Xbit_r207_c7 bl[7] br[7] wl[207] vdd gnd cell_6t
Xbit_r208_c7 bl[7] br[7] wl[208] vdd gnd cell_6t
Xbit_r209_c7 bl[7] br[7] wl[209] vdd gnd cell_6t
Xbit_r210_c7 bl[7] br[7] wl[210] vdd gnd cell_6t
Xbit_r211_c7 bl[7] br[7] wl[211] vdd gnd cell_6t
Xbit_r212_c7 bl[7] br[7] wl[212] vdd gnd cell_6t
Xbit_r213_c7 bl[7] br[7] wl[213] vdd gnd cell_6t
Xbit_r214_c7 bl[7] br[7] wl[214] vdd gnd cell_6t
Xbit_r215_c7 bl[7] br[7] wl[215] vdd gnd cell_6t
Xbit_r216_c7 bl[7] br[7] wl[216] vdd gnd cell_6t
Xbit_r217_c7 bl[7] br[7] wl[217] vdd gnd cell_6t
Xbit_r218_c7 bl[7] br[7] wl[218] vdd gnd cell_6t
Xbit_r219_c7 bl[7] br[7] wl[219] vdd gnd cell_6t
Xbit_r220_c7 bl[7] br[7] wl[220] vdd gnd cell_6t
Xbit_r221_c7 bl[7] br[7] wl[221] vdd gnd cell_6t
Xbit_r222_c7 bl[7] br[7] wl[222] vdd gnd cell_6t
Xbit_r223_c7 bl[7] br[7] wl[223] vdd gnd cell_6t
Xbit_r224_c7 bl[7] br[7] wl[224] vdd gnd cell_6t
Xbit_r225_c7 bl[7] br[7] wl[225] vdd gnd cell_6t
Xbit_r226_c7 bl[7] br[7] wl[226] vdd gnd cell_6t
Xbit_r227_c7 bl[7] br[7] wl[227] vdd gnd cell_6t
Xbit_r228_c7 bl[7] br[7] wl[228] vdd gnd cell_6t
Xbit_r229_c7 bl[7] br[7] wl[229] vdd gnd cell_6t
Xbit_r230_c7 bl[7] br[7] wl[230] vdd gnd cell_6t
Xbit_r231_c7 bl[7] br[7] wl[231] vdd gnd cell_6t
Xbit_r232_c7 bl[7] br[7] wl[232] vdd gnd cell_6t
Xbit_r233_c7 bl[7] br[7] wl[233] vdd gnd cell_6t
Xbit_r234_c7 bl[7] br[7] wl[234] vdd gnd cell_6t
Xbit_r235_c7 bl[7] br[7] wl[235] vdd gnd cell_6t
Xbit_r236_c7 bl[7] br[7] wl[236] vdd gnd cell_6t
Xbit_r237_c7 bl[7] br[7] wl[237] vdd gnd cell_6t
Xbit_r238_c7 bl[7] br[7] wl[238] vdd gnd cell_6t
Xbit_r239_c7 bl[7] br[7] wl[239] vdd gnd cell_6t
Xbit_r240_c7 bl[7] br[7] wl[240] vdd gnd cell_6t
Xbit_r241_c7 bl[7] br[7] wl[241] vdd gnd cell_6t
Xbit_r242_c7 bl[7] br[7] wl[242] vdd gnd cell_6t
Xbit_r243_c7 bl[7] br[7] wl[243] vdd gnd cell_6t
Xbit_r244_c7 bl[7] br[7] wl[244] vdd gnd cell_6t
Xbit_r245_c7 bl[7] br[7] wl[245] vdd gnd cell_6t
Xbit_r246_c7 bl[7] br[7] wl[246] vdd gnd cell_6t
Xbit_r247_c7 bl[7] br[7] wl[247] vdd gnd cell_6t
Xbit_r248_c7 bl[7] br[7] wl[248] vdd gnd cell_6t
Xbit_r249_c7 bl[7] br[7] wl[249] vdd gnd cell_6t
Xbit_r250_c7 bl[7] br[7] wl[250] vdd gnd cell_6t
Xbit_r251_c7 bl[7] br[7] wl[251] vdd gnd cell_6t
Xbit_r252_c7 bl[7] br[7] wl[252] vdd gnd cell_6t
Xbit_r253_c7 bl[7] br[7] wl[253] vdd gnd cell_6t
Xbit_r254_c7 bl[7] br[7] wl[254] vdd gnd cell_6t
Xbit_r255_c7 bl[7] br[7] wl[255] vdd gnd cell_6t
Xbit_r0_c8 bl[8] br[8] wl[0] vdd gnd cell_6t
Xbit_r1_c8 bl[8] br[8] wl[1] vdd gnd cell_6t
Xbit_r2_c8 bl[8] br[8] wl[2] vdd gnd cell_6t
Xbit_r3_c8 bl[8] br[8] wl[3] vdd gnd cell_6t
Xbit_r4_c8 bl[8] br[8] wl[4] vdd gnd cell_6t
Xbit_r5_c8 bl[8] br[8] wl[5] vdd gnd cell_6t
Xbit_r6_c8 bl[8] br[8] wl[6] vdd gnd cell_6t
Xbit_r7_c8 bl[8] br[8] wl[7] vdd gnd cell_6t
Xbit_r8_c8 bl[8] br[8] wl[8] vdd gnd cell_6t
Xbit_r9_c8 bl[8] br[8] wl[9] vdd gnd cell_6t
Xbit_r10_c8 bl[8] br[8] wl[10] vdd gnd cell_6t
Xbit_r11_c8 bl[8] br[8] wl[11] vdd gnd cell_6t
Xbit_r12_c8 bl[8] br[8] wl[12] vdd gnd cell_6t
Xbit_r13_c8 bl[8] br[8] wl[13] vdd gnd cell_6t
Xbit_r14_c8 bl[8] br[8] wl[14] vdd gnd cell_6t
Xbit_r15_c8 bl[8] br[8] wl[15] vdd gnd cell_6t
Xbit_r16_c8 bl[8] br[8] wl[16] vdd gnd cell_6t
Xbit_r17_c8 bl[8] br[8] wl[17] vdd gnd cell_6t
Xbit_r18_c8 bl[8] br[8] wl[18] vdd gnd cell_6t
Xbit_r19_c8 bl[8] br[8] wl[19] vdd gnd cell_6t
Xbit_r20_c8 bl[8] br[8] wl[20] vdd gnd cell_6t
Xbit_r21_c8 bl[8] br[8] wl[21] vdd gnd cell_6t
Xbit_r22_c8 bl[8] br[8] wl[22] vdd gnd cell_6t
Xbit_r23_c8 bl[8] br[8] wl[23] vdd gnd cell_6t
Xbit_r24_c8 bl[8] br[8] wl[24] vdd gnd cell_6t
Xbit_r25_c8 bl[8] br[8] wl[25] vdd gnd cell_6t
Xbit_r26_c8 bl[8] br[8] wl[26] vdd gnd cell_6t
Xbit_r27_c8 bl[8] br[8] wl[27] vdd gnd cell_6t
Xbit_r28_c8 bl[8] br[8] wl[28] vdd gnd cell_6t
Xbit_r29_c8 bl[8] br[8] wl[29] vdd gnd cell_6t
Xbit_r30_c8 bl[8] br[8] wl[30] vdd gnd cell_6t
Xbit_r31_c8 bl[8] br[8] wl[31] vdd gnd cell_6t
Xbit_r32_c8 bl[8] br[8] wl[32] vdd gnd cell_6t
Xbit_r33_c8 bl[8] br[8] wl[33] vdd gnd cell_6t
Xbit_r34_c8 bl[8] br[8] wl[34] vdd gnd cell_6t
Xbit_r35_c8 bl[8] br[8] wl[35] vdd gnd cell_6t
Xbit_r36_c8 bl[8] br[8] wl[36] vdd gnd cell_6t
Xbit_r37_c8 bl[8] br[8] wl[37] vdd gnd cell_6t
Xbit_r38_c8 bl[8] br[8] wl[38] vdd gnd cell_6t
Xbit_r39_c8 bl[8] br[8] wl[39] vdd gnd cell_6t
Xbit_r40_c8 bl[8] br[8] wl[40] vdd gnd cell_6t
Xbit_r41_c8 bl[8] br[8] wl[41] vdd gnd cell_6t
Xbit_r42_c8 bl[8] br[8] wl[42] vdd gnd cell_6t
Xbit_r43_c8 bl[8] br[8] wl[43] vdd gnd cell_6t
Xbit_r44_c8 bl[8] br[8] wl[44] vdd gnd cell_6t
Xbit_r45_c8 bl[8] br[8] wl[45] vdd gnd cell_6t
Xbit_r46_c8 bl[8] br[8] wl[46] vdd gnd cell_6t
Xbit_r47_c8 bl[8] br[8] wl[47] vdd gnd cell_6t
Xbit_r48_c8 bl[8] br[8] wl[48] vdd gnd cell_6t
Xbit_r49_c8 bl[8] br[8] wl[49] vdd gnd cell_6t
Xbit_r50_c8 bl[8] br[8] wl[50] vdd gnd cell_6t
Xbit_r51_c8 bl[8] br[8] wl[51] vdd gnd cell_6t
Xbit_r52_c8 bl[8] br[8] wl[52] vdd gnd cell_6t
Xbit_r53_c8 bl[8] br[8] wl[53] vdd gnd cell_6t
Xbit_r54_c8 bl[8] br[8] wl[54] vdd gnd cell_6t
Xbit_r55_c8 bl[8] br[8] wl[55] vdd gnd cell_6t
Xbit_r56_c8 bl[8] br[8] wl[56] vdd gnd cell_6t
Xbit_r57_c8 bl[8] br[8] wl[57] vdd gnd cell_6t
Xbit_r58_c8 bl[8] br[8] wl[58] vdd gnd cell_6t
Xbit_r59_c8 bl[8] br[8] wl[59] vdd gnd cell_6t
Xbit_r60_c8 bl[8] br[8] wl[60] vdd gnd cell_6t
Xbit_r61_c8 bl[8] br[8] wl[61] vdd gnd cell_6t
Xbit_r62_c8 bl[8] br[8] wl[62] vdd gnd cell_6t
Xbit_r63_c8 bl[8] br[8] wl[63] vdd gnd cell_6t
Xbit_r64_c8 bl[8] br[8] wl[64] vdd gnd cell_6t
Xbit_r65_c8 bl[8] br[8] wl[65] vdd gnd cell_6t
Xbit_r66_c8 bl[8] br[8] wl[66] vdd gnd cell_6t
Xbit_r67_c8 bl[8] br[8] wl[67] vdd gnd cell_6t
Xbit_r68_c8 bl[8] br[8] wl[68] vdd gnd cell_6t
Xbit_r69_c8 bl[8] br[8] wl[69] vdd gnd cell_6t
Xbit_r70_c8 bl[8] br[8] wl[70] vdd gnd cell_6t
Xbit_r71_c8 bl[8] br[8] wl[71] vdd gnd cell_6t
Xbit_r72_c8 bl[8] br[8] wl[72] vdd gnd cell_6t
Xbit_r73_c8 bl[8] br[8] wl[73] vdd gnd cell_6t
Xbit_r74_c8 bl[8] br[8] wl[74] vdd gnd cell_6t
Xbit_r75_c8 bl[8] br[8] wl[75] vdd gnd cell_6t
Xbit_r76_c8 bl[8] br[8] wl[76] vdd gnd cell_6t
Xbit_r77_c8 bl[8] br[8] wl[77] vdd gnd cell_6t
Xbit_r78_c8 bl[8] br[8] wl[78] vdd gnd cell_6t
Xbit_r79_c8 bl[8] br[8] wl[79] vdd gnd cell_6t
Xbit_r80_c8 bl[8] br[8] wl[80] vdd gnd cell_6t
Xbit_r81_c8 bl[8] br[8] wl[81] vdd gnd cell_6t
Xbit_r82_c8 bl[8] br[8] wl[82] vdd gnd cell_6t
Xbit_r83_c8 bl[8] br[8] wl[83] vdd gnd cell_6t
Xbit_r84_c8 bl[8] br[8] wl[84] vdd gnd cell_6t
Xbit_r85_c8 bl[8] br[8] wl[85] vdd gnd cell_6t
Xbit_r86_c8 bl[8] br[8] wl[86] vdd gnd cell_6t
Xbit_r87_c8 bl[8] br[8] wl[87] vdd gnd cell_6t
Xbit_r88_c8 bl[8] br[8] wl[88] vdd gnd cell_6t
Xbit_r89_c8 bl[8] br[8] wl[89] vdd gnd cell_6t
Xbit_r90_c8 bl[8] br[8] wl[90] vdd gnd cell_6t
Xbit_r91_c8 bl[8] br[8] wl[91] vdd gnd cell_6t
Xbit_r92_c8 bl[8] br[8] wl[92] vdd gnd cell_6t
Xbit_r93_c8 bl[8] br[8] wl[93] vdd gnd cell_6t
Xbit_r94_c8 bl[8] br[8] wl[94] vdd gnd cell_6t
Xbit_r95_c8 bl[8] br[8] wl[95] vdd gnd cell_6t
Xbit_r96_c8 bl[8] br[8] wl[96] vdd gnd cell_6t
Xbit_r97_c8 bl[8] br[8] wl[97] vdd gnd cell_6t
Xbit_r98_c8 bl[8] br[8] wl[98] vdd gnd cell_6t
Xbit_r99_c8 bl[8] br[8] wl[99] vdd gnd cell_6t
Xbit_r100_c8 bl[8] br[8] wl[100] vdd gnd cell_6t
Xbit_r101_c8 bl[8] br[8] wl[101] vdd gnd cell_6t
Xbit_r102_c8 bl[8] br[8] wl[102] vdd gnd cell_6t
Xbit_r103_c8 bl[8] br[8] wl[103] vdd gnd cell_6t
Xbit_r104_c8 bl[8] br[8] wl[104] vdd gnd cell_6t
Xbit_r105_c8 bl[8] br[8] wl[105] vdd gnd cell_6t
Xbit_r106_c8 bl[8] br[8] wl[106] vdd gnd cell_6t
Xbit_r107_c8 bl[8] br[8] wl[107] vdd gnd cell_6t
Xbit_r108_c8 bl[8] br[8] wl[108] vdd gnd cell_6t
Xbit_r109_c8 bl[8] br[8] wl[109] vdd gnd cell_6t
Xbit_r110_c8 bl[8] br[8] wl[110] vdd gnd cell_6t
Xbit_r111_c8 bl[8] br[8] wl[111] vdd gnd cell_6t
Xbit_r112_c8 bl[8] br[8] wl[112] vdd gnd cell_6t
Xbit_r113_c8 bl[8] br[8] wl[113] vdd gnd cell_6t
Xbit_r114_c8 bl[8] br[8] wl[114] vdd gnd cell_6t
Xbit_r115_c8 bl[8] br[8] wl[115] vdd gnd cell_6t
Xbit_r116_c8 bl[8] br[8] wl[116] vdd gnd cell_6t
Xbit_r117_c8 bl[8] br[8] wl[117] vdd gnd cell_6t
Xbit_r118_c8 bl[8] br[8] wl[118] vdd gnd cell_6t
Xbit_r119_c8 bl[8] br[8] wl[119] vdd gnd cell_6t
Xbit_r120_c8 bl[8] br[8] wl[120] vdd gnd cell_6t
Xbit_r121_c8 bl[8] br[8] wl[121] vdd gnd cell_6t
Xbit_r122_c8 bl[8] br[8] wl[122] vdd gnd cell_6t
Xbit_r123_c8 bl[8] br[8] wl[123] vdd gnd cell_6t
Xbit_r124_c8 bl[8] br[8] wl[124] vdd gnd cell_6t
Xbit_r125_c8 bl[8] br[8] wl[125] vdd gnd cell_6t
Xbit_r126_c8 bl[8] br[8] wl[126] vdd gnd cell_6t
Xbit_r127_c8 bl[8] br[8] wl[127] vdd gnd cell_6t
Xbit_r128_c8 bl[8] br[8] wl[128] vdd gnd cell_6t
Xbit_r129_c8 bl[8] br[8] wl[129] vdd gnd cell_6t
Xbit_r130_c8 bl[8] br[8] wl[130] vdd gnd cell_6t
Xbit_r131_c8 bl[8] br[8] wl[131] vdd gnd cell_6t
Xbit_r132_c8 bl[8] br[8] wl[132] vdd gnd cell_6t
Xbit_r133_c8 bl[8] br[8] wl[133] vdd gnd cell_6t
Xbit_r134_c8 bl[8] br[8] wl[134] vdd gnd cell_6t
Xbit_r135_c8 bl[8] br[8] wl[135] vdd gnd cell_6t
Xbit_r136_c8 bl[8] br[8] wl[136] vdd gnd cell_6t
Xbit_r137_c8 bl[8] br[8] wl[137] vdd gnd cell_6t
Xbit_r138_c8 bl[8] br[8] wl[138] vdd gnd cell_6t
Xbit_r139_c8 bl[8] br[8] wl[139] vdd gnd cell_6t
Xbit_r140_c8 bl[8] br[8] wl[140] vdd gnd cell_6t
Xbit_r141_c8 bl[8] br[8] wl[141] vdd gnd cell_6t
Xbit_r142_c8 bl[8] br[8] wl[142] vdd gnd cell_6t
Xbit_r143_c8 bl[8] br[8] wl[143] vdd gnd cell_6t
Xbit_r144_c8 bl[8] br[8] wl[144] vdd gnd cell_6t
Xbit_r145_c8 bl[8] br[8] wl[145] vdd gnd cell_6t
Xbit_r146_c8 bl[8] br[8] wl[146] vdd gnd cell_6t
Xbit_r147_c8 bl[8] br[8] wl[147] vdd gnd cell_6t
Xbit_r148_c8 bl[8] br[8] wl[148] vdd gnd cell_6t
Xbit_r149_c8 bl[8] br[8] wl[149] vdd gnd cell_6t
Xbit_r150_c8 bl[8] br[8] wl[150] vdd gnd cell_6t
Xbit_r151_c8 bl[8] br[8] wl[151] vdd gnd cell_6t
Xbit_r152_c8 bl[8] br[8] wl[152] vdd gnd cell_6t
Xbit_r153_c8 bl[8] br[8] wl[153] vdd gnd cell_6t
Xbit_r154_c8 bl[8] br[8] wl[154] vdd gnd cell_6t
Xbit_r155_c8 bl[8] br[8] wl[155] vdd gnd cell_6t
Xbit_r156_c8 bl[8] br[8] wl[156] vdd gnd cell_6t
Xbit_r157_c8 bl[8] br[8] wl[157] vdd gnd cell_6t
Xbit_r158_c8 bl[8] br[8] wl[158] vdd gnd cell_6t
Xbit_r159_c8 bl[8] br[8] wl[159] vdd gnd cell_6t
Xbit_r160_c8 bl[8] br[8] wl[160] vdd gnd cell_6t
Xbit_r161_c8 bl[8] br[8] wl[161] vdd gnd cell_6t
Xbit_r162_c8 bl[8] br[8] wl[162] vdd gnd cell_6t
Xbit_r163_c8 bl[8] br[8] wl[163] vdd gnd cell_6t
Xbit_r164_c8 bl[8] br[8] wl[164] vdd gnd cell_6t
Xbit_r165_c8 bl[8] br[8] wl[165] vdd gnd cell_6t
Xbit_r166_c8 bl[8] br[8] wl[166] vdd gnd cell_6t
Xbit_r167_c8 bl[8] br[8] wl[167] vdd gnd cell_6t
Xbit_r168_c8 bl[8] br[8] wl[168] vdd gnd cell_6t
Xbit_r169_c8 bl[8] br[8] wl[169] vdd gnd cell_6t
Xbit_r170_c8 bl[8] br[8] wl[170] vdd gnd cell_6t
Xbit_r171_c8 bl[8] br[8] wl[171] vdd gnd cell_6t
Xbit_r172_c8 bl[8] br[8] wl[172] vdd gnd cell_6t
Xbit_r173_c8 bl[8] br[8] wl[173] vdd gnd cell_6t
Xbit_r174_c8 bl[8] br[8] wl[174] vdd gnd cell_6t
Xbit_r175_c8 bl[8] br[8] wl[175] vdd gnd cell_6t
Xbit_r176_c8 bl[8] br[8] wl[176] vdd gnd cell_6t
Xbit_r177_c8 bl[8] br[8] wl[177] vdd gnd cell_6t
Xbit_r178_c8 bl[8] br[8] wl[178] vdd gnd cell_6t
Xbit_r179_c8 bl[8] br[8] wl[179] vdd gnd cell_6t
Xbit_r180_c8 bl[8] br[8] wl[180] vdd gnd cell_6t
Xbit_r181_c8 bl[8] br[8] wl[181] vdd gnd cell_6t
Xbit_r182_c8 bl[8] br[8] wl[182] vdd gnd cell_6t
Xbit_r183_c8 bl[8] br[8] wl[183] vdd gnd cell_6t
Xbit_r184_c8 bl[8] br[8] wl[184] vdd gnd cell_6t
Xbit_r185_c8 bl[8] br[8] wl[185] vdd gnd cell_6t
Xbit_r186_c8 bl[8] br[8] wl[186] vdd gnd cell_6t
Xbit_r187_c8 bl[8] br[8] wl[187] vdd gnd cell_6t
Xbit_r188_c8 bl[8] br[8] wl[188] vdd gnd cell_6t
Xbit_r189_c8 bl[8] br[8] wl[189] vdd gnd cell_6t
Xbit_r190_c8 bl[8] br[8] wl[190] vdd gnd cell_6t
Xbit_r191_c8 bl[8] br[8] wl[191] vdd gnd cell_6t
Xbit_r192_c8 bl[8] br[8] wl[192] vdd gnd cell_6t
Xbit_r193_c8 bl[8] br[8] wl[193] vdd gnd cell_6t
Xbit_r194_c8 bl[8] br[8] wl[194] vdd gnd cell_6t
Xbit_r195_c8 bl[8] br[8] wl[195] vdd gnd cell_6t
Xbit_r196_c8 bl[8] br[8] wl[196] vdd gnd cell_6t
Xbit_r197_c8 bl[8] br[8] wl[197] vdd gnd cell_6t
Xbit_r198_c8 bl[8] br[8] wl[198] vdd gnd cell_6t
Xbit_r199_c8 bl[8] br[8] wl[199] vdd gnd cell_6t
Xbit_r200_c8 bl[8] br[8] wl[200] vdd gnd cell_6t
Xbit_r201_c8 bl[8] br[8] wl[201] vdd gnd cell_6t
Xbit_r202_c8 bl[8] br[8] wl[202] vdd gnd cell_6t
Xbit_r203_c8 bl[8] br[8] wl[203] vdd gnd cell_6t
Xbit_r204_c8 bl[8] br[8] wl[204] vdd gnd cell_6t
Xbit_r205_c8 bl[8] br[8] wl[205] vdd gnd cell_6t
Xbit_r206_c8 bl[8] br[8] wl[206] vdd gnd cell_6t
Xbit_r207_c8 bl[8] br[8] wl[207] vdd gnd cell_6t
Xbit_r208_c8 bl[8] br[8] wl[208] vdd gnd cell_6t
Xbit_r209_c8 bl[8] br[8] wl[209] vdd gnd cell_6t
Xbit_r210_c8 bl[8] br[8] wl[210] vdd gnd cell_6t
Xbit_r211_c8 bl[8] br[8] wl[211] vdd gnd cell_6t
Xbit_r212_c8 bl[8] br[8] wl[212] vdd gnd cell_6t
Xbit_r213_c8 bl[8] br[8] wl[213] vdd gnd cell_6t
Xbit_r214_c8 bl[8] br[8] wl[214] vdd gnd cell_6t
Xbit_r215_c8 bl[8] br[8] wl[215] vdd gnd cell_6t
Xbit_r216_c8 bl[8] br[8] wl[216] vdd gnd cell_6t
Xbit_r217_c8 bl[8] br[8] wl[217] vdd gnd cell_6t
Xbit_r218_c8 bl[8] br[8] wl[218] vdd gnd cell_6t
Xbit_r219_c8 bl[8] br[8] wl[219] vdd gnd cell_6t
Xbit_r220_c8 bl[8] br[8] wl[220] vdd gnd cell_6t
Xbit_r221_c8 bl[8] br[8] wl[221] vdd gnd cell_6t
Xbit_r222_c8 bl[8] br[8] wl[222] vdd gnd cell_6t
Xbit_r223_c8 bl[8] br[8] wl[223] vdd gnd cell_6t
Xbit_r224_c8 bl[8] br[8] wl[224] vdd gnd cell_6t
Xbit_r225_c8 bl[8] br[8] wl[225] vdd gnd cell_6t
Xbit_r226_c8 bl[8] br[8] wl[226] vdd gnd cell_6t
Xbit_r227_c8 bl[8] br[8] wl[227] vdd gnd cell_6t
Xbit_r228_c8 bl[8] br[8] wl[228] vdd gnd cell_6t
Xbit_r229_c8 bl[8] br[8] wl[229] vdd gnd cell_6t
Xbit_r230_c8 bl[8] br[8] wl[230] vdd gnd cell_6t
Xbit_r231_c8 bl[8] br[8] wl[231] vdd gnd cell_6t
Xbit_r232_c8 bl[8] br[8] wl[232] vdd gnd cell_6t
Xbit_r233_c8 bl[8] br[8] wl[233] vdd gnd cell_6t
Xbit_r234_c8 bl[8] br[8] wl[234] vdd gnd cell_6t
Xbit_r235_c8 bl[8] br[8] wl[235] vdd gnd cell_6t
Xbit_r236_c8 bl[8] br[8] wl[236] vdd gnd cell_6t
Xbit_r237_c8 bl[8] br[8] wl[237] vdd gnd cell_6t
Xbit_r238_c8 bl[8] br[8] wl[238] vdd gnd cell_6t
Xbit_r239_c8 bl[8] br[8] wl[239] vdd gnd cell_6t
Xbit_r240_c8 bl[8] br[8] wl[240] vdd gnd cell_6t
Xbit_r241_c8 bl[8] br[8] wl[241] vdd gnd cell_6t
Xbit_r242_c8 bl[8] br[8] wl[242] vdd gnd cell_6t
Xbit_r243_c8 bl[8] br[8] wl[243] vdd gnd cell_6t
Xbit_r244_c8 bl[8] br[8] wl[244] vdd gnd cell_6t
Xbit_r245_c8 bl[8] br[8] wl[245] vdd gnd cell_6t
Xbit_r246_c8 bl[8] br[8] wl[246] vdd gnd cell_6t
Xbit_r247_c8 bl[8] br[8] wl[247] vdd gnd cell_6t
Xbit_r248_c8 bl[8] br[8] wl[248] vdd gnd cell_6t
Xbit_r249_c8 bl[8] br[8] wl[249] vdd gnd cell_6t
Xbit_r250_c8 bl[8] br[8] wl[250] vdd gnd cell_6t
Xbit_r251_c8 bl[8] br[8] wl[251] vdd gnd cell_6t
Xbit_r252_c8 bl[8] br[8] wl[252] vdd gnd cell_6t
Xbit_r253_c8 bl[8] br[8] wl[253] vdd gnd cell_6t
Xbit_r254_c8 bl[8] br[8] wl[254] vdd gnd cell_6t
Xbit_r255_c8 bl[8] br[8] wl[255] vdd gnd cell_6t
Xbit_r0_c9 bl[9] br[9] wl[0] vdd gnd cell_6t
Xbit_r1_c9 bl[9] br[9] wl[1] vdd gnd cell_6t
Xbit_r2_c9 bl[9] br[9] wl[2] vdd gnd cell_6t
Xbit_r3_c9 bl[9] br[9] wl[3] vdd gnd cell_6t
Xbit_r4_c9 bl[9] br[9] wl[4] vdd gnd cell_6t
Xbit_r5_c9 bl[9] br[9] wl[5] vdd gnd cell_6t
Xbit_r6_c9 bl[9] br[9] wl[6] vdd gnd cell_6t
Xbit_r7_c9 bl[9] br[9] wl[7] vdd gnd cell_6t
Xbit_r8_c9 bl[9] br[9] wl[8] vdd gnd cell_6t
Xbit_r9_c9 bl[9] br[9] wl[9] vdd gnd cell_6t
Xbit_r10_c9 bl[9] br[9] wl[10] vdd gnd cell_6t
Xbit_r11_c9 bl[9] br[9] wl[11] vdd gnd cell_6t
Xbit_r12_c9 bl[9] br[9] wl[12] vdd gnd cell_6t
Xbit_r13_c9 bl[9] br[9] wl[13] vdd gnd cell_6t
Xbit_r14_c9 bl[9] br[9] wl[14] vdd gnd cell_6t
Xbit_r15_c9 bl[9] br[9] wl[15] vdd gnd cell_6t
Xbit_r16_c9 bl[9] br[9] wl[16] vdd gnd cell_6t
Xbit_r17_c9 bl[9] br[9] wl[17] vdd gnd cell_6t
Xbit_r18_c9 bl[9] br[9] wl[18] vdd gnd cell_6t
Xbit_r19_c9 bl[9] br[9] wl[19] vdd gnd cell_6t
Xbit_r20_c9 bl[9] br[9] wl[20] vdd gnd cell_6t
Xbit_r21_c9 bl[9] br[9] wl[21] vdd gnd cell_6t
Xbit_r22_c9 bl[9] br[9] wl[22] vdd gnd cell_6t
Xbit_r23_c9 bl[9] br[9] wl[23] vdd gnd cell_6t
Xbit_r24_c9 bl[9] br[9] wl[24] vdd gnd cell_6t
Xbit_r25_c9 bl[9] br[9] wl[25] vdd gnd cell_6t
Xbit_r26_c9 bl[9] br[9] wl[26] vdd gnd cell_6t
Xbit_r27_c9 bl[9] br[9] wl[27] vdd gnd cell_6t
Xbit_r28_c9 bl[9] br[9] wl[28] vdd gnd cell_6t
Xbit_r29_c9 bl[9] br[9] wl[29] vdd gnd cell_6t
Xbit_r30_c9 bl[9] br[9] wl[30] vdd gnd cell_6t
Xbit_r31_c9 bl[9] br[9] wl[31] vdd gnd cell_6t
Xbit_r32_c9 bl[9] br[9] wl[32] vdd gnd cell_6t
Xbit_r33_c9 bl[9] br[9] wl[33] vdd gnd cell_6t
Xbit_r34_c9 bl[9] br[9] wl[34] vdd gnd cell_6t
Xbit_r35_c9 bl[9] br[9] wl[35] vdd gnd cell_6t
Xbit_r36_c9 bl[9] br[9] wl[36] vdd gnd cell_6t
Xbit_r37_c9 bl[9] br[9] wl[37] vdd gnd cell_6t
Xbit_r38_c9 bl[9] br[9] wl[38] vdd gnd cell_6t
Xbit_r39_c9 bl[9] br[9] wl[39] vdd gnd cell_6t
Xbit_r40_c9 bl[9] br[9] wl[40] vdd gnd cell_6t
Xbit_r41_c9 bl[9] br[9] wl[41] vdd gnd cell_6t
Xbit_r42_c9 bl[9] br[9] wl[42] vdd gnd cell_6t
Xbit_r43_c9 bl[9] br[9] wl[43] vdd gnd cell_6t
Xbit_r44_c9 bl[9] br[9] wl[44] vdd gnd cell_6t
Xbit_r45_c9 bl[9] br[9] wl[45] vdd gnd cell_6t
Xbit_r46_c9 bl[9] br[9] wl[46] vdd gnd cell_6t
Xbit_r47_c9 bl[9] br[9] wl[47] vdd gnd cell_6t
Xbit_r48_c9 bl[9] br[9] wl[48] vdd gnd cell_6t
Xbit_r49_c9 bl[9] br[9] wl[49] vdd gnd cell_6t
Xbit_r50_c9 bl[9] br[9] wl[50] vdd gnd cell_6t
Xbit_r51_c9 bl[9] br[9] wl[51] vdd gnd cell_6t
Xbit_r52_c9 bl[9] br[9] wl[52] vdd gnd cell_6t
Xbit_r53_c9 bl[9] br[9] wl[53] vdd gnd cell_6t
Xbit_r54_c9 bl[9] br[9] wl[54] vdd gnd cell_6t
Xbit_r55_c9 bl[9] br[9] wl[55] vdd gnd cell_6t
Xbit_r56_c9 bl[9] br[9] wl[56] vdd gnd cell_6t
Xbit_r57_c9 bl[9] br[9] wl[57] vdd gnd cell_6t
Xbit_r58_c9 bl[9] br[9] wl[58] vdd gnd cell_6t
Xbit_r59_c9 bl[9] br[9] wl[59] vdd gnd cell_6t
Xbit_r60_c9 bl[9] br[9] wl[60] vdd gnd cell_6t
Xbit_r61_c9 bl[9] br[9] wl[61] vdd gnd cell_6t
Xbit_r62_c9 bl[9] br[9] wl[62] vdd gnd cell_6t
Xbit_r63_c9 bl[9] br[9] wl[63] vdd gnd cell_6t
Xbit_r64_c9 bl[9] br[9] wl[64] vdd gnd cell_6t
Xbit_r65_c9 bl[9] br[9] wl[65] vdd gnd cell_6t
Xbit_r66_c9 bl[9] br[9] wl[66] vdd gnd cell_6t
Xbit_r67_c9 bl[9] br[9] wl[67] vdd gnd cell_6t
Xbit_r68_c9 bl[9] br[9] wl[68] vdd gnd cell_6t
Xbit_r69_c9 bl[9] br[9] wl[69] vdd gnd cell_6t
Xbit_r70_c9 bl[9] br[9] wl[70] vdd gnd cell_6t
Xbit_r71_c9 bl[9] br[9] wl[71] vdd gnd cell_6t
Xbit_r72_c9 bl[9] br[9] wl[72] vdd gnd cell_6t
Xbit_r73_c9 bl[9] br[9] wl[73] vdd gnd cell_6t
Xbit_r74_c9 bl[9] br[9] wl[74] vdd gnd cell_6t
Xbit_r75_c9 bl[9] br[9] wl[75] vdd gnd cell_6t
Xbit_r76_c9 bl[9] br[9] wl[76] vdd gnd cell_6t
Xbit_r77_c9 bl[9] br[9] wl[77] vdd gnd cell_6t
Xbit_r78_c9 bl[9] br[9] wl[78] vdd gnd cell_6t
Xbit_r79_c9 bl[9] br[9] wl[79] vdd gnd cell_6t
Xbit_r80_c9 bl[9] br[9] wl[80] vdd gnd cell_6t
Xbit_r81_c9 bl[9] br[9] wl[81] vdd gnd cell_6t
Xbit_r82_c9 bl[9] br[9] wl[82] vdd gnd cell_6t
Xbit_r83_c9 bl[9] br[9] wl[83] vdd gnd cell_6t
Xbit_r84_c9 bl[9] br[9] wl[84] vdd gnd cell_6t
Xbit_r85_c9 bl[9] br[9] wl[85] vdd gnd cell_6t
Xbit_r86_c9 bl[9] br[9] wl[86] vdd gnd cell_6t
Xbit_r87_c9 bl[9] br[9] wl[87] vdd gnd cell_6t
Xbit_r88_c9 bl[9] br[9] wl[88] vdd gnd cell_6t
Xbit_r89_c9 bl[9] br[9] wl[89] vdd gnd cell_6t
Xbit_r90_c9 bl[9] br[9] wl[90] vdd gnd cell_6t
Xbit_r91_c9 bl[9] br[9] wl[91] vdd gnd cell_6t
Xbit_r92_c9 bl[9] br[9] wl[92] vdd gnd cell_6t
Xbit_r93_c9 bl[9] br[9] wl[93] vdd gnd cell_6t
Xbit_r94_c9 bl[9] br[9] wl[94] vdd gnd cell_6t
Xbit_r95_c9 bl[9] br[9] wl[95] vdd gnd cell_6t
Xbit_r96_c9 bl[9] br[9] wl[96] vdd gnd cell_6t
Xbit_r97_c9 bl[9] br[9] wl[97] vdd gnd cell_6t
Xbit_r98_c9 bl[9] br[9] wl[98] vdd gnd cell_6t
Xbit_r99_c9 bl[9] br[9] wl[99] vdd gnd cell_6t
Xbit_r100_c9 bl[9] br[9] wl[100] vdd gnd cell_6t
Xbit_r101_c9 bl[9] br[9] wl[101] vdd gnd cell_6t
Xbit_r102_c9 bl[9] br[9] wl[102] vdd gnd cell_6t
Xbit_r103_c9 bl[9] br[9] wl[103] vdd gnd cell_6t
Xbit_r104_c9 bl[9] br[9] wl[104] vdd gnd cell_6t
Xbit_r105_c9 bl[9] br[9] wl[105] vdd gnd cell_6t
Xbit_r106_c9 bl[9] br[9] wl[106] vdd gnd cell_6t
Xbit_r107_c9 bl[9] br[9] wl[107] vdd gnd cell_6t
Xbit_r108_c9 bl[9] br[9] wl[108] vdd gnd cell_6t
Xbit_r109_c9 bl[9] br[9] wl[109] vdd gnd cell_6t
Xbit_r110_c9 bl[9] br[9] wl[110] vdd gnd cell_6t
Xbit_r111_c9 bl[9] br[9] wl[111] vdd gnd cell_6t
Xbit_r112_c9 bl[9] br[9] wl[112] vdd gnd cell_6t
Xbit_r113_c9 bl[9] br[9] wl[113] vdd gnd cell_6t
Xbit_r114_c9 bl[9] br[9] wl[114] vdd gnd cell_6t
Xbit_r115_c9 bl[9] br[9] wl[115] vdd gnd cell_6t
Xbit_r116_c9 bl[9] br[9] wl[116] vdd gnd cell_6t
Xbit_r117_c9 bl[9] br[9] wl[117] vdd gnd cell_6t
Xbit_r118_c9 bl[9] br[9] wl[118] vdd gnd cell_6t
Xbit_r119_c9 bl[9] br[9] wl[119] vdd gnd cell_6t
Xbit_r120_c9 bl[9] br[9] wl[120] vdd gnd cell_6t
Xbit_r121_c9 bl[9] br[9] wl[121] vdd gnd cell_6t
Xbit_r122_c9 bl[9] br[9] wl[122] vdd gnd cell_6t
Xbit_r123_c9 bl[9] br[9] wl[123] vdd gnd cell_6t
Xbit_r124_c9 bl[9] br[9] wl[124] vdd gnd cell_6t
Xbit_r125_c9 bl[9] br[9] wl[125] vdd gnd cell_6t
Xbit_r126_c9 bl[9] br[9] wl[126] vdd gnd cell_6t
Xbit_r127_c9 bl[9] br[9] wl[127] vdd gnd cell_6t
Xbit_r128_c9 bl[9] br[9] wl[128] vdd gnd cell_6t
Xbit_r129_c9 bl[9] br[9] wl[129] vdd gnd cell_6t
Xbit_r130_c9 bl[9] br[9] wl[130] vdd gnd cell_6t
Xbit_r131_c9 bl[9] br[9] wl[131] vdd gnd cell_6t
Xbit_r132_c9 bl[9] br[9] wl[132] vdd gnd cell_6t
Xbit_r133_c9 bl[9] br[9] wl[133] vdd gnd cell_6t
Xbit_r134_c9 bl[9] br[9] wl[134] vdd gnd cell_6t
Xbit_r135_c9 bl[9] br[9] wl[135] vdd gnd cell_6t
Xbit_r136_c9 bl[9] br[9] wl[136] vdd gnd cell_6t
Xbit_r137_c9 bl[9] br[9] wl[137] vdd gnd cell_6t
Xbit_r138_c9 bl[9] br[9] wl[138] vdd gnd cell_6t
Xbit_r139_c9 bl[9] br[9] wl[139] vdd gnd cell_6t
Xbit_r140_c9 bl[9] br[9] wl[140] vdd gnd cell_6t
Xbit_r141_c9 bl[9] br[9] wl[141] vdd gnd cell_6t
Xbit_r142_c9 bl[9] br[9] wl[142] vdd gnd cell_6t
Xbit_r143_c9 bl[9] br[9] wl[143] vdd gnd cell_6t
Xbit_r144_c9 bl[9] br[9] wl[144] vdd gnd cell_6t
Xbit_r145_c9 bl[9] br[9] wl[145] vdd gnd cell_6t
Xbit_r146_c9 bl[9] br[9] wl[146] vdd gnd cell_6t
Xbit_r147_c9 bl[9] br[9] wl[147] vdd gnd cell_6t
Xbit_r148_c9 bl[9] br[9] wl[148] vdd gnd cell_6t
Xbit_r149_c9 bl[9] br[9] wl[149] vdd gnd cell_6t
Xbit_r150_c9 bl[9] br[9] wl[150] vdd gnd cell_6t
Xbit_r151_c9 bl[9] br[9] wl[151] vdd gnd cell_6t
Xbit_r152_c9 bl[9] br[9] wl[152] vdd gnd cell_6t
Xbit_r153_c9 bl[9] br[9] wl[153] vdd gnd cell_6t
Xbit_r154_c9 bl[9] br[9] wl[154] vdd gnd cell_6t
Xbit_r155_c9 bl[9] br[9] wl[155] vdd gnd cell_6t
Xbit_r156_c9 bl[9] br[9] wl[156] vdd gnd cell_6t
Xbit_r157_c9 bl[9] br[9] wl[157] vdd gnd cell_6t
Xbit_r158_c9 bl[9] br[9] wl[158] vdd gnd cell_6t
Xbit_r159_c9 bl[9] br[9] wl[159] vdd gnd cell_6t
Xbit_r160_c9 bl[9] br[9] wl[160] vdd gnd cell_6t
Xbit_r161_c9 bl[9] br[9] wl[161] vdd gnd cell_6t
Xbit_r162_c9 bl[9] br[9] wl[162] vdd gnd cell_6t
Xbit_r163_c9 bl[9] br[9] wl[163] vdd gnd cell_6t
Xbit_r164_c9 bl[9] br[9] wl[164] vdd gnd cell_6t
Xbit_r165_c9 bl[9] br[9] wl[165] vdd gnd cell_6t
Xbit_r166_c9 bl[9] br[9] wl[166] vdd gnd cell_6t
Xbit_r167_c9 bl[9] br[9] wl[167] vdd gnd cell_6t
Xbit_r168_c9 bl[9] br[9] wl[168] vdd gnd cell_6t
Xbit_r169_c9 bl[9] br[9] wl[169] vdd gnd cell_6t
Xbit_r170_c9 bl[9] br[9] wl[170] vdd gnd cell_6t
Xbit_r171_c9 bl[9] br[9] wl[171] vdd gnd cell_6t
Xbit_r172_c9 bl[9] br[9] wl[172] vdd gnd cell_6t
Xbit_r173_c9 bl[9] br[9] wl[173] vdd gnd cell_6t
Xbit_r174_c9 bl[9] br[9] wl[174] vdd gnd cell_6t
Xbit_r175_c9 bl[9] br[9] wl[175] vdd gnd cell_6t
Xbit_r176_c9 bl[9] br[9] wl[176] vdd gnd cell_6t
Xbit_r177_c9 bl[9] br[9] wl[177] vdd gnd cell_6t
Xbit_r178_c9 bl[9] br[9] wl[178] vdd gnd cell_6t
Xbit_r179_c9 bl[9] br[9] wl[179] vdd gnd cell_6t
Xbit_r180_c9 bl[9] br[9] wl[180] vdd gnd cell_6t
Xbit_r181_c9 bl[9] br[9] wl[181] vdd gnd cell_6t
Xbit_r182_c9 bl[9] br[9] wl[182] vdd gnd cell_6t
Xbit_r183_c9 bl[9] br[9] wl[183] vdd gnd cell_6t
Xbit_r184_c9 bl[9] br[9] wl[184] vdd gnd cell_6t
Xbit_r185_c9 bl[9] br[9] wl[185] vdd gnd cell_6t
Xbit_r186_c9 bl[9] br[9] wl[186] vdd gnd cell_6t
Xbit_r187_c9 bl[9] br[9] wl[187] vdd gnd cell_6t
Xbit_r188_c9 bl[9] br[9] wl[188] vdd gnd cell_6t
Xbit_r189_c9 bl[9] br[9] wl[189] vdd gnd cell_6t
Xbit_r190_c9 bl[9] br[9] wl[190] vdd gnd cell_6t
Xbit_r191_c9 bl[9] br[9] wl[191] vdd gnd cell_6t
Xbit_r192_c9 bl[9] br[9] wl[192] vdd gnd cell_6t
Xbit_r193_c9 bl[9] br[9] wl[193] vdd gnd cell_6t
Xbit_r194_c9 bl[9] br[9] wl[194] vdd gnd cell_6t
Xbit_r195_c9 bl[9] br[9] wl[195] vdd gnd cell_6t
Xbit_r196_c9 bl[9] br[9] wl[196] vdd gnd cell_6t
Xbit_r197_c9 bl[9] br[9] wl[197] vdd gnd cell_6t
Xbit_r198_c9 bl[9] br[9] wl[198] vdd gnd cell_6t
Xbit_r199_c9 bl[9] br[9] wl[199] vdd gnd cell_6t
Xbit_r200_c9 bl[9] br[9] wl[200] vdd gnd cell_6t
Xbit_r201_c9 bl[9] br[9] wl[201] vdd gnd cell_6t
Xbit_r202_c9 bl[9] br[9] wl[202] vdd gnd cell_6t
Xbit_r203_c9 bl[9] br[9] wl[203] vdd gnd cell_6t
Xbit_r204_c9 bl[9] br[9] wl[204] vdd gnd cell_6t
Xbit_r205_c9 bl[9] br[9] wl[205] vdd gnd cell_6t
Xbit_r206_c9 bl[9] br[9] wl[206] vdd gnd cell_6t
Xbit_r207_c9 bl[9] br[9] wl[207] vdd gnd cell_6t
Xbit_r208_c9 bl[9] br[9] wl[208] vdd gnd cell_6t
Xbit_r209_c9 bl[9] br[9] wl[209] vdd gnd cell_6t
Xbit_r210_c9 bl[9] br[9] wl[210] vdd gnd cell_6t
Xbit_r211_c9 bl[9] br[9] wl[211] vdd gnd cell_6t
Xbit_r212_c9 bl[9] br[9] wl[212] vdd gnd cell_6t
Xbit_r213_c9 bl[9] br[9] wl[213] vdd gnd cell_6t
Xbit_r214_c9 bl[9] br[9] wl[214] vdd gnd cell_6t
Xbit_r215_c9 bl[9] br[9] wl[215] vdd gnd cell_6t
Xbit_r216_c9 bl[9] br[9] wl[216] vdd gnd cell_6t
Xbit_r217_c9 bl[9] br[9] wl[217] vdd gnd cell_6t
Xbit_r218_c9 bl[9] br[9] wl[218] vdd gnd cell_6t
Xbit_r219_c9 bl[9] br[9] wl[219] vdd gnd cell_6t
Xbit_r220_c9 bl[9] br[9] wl[220] vdd gnd cell_6t
Xbit_r221_c9 bl[9] br[9] wl[221] vdd gnd cell_6t
Xbit_r222_c9 bl[9] br[9] wl[222] vdd gnd cell_6t
Xbit_r223_c9 bl[9] br[9] wl[223] vdd gnd cell_6t
Xbit_r224_c9 bl[9] br[9] wl[224] vdd gnd cell_6t
Xbit_r225_c9 bl[9] br[9] wl[225] vdd gnd cell_6t
Xbit_r226_c9 bl[9] br[9] wl[226] vdd gnd cell_6t
Xbit_r227_c9 bl[9] br[9] wl[227] vdd gnd cell_6t
Xbit_r228_c9 bl[9] br[9] wl[228] vdd gnd cell_6t
Xbit_r229_c9 bl[9] br[9] wl[229] vdd gnd cell_6t
Xbit_r230_c9 bl[9] br[9] wl[230] vdd gnd cell_6t
Xbit_r231_c9 bl[9] br[9] wl[231] vdd gnd cell_6t
Xbit_r232_c9 bl[9] br[9] wl[232] vdd gnd cell_6t
Xbit_r233_c9 bl[9] br[9] wl[233] vdd gnd cell_6t
Xbit_r234_c9 bl[9] br[9] wl[234] vdd gnd cell_6t
Xbit_r235_c9 bl[9] br[9] wl[235] vdd gnd cell_6t
Xbit_r236_c9 bl[9] br[9] wl[236] vdd gnd cell_6t
Xbit_r237_c9 bl[9] br[9] wl[237] vdd gnd cell_6t
Xbit_r238_c9 bl[9] br[9] wl[238] vdd gnd cell_6t
Xbit_r239_c9 bl[9] br[9] wl[239] vdd gnd cell_6t
Xbit_r240_c9 bl[9] br[9] wl[240] vdd gnd cell_6t
Xbit_r241_c9 bl[9] br[9] wl[241] vdd gnd cell_6t
Xbit_r242_c9 bl[9] br[9] wl[242] vdd gnd cell_6t
Xbit_r243_c9 bl[9] br[9] wl[243] vdd gnd cell_6t
Xbit_r244_c9 bl[9] br[9] wl[244] vdd gnd cell_6t
Xbit_r245_c9 bl[9] br[9] wl[245] vdd gnd cell_6t
Xbit_r246_c9 bl[9] br[9] wl[246] vdd gnd cell_6t
Xbit_r247_c9 bl[9] br[9] wl[247] vdd gnd cell_6t
Xbit_r248_c9 bl[9] br[9] wl[248] vdd gnd cell_6t
Xbit_r249_c9 bl[9] br[9] wl[249] vdd gnd cell_6t
Xbit_r250_c9 bl[9] br[9] wl[250] vdd gnd cell_6t
Xbit_r251_c9 bl[9] br[9] wl[251] vdd gnd cell_6t
Xbit_r252_c9 bl[9] br[9] wl[252] vdd gnd cell_6t
Xbit_r253_c9 bl[9] br[9] wl[253] vdd gnd cell_6t
Xbit_r254_c9 bl[9] br[9] wl[254] vdd gnd cell_6t
Xbit_r255_c9 bl[9] br[9] wl[255] vdd gnd cell_6t
Xbit_r0_c10 bl[10] br[10] wl[0] vdd gnd cell_6t
Xbit_r1_c10 bl[10] br[10] wl[1] vdd gnd cell_6t
Xbit_r2_c10 bl[10] br[10] wl[2] vdd gnd cell_6t
Xbit_r3_c10 bl[10] br[10] wl[3] vdd gnd cell_6t
Xbit_r4_c10 bl[10] br[10] wl[4] vdd gnd cell_6t
Xbit_r5_c10 bl[10] br[10] wl[5] vdd gnd cell_6t
Xbit_r6_c10 bl[10] br[10] wl[6] vdd gnd cell_6t
Xbit_r7_c10 bl[10] br[10] wl[7] vdd gnd cell_6t
Xbit_r8_c10 bl[10] br[10] wl[8] vdd gnd cell_6t
Xbit_r9_c10 bl[10] br[10] wl[9] vdd gnd cell_6t
Xbit_r10_c10 bl[10] br[10] wl[10] vdd gnd cell_6t
Xbit_r11_c10 bl[10] br[10] wl[11] vdd gnd cell_6t
Xbit_r12_c10 bl[10] br[10] wl[12] vdd gnd cell_6t
Xbit_r13_c10 bl[10] br[10] wl[13] vdd gnd cell_6t
Xbit_r14_c10 bl[10] br[10] wl[14] vdd gnd cell_6t
Xbit_r15_c10 bl[10] br[10] wl[15] vdd gnd cell_6t
Xbit_r16_c10 bl[10] br[10] wl[16] vdd gnd cell_6t
Xbit_r17_c10 bl[10] br[10] wl[17] vdd gnd cell_6t
Xbit_r18_c10 bl[10] br[10] wl[18] vdd gnd cell_6t
Xbit_r19_c10 bl[10] br[10] wl[19] vdd gnd cell_6t
Xbit_r20_c10 bl[10] br[10] wl[20] vdd gnd cell_6t
Xbit_r21_c10 bl[10] br[10] wl[21] vdd gnd cell_6t
Xbit_r22_c10 bl[10] br[10] wl[22] vdd gnd cell_6t
Xbit_r23_c10 bl[10] br[10] wl[23] vdd gnd cell_6t
Xbit_r24_c10 bl[10] br[10] wl[24] vdd gnd cell_6t
Xbit_r25_c10 bl[10] br[10] wl[25] vdd gnd cell_6t
Xbit_r26_c10 bl[10] br[10] wl[26] vdd gnd cell_6t
Xbit_r27_c10 bl[10] br[10] wl[27] vdd gnd cell_6t
Xbit_r28_c10 bl[10] br[10] wl[28] vdd gnd cell_6t
Xbit_r29_c10 bl[10] br[10] wl[29] vdd gnd cell_6t
Xbit_r30_c10 bl[10] br[10] wl[30] vdd gnd cell_6t
Xbit_r31_c10 bl[10] br[10] wl[31] vdd gnd cell_6t
Xbit_r32_c10 bl[10] br[10] wl[32] vdd gnd cell_6t
Xbit_r33_c10 bl[10] br[10] wl[33] vdd gnd cell_6t
Xbit_r34_c10 bl[10] br[10] wl[34] vdd gnd cell_6t
Xbit_r35_c10 bl[10] br[10] wl[35] vdd gnd cell_6t
Xbit_r36_c10 bl[10] br[10] wl[36] vdd gnd cell_6t
Xbit_r37_c10 bl[10] br[10] wl[37] vdd gnd cell_6t
Xbit_r38_c10 bl[10] br[10] wl[38] vdd gnd cell_6t
Xbit_r39_c10 bl[10] br[10] wl[39] vdd gnd cell_6t
Xbit_r40_c10 bl[10] br[10] wl[40] vdd gnd cell_6t
Xbit_r41_c10 bl[10] br[10] wl[41] vdd gnd cell_6t
Xbit_r42_c10 bl[10] br[10] wl[42] vdd gnd cell_6t
Xbit_r43_c10 bl[10] br[10] wl[43] vdd gnd cell_6t
Xbit_r44_c10 bl[10] br[10] wl[44] vdd gnd cell_6t
Xbit_r45_c10 bl[10] br[10] wl[45] vdd gnd cell_6t
Xbit_r46_c10 bl[10] br[10] wl[46] vdd gnd cell_6t
Xbit_r47_c10 bl[10] br[10] wl[47] vdd gnd cell_6t
Xbit_r48_c10 bl[10] br[10] wl[48] vdd gnd cell_6t
Xbit_r49_c10 bl[10] br[10] wl[49] vdd gnd cell_6t
Xbit_r50_c10 bl[10] br[10] wl[50] vdd gnd cell_6t
Xbit_r51_c10 bl[10] br[10] wl[51] vdd gnd cell_6t
Xbit_r52_c10 bl[10] br[10] wl[52] vdd gnd cell_6t
Xbit_r53_c10 bl[10] br[10] wl[53] vdd gnd cell_6t
Xbit_r54_c10 bl[10] br[10] wl[54] vdd gnd cell_6t
Xbit_r55_c10 bl[10] br[10] wl[55] vdd gnd cell_6t
Xbit_r56_c10 bl[10] br[10] wl[56] vdd gnd cell_6t
Xbit_r57_c10 bl[10] br[10] wl[57] vdd gnd cell_6t
Xbit_r58_c10 bl[10] br[10] wl[58] vdd gnd cell_6t
Xbit_r59_c10 bl[10] br[10] wl[59] vdd gnd cell_6t
Xbit_r60_c10 bl[10] br[10] wl[60] vdd gnd cell_6t
Xbit_r61_c10 bl[10] br[10] wl[61] vdd gnd cell_6t
Xbit_r62_c10 bl[10] br[10] wl[62] vdd gnd cell_6t
Xbit_r63_c10 bl[10] br[10] wl[63] vdd gnd cell_6t
Xbit_r64_c10 bl[10] br[10] wl[64] vdd gnd cell_6t
Xbit_r65_c10 bl[10] br[10] wl[65] vdd gnd cell_6t
Xbit_r66_c10 bl[10] br[10] wl[66] vdd gnd cell_6t
Xbit_r67_c10 bl[10] br[10] wl[67] vdd gnd cell_6t
Xbit_r68_c10 bl[10] br[10] wl[68] vdd gnd cell_6t
Xbit_r69_c10 bl[10] br[10] wl[69] vdd gnd cell_6t
Xbit_r70_c10 bl[10] br[10] wl[70] vdd gnd cell_6t
Xbit_r71_c10 bl[10] br[10] wl[71] vdd gnd cell_6t
Xbit_r72_c10 bl[10] br[10] wl[72] vdd gnd cell_6t
Xbit_r73_c10 bl[10] br[10] wl[73] vdd gnd cell_6t
Xbit_r74_c10 bl[10] br[10] wl[74] vdd gnd cell_6t
Xbit_r75_c10 bl[10] br[10] wl[75] vdd gnd cell_6t
Xbit_r76_c10 bl[10] br[10] wl[76] vdd gnd cell_6t
Xbit_r77_c10 bl[10] br[10] wl[77] vdd gnd cell_6t
Xbit_r78_c10 bl[10] br[10] wl[78] vdd gnd cell_6t
Xbit_r79_c10 bl[10] br[10] wl[79] vdd gnd cell_6t
Xbit_r80_c10 bl[10] br[10] wl[80] vdd gnd cell_6t
Xbit_r81_c10 bl[10] br[10] wl[81] vdd gnd cell_6t
Xbit_r82_c10 bl[10] br[10] wl[82] vdd gnd cell_6t
Xbit_r83_c10 bl[10] br[10] wl[83] vdd gnd cell_6t
Xbit_r84_c10 bl[10] br[10] wl[84] vdd gnd cell_6t
Xbit_r85_c10 bl[10] br[10] wl[85] vdd gnd cell_6t
Xbit_r86_c10 bl[10] br[10] wl[86] vdd gnd cell_6t
Xbit_r87_c10 bl[10] br[10] wl[87] vdd gnd cell_6t
Xbit_r88_c10 bl[10] br[10] wl[88] vdd gnd cell_6t
Xbit_r89_c10 bl[10] br[10] wl[89] vdd gnd cell_6t
Xbit_r90_c10 bl[10] br[10] wl[90] vdd gnd cell_6t
Xbit_r91_c10 bl[10] br[10] wl[91] vdd gnd cell_6t
Xbit_r92_c10 bl[10] br[10] wl[92] vdd gnd cell_6t
Xbit_r93_c10 bl[10] br[10] wl[93] vdd gnd cell_6t
Xbit_r94_c10 bl[10] br[10] wl[94] vdd gnd cell_6t
Xbit_r95_c10 bl[10] br[10] wl[95] vdd gnd cell_6t
Xbit_r96_c10 bl[10] br[10] wl[96] vdd gnd cell_6t
Xbit_r97_c10 bl[10] br[10] wl[97] vdd gnd cell_6t
Xbit_r98_c10 bl[10] br[10] wl[98] vdd gnd cell_6t
Xbit_r99_c10 bl[10] br[10] wl[99] vdd gnd cell_6t
Xbit_r100_c10 bl[10] br[10] wl[100] vdd gnd cell_6t
Xbit_r101_c10 bl[10] br[10] wl[101] vdd gnd cell_6t
Xbit_r102_c10 bl[10] br[10] wl[102] vdd gnd cell_6t
Xbit_r103_c10 bl[10] br[10] wl[103] vdd gnd cell_6t
Xbit_r104_c10 bl[10] br[10] wl[104] vdd gnd cell_6t
Xbit_r105_c10 bl[10] br[10] wl[105] vdd gnd cell_6t
Xbit_r106_c10 bl[10] br[10] wl[106] vdd gnd cell_6t
Xbit_r107_c10 bl[10] br[10] wl[107] vdd gnd cell_6t
Xbit_r108_c10 bl[10] br[10] wl[108] vdd gnd cell_6t
Xbit_r109_c10 bl[10] br[10] wl[109] vdd gnd cell_6t
Xbit_r110_c10 bl[10] br[10] wl[110] vdd gnd cell_6t
Xbit_r111_c10 bl[10] br[10] wl[111] vdd gnd cell_6t
Xbit_r112_c10 bl[10] br[10] wl[112] vdd gnd cell_6t
Xbit_r113_c10 bl[10] br[10] wl[113] vdd gnd cell_6t
Xbit_r114_c10 bl[10] br[10] wl[114] vdd gnd cell_6t
Xbit_r115_c10 bl[10] br[10] wl[115] vdd gnd cell_6t
Xbit_r116_c10 bl[10] br[10] wl[116] vdd gnd cell_6t
Xbit_r117_c10 bl[10] br[10] wl[117] vdd gnd cell_6t
Xbit_r118_c10 bl[10] br[10] wl[118] vdd gnd cell_6t
Xbit_r119_c10 bl[10] br[10] wl[119] vdd gnd cell_6t
Xbit_r120_c10 bl[10] br[10] wl[120] vdd gnd cell_6t
Xbit_r121_c10 bl[10] br[10] wl[121] vdd gnd cell_6t
Xbit_r122_c10 bl[10] br[10] wl[122] vdd gnd cell_6t
Xbit_r123_c10 bl[10] br[10] wl[123] vdd gnd cell_6t
Xbit_r124_c10 bl[10] br[10] wl[124] vdd gnd cell_6t
Xbit_r125_c10 bl[10] br[10] wl[125] vdd gnd cell_6t
Xbit_r126_c10 bl[10] br[10] wl[126] vdd gnd cell_6t
Xbit_r127_c10 bl[10] br[10] wl[127] vdd gnd cell_6t
Xbit_r128_c10 bl[10] br[10] wl[128] vdd gnd cell_6t
Xbit_r129_c10 bl[10] br[10] wl[129] vdd gnd cell_6t
Xbit_r130_c10 bl[10] br[10] wl[130] vdd gnd cell_6t
Xbit_r131_c10 bl[10] br[10] wl[131] vdd gnd cell_6t
Xbit_r132_c10 bl[10] br[10] wl[132] vdd gnd cell_6t
Xbit_r133_c10 bl[10] br[10] wl[133] vdd gnd cell_6t
Xbit_r134_c10 bl[10] br[10] wl[134] vdd gnd cell_6t
Xbit_r135_c10 bl[10] br[10] wl[135] vdd gnd cell_6t
Xbit_r136_c10 bl[10] br[10] wl[136] vdd gnd cell_6t
Xbit_r137_c10 bl[10] br[10] wl[137] vdd gnd cell_6t
Xbit_r138_c10 bl[10] br[10] wl[138] vdd gnd cell_6t
Xbit_r139_c10 bl[10] br[10] wl[139] vdd gnd cell_6t
Xbit_r140_c10 bl[10] br[10] wl[140] vdd gnd cell_6t
Xbit_r141_c10 bl[10] br[10] wl[141] vdd gnd cell_6t
Xbit_r142_c10 bl[10] br[10] wl[142] vdd gnd cell_6t
Xbit_r143_c10 bl[10] br[10] wl[143] vdd gnd cell_6t
Xbit_r144_c10 bl[10] br[10] wl[144] vdd gnd cell_6t
Xbit_r145_c10 bl[10] br[10] wl[145] vdd gnd cell_6t
Xbit_r146_c10 bl[10] br[10] wl[146] vdd gnd cell_6t
Xbit_r147_c10 bl[10] br[10] wl[147] vdd gnd cell_6t
Xbit_r148_c10 bl[10] br[10] wl[148] vdd gnd cell_6t
Xbit_r149_c10 bl[10] br[10] wl[149] vdd gnd cell_6t
Xbit_r150_c10 bl[10] br[10] wl[150] vdd gnd cell_6t
Xbit_r151_c10 bl[10] br[10] wl[151] vdd gnd cell_6t
Xbit_r152_c10 bl[10] br[10] wl[152] vdd gnd cell_6t
Xbit_r153_c10 bl[10] br[10] wl[153] vdd gnd cell_6t
Xbit_r154_c10 bl[10] br[10] wl[154] vdd gnd cell_6t
Xbit_r155_c10 bl[10] br[10] wl[155] vdd gnd cell_6t
Xbit_r156_c10 bl[10] br[10] wl[156] vdd gnd cell_6t
Xbit_r157_c10 bl[10] br[10] wl[157] vdd gnd cell_6t
Xbit_r158_c10 bl[10] br[10] wl[158] vdd gnd cell_6t
Xbit_r159_c10 bl[10] br[10] wl[159] vdd gnd cell_6t
Xbit_r160_c10 bl[10] br[10] wl[160] vdd gnd cell_6t
Xbit_r161_c10 bl[10] br[10] wl[161] vdd gnd cell_6t
Xbit_r162_c10 bl[10] br[10] wl[162] vdd gnd cell_6t
Xbit_r163_c10 bl[10] br[10] wl[163] vdd gnd cell_6t
Xbit_r164_c10 bl[10] br[10] wl[164] vdd gnd cell_6t
Xbit_r165_c10 bl[10] br[10] wl[165] vdd gnd cell_6t
Xbit_r166_c10 bl[10] br[10] wl[166] vdd gnd cell_6t
Xbit_r167_c10 bl[10] br[10] wl[167] vdd gnd cell_6t
Xbit_r168_c10 bl[10] br[10] wl[168] vdd gnd cell_6t
Xbit_r169_c10 bl[10] br[10] wl[169] vdd gnd cell_6t
Xbit_r170_c10 bl[10] br[10] wl[170] vdd gnd cell_6t
Xbit_r171_c10 bl[10] br[10] wl[171] vdd gnd cell_6t
Xbit_r172_c10 bl[10] br[10] wl[172] vdd gnd cell_6t
Xbit_r173_c10 bl[10] br[10] wl[173] vdd gnd cell_6t
Xbit_r174_c10 bl[10] br[10] wl[174] vdd gnd cell_6t
Xbit_r175_c10 bl[10] br[10] wl[175] vdd gnd cell_6t
Xbit_r176_c10 bl[10] br[10] wl[176] vdd gnd cell_6t
Xbit_r177_c10 bl[10] br[10] wl[177] vdd gnd cell_6t
Xbit_r178_c10 bl[10] br[10] wl[178] vdd gnd cell_6t
Xbit_r179_c10 bl[10] br[10] wl[179] vdd gnd cell_6t
Xbit_r180_c10 bl[10] br[10] wl[180] vdd gnd cell_6t
Xbit_r181_c10 bl[10] br[10] wl[181] vdd gnd cell_6t
Xbit_r182_c10 bl[10] br[10] wl[182] vdd gnd cell_6t
Xbit_r183_c10 bl[10] br[10] wl[183] vdd gnd cell_6t
Xbit_r184_c10 bl[10] br[10] wl[184] vdd gnd cell_6t
Xbit_r185_c10 bl[10] br[10] wl[185] vdd gnd cell_6t
Xbit_r186_c10 bl[10] br[10] wl[186] vdd gnd cell_6t
Xbit_r187_c10 bl[10] br[10] wl[187] vdd gnd cell_6t
Xbit_r188_c10 bl[10] br[10] wl[188] vdd gnd cell_6t
Xbit_r189_c10 bl[10] br[10] wl[189] vdd gnd cell_6t
Xbit_r190_c10 bl[10] br[10] wl[190] vdd gnd cell_6t
Xbit_r191_c10 bl[10] br[10] wl[191] vdd gnd cell_6t
Xbit_r192_c10 bl[10] br[10] wl[192] vdd gnd cell_6t
Xbit_r193_c10 bl[10] br[10] wl[193] vdd gnd cell_6t
Xbit_r194_c10 bl[10] br[10] wl[194] vdd gnd cell_6t
Xbit_r195_c10 bl[10] br[10] wl[195] vdd gnd cell_6t
Xbit_r196_c10 bl[10] br[10] wl[196] vdd gnd cell_6t
Xbit_r197_c10 bl[10] br[10] wl[197] vdd gnd cell_6t
Xbit_r198_c10 bl[10] br[10] wl[198] vdd gnd cell_6t
Xbit_r199_c10 bl[10] br[10] wl[199] vdd gnd cell_6t
Xbit_r200_c10 bl[10] br[10] wl[200] vdd gnd cell_6t
Xbit_r201_c10 bl[10] br[10] wl[201] vdd gnd cell_6t
Xbit_r202_c10 bl[10] br[10] wl[202] vdd gnd cell_6t
Xbit_r203_c10 bl[10] br[10] wl[203] vdd gnd cell_6t
Xbit_r204_c10 bl[10] br[10] wl[204] vdd gnd cell_6t
Xbit_r205_c10 bl[10] br[10] wl[205] vdd gnd cell_6t
Xbit_r206_c10 bl[10] br[10] wl[206] vdd gnd cell_6t
Xbit_r207_c10 bl[10] br[10] wl[207] vdd gnd cell_6t
Xbit_r208_c10 bl[10] br[10] wl[208] vdd gnd cell_6t
Xbit_r209_c10 bl[10] br[10] wl[209] vdd gnd cell_6t
Xbit_r210_c10 bl[10] br[10] wl[210] vdd gnd cell_6t
Xbit_r211_c10 bl[10] br[10] wl[211] vdd gnd cell_6t
Xbit_r212_c10 bl[10] br[10] wl[212] vdd gnd cell_6t
Xbit_r213_c10 bl[10] br[10] wl[213] vdd gnd cell_6t
Xbit_r214_c10 bl[10] br[10] wl[214] vdd gnd cell_6t
Xbit_r215_c10 bl[10] br[10] wl[215] vdd gnd cell_6t
Xbit_r216_c10 bl[10] br[10] wl[216] vdd gnd cell_6t
Xbit_r217_c10 bl[10] br[10] wl[217] vdd gnd cell_6t
Xbit_r218_c10 bl[10] br[10] wl[218] vdd gnd cell_6t
Xbit_r219_c10 bl[10] br[10] wl[219] vdd gnd cell_6t
Xbit_r220_c10 bl[10] br[10] wl[220] vdd gnd cell_6t
Xbit_r221_c10 bl[10] br[10] wl[221] vdd gnd cell_6t
Xbit_r222_c10 bl[10] br[10] wl[222] vdd gnd cell_6t
Xbit_r223_c10 bl[10] br[10] wl[223] vdd gnd cell_6t
Xbit_r224_c10 bl[10] br[10] wl[224] vdd gnd cell_6t
Xbit_r225_c10 bl[10] br[10] wl[225] vdd gnd cell_6t
Xbit_r226_c10 bl[10] br[10] wl[226] vdd gnd cell_6t
Xbit_r227_c10 bl[10] br[10] wl[227] vdd gnd cell_6t
Xbit_r228_c10 bl[10] br[10] wl[228] vdd gnd cell_6t
Xbit_r229_c10 bl[10] br[10] wl[229] vdd gnd cell_6t
Xbit_r230_c10 bl[10] br[10] wl[230] vdd gnd cell_6t
Xbit_r231_c10 bl[10] br[10] wl[231] vdd gnd cell_6t
Xbit_r232_c10 bl[10] br[10] wl[232] vdd gnd cell_6t
Xbit_r233_c10 bl[10] br[10] wl[233] vdd gnd cell_6t
Xbit_r234_c10 bl[10] br[10] wl[234] vdd gnd cell_6t
Xbit_r235_c10 bl[10] br[10] wl[235] vdd gnd cell_6t
Xbit_r236_c10 bl[10] br[10] wl[236] vdd gnd cell_6t
Xbit_r237_c10 bl[10] br[10] wl[237] vdd gnd cell_6t
Xbit_r238_c10 bl[10] br[10] wl[238] vdd gnd cell_6t
Xbit_r239_c10 bl[10] br[10] wl[239] vdd gnd cell_6t
Xbit_r240_c10 bl[10] br[10] wl[240] vdd gnd cell_6t
Xbit_r241_c10 bl[10] br[10] wl[241] vdd gnd cell_6t
Xbit_r242_c10 bl[10] br[10] wl[242] vdd gnd cell_6t
Xbit_r243_c10 bl[10] br[10] wl[243] vdd gnd cell_6t
Xbit_r244_c10 bl[10] br[10] wl[244] vdd gnd cell_6t
Xbit_r245_c10 bl[10] br[10] wl[245] vdd gnd cell_6t
Xbit_r246_c10 bl[10] br[10] wl[246] vdd gnd cell_6t
Xbit_r247_c10 bl[10] br[10] wl[247] vdd gnd cell_6t
Xbit_r248_c10 bl[10] br[10] wl[248] vdd gnd cell_6t
Xbit_r249_c10 bl[10] br[10] wl[249] vdd gnd cell_6t
Xbit_r250_c10 bl[10] br[10] wl[250] vdd gnd cell_6t
Xbit_r251_c10 bl[10] br[10] wl[251] vdd gnd cell_6t
Xbit_r252_c10 bl[10] br[10] wl[252] vdd gnd cell_6t
Xbit_r253_c10 bl[10] br[10] wl[253] vdd gnd cell_6t
Xbit_r254_c10 bl[10] br[10] wl[254] vdd gnd cell_6t
Xbit_r255_c10 bl[10] br[10] wl[255] vdd gnd cell_6t
Xbit_r0_c11 bl[11] br[11] wl[0] vdd gnd cell_6t
Xbit_r1_c11 bl[11] br[11] wl[1] vdd gnd cell_6t
Xbit_r2_c11 bl[11] br[11] wl[2] vdd gnd cell_6t
Xbit_r3_c11 bl[11] br[11] wl[3] vdd gnd cell_6t
Xbit_r4_c11 bl[11] br[11] wl[4] vdd gnd cell_6t
Xbit_r5_c11 bl[11] br[11] wl[5] vdd gnd cell_6t
Xbit_r6_c11 bl[11] br[11] wl[6] vdd gnd cell_6t
Xbit_r7_c11 bl[11] br[11] wl[7] vdd gnd cell_6t
Xbit_r8_c11 bl[11] br[11] wl[8] vdd gnd cell_6t
Xbit_r9_c11 bl[11] br[11] wl[9] vdd gnd cell_6t
Xbit_r10_c11 bl[11] br[11] wl[10] vdd gnd cell_6t
Xbit_r11_c11 bl[11] br[11] wl[11] vdd gnd cell_6t
Xbit_r12_c11 bl[11] br[11] wl[12] vdd gnd cell_6t
Xbit_r13_c11 bl[11] br[11] wl[13] vdd gnd cell_6t
Xbit_r14_c11 bl[11] br[11] wl[14] vdd gnd cell_6t
Xbit_r15_c11 bl[11] br[11] wl[15] vdd gnd cell_6t
Xbit_r16_c11 bl[11] br[11] wl[16] vdd gnd cell_6t
Xbit_r17_c11 bl[11] br[11] wl[17] vdd gnd cell_6t
Xbit_r18_c11 bl[11] br[11] wl[18] vdd gnd cell_6t
Xbit_r19_c11 bl[11] br[11] wl[19] vdd gnd cell_6t
Xbit_r20_c11 bl[11] br[11] wl[20] vdd gnd cell_6t
Xbit_r21_c11 bl[11] br[11] wl[21] vdd gnd cell_6t
Xbit_r22_c11 bl[11] br[11] wl[22] vdd gnd cell_6t
Xbit_r23_c11 bl[11] br[11] wl[23] vdd gnd cell_6t
Xbit_r24_c11 bl[11] br[11] wl[24] vdd gnd cell_6t
Xbit_r25_c11 bl[11] br[11] wl[25] vdd gnd cell_6t
Xbit_r26_c11 bl[11] br[11] wl[26] vdd gnd cell_6t
Xbit_r27_c11 bl[11] br[11] wl[27] vdd gnd cell_6t
Xbit_r28_c11 bl[11] br[11] wl[28] vdd gnd cell_6t
Xbit_r29_c11 bl[11] br[11] wl[29] vdd gnd cell_6t
Xbit_r30_c11 bl[11] br[11] wl[30] vdd gnd cell_6t
Xbit_r31_c11 bl[11] br[11] wl[31] vdd gnd cell_6t
Xbit_r32_c11 bl[11] br[11] wl[32] vdd gnd cell_6t
Xbit_r33_c11 bl[11] br[11] wl[33] vdd gnd cell_6t
Xbit_r34_c11 bl[11] br[11] wl[34] vdd gnd cell_6t
Xbit_r35_c11 bl[11] br[11] wl[35] vdd gnd cell_6t
Xbit_r36_c11 bl[11] br[11] wl[36] vdd gnd cell_6t
Xbit_r37_c11 bl[11] br[11] wl[37] vdd gnd cell_6t
Xbit_r38_c11 bl[11] br[11] wl[38] vdd gnd cell_6t
Xbit_r39_c11 bl[11] br[11] wl[39] vdd gnd cell_6t
Xbit_r40_c11 bl[11] br[11] wl[40] vdd gnd cell_6t
Xbit_r41_c11 bl[11] br[11] wl[41] vdd gnd cell_6t
Xbit_r42_c11 bl[11] br[11] wl[42] vdd gnd cell_6t
Xbit_r43_c11 bl[11] br[11] wl[43] vdd gnd cell_6t
Xbit_r44_c11 bl[11] br[11] wl[44] vdd gnd cell_6t
Xbit_r45_c11 bl[11] br[11] wl[45] vdd gnd cell_6t
Xbit_r46_c11 bl[11] br[11] wl[46] vdd gnd cell_6t
Xbit_r47_c11 bl[11] br[11] wl[47] vdd gnd cell_6t
Xbit_r48_c11 bl[11] br[11] wl[48] vdd gnd cell_6t
Xbit_r49_c11 bl[11] br[11] wl[49] vdd gnd cell_6t
Xbit_r50_c11 bl[11] br[11] wl[50] vdd gnd cell_6t
Xbit_r51_c11 bl[11] br[11] wl[51] vdd gnd cell_6t
Xbit_r52_c11 bl[11] br[11] wl[52] vdd gnd cell_6t
Xbit_r53_c11 bl[11] br[11] wl[53] vdd gnd cell_6t
Xbit_r54_c11 bl[11] br[11] wl[54] vdd gnd cell_6t
Xbit_r55_c11 bl[11] br[11] wl[55] vdd gnd cell_6t
Xbit_r56_c11 bl[11] br[11] wl[56] vdd gnd cell_6t
Xbit_r57_c11 bl[11] br[11] wl[57] vdd gnd cell_6t
Xbit_r58_c11 bl[11] br[11] wl[58] vdd gnd cell_6t
Xbit_r59_c11 bl[11] br[11] wl[59] vdd gnd cell_6t
Xbit_r60_c11 bl[11] br[11] wl[60] vdd gnd cell_6t
Xbit_r61_c11 bl[11] br[11] wl[61] vdd gnd cell_6t
Xbit_r62_c11 bl[11] br[11] wl[62] vdd gnd cell_6t
Xbit_r63_c11 bl[11] br[11] wl[63] vdd gnd cell_6t
Xbit_r64_c11 bl[11] br[11] wl[64] vdd gnd cell_6t
Xbit_r65_c11 bl[11] br[11] wl[65] vdd gnd cell_6t
Xbit_r66_c11 bl[11] br[11] wl[66] vdd gnd cell_6t
Xbit_r67_c11 bl[11] br[11] wl[67] vdd gnd cell_6t
Xbit_r68_c11 bl[11] br[11] wl[68] vdd gnd cell_6t
Xbit_r69_c11 bl[11] br[11] wl[69] vdd gnd cell_6t
Xbit_r70_c11 bl[11] br[11] wl[70] vdd gnd cell_6t
Xbit_r71_c11 bl[11] br[11] wl[71] vdd gnd cell_6t
Xbit_r72_c11 bl[11] br[11] wl[72] vdd gnd cell_6t
Xbit_r73_c11 bl[11] br[11] wl[73] vdd gnd cell_6t
Xbit_r74_c11 bl[11] br[11] wl[74] vdd gnd cell_6t
Xbit_r75_c11 bl[11] br[11] wl[75] vdd gnd cell_6t
Xbit_r76_c11 bl[11] br[11] wl[76] vdd gnd cell_6t
Xbit_r77_c11 bl[11] br[11] wl[77] vdd gnd cell_6t
Xbit_r78_c11 bl[11] br[11] wl[78] vdd gnd cell_6t
Xbit_r79_c11 bl[11] br[11] wl[79] vdd gnd cell_6t
Xbit_r80_c11 bl[11] br[11] wl[80] vdd gnd cell_6t
Xbit_r81_c11 bl[11] br[11] wl[81] vdd gnd cell_6t
Xbit_r82_c11 bl[11] br[11] wl[82] vdd gnd cell_6t
Xbit_r83_c11 bl[11] br[11] wl[83] vdd gnd cell_6t
Xbit_r84_c11 bl[11] br[11] wl[84] vdd gnd cell_6t
Xbit_r85_c11 bl[11] br[11] wl[85] vdd gnd cell_6t
Xbit_r86_c11 bl[11] br[11] wl[86] vdd gnd cell_6t
Xbit_r87_c11 bl[11] br[11] wl[87] vdd gnd cell_6t
Xbit_r88_c11 bl[11] br[11] wl[88] vdd gnd cell_6t
Xbit_r89_c11 bl[11] br[11] wl[89] vdd gnd cell_6t
Xbit_r90_c11 bl[11] br[11] wl[90] vdd gnd cell_6t
Xbit_r91_c11 bl[11] br[11] wl[91] vdd gnd cell_6t
Xbit_r92_c11 bl[11] br[11] wl[92] vdd gnd cell_6t
Xbit_r93_c11 bl[11] br[11] wl[93] vdd gnd cell_6t
Xbit_r94_c11 bl[11] br[11] wl[94] vdd gnd cell_6t
Xbit_r95_c11 bl[11] br[11] wl[95] vdd gnd cell_6t
Xbit_r96_c11 bl[11] br[11] wl[96] vdd gnd cell_6t
Xbit_r97_c11 bl[11] br[11] wl[97] vdd gnd cell_6t
Xbit_r98_c11 bl[11] br[11] wl[98] vdd gnd cell_6t
Xbit_r99_c11 bl[11] br[11] wl[99] vdd gnd cell_6t
Xbit_r100_c11 bl[11] br[11] wl[100] vdd gnd cell_6t
Xbit_r101_c11 bl[11] br[11] wl[101] vdd gnd cell_6t
Xbit_r102_c11 bl[11] br[11] wl[102] vdd gnd cell_6t
Xbit_r103_c11 bl[11] br[11] wl[103] vdd gnd cell_6t
Xbit_r104_c11 bl[11] br[11] wl[104] vdd gnd cell_6t
Xbit_r105_c11 bl[11] br[11] wl[105] vdd gnd cell_6t
Xbit_r106_c11 bl[11] br[11] wl[106] vdd gnd cell_6t
Xbit_r107_c11 bl[11] br[11] wl[107] vdd gnd cell_6t
Xbit_r108_c11 bl[11] br[11] wl[108] vdd gnd cell_6t
Xbit_r109_c11 bl[11] br[11] wl[109] vdd gnd cell_6t
Xbit_r110_c11 bl[11] br[11] wl[110] vdd gnd cell_6t
Xbit_r111_c11 bl[11] br[11] wl[111] vdd gnd cell_6t
Xbit_r112_c11 bl[11] br[11] wl[112] vdd gnd cell_6t
Xbit_r113_c11 bl[11] br[11] wl[113] vdd gnd cell_6t
Xbit_r114_c11 bl[11] br[11] wl[114] vdd gnd cell_6t
Xbit_r115_c11 bl[11] br[11] wl[115] vdd gnd cell_6t
Xbit_r116_c11 bl[11] br[11] wl[116] vdd gnd cell_6t
Xbit_r117_c11 bl[11] br[11] wl[117] vdd gnd cell_6t
Xbit_r118_c11 bl[11] br[11] wl[118] vdd gnd cell_6t
Xbit_r119_c11 bl[11] br[11] wl[119] vdd gnd cell_6t
Xbit_r120_c11 bl[11] br[11] wl[120] vdd gnd cell_6t
Xbit_r121_c11 bl[11] br[11] wl[121] vdd gnd cell_6t
Xbit_r122_c11 bl[11] br[11] wl[122] vdd gnd cell_6t
Xbit_r123_c11 bl[11] br[11] wl[123] vdd gnd cell_6t
Xbit_r124_c11 bl[11] br[11] wl[124] vdd gnd cell_6t
Xbit_r125_c11 bl[11] br[11] wl[125] vdd gnd cell_6t
Xbit_r126_c11 bl[11] br[11] wl[126] vdd gnd cell_6t
Xbit_r127_c11 bl[11] br[11] wl[127] vdd gnd cell_6t
Xbit_r128_c11 bl[11] br[11] wl[128] vdd gnd cell_6t
Xbit_r129_c11 bl[11] br[11] wl[129] vdd gnd cell_6t
Xbit_r130_c11 bl[11] br[11] wl[130] vdd gnd cell_6t
Xbit_r131_c11 bl[11] br[11] wl[131] vdd gnd cell_6t
Xbit_r132_c11 bl[11] br[11] wl[132] vdd gnd cell_6t
Xbit_r133_c11 bl[11] br[11] wl[133] vdd gnd cell_6t
Xbit_r134_c11 bl[11] br[11] wl[134] vdd gnd cell_6t
Xbit_r135_c11 bl[11] br[11] wl[135] vdd gnd cell_6t
Xbit_r136_c11 bl[11] br[11] wl[136] vdd gnd cell_6t
Xbit_r137_c11 bl[11] br[11] wl[137] vdd gnd cell_6t
Xbit_r138_c11 bl[11] br[11] wl[138] vdd gnd cell_6t
Xbit_r139_c11 bl[11] br[11] wl[139] vdd gnd cell_6t
Xbit_r140_c11 bl[11] br[11] wl[140] vdd gnd cell_6t
Xbit_r141_c11 bl[11] br[11] wl[141] vdd gnd cell_6t
Xbit_r142_c11 bl[11] br[11] wl[142] vdd gnd cell_6t
Xbit_r143_c11 bl[11] br[11] wl[143] vdd gnd cell_6t
Xbit_r144_c11 bl[11] br[11] wl[144] vdd gnd cell_6t
Xbit_r145_c11 bl[11] br[11] wl[145] vdd gnd cell_6t
Xbit_r146_c11 bl[11] br[11] wl[146] vdd gnd cell_6t
Xbit_r147_c11 bl[11] br[11] wl[147] vdd gnd cell_6t
Xbit_r148_c11 bl[11] br[11] wl[148] vdd gnd cell_6t
Xbit_r149_c11 bl[11] br[11] wl[149] vdd gnd cell_6t
Xbit_r150_c11 bl[11] br[11] wl[150] vdd gnd cell_6t
Xbit_r151_c11 bl[11] br[11] wl[151] vdd gnd cell_6t
Xbit_r152_c11 bl[11] br[11] wl[152] vdd gnd cell_6t
Xbit_r153_c11 bl[11] br[11] wl[153] vdd gnd cell_6t
Xbit_r154_c11 bl[11] br[11] wl[154] vdd gnd cell_6t
Xbit_r155_c11 bl[11] br[11] wl[155] vdd gnd cell_6t
Xbit_r156_c11 bl[11] br[11] wl[156] vdd gnd cell_6t
Xbit_r157_c11 bl[11] br[11] wl[157] vdd gnd cell_6t
Xbit_r158_c11 bl[11] br[11] wl[158] vdd gnd cell_6t
Xbit_r159_c11 bl[11] br[11] wl[159] vdd gnd cell_6t
Xbit_r160_c11 bl[11] br[11] wl[160] vdd gnd cell_6t
Xbit_r161_c11 bl[11] br[11] wl[161] vdd gnd cell_6t
Xbit_r162_c11 bl[11] br[11] wl[162] vdd gnd cell_6t
Xbit_r163_c11 bl[11] br[11] wl[163] vdd gnd cell_6t
Xbit_r164_c11 bl[11] br[11] wl[164] vdd gnd cell_6t
Xbit_r165_c11 bl[11] br[11] wl[165] vdd gnd cell_6t
Xbit_r166_c11 bl[11] br[11] wl[166] vdd gnd cell_6t
Xbit_r167_c11 bl[11] br[11] wl[167] vdd gnd cell_6t
Xbit_r168_c11 bl[11] br[11] wl[168] vdd gnd cell_6t
Xbit_r169_c11 bl[11] br[11] wl[169] vdd gnd cell_6t
Xbit_r170_c11 bl[11] br[11] wl[170] vdd gnd cell_6t
Xbit_r171_c11 bl[11] br[11] wl[171] vdd gnd cell_6t
Xbit_r172_c11 bl[11] br[11] wl[172] vdd gnd cell_6t
Xbit_r173_c11 bl[11] br[11] wl[173] vdd gnd cell_6t
Xbit_r174_c11 bl[11] br[11] wl[174] vdd gnd cell_6t
Xbit_r175_c11 bl[11] br[11] wl[175] vdd gnd cell_6t
Xbit_r176_c11 bl[11] br[11] wl[176] vdd gnd cell_6t
Xbit_r177_c11 bl[11] br[11] wl[177] vdd gnd cell_6t
Xbit_r178_c11 bl[11] br[11] wl[178] vdd gnd cell_6t
Xbit_r179_c11 bl[11] br[11] wl[179] vdd gnd cell_6t
Xbit_r180_c11 bl[11] br[11] wl[180] vdd gnd cell_6t
Xbit_r181_c11 bl[11] br[11] wl[181] vdd gnd cell_6t
Xbit_r182_c11 bl[11] br[11] wl[182] vdd gnd cell_6t
Xbit_r183_c11 bl[11] br[11] wl[183] vdd gnd cell_6t
Xbit_r184_c11 bl[11] br[11] wl[184] vdd gnd cell_6t
Xbit_r185_c11 bl[11] br[11] wl[185] vdd gnd cell_6t
Xbit_r186_c11 bl[11] br[11] wl[186] vdd gnd cell_6t
Xbit_r187_c11 bl[11] br[11] wl[187] vdd gnd cell_6t
Xbit_r188_c11 bl[11] br[11] wl[188] vdd gnd cell_6t
Xbit_r189_c11 bl[11] br[11] wl[189] vdd gnd cell_6t
Xbit_r190_c11 bl[11] br[11] wl[190] vdd gnd cell_6t
Xbit_r191_c11 bl[11] br[11] wl[191] vdd gnd cell_6t
Xbit_r192_c11 bl[11] br[11] wl[192] vdd gnd cell_6t
Xbit_r193_c11 bl[11] br[11] wl[193] vdd gnd cell_6t
Xbit_r194_c11 bl[11] br[11] wl[194] vdd gnd cell_6t
Xbit_r195_c11 bl[11] br[11] wl[195] vdd gnd cell_6t
Xbit_r196_c11 bl[11] br[11] wl[196] vdd gnd cell_6t
Xbit_r197_c11 bl[11] br[11] wl[197] vdd gnd cell_6t
Xbit_r198_c11 bl[11] br[11] wl[198] vdd gnd cell_6t
Xbit_r199_c11 bl[11] br[11] wl[199] vdd gnd cell_6t
Xbit_r200_c11 bl[11] br[11] wl[200] vdd gnd cell_6t
Xbit_r201_c11 bl[11] br[11] wl[201] vdd gnd cell_6t
Xbit_r202_c11 bl[11] br[11] wl[202] vdd gnd cell_6t
Xbit_r203_c11 bl[11] br[11] wl[203] vdd gnd cell_6t
Xbit_r204_c11 bl[11] br[11] wl[204] vdd gnd cell_6t
Xbit_r205_c11 bl[11] br[11] wl[205] vdd gnd cell_6t
Xbit_r206_c11 bl[11] br[11] wl[206] vdd gnd cell_6t
Xbit_r207_c11 bl[11] br[11] wl[207] vdd gnd cell_6t
Xbit_r208_c11 bl[11] br[11] wl[208] vdd gnd cell_6t
Xbit_r209_c11 bl[11] br[11] wl[209] vdd gnd cell_6t
Xbit_r210_c11 bl[11] br[11] wl[210] vdd gnd cell_6t
Xbit_r211_c11 bl[11] br[11] wl[211] vdd gnd cell_6t
Xbit_r212_c11 bl[11] br[11] wl[212] vdd gnd cell_6t
Xbit_r213_c11 bl[11] br[11] wl[213] vdd gnd cell_6t
Xbit_r214_c11 bl[11] br[11] wl[214] vdd gnd cell_6t
Xbit_r215_c11 bl[11] br[11] wl[215] vdd gnd cell_6t
Xbit_r216_c11 bl[11] br[11] wl[216] vdd gnd cell_6t
Xbit_r217_c11 bl[11] br[11] wl[217] vdd gnd cell_6t
Xbit_r218_c11 bl[11] br[11] wl[218] vdd gnd cell_6t
Xbit_r219_c11 bl[11] br[11] wl[219] vdd gnd cell_6t
Xbit_r220_c11 bl[11] br[11] wl[220] vdd gnd cell_6t
Xbit_r221_c11 bl[11] br[11] wl[221] vdd gnd cell_6t
Xbit_r222_c11 bl[11] br[11] wl[222] vdd gnd cell_6t
Xbit_r223_c11 bl[11] br[11] wl[223] vdd gnd cell_6t
Xbit_r224_c11 bl[11] br[11] wl[224] vdd gnd cell_6t
Xbit_r225_c11 bl[11] br[11] wl[225] vdd gnd cell_6t
Xbit_r226_c11 bl[11] br[11] wl[226] vdd gnd cell_6t
Xbit_r227_c11 bl[11] br[11] wl[227] vdd gnd cell_6t
Xbit_r228_c11 bl[11] br[11] wl[228] vdd gnd cell_6t
Xbit_r229_c11 bl[11] br[11] wl[229] vdd gnd cell_6t
Xbit_r230_c11 bl[11] br[11] wl[230] vdd gnd cell_6t
Xbit_r231_c11 bl[11] br[11] wl[231] vdd gnd cell_6t
Xbit_r232_c11 bl[11] br[11] wl[232] vdd gnd cell_6t
Xbit_r233_c11 bl[11] br[11] wl[233] vdd gnd cell_6t
Xbit_r234_c11 bl[11] br[11] wl[234] vdd gnd cell_6t
Xbit_r235_c11 bl[11] br[11] wl[235] vdd gnd cell_6t
Xbit_r236_c11 bl[11] br[11] wl[236] vdd gnd cell_6t
Xbit_r237_c11 bl[11] br[11] wl[237] vdd gnd cell_6t
Xbit_r238_c11 bl[11] br[11] wl[238] vdd gnd cell_6t
Xbit_r239_c11 bl[11] br[11] wl[239] vdd gnd cell_6t
Xbit_r240_c11 bl[11] br[11] wl[240] vdd gnd cell_6t
Xbit_r241_c11 bl[11] br[11] wl[241] vdd gnd cell_6t
Xbit_r242_c11 bl[11] br[11] wl[242] vdd gnd cell_6t
Xbit_r243_c11 bl[11] br[11] wl[243] vdd gnd cell_6t
Xbit_r244_c11 bl[11] br[11] wl[244] vdd gnd cell_6t
Xbit_r245_c11 bl[11] br[11] wl[245] vdd gnd cell_6t
Xbit_r246_c11 bl[11] br[11] wl[246] vdd gnd cell_6t
Xbit_r247_c11 bl[11] br[11] wl[247] vdd gnd cell_6t
Xbit_r248_c11 bl[11] br[11] wl[248] vdd gnd cell_6t
Xbit_r249_c11 bl[11] br[11] wl[249] vdd gnd cell_6t
Xbit_r250_c11 bl[11] br[11] wl[250] vdd gnd cell_6t
Xbit_r251_c11 bl[11] br[11] wl[251] vdd gnd cell_6t
Xbit_r252_c11 bl[11] br[11] wl[252] vdd gnd cell_6t
Xbit_r253_c11 bl[11] br[11] wl[253] vdd gnd cell_6t
Xbit_r254_c11 bl[11] br[11] wl[254] vdd gnd cell_6t
Xbit_r255_c11 bl[11] br[11] wl[255] vdd gnd cell_6t
Xbit_r0_c12 bl[12] br[12] wl[0] vdd gnd cell_6t
Xbit_r1_c12 bl[12] br[12] wl[1] vdd gnd cell_6t
Xbit_r2_c12 bl[12] br[12] wl[2] vdd gnd cell_6t
Xbit_r3_c12 bl[12] br[12] wl[3] vdd gnd cell_6t
Xbit_r4_c12 bl[12] br[12] wl[4] vdd gnd cell_6t
Xbit_r5_c12 bl[12] br[12] wl[5] vdd gnd cell_6t
Xbit_r6_c12 bl[12] br[12] wl[6] vdd gnd cell_6t
Xbit_r7_c12 bl[12] br[12] wl[7] vdd gnd cell_6t
Xbit_r8_c12 bl[12] br[12] wl[8] vdd gnd cell_6t
Xbit_r9_c12 bl[12] br[12] wl[9] vdd gnd cell_6t
Xbit_r10_c12 bl[12] br[12] wl[10] vdd gnd cell_6t
Xbit_r11_c12 bl[12] br[12] wl[11] vdd gnd cell_6t
Xbit_r12_c12 bl[12] br[12] wl[12] vdd gnd cell_6t
Xbit_r13_c12 bl[12] br[12] wl[13] vdd gnd cell_6t
Xbit_r14_c12 bl[12] br[12] wl[14] vdd gnd cell_6t
Xbit_r15_c12 bl[12] br[12] wl[15] vdd gnd cell_6t
Xbit_r16_c12 bl[12] br[12] wl[16] vdd gnd cell_6t
Xbit_r17_c12 bl[12] br[12] wl[17] vdd gnd cell_6t
Xbit_r18_c12 bl[12] br[12] wl[18] vdd gnd cell_6t
Xbit_r19_c12 bl[12] br[12] wl[19] vdd gnd cell_6t
Xbit_r20_c12 bl[12] br[12] wl[20] vdd gnd cell_6t
Xbit_r21_c12 bl[12] br[12] wl[21] vdd gnd cell_6t
Xbit_r22_c12 bl[12] br[12] wl[22] vdd gnd cell_6t
Xbit_r23_c12 bl[12] br[12] wl[23] vdd gnd cell_6t
Xbit_r24_c12 bl[12] br[12] wl[24] vdd gnd cell_6t
Xbit_r25_c12 bl[12] br[12] wl[25] vdd gnd cell_6t
Xbit_r26_c12 bl[12] br[12] wl[26] vdd gnd cell_6t
Xbit_r27_c12 bl[12] br[12] wl[27] vdd gnd cell_6t
Xbit_r28_c12 bl[12] br[12] wl[28] vdd gnd cell_6t
Xbit_r29_c12 bl[12] br[12] wl[29] vdd gnd cell_6t
Xbit_r30_c12 bl[12] br[12] wl[30] vdd gnd cell_6t
Xbit_r31_c12 bl[12] br[12] wl[31] vdd gnd cell_6t
Xbit_r32_c12 bl[12] br[12] wl[32] vdd gnd cell_6t
Xbit_r33_c12 bl[12] br[12] wl[33] vdd gnd cell_6t
Xbit_r34_c12 bl[12] br[12] wl[34] vdd gnd cell_6t
Xbit_r35_c12 bl[12] br[12] wl[35] vdd gnd cell_6t
Xbit_r36_c12 bl[12] br[12] wl[36] vdd gnd cell_6t
Xbit_r37_c12 bl[12] br[12] wl[37] vdd gnd cell_6t
Xbit_r38_c12 bl[12] br[12] wl[38] vdd gnd cell_6t
Xbit_r39_c12 bl[12] br[12] wl[39] vdd gnd cell_6t
Xbit_r40_c12 bl[12] br[12] wl[40] vdd gnd cell_6t
Xbit_r41_c12 bl[12] br[12] wl[41] vdd gnd cell_6t
Xbit_r42_c12 bl[12] br[12] wl[42] vdd gnd cell_6t
Xbit_r43_c12 bl[12] br[12] wl[43] vdd gnd cell_6t
Xbit_r44_c12 bl[12] br[12] wl[44] vdd gnd cell_6t
Xbit_r45_c12 bl[12] br[12] wl[45] vdd gnd cell_6t
Xbit_r46_c12 bl[12] br[12] wl[46] vdd gnd cell_6t
Xbit_r47_c12 bl[12] br[12] wl[47] vdd gnd cell_6t
Xbit_r48_c12 bl[12] br[12] wl[48] vdd gnd cell_6t
Xbit_r49_c12 bl[12] br[12] wl[49] vdd gnd cell_6t
Xbit_r50_c12 bl[12] br[12] wl[50] vdd gnd cell_6t
Xbit_r51_c12 bl[12] br[12] wl[51] vdd gnd cell_6t
Xbit_r52_c12 bl[12] br[12] wl[52] vdd gnd cell_6t
Xbit_r53_c12 bl[12] br[12] wl[53] vdd gnd cell_6t
Xbit_r54_c12 bl[12] br[12] wl[54] vdd gnd cell_6t
Xbit_r55_c12 bl[12] br[12] wl[55] vdd gnd cell_6t
Xbit_r56_c12 bl[12] br[12] wl[56] vdd gnd cell_6t
Xbit_r57_c12 bl[12] br[12] wl[57] vdd gnd cell_6t
Xbit_r58_c12 bl[12] br[12] wl[58] vdd gnd cell_6t
Xbit_r59_c12 bl[12] br[12] wl[59] vdd gnd cell_6t
Xbit_r60_c12 bl[12] br[12] wl[60] vdd gnd cell_6t
Xbit_r61_c12 bl[12] br[12] wl[61] vdd gnd cell_6t
Xbit_r62_c12 bl[12] br[12] wl[62] vdd gnd cell_6t
Xbit_r63_c12 bl[12] br[12] wl[63] vdd gnd cell_6t
Xbit_r64_c12 bl[12] br[12] wl[64] vdd gnd cell_6t
Xbit_r65_c12 bl[12] br[12] wl[65] vdd gnd cell_6t
Xbit_r66_c12 bl[12] br[12] wl[66] vdd gnd cell_6t
Xbit_r67_c12 bl[12] br[12] wl[67] vdd gnd cell_6t
Xbit_r68_c12 bl[12] br[12] wl[68] vdd gnd cell_6t
Xbit_r69_c12 bl[12] br[12] wl[69] vdd gnd cell_6t
Xbit_r70_c12 bl[12] br[12] wl[70] vdd gnd cell_6t
Xbit_r71_c12 bl[12] br[12] wl[71] vdd gnd cell_6t
Xbit_r72_c12 bl[12] br[12] wl[72] vdd gnd cell_6t
Xbit_r73_c12 bl[12] br[12] wl[73] vdd gnd cell_6t
Xbit_r74_c12 bl[12] br[12] wl[74] vdd gnd cell_6t
Xbit_r75_c12 bl[12] br[12] wl[75] vdd gnd cell_6t
Xbit_r76_c12 bl[12] br[12] wl[76] vdd gnd cell_6t
Xbit_r77_c12 bl[12] br[12] wl[77] vdd gnd cell_6t
Xbit_r78_c12 bl[12] br[12] wl[78] vdd gnd cell_6t
Xbit_r79_c12 bl[12] br[12] wl[79] vdd gnd cell_6t
Xbit_r80_c12 bl[12] br[12] wl[80] vdd gnd cell_6t
Xbit_r81_c12 bl[12] br[12] wl[81] vdd gnd cell_6t
Xbit_r82_c12 bl[12] br[12] wl[82] vdd gnd cell_6t
Xbit_r83_c12 bl[12] br[12] wl[83] vdd gnd cell_6t
Xbit_r84_c12 bl[12] br[12] wl[84] vdd gnd cell_6t
Xbit_r85_c12 bl[12] br[12] wl[85] vdd gnd cell_6t
Xbit_r86_c12 bl[12] br[12] wl[86] vdd gnd cell_6t
Xbit_r87_c12 bl[12] br[12] wl[87] vdd gnd cell_6t
Xbit_r88_c12 bl[12] br[12] wl[88] vdd gnd cell_6t
Xbit_r89_c12 bl[12] br[12] wl[89] vdd gnd cell_6t
Xbit_r90_c12 bl[12] br[12] wl[90] vdd gnd cell_6t
Xbit_r91_c12 bl[12] br[12] wl[91] vdd gnd cell_6t
Xbit_r92_c12 bl[12] br[12] wl[92] vdd gnd cell_6t
Xbit_r93_c12 bl[12] br[12] wl[93] vdd gnd cell_6t
Xbit_r94_c12 bl[12] br[12] wl[94] vdd gnd cell_6t
Xbit_r95_c12 bl[12] br[12] wl[95] vdd gnd cell_6t
Xbit_r96_c12 bl[12] br[12] wl[96] vdd gnd cell_6t
Xbit_r97_c12 bl[12] br[12] wl[97] vdd gnd cell_6t
Xbit_r98_c12 bl[12] br[12] wl[98] vdd gnd cell_6t
Xbit_r99_c12 bl[12] br[12] wl[99] vdd gnd cell_6t
Xbit_r100_c12 bl[12] br[12] wl[100] vdd gnd cell_6t
Xbit_r101_c12 bl[12] br[12] wl[101] vdd gnd cell_6t
Xbit_r102_c12 bl[12] br[12] wl[102] vdd gnd cell_6t
Xbit_r103_c12 bl[12] br[12] wl[103] vdd gnd cell_6t
Xbit_r104_c12 bl[12] br[12] wl[104] vdd gnd cell_6t
Xbit_r105_c12 bl[12] br[12] wl[105] vdd gnd cell_6t
Xbit_r106_c12 bl[12] br[12] wl[106] vdd gnd cell_6t
Xbit_r107_c12 bl[12] br[12] wl[107] vdd gnd cell_6t
Xbit_r108_c12 bl[12] br[12] wl[108] vdd gnd cell_6t
Xbit_r109_c12 bl[12] br[12] wl[109] vdd gnd cell_6t
Xbit_r110_c12 bl[12] br[12] wl[110] vdd gnd cell_6t
Xbit_r111_c12 bl[12] br[12] wl[111] vdd gnd cell_6t
Xbit_r112_c12 bl[12] br[12] wl[112] vdd gnd cell_6t
Xbit_r113_c12 bl[12] br[12] wl[113] vdd gnd cell_6t
Xbit_r114_c12 bl[12] br[12] wl[114] vdd gnd cell_6t
Xbit_r115_c12 bl[12] br[12] wl[115] vdd gnd cell_6t
Xbit_r116_c12 bl[12] br[12] wl[116] vdd gnd cell_6t
Xbit_r117_c12 bl[12] br[12] wl[117] vdd gnd cell_6t
Xbit_r118_c12 bl[12] br[12] wl[118] vdd gnd cell_6t
Xbit_r119_c12 bl[12] br[12] wl[119] vdd gnd cell_6t
Xbit_r120_c12 bl[12] br[12] wl[120] vdd gnd cell_6t
Xbit_r121_c12 bl[12] br[12] wl[121] vdd gnd cell_6t
Xbit_r122_c12 bl[12] br[12] wl[122] vdd gnd cell_6t
Xbit_r123_c12 bl[12] br[12] wl[123] vdd gnd cell_6t
Xbit_r124_c12 bl[12] br[12] wl[124] vdd gnd cell_6t
Xbit_r125_c12 bl[12] br[12] wl[125] vdd gnd cell_6t
Xbit_r126_c12 bl[12] br[12] wl[126] vdd gnd cell_6t
Xbit_r127_c12 bl[12] br[12] wl[127] vdd gnd cell_6t
Xbit_r128_c12 bl[12] br[12] wl[128] vdd gnd cell_6t
Xbit_r129_c12 bl[12] br[12] wl[129] vdd gnd cell_6t
Xbit_r130_c12 bl[12] br[12] wl[130] vdd gnd cell_6t
Xbit_r131_c12 bl[12] br[12] wl[131] vdd gnd cell_6t
Xbit_r132_c12 bl[12] br[12] wl[132] vdd gnd cell_6t
Xbit_r133_c12 bl[12] br[12] wl[133] vdd gnd cell_6t
Xbit_r134_c12 bl[12] br[12] wl[134] vdd gnd cell_6t
Xbit_r135_c12 bl[12] br[12] wl[135] vdd gnd cell_6t
Xbit_r136_c12 bl[12] br[12] wl[136] vdd gnd cell_6t
Xbit_r137_c12 bl[12] br[12] wl[137] vdd gnd cell_6t
Xbit_r138_c12 bl[12] br[12] wl[138] vdd gnd cell_6t
Xbit_r139_c12 bl[12] br[12] wl[139] vdd gnd cell_6t
Xbit_r140_c12 bl[12] br[12] wl[140] vdd gnd cell_6t
Xbit_r141_c12 bl[12] br[12] wl[141] vdd gnd cell_6t
Xbit_r142_c12 bl[12] br[12] wl[142] vdd gnd cell_6t
Xbit_r143_c12 bl[12] br[12] wl[143] vdd gnd cell_6t
Xbit_r144_c12 bl[12] br[12] wl[144] vdd gnd cell_6t
Xbit_r145_c12 bl[12] br[12] wl[145] vdd gnd cell_6t
Xbit_r146_c12 bl[12] br[12] wl[146] vdd gnd cell_6t
Xbit_r147_c12 bl[12] br[12] wl[147] vdd gnd cell_6t
Xbit_r148_c12 bl[12] br[12] wl[148] vdd gnd cell_6t
Xbit_r149_c12 bl[12] br[12] wl[149] vdd gnd cell_6t
Xbit_r150_c12 bl[12] br[12] wl[150] vdd gnd cell_6t
Xbit_r151_c12 bl[12] br[12] wl[151] vdd gnd cell_6t
Xbit_r152_c12 bl[12] br[12] wl[152] vdd gnd cell_6t
Xbit_r153_c12 bl[12] br[12] wl[153] vdd gnd cell_6t
Xbit_r154_c12 bl[12] br[12] wl[154] vdd gnd cell_6t
Xbit_r155_c12 bl[12] br[12] wl[155] vdd gnd cell_6t
Xbit_r156_c12 bl[12] br[12] wl[156] vdd gnd cell_6t
Xbit_r157_c12 bl[12] br[12] wl[157] vdd gnd cell_6t
Xbit_r158_c12 bl[12] br[12] wl[158] vdd gnd cell_6t
Xbit_r159_c12 bl[12] br[12] wl[159] vdd gnd cell_6t
Xbit_r160_c12 bl[12] br[12] wl[160] vdd gnd cell_6t
Xbit_r161_c12 bl[12] br[12] wl[161] vdd gnd cell_6t
Xbit_r162_c12 bl[12] br[12] wl[162] vdd gnd cell_6t
Xbit_r163_c12 bl[12] br[12] wl[163] vdd gnd cell_6t
Xbit_r164_c12 bl[12] br[12] wl[164] vdd gnd cell_6t
Xbit_r165_c12 bl[12] br[12] wl[165] vdd gnd cell_6t
Xbit_r166_c12 bl[12] br[12] wl[166] vdd gnd cell_6t
Xbit_r167_c12 bl[12] br[12] wl[167] vdd gnd cell_6t
Xbit_r168_c12 bl[12] br[12] wl[168] vdd gnd cell_6t
Xbit_r169_c12 bl[12] br[12] wl[169] vdd gnd cell_6t
Xbit_r170_c12 bl[12] br[12] wl[170] vdd gnd cell_6t
Xbit_r171_c12 bl[12] br[12] wl[171] vdd gnd cell_6t
Xbit_r172_c12 bl[12] br[12] wl[172] vdd gnd cell_6t
Xbit_r173_c12 bl[12] br[12] wl[173] vdd gnd cell_6t
Xbit_r174_c12 bl[12] br[12] wl[174] vdd gnd cell_6t
Xbit_r175_c12 bl[12] br[12] wl[175] vdd gnd cell_6t
Xbit_r176_c12 bl[12] br[12] wl[176] vdd gnd cell_6t
Xbit_r177_c12 bl[12] br[12] wl[177] vdd gnd cell_6t
Xbit_r178_c12 bl[12] br[12] wl[178] vdd gnd cell_6t
Xbit_r179_c12 bl[12] br[12] wl[179] vdd gnd cell_6t
Xbit_r180_c12 bl[12] br[12] wl[180] vdd gnd cell_6t
Xbit_r181_c12 bl[12] br[12] wl[181] vdd gnd cell_6t
Xbit_r182_c12 bl[12] br[12] wl[182] vdd gnd cell_6t
Xbit_r183_c12 bl[12] br[12] wl[183] vdd gnd cell_6t
Xbit_r184_c12 bl[12] br[12] wl[184] vdd gnd cell_6t
Xbit_r185_c12 bl[12] br[12] wl[185] vdd gnd cell_6t
Xbit_r186_c12 bl[12] br[12] wl[186] vdd gnd cell_6t
Xbit_r187_c12 bl[12] br[12] wl[187] vdd gnd cell_6t
Xbit_r188_c12 bl[12] br[12] wl[188] vdd gnd cell_6t
Xbit_r189_c12 bl[12] br[12] wl[189] vdd gnd cell_6t
Xbit_r190_c12 bl[12] br[12] wl[190] vdd gnd cell_6t
Xbit_r191_c12 bl[12] br[12] wl[191] vdd gnd cell_6t
Xbit_r192_c12 bl[12] br[12] wl[192] vdd gnd cell_6t
Xbit_r193_c12 bl[12] br[12] wl[193] vdd gnd cell_6t
Xbit_r194_c12 bl[12] br[12] wl[194] vdd gnd cell_6t
Xbit_r195_c12 bl[12] br[12] wl[195] vdd gnd cell_6t
Xbit_r196_c12 bl[12] br[12] wl[196] vdd gnd cell_6t
Xbit_r197_c12 bl[12] br[12] wl[197] vdd gnd cell_6t
Xbit_r198_c12 bl[12] br[12] wl[198] vdd gnd cell_6t
Xbit_r199_c12 bl[12] br[12] wl[199] vdd gnd cell_6t
Xbit_r200_c12 bl[12] br[12] wl[200] vdd gnd cell_6t
Xbit_r201_c12 bl[12] br[12] wl[201] vdd gnd cell_6t
Xbit_r202_c12 bl[12] br[12] wl[202] vdd gnd cell_6t
Xbit_r203_c12 bl[12] br[12] wl[203] vdd gnd cell_6t
Xbit_r204_c12 bl[12] br[12] wl[204] vdd gnd cell_6t
Xbit_r205_c12 bl[12] br[12] wl[205] vdd gnd cell_6t
Xbit_r206_c12 bl[12] br[12] wl[206] vdd gnd cell_6t
Xbit_r207_c12 bl[12] br[12] wl[207] vdd gnd cell_6t
Xbit_r208_c12 bl[12] br[12] wl[208] vdd gnd cell_6t
Xbit_r209_c12 bl[12] br[12] wl[209] vdd gnd cell_6t
Xbit_r210_c12 bl[12] br[12] wl[210] vdd gnd cell_6t
Xbit_r211_c12 bl[12] br[12] wl[211] vdd gnd cell_6t
Xbit_r212_c12 bl[12] br[12] wl[212] vdd gnd cell_6t
Xbit_r213_c12 bl[12] br[12] wl[213] vdd gnd cell_6t
Xbit_r214_c12 bl[12] br[12] wl[214] vdd gnd cell_6t
Xbit_r215_c12 bl[12] br[12] wl[215] vdd gnd cell_6t
Xbit_r216_c12 bl[12] br[12] wl[216] vdd gnd cell_6t
Xbit_r217_c12 bl[12] br[12] wl[217] vdd gnd cell_6t
Xbit_r218_c12 bl[12] br[12] wl[218] vdd gnd cell_6t
Xbit_r219_c12 bl[12] br[12] wl[219] vdd gnd cell_6t
Xbit_r220_c12 bl[12] br[12] wl[220] vdd gnd cell_6t
Xbit_r221_c12 bl[12] br[12] wl[221] vdd gnd cell_6t
Xbit_r222_c12 bl[12] br[12] wl[222] vdd gnd cell_6t
Xbit_r223_c12 bl[12] br[12] wl[223] vdd gnd cell_6t
Xbit_r224_c12 bl[12] br[12] wl[224] vdd gnd cell_6t
Xbit_r225_c12 bl[12] br[12] wl[225] vdd gnd cell_6t
Xbit_r226_c12 bl[12] br[12] wl[226] vdd gnd cell_6t
Xbit_r227_c12 bl[12] br[12] wl[227] vdd gnd cell_6t
Xbit_r228_c12 bl[12] br[12] wl[228] vdd gnd cell_6t
Xbit_r229_c12 bl[12] br[12] wl[229] vdd gnd cell_6t
Xbit_r230_c12 bl[12] br[12] wl[230] vdd gnd cell_6t
Xbit_r231_c12 bl[12] br[12] wl[231] vdd gnd cell_6t
Xbit_r232_c12 bl[12] br[12] wl[232] vdd gnd cell_6t
Xbit_r233_c12 bl[12] br[12] wl[233] vdd gnd cell_6t
Xbit_r234_c12 bl[12] br[12] wl[234] vdd gnd cell_6t
Xbit_r235_c12 bl[12] br[12] wl[235] vdd gnd cell_6t
Xbit_r236_c12 bl[12] br[12] wl[236] vdd gnd cell_6t
Xbit_r237_c12 bl[12] br[12] wl[237] vdd gnd cell_6t
Xbit_r238_c12 bl[12] br[12] wl[238] vdd gnd cell_6t
Xbit_r239_c12 bl[12] br[12] wl[239] vdd gnd cell_6t
Xbit_r240_c12 bl[12] br[12] wl[240] vdd gnd cell_6t
Xbit_r241_c12 bl[12] br[12] wl[241] vdd gnd cell_6t
Xbit_r242_c12 bl[12] br[12] wl[242] vdd gnd cell_6t
Xbit_r243_c12 bl[12] br[12] wl[243] vdd gnd cell_6t
Xbit_r244_c12 bl[12] br[12] wl[244] vdd gnd cell_6t
Xbit_r245_c12 bl[12] br[12] wl[245] vdd gnd cell_6t
Xbit_r246_c12 bl[12] br[12] wl[246] vdd gnd cell_6t
Xbit_r247_c12 bl[12] br[12] wl[247] vdd gnd cell_6t
Xbit_r248_c12 bl[12] br[12] wl[248] vdd gnd cell_6t
Xbit_r249_c12 bl[12] br[12] wl[249] vdd gnd cell_6t
Xbit_r250_c12 bl[12] br[12] wl[250] vdd gnd cell_6t
Xbit_r251_c12 bl[12] br[12] wl[251] vdd gnd cell_6t
Xbit_r252_c12 bl[12] br[12] wl[252] vdd gnd cell_6t
Xbit_r253_c12 bl[12] br[12] wl[253] vdd gnd cell_6t
Xbit_r254_c12 bl[12] br[12] wl[254] vdd gnd cell_6t
Xbit_r255_c12 bl[12] br[12] wl[255] vdd gnd cell_6t
Xbit_r0_c13 bl[13] br[13] wl[0] vdd gnd cell_6t
Xbit_r1_c13 bl[13] br[13] wl[1] vdd gnd cell_6t
Xbit_r2_c13 bl[13] br[13] wl[2] vdd gnd cell_6t
Xbit_r3_c13 bl[13] br[13] wl[3] vdd gnd cell_6t
Xbit_r4_c13 bl[13] br[13] wl[4] vdd gnd cell_6t
Xbit_r5_c13 bl[13] br[13] wl[5] vdd gnd cell_6t
Xbit_r6_c13 bl[13] br[13] wl[6] vdd gnd cell_6t
Xbit_r7_c13 bl[13] br[13] wl[7] vdd gnd cell_6t
Xbit_r8_c13 bl[13] br[13] wl[8] vdd gnd cell_6t
Xbit_r9_c13 bl[13] br[13] wl[9] vdd gnd cell_6t
Xbit_r10_c13 bl[13] br[13] wl[10] vdd gnd cell_6t
Xbit_r11_c13 bl[13] br[13] wl[11] vdd gnd cell_6t
Xbit_r12_c13 bl[13] br[13] wl[12] vdd gnd cell_6t
Xbit_r13_c13 bl[13] br[13] wl[13] vdd gnd cell_6t
Xbit_r14_c13 bl[13] br[13] wl[14] vdd gnd cell_6t
Xbit_r15_c13 bl[13] br[13] wl[15] vdd gnd cell_6t
Xbit_r16_c13 bl[13] br[13] wl[16] vdd gnd cell_6t
Xbit_r17_c13 bl[13] br[13] wl[17] vdd gnd cell_6t
Xbit_r18_c13 bl[13] br[13] wl[18] vdd gnd cell_6t
Xbit_r19_c13 bl[13] br[13] wl[19] vdd gnd cell_6t
Xbit_r20_c13 bl[13] br[13] wl[20] vdd gnd cell_6t
Xbit_r21_c13 bl[13] br[13] wl[21] vdd gnd cell_6t
Xbit_r22_c13 bl[13] br[13] wl[22] vdd gnd cell_6t
Xbit_r23_c13 bl[13] br[13] wl[23] vdd gnd cell_6t
Xbit_r24_c13 bl[13] br[13] wl[24] vdd gnd cell_6t
Xbit_r25_c13 bl[13] br[13] wl[25] vdd gnd cell_6t
Xbit_r26_c13 bl[13] br[13] wl[26] vdd gnd cell_6t
Xbit_r27_c13 bl[13] br[13] wl[27] vdd gnd cell_6t
Xbit_r28_c13 bl[13] br[13] wl[28] vdd gnd cell_6t
Xbit_r29_c13 bl[13] br[13] wl[29] vdd gnd cell_6t
Xbit_r30_c13 bl[13] br[13] wl[30] vdd gnd cell_6t
Xbit_r31_c13 bl[13] br[13] wl[31] vdd gnd cell_6t
Xbit_r32_c13 bl[13] br[13] wl[32] vdd gnd cell_6t
Xbit_r33_c13 bl[13] br[13] wl[33] vdd gnd cell_6t
Xbit_r34_c13 bl[13] br[13] wl[34] vdd gnd cell_6t
Xbit_r35_c13 bl[13] br[13] wl[35] vdd gnd cell_6t
Xbit_r36_c13 bl[13] br[13] wl[36] vdd gnd cell_6t
Xbit_r37_c13 bl[13] br[13] wl[37] vdd gnd cell_6t
Xbit_r38_c13 bl[13] br[13] wl[38] vdd gnd cell_6t
Xbit_r39_c13 bl[13] br[13] wl[39] vdd gnd cell_6t
Xbit_r40_c13 bl[13] br[13] wl[40] vdd gnd cell_6t
Xbit_r41_c13 bl[13] br[13] wl[41] vdd gnd cell_6t
Xbit_r42_c13 bl[13] br[13] wl[42] vdd gnd cell_6t
Xbit_r43_c13 bl[13] br[13] wl[43] vdd gnd cell_6t
Xbit_r44_c13 bl[13] br[13] wl[44] vdd gnd cell_6t
Xbit_r45_c13 bl[13] br[13] wl[45] vdd gnd cell_6t
Xbit_r46_c13 bl[13] br[13] wl[46] vdd gnd cell_6t
Xbit_r47_c13 bl[13] br[13] wl[47] vdd gnd cell_6t
Xbit_r48_c13 bl[13] br[13] wl[48] vdd gnd cell_6t
Xbit_r49_c13 bl[13] br[13] wl[49] vdd gnd cell_6t
Xbit_r50_c13 bl[13] br[13] wl[50] vdd gnd cell_6t
Xbit_r51_c13 bl[13] br[13] wl[51] vdd gnd cell_6t
Xbit_r52_c13 bl[13] br[13] wl[52] vdd gnd cell_6t
Xbit_r53_c13 bl[13] br[13] wl[53] vdd gnd cell_6t
Xbit_r54_c13 bl[13] br[13] wl[54] vdd gnd cell_6t
Xbit_r55_c13 bl[13] br[13] wl[55] vdd gnd cell_6t
Xbit_r56_c13 bl[13] br[13] wl[56] vdd gnd cell_6t
Xbit_r57_c13 bl[13] br[13] wl[57] vdd gnd cell_6t
Xbit_r58_c13 bl[13] br[13] wl[58] vdd gnd cell_6t
Xbit_r59_c13 bl[13] br[13] wl[59] vdd gnd cell_6t
Xbit_r60_c13 bl[13] br[13] wl[60] vdd gnd cell_6t
Xbit_r61_c13 bl[13] br[13] wl[61] vdd gnd cell_6t
Xbit_r62_c13 bl[13] br[13] wl[62] vdd gnd cell_6t
Xbit_r63_c13 bl[13] br[13] wl[63] vdd gnd cell_6t
Xbit_r64_c13 bl[13] br[13] wl[64] vdd gnd cell_6t
Xbit_r65_c13 bl[13] br[13] wl[65] vdd gnd cell_6t
Xbit_r66_c13 bl[13] br[13] wl[66] vdd gnd cell_6t
Xbit_r67_c13 bl[13] br[13] wl[67] vdd gnd cell_6t
Xbit_r68_c13 bl[13] br[13] wl[68] vdd gnd cell_6t
Xbit_r69_c13 bl[13] br[13] wl[69] vdd gnd cell_6t
Xbit_r70_c13 bl[13] br[13] wl[70] vdd gnd cell_6t
Xbit_r71_c13 bl[13] br[13] wl[71] vdd gnd cell_6t
Xbit_r72_c13 bl[13] br[13] wl[72] vdd gnd cell_6t
Xbit_r73_c13 bl[13] br[13] wl[73] vdd gnd cell_6t
Xbit_r74_c13 bl[13] br[13] wl[74] vdd gnd cell_6t
Xbit_r75_c13 bl[13] br[13] wl[75] vdd gnd cell_6t
Xbit_r76_c13 bl[13] br[13] wl[76] vdd gnd cell_6t
Xbit_r77_c13 bl[13] br[13] wl[77] vdd gnd cell_6t
Xbit_r78_c13 bl[13] br[13] wl[78] vdd gnd cell_6t
Xbit_r79_c13 bl[13] br[13] wl[79] vdd gnd cell_6t
Xbit_r80_c13 bl[13] br[13] wl[80] vdd gnd cell_6t
Xbit_r81_c13 bl[13] br[13] wl[81] vdd gnd cell_6t
Xbit_r82_c13 bl[13] br[13] wl[82] vdd gnd cell_6t
Xbit_r83_c13 bl[13] br[13] wl[83] vdd gnd cell_6t
Xbit_r84_c13 bl[13] br[13] wl[84] vdd gnd cell_6t
Xbit_r85_c13 bl[13] br[13] wl[85] vdd gnd cell_6t
Xbit_r86_c13 bl[13] br[13] wl[86] vdd gnd cell_6t
Xbit_r87_c13 bl[13] br[13] wl[87] vdd gnd cell_6t
Xbit_r88_c13 bl[13] br[13] wl[88] vdd gnd cell_6t
Xbit_r89_c13 bl[13] br[13] wl[89] vdd gnd cell_6t
Xbit_r90_c13 bl[13] br[13] wl[90] vdd gnd cell_6t
Xbit_r91_c13 bl[13] br[13] wl[91] vdd gnd cell_6t
Xbit_r92_c13 bl[13] br[13] wl[92] vdd gnd cell_6t
Xbit_r93_c13 bl[13] br[13] wl[93] vdd gnd cell_6t
Xbit_r94_c13 bl[13] br[13] wl[94] vdd gnd cell_6t
Xbit_r95_c13 bl[13] br[13] wl[95] vdd gnd cell_6t
Xbit_r96_c13 bl[13] br[13] wl[96] vdd gnd cell_6t
Xbit_r97_c13 bl[13] br[13] wl[97] vdd gnd cell_6t
Xbit_r98_c13 bl[13] br[13] wl[98] vdd gnd cell_6t
Xbit_r99_c13 bl[13] br[13] wl[99] vdd gnd cell_6t
Xbit_r100_c13 bl[13] br[13] wl[100] vdd gnd cell_6t
Xbit_r101_c13 bl[13] br[13] wl[101] vdd gnd cell_6t
Xbit_r102_c13 bl[13] br[13] wl[102] vdd gnd cell_6t
Xbit_r103_c13 bl[13] br[13] wl[103] vdd gnd cell_6t
Xbit_r104_c13 bl[13] br[13] wl[104] vdd gnd cell_6t
Xbit_r105_c13 bl[13] br[13] wl[105] vdd gnd cell_6t
Xbit_r106_c13 bl[13] br[13] wl[106] vdd gnd cell_6t
Xbit_r107_c13 bl[13] br[13] wl[107] vdd gnd cell_6t
Xbit_r108_c13 bl[13] br[13] wl[108] vdd gnd cell_6t
Xbit_r109_c13 bl[13] br[13] wl[109] vdd gnd cell_6t
Xbit_r110_c13 bl[13] br[13] wl[110] vdd gnd cell_6t
Xbit_r111_c13 bl[13] br[13] wl[111] vdd gnd cell_6t
Xbit_r112_c13 bl[13] br[13] wl[112] vdd gnd cell_6t
Xbit_r113_c13 bl[13] br[13] wl[113] vdd gnd cell_6t
Xbit_r114_c13 bl[13] br[13] wl[114] vdd gnd cell_6t
Xbit_r115_c13 bl[13] br[13] wl[115] vdd gnd cell_6t
Xbit_r116_c13 bl[13] br[13] wl[116] vdd gnd cell_6t
Xbit_r117_c13 bl[13] br[13] wl[117] vdd gnd cell_6t
Xbit_r118_c13 bl[13] br[13] wl[118] vdd gnd cell_6t
Xbit_r119_c13 bl[13] br[13] wl[119] vdd gnd cell_6t
Xbit_r120_c13 bl[13] br[13] wl[120] vdd gnd cell_6t
Xbit_r121_c13 bl[13] br[13] wl[121] vdd gnd cell_6t
Xbit_r122_c13 bl[13] br[13] wl[122] vdd gnd cell_6t
Xbit_r123_c13 bl[13] br[13] wl[123] vdd gnd cell_6t
Xbit_r124_c13 bl[13] br[13] wl[124] vdd gnd cell_6t
Xbit_r125_c13 bl[13] br[13] wl[125] vdd gnd cell_6t
Xbit_r126_c13 bl[13] br[13] wl[126] vdd gnd cell_6t
Xbit_r127_c13 bl[13] br[13] wl[127] vdd gnd cell_6t
Xbit_r128_c13 bl[13] br[13] wl[128] vdd gnd cell_6t
Xbit_r129_c13 bl[13] br[13] wl[129] vdd gnd cell_6t
Xbit_r130_c13 bl[13] br[13] wl[130] vdd gnd cell_6t
Xbit_r131_c13 bl[13] br[13] wl[131] vdd gnd cell_6t
Xbit_r132_c13 bl[13] br[13] wl[132] vdd gnd cell_6t
Xbit_r133_c13 bl[13] br[13] wl[133] vdd gnd cell_6t
Xbit_r134_c13 bl[13] br[13] wl[134] vdd gnd cell_6t
Xbit_r135_c13 bl[13] br[13] wl[135] vdd gnd cell_6t
Xbit_r136_c13 bl[13] br[13] wl[136] vdd gnd cell_6t
Xbit_r137_c13 bl[13] br[13] wl[137] vdd gnd cell_6t
Xbit_r138_c13 bl[13] br[13] wl[138] vdd gnd cell_6t
Xbit_r139_c13 bl[13] br[13] wl[139] vdd gnd cell_6t
Xbit_r140_c13 bl[13] br[13] wl[140] vdd gnd cell_6t
Xbit_r141_c13 bl[13] br[13] wl[141] vdd gnd cell_6t
Xbit_r142_c13 bl[13] br[13] wl[142] vdd gnd cell_6t
Xbit_r143_c13 bl[13] br[13] wl[143] vdd gnd cell_6t
Xbit_r144_c13 bl[13] br[13] wl[144] vdd gnd cell_6t
Xbit_r145_c13 bl[13] br[13] wl[145] vdd gnd cell_6t
Xbit_r146_c13 bl[13] br[13] wl[146] vdd gnd cell_6t
Xbit_r147_c13 bl[13] br[13] wl[147] vdd gnd cell_6t
Xbit_r148_c13 bl[13] br[13] wl[148] vdd gnd cell_6t
Xbit_r149_c13 bl[13] br[13] wl[149] vdd gnd cell_6t
Xbit_r150_c13 bl[13] br[13] wl[150] vdd gnd cell_6t
Xbit_r151_c13 bl[13] br[13] wl[151] vdd gnd cell_6t
Xbit_r152_c13 bl[13] br[13] wl[152] vdd gnd cell_6t
Xbit_r153_c13 bl[13] br[13] wl[153] vdd gnd cell_6t
Xbit_r154_c13 bl[13] br[13] wl[154] vdd gnd cell_6t
Xbit_r155_c13 bl[13] br[13] wl[155] vdd gnd cell_6t
Xbit_r156_c13 bl[13] br[13] wl[156] vdd gnd cell_6t
Xbit_r157_c13 bl[13] br[13] wl[157] vdd gnd cell_6t
Xbit_r158_c13 bl[13] br[13] wl[158] vdd gnd cell_6t
Xbit_r159_c13 bl[13] br[13] wl[159] vdd gnd cell_6t
Xbit_r160_c13 bl[13] br[13] wl[160] vdd gnd cell_6t
Xbit_r161_c13 bl[13] br[13] wl[161] vdd gnd cell_6t
Xbit_r162_c13 bl[13] br[13] wl[162] vdd gnd cell_6t
Xbit_r163_c13 bl[13] br[13] wl[163] vdd gnd cell_6t
Xbit_r164_c13 bl[13] br[13] wl[164] vdd gnd cell_6t
Xbit_r165_c13 bl[13] br[13] wl[165] vdd gnd cell_6t
Xbit_r166_c13 bl[13] br[13] wl[166] vdd gnd cell_6t
Xbit_r167_c13 bl[13] br[13] wl[167] vdd gnd cell_6t
Xbit_r168_c13 bl[13] br[13] wl[168] vdd gnd cell_6t
Xbit_r169_c13 bl[13] br[13] wl[169] vdd gnd cell_6t
Xbit_r170_c13 bl[13] br[13] wl[170] vdd gnd cell_6t
Xbit_r171_c13 bl[13] br[13] wl[171] vdd gnd cell_6t
Xbit_r172_c13 bl[13] br[13] wl[172] vdd gnd cell_6t
Xbit_r173_c13 bl[13] br[13] wl[173] vdd gnd cell_6t
Xbit_r174_c13 bl[13] br[13] wl[174] vdd gnd cell_6t
Xbit_r175_c13 bl[13] br[13] wl[175] vdd gnd cell_6t
Xbit_r176_c13 bl[13] br[13] wl[176] vdd gnd cell_6t
Xbit_r177_c13 bl[13] br[13] wl[177] vdd gnd cell_6t
Xbit_r178_c13 bl[13] br[13] wl[178] vdd gnd cell_6t
Xbit_r179_c13 bl[13] br[13] wl[179] vdd gnd cell_6t
Xbit_r180_c13 bl[13] br[13] wl[180] vdd gnd cell_6t
Xbit_r181_c13 bl[13] br[13] wl[181] vdd gnd cell_6t
Xbit_r182_c13 bl[13] br[13] wl[182] vdd gnd cell_6t
Xbit_r183_c13 bl[13] br[13] wl[183] vdd gnd cell_6t
Xbit_r184_c13 bl[13] br[13] wl[184] vdd gnd cell_6t
Xbit_r185_c13 bl[13] br[13] wl[185] vdd gnd cell_6t
Xbit_r186_c13 bl[13] br[13] wl[186] vdd gnd cell_6t
Xbit_r187_c13 bl[13] br[13] wl[187] vdd gnd cell_6t
Xbit_r188_c13 bl[13] br[13] wl[188] vdd gnd cell_6t
Xbit_r189_c13 bl[13] br[13] wl[189] vdd gnd cell_6t
Xbit_r190_c13 bl[13] br[13] wl[190] vdd gnd cell_6t
Xbit_r191_c13 bl[13] br[13] wl[191] vdd gnd cell_6t
Xbit_r192_c13 bl[13] br[13] wl[192] vdd gnd cell_6t
Xbit_r193_c13 bl[13] br[13] wl[193] vdd gnd cell_6t
Xbit_r194_c13 bl[13] br[13] wl[194] vdd gnd cell_6t
Xbit_r195_c13 bl[13] br[13] wl[195] vdd gnd cell_6t
Xbit_r196_c13 bl[13] br[13] wl[196] vdd gnd cell_6t
Xbit_r197_c13 bl[13] br[13] wl[197] vdd gnd cell_6t
Xbit_r198_c13 bl[13] br[13] wl[198] vdd gnd cell_6t
Xbit_r199_c13 bl[13] br[13] wl[199] vdd gnd cell_6t
Xbit_r200_c13 bl[13] br[13] wl[200] vdd gnd cell_6t
Xbit_r201_c13 bl[13] br[13] wl[201] vdd gnd cell_6t
Xbit_r202_c13 bl[13] br[13] wl[202] vdd gnd cell_6t
Xbit_r203_c13 bl[13] br[13] wl[203] vdd gnd cell_6t
Xbit_r204_c13 bl[13] br[13] wl[204] vdd gnd cell_6t
Xbit_r205_c13 bl[13] br[13] wl[205] vdd gnd cell_6t
Xbit_r206_c13 bl[13] br[13] wl[206] vdd gnd cell_6t
Xbit_r207_c13 bl[13] br[13] wl[207] vdd gnd cell_6t
Xbit_r208_c13 bl[13] br[13] wl[208] vdd gnd cell_6t
Xbit_r209_c13 bl[13] br[13] wl[209] vdd gnd cell_6t
Xbit_r210_c13 bl[13] br[13] wl[210] vdd gnd cell_6t
Xbit_r211_c13 bl[13] br[13] wl[211] vdd gnd cell_6t
Xbit_r212_c13 bl[13] br[13] wl[212] vdd gnd cell_6t
Xbit_r213_c13 bl[13] br[13] wl[213] vdd gnd cell_6t
Xbit_r214_c13 bl[13] br[13] wl[214] vdd gnd cell_6t
Xbit_r215_c13 bl[13] br[13] wl[215] vdd gnd cell_6t
Xbit_r216_c13 bl[13] br[13] wl[216] vdd gnd cell_6t
Xbit_r217_c13 bl[13] br[13] wl[217] vdd gnd cell_6t
Xbit_r218_c13 bl[13] br[13] wl[218] vdd gnd cell_6t
Xbit_r219_c13 bl[13] br[13] wl[219] vdd gnd cell_6t
Xbit_r220_c13 bl[13] br[13] wl[220] vdd gnd cell_6t
Xbit_r221_c13 bl[13] br[13] wl[221] vdd gnd cell_6t
Xbit_r222_c13 bl[13] br[13] wl[222] vdd gnd cell_6t
Xbit_r223_c13 bl[13] br[13] wl[223] vdd gnd cell_6t
Xbit_r224_c13 bl[13] br[13] wl[224] vdd gnd cell_6t
Xbit_r225_c13 bl[13] br[13] wl[225] vdd gnd cell_6t
Xbit_r226_c13 bl[13] br[13] wl[226] vdd gnd cell_6t
Xbit_r227_c13 bl[13] br[13] wl[227] vdd gnd cell_6t
Xbit_r228_c13 bl[13] br[13] wl[228] vdd gnd cell_6t
Xbit_r229_c13 bl[13] br[13] wl[229] vdd gnd cell_6t
Xbit_r230_c13 bl[13] br[13] wl[230] vdd gnd cell_6t
Xbit_r231_c13 bl[13] br[13] wl[231] vdd gnd cell_6t
Xbit_r232_c13 bl[13] br[13] wl[232] vdd gnd cell_6t
Xbit_r233_c13 bl[13] br[13] wl[233] vdd gnd cell_6t
Xbit_r234_c13 bl[13] br[13] wl[234] vdd gnd cell_6t
Xbit_r235_c13 bl[13] br[13] wl[235] vdd gnd cell_6t
Xbit_r236_c13 bl[13] br[13] wl[236] vdd gnd cell_6t
Xbit_r237_c13 bl[13] br[13] wl[237] vdd gnd cell_6t
Xbit_r238_c13 bl[13] br[13] wl[238] vdd gnd cell_6t
Xbit_r239_c13 bl[13] br[13] wl[239] vdd gnd cell_6t
Xbit_r240_c13 bl[13] br[13] wl[240] vdd gnd cell_6t
Xbit_r241_c13 bl[13] br[13] wl[241] vdd gnd cell_6t
Xbit_r242_c13 bl[13] br[13] wl[242] vdd gnd cell_6t
Xbit_r243_c13 bl[13] br[13] wl[243] vdd gnd cell_6t
Xbit_r244_c13 bl[13] br[13] wl[244] vdd gnd cell_6t
Xbit_r245_c13 bl[13] br[13] wl[245] vdd gnd cell_6t
Xbit_r246_c13 bl[13] br[13] wl[246] vdd gnd cell_6t
Xbit_r247_c13 bl[13] br[13] wl[247] vdd gnd cell_6t
Xbit_r248_c13 bl[13] br[13] wl[248] vdd gnd cell_6t
Xbit_r249_c13 bl[13] br[13] wl[249] vdd gnd cell_6t
Xbit_r250_c13 bl[13] br[13] wl[250] vdd gnd cell_6t
Xbit_r251_c13 bl[13] br[13] wl[251] vdd gnd cell_6t
Xbit_r252_c13 bl[13] br[13] wl[252] vdd gnd cell_6t
Xbit_r253_c13 bl[13] br[13] wl[253] vdd gnd cell_6t
Xbit_r254_c13 bl[13] br[13] wl[254] vdd gnd cell_6t
Xbit_r255_c13 bl[13] br[13] wl[255] vdd gnd cell_6t
Xbit_r0_c14 bl[14] br[14] wl[0] vdd gnd cell_6t
Xbit_r1_c14 bl[14] br[14] wl[1] vdd gnd cell_6t
Xbit_r2_c14 bl[14] br[14] wl[2] vdd gnd cell_6t
Xbit_r3_c14 bl[14] br[14] wl[3] vdd gnd cell_6t
Xbit_r4_c14 bl[14] br[14] wl[4] vdd gnd cell_6t
Xbit_r5_c14 bl[14] br[14] wl[5] vdd gnd cell_6t
Xbit_r6_c14 bl[14] br[14] wl[6] vdd gnd cell_6t
Xbit_r7_c14 bl[14] br[14] wl[7] vdd gnd cell_6t
Xbit_r8_c14 bl[14] br[14] wl[8] vdd gnd cell_6t
Xbit_r9_c14 bl[14] br[14] wl[9] vdd gnd cell_6t
Xbit_r10_c14 bl[14] br[14] wl[10] vdd gnd cell_6t
Xbit_r11_c14 bl[14] br[14] wl[11] vdd gnd cell_6t
Xbit_r12_c14 bl[14] br[14] wl[12] vdd gnd cell_6t
Xbit_r13_c14 bl[14] br[14] wl[13] vdd gnd cell_6t
Xbit_r14_c14 bl[14] br[14] wl[14] vdd gnd cell_6t
Xbit_r15_c14 bl[14] br[14] wl[15] vdd gnd cell_6t
Xbit_r16_c14 bl[14] br[14] wl[16] vdd gnd cell_6t
Xbit_r17_c14 bl[14] br[14] wl[17] vdd gnd cell_6t
Xbit_r18_c14 bl[14] br[14] wl[18] vdd gnd cell_6t
Xbit_r19_c14 bl[14] br[14] wl[19] vdd gnd cell_6t
Xbit_r20_c14 bl[14] br[14] wl[20] vdd gnd cell_6t
Xbit_r21_c14 bl[14] br[14] wl[21] vdd gnd cell_6t
Xbit_r22_c14 bl[14] br[14] wl[22] vdd gnd cell_6t
Xbit_r23_c14 bl[14] br[14] wl[23] vdd gnd cell_6t
Xbit_r24_c14 bl[14] br[14] wl[24] vdd gnd cell_6t
Xbit_r25_c14 bl[14] br[14] wl[25] vdd gnd cell_6t
Xbit_r26_c14 bl[14] br[14] wl[26] vdd gnd cell_6t
Xbit_r27_c14 bl[14] br[14] wl[27] vdd gnd cell_6t
Xbit_r28_c14 bl[14] br[14] wl[28] vdd gnd cell_6t
Xbit_r29_c14 bl[14] br[14] wl[29] vdd gnd cell_6t
Xbit_r30_c14 bl[14] br[14] wl[30] vdd gnd cell_6t
Xbit_r31_c14 bl[14] br[14] wl[31] vdd gnd cell_6t
Xbit_r32_c14 bl[14] br[14] wl[32] vdd gnd cell_6t
Xbit_r33_c14 bl[14] br[14] wl[33] vdd gnd cell_6t
Xbit_r34_c14 bl[14] br[14] wl[34] vdd gnd cell_6t
Xbit_r35_c14 bl[14] br[14] wl[35] vdd gnd cell_6t
Xbit_r36_c14 bl[14] br[14] wl[36] vdd gnd cell_6t
Xbit_r37_c14 bl[14] br[14] wl[37] vdd gnd cell_6t
Xbit_r38_c14 bl[14] br[14] wl[38] vdd gnd cell_6t
Xbit_r39_c14 bl[14] br[14] wl[39] vdd gnd cell_6t
Xbit_r40_c14 bl[14] br[14] wl[40] vdd gnd cell_6t
Xbit_r41_c14 bl[14] br[14] wl[41] vdd gnd cell_6t
Xbit_r42_c14 bl[14] br[14] wl[42] vdd gnd cell_6t
Xbit_r43_c14 bl[14] br[14] wl[43] vdd gnd cell_6t
Xbit_r44_c14 bl[14] br[14] wl[44] vdd gnd cell_6t
Xbit_r45_c14 bl[14] br[14] wl[45] vdd gnd cell_6t
Xbit_r46_c14 bl[14] br[14] wl[46] vdd gnd cell_6t
Xbit_r47_c14 bl[14] br[14] wl[47] vdd gnd cell_6t
Xbit_r48_c14 bl[14] br[14] wl[48] vdd gnd cell_6t
Xbit_r49_c14 bl[14] br[14] wl[49] vdd gnd cell_6t
Xbit_r50_c14 bl[14] br[14] wl[50] vdd gnd cell_6t
Xbit_r51_c14 bl[14] br[14] wl[51] vdd gnd cell_6t
Xbit_r52_c14 bl[14] br[14] wl[52] vdd gnd cell_6t
Xbit_r53_c14 bl[14] br[14] wl[53] vdd gnd cell_6t
Xbit_r54_c14 bl[14] br[14] wl[54] vdd gnd cell_6t
Xbit_r55_c14 bl[14] br[14] wl[55] vdd gnd cell_6t
Xbit_r56_c14 bl[14] br[14] wl[56] vdd gnd cell_6t
Xbit_r57_c14 bl[14] br[14] wl[57] vdd gnd cell_6t
Xbit_r58_c14 bl[14] br[14] wl[58] vdd gnd cell_6t
Xbit_r59_c14 bl[14] br[14] wl[59] vdd gnd cell_6t
Xbit_r60_c14 bl[14] br[14] wl[60] vdd gnd cell_6t
Xbit_r61_c14 bl[14] br[14] wl[61] vdd gnd cell_6t
Xbit_r62_c14 bl[14] br[14] wl[62] vdd gnd cell_6t
Xbit_r63_c14 bl[14] br[14] wl[63] vdd gnd cell_6t
Xbit_r64_c14 bl[14] br[14] wl[64] vdd gnd cell_6t
Xbit_r65_c14 bl[14] br[14] wl[65] vdd gnd cell_6t
Xbit_r66_c14 bl[14] br[14] wl[66] vdd gnd cell_6t
Xbit_r67_c14 bl[14] br[14] wl[67] vdd gnd cell_6t
Xbit_r68_c14 bl[14] br[14] wl[68] vdd gnd cell_6t
Xbit_r69_c14 bl[14] br[14] wl[69] vdd gnd cell_6t
Xbit_r70_c14 bl[14] br[14] wl[70] vdd gnd cell_6t
Xbit_r71_c14 bl[14] br[14] wl[71] vdd gnd cell_6t
Xbit_r72_c14 bl[14] br[14] wl[72] vdd gnd cell_6t
Xbit_r73_c14 bl[14] br[14] wl[73] vdd gnd cell_6t
Xbit_r74_c14 bl[14] br[14] wl[74] vdd gnd cell_6t
Xbit_r75_c14 bl[14] br[14] wl[75] vdd gnd cell_6t
Xbit_r76_c14 bl[14] br[14] wl[76] vdd gnd cell_6t
Xbit_r77_c14 bl[14] br[14] wl[77] vdd gnd cell_6t
Xbit_r78_c14 bl[14] br[14] wl[78] vdd gnd cell_6t
Xbit_r79_c14 bl[14] br[14] wl[79] vdd gnd cell_6t
Xbit_r80_c14 bl[14] br[14] wl[80] vdd gnd cell_6t
Xbit_r81_c14 bl[14] br[14] wl[81] vdd gnd cell_6t
Xbit_r82_c14 bl[14] br[14] wl[82] vdd gnd cell_6t
Xbit_r83_c14 bl[14] br[14] wl[83] vdd gnd cell_6t
Xbit_r84_c14 bl[14] br[14] wl[84] vdd gnd cell_6t
Xbit_r85_c14 bl[14] br[14] wl[85] vdd gnd cell_6t
Xbit_r86_c14 bl[14] br[14] wl[86] vdd gnd cell_6t
Xbit_r87_c14 bl[14] br[14] wl[87] vdd gnd cell_6t
Xbit_r88_c14 bl[14] br[14] wl[88] vdd gnd cell_6t
Xbit_r89_c14 bl[14] br[14] wl[89] vdd gnd cell_6t
Xbit_r90_c14 bl[14] br[14] wl[90] vdd gnd cell_6t
Xbit_r91_c14 bl[14] br[14] wl[91] vdd gnd cell_6t
Xbit_r92_c14 bl[14] br[14] wl[92] vdd gnd cell_6t
Xbit_r93_c14 bl[14] br[14] wl[93] vdd gnd cell_6t
Xbit_r94_c14 bl[14] br[14] wl[94] vdd gnd cell_6t
Xbit_r95_c14 bl[14] br[14] wl[95] vdd gnd cell_6t
Xbit_r96_c14 bl[14] br[14] wl[96] vdd gnd cell_6t
Xbit_r97_c14 bl[14] br[14] wl[97] vdd gnd cell_6t
Xbit_r98_c14 bl[14] br[14] wl[98] vdd gnd cell_6t
Xbit_r99_c14 bl[14] br[14] wl[99] vdd gnd cell_6t
Xbit_r100_c14 bl[14] br[14] wl[100] vdd gnd cell_6t
Xbit_r101_c14 bl[14] br[14] wl[101] vdd gnd cell_6t
Xbit_r102_c14 bl[14] br[14] wl[102] vdd gnd cell_6t
Xbit_r103_c14 bl[14] br[14] wl[103] vdd gnd cell_6t
Xbit_r104_c14 bl[14] br[14] wl[104] vdd gnd cell_6t
Xbit_r105_c14 bl[14] br[14] wl[105] vdd gnd cell_6t
Xbit_r106_c14 bl[14] br[14] wl[106] vdd gnd cell_6t
Xbit_r107_c14 bl[14] br[14] wl[107] vdd gnd cell_6t
Xbit_r108_c14 bl[14] br[14] wl[108] vdd gnd cell_6t
Xbit_r109_c14 bl[14] br[14] wl[109] vdd gnd cell_6t
Xbit_r110_c14 bl[14] br[14] wl[110] vdd gnd cell_6t
Xbit_r111_c14 bl[14] br[14] wl[111] vdd gnd cell_6t
Xbit_r112_c14 bl[14] br[14] wl[112] vdd gnd cell_6t
Xbit_r113_c14 bl[14] br[14] wl[113] vdd gnd cell_6t
Xbit_r114_c14 bl[14] br[14] wl[114] vdd gnd cell_6t
Xbit_r115_c14 bl[14] br[14] wl[115] vdd gnd cell_6t
Xbit_r116_c14 bl[14] br[14] wl[116] vdd gnd cell_6t
Xbit_r117_c14 bl[14] br[14] wl[117] vdd gnd cell_6t
Xbit_r118_c14 bl[14] br[14] wl[118] vdd gnd cell_6t
Xbit_r119_c14 bl[14] br[14] wl[119] vdd gnd cell_6t
Xbit_r120_c14 bl[14] br[14] wl[120] vdd gnd cell_6t
Xbit_r121_c14 bl[14] br[14] wl[121] vdd gnd cell_6t
Xbit_r122_c14 bl[14] br[14] wl[122] vdd gnd cell_6t
Xbit_r123_c14 bl[14] br[14] wl[123] vdd gnd cell_6t
Xbit_r124_c14 bl[14] br[14] wl[124] vdd gnd cell_6t
Xbit_r125_c14 bl[14] br[14] wl[125] vdd gnd cell_6t
Xbit_r126_c14 bl[14] br[14] wl[126] vdd gnd cell_6t
Xbit_r127_c14 bl[14] br[14] wl[127] vdd gnd cell_6t
Xbit_r128_c14 bl[14] br[14] wl[128] vdd gnd cell_6t
Xbit_r129_c14 bl[14] br[14] wl[129] vdd gnd cell_6t
Xbit_r130_c14 bl[14] br[14] wl[130] vdd gnd cell_6t
Xbit_r131_c14 bl[14] br[14] wl[131] vdd gnd cell_6t
Xbit_r132_c14 bl[14] br[14] wl[132] vdd gnd cell_6t
Xbit_r133_c14 bl[14] br[14] wl[133] vdd gnd cell_6t
Xbit_r134_c14 bl[14] br[14] wl[134] vdd gnd cell_6t
Xbit_r135_c14 bl[14] br[14] wl[135] vdd gnd cell_6t
Xbit_r136_c14 bl[14] br[14] wl[136] vdd gnd cell_6t
Xbit_r137_c14 bl[14] br[14] wl[137] vdd gnd cell_6t
Xbit_r138_c14 bl[14] br[14] wl[138] vdd gnd cell_6t
Xbit_r139_c14 bl[14] br[14] wl[139] vdd gnd cell_6t
Xbit_r140_c14 bl[14] br[14] wl[140] vdd gnd cell_6t
Xbit_r141_c14 bl[14] br[14] wl[141] vdd gnd cell_6t
Xbit_r142_c14 bl[14] br[14] wl[142] vdd gnd cell_6t
Xbit_r143_c14 bl[14] br[14] wl[143] vdd gnd cell_6t
Xbit_r144_c14 bl[14] br[14] wl[144] vdd gnd cell_6t
Xbit_r145_c14 bl[14] br[14] wl[145] vdd gnd cell_6t
Xbit_r146_c14 bl[14] br[14] wl[146] vdd gnd cell_6t
Xbit_r147_c14 bl[14] br[14] wl[147] vdd gnd cell_6t
Xbit_r148_c14 bl[14] br[14] wl[148] vdd gnd cell_6t
Xbit_r149_c14 bl[14] br[14] wl[149] vdd gnd cell_6t
Xbit_r150_c14 bl[14] br[14] wl[150] vdd gnd cell_6t
Xbit_r151_c14 bl[14] br[14] wl[151] vdd gnd cell_6t
Xbit_r152_c14 bl[14] br[14] wl[152] vdd gnd cell_6t
Xbit_r153_c14 bl[14] br[14] wl[153] vdd gnd cell_6t
Xbit_r154_c14 bl[14] br[14] wl[154] vdd gnd cell_6t
Xbit_r155_c14 bl[14] br[14] wl[155] vdd gnd cell_6t
Xbit_r156_c14 bl[14] br[14] wl[156] vdd gnd cell_6t
Xbit_r157_c14 bl[14] br[14] wl[157] vdd gnd cell_6t
Xbit_r158_c14 bl[14] br[14] wl[158] vdd gnd cell_6t
Xbit_r159_c14 bl[14] br[14] wl[159] vdd gnd cell_6t
Xbit_r160_c14 bl[14] br[14] wl[160] vdd gnd cell_6t
Xbit_r161_c14 bl[14] br[14] wl[161] vdd gnd cell_6t
Xbit_r162_c14 bl[14] br[14] wl[162] vdd gnd cell_6t
Xbit_r163_c14 bl[14] br[14] wl[163] vdd gnd cell_6t
Xbit_r164_c14 bl[14] br[14] wl[164] vdd gnd cell_6t
Xbit_r165_c14 bl[14] br[14] wl[165] vdd gnd cell_6t
Xbit_r166_c14 bl[14] br[14] wl[166] vdd gnd cell_6t
Xbit_r167_c14 bl[14] br[14] wl[167] vdd gnd cell_6t
Xbit_r168_c14 bl[14] br[14] wl[168] vdd gnd cell_6t
Xbit_r169_c14 bl[14] br[14] wl[169] vdd gnd cell_6t
Xbit_r170_c14 bl[14] br[14] wl[170] vdd gnd cell_6t
Xbit_r171_c14 bl[14] br[14] wl[171] vdd gnd cell_6t
Xbit_r172_c14 bl[14] br[14] wl[172] vdd gnd cell_6t
Xbit_r173_c14 bl[14] br[14] wl[173] vdd gnd cell_6t
Xbit_r174_c14 bl[14] br[14] wl[174] vdd gnd cell_6t
Xbit_r175_c14 bl[14] br[14] wl[175] vdd gnd cell_6t
Xbit_r176_c14 bl[14] br[14] wl[176] vdd gnd cell_6t
Xbit_r177_c14 bl[14] br[14] wl[177] vdd gnd cell_6t
Xbit_r178_c14 bl[14] br[14] wl[178] vdd gnd cell_6t
Xbit_r179_c14 bl[14] br[14] wl[179] vdd gnd cell_6t
Xbit_r180_c14 bl[14] br[14] wl[180] vdd gnd cell_6t
Xbit_r181_c14 bl[14] br[14] wl[181] vdd gnd cell_6t
Xbit_r182_c14 bl[14] br[14] wl[182] vdd gnd cell_6t
Xbit_r183_c14 bl[14] br[14] wl[183] vdd gnd cell_6t
Xbit_r184_c14 bl[14] br[14] wl[184] vdd gnd cell_6t
Xbit_r185_c14 bl[14] br[14] wl[185] vdd gnd cell_6t
Xbit_r186_c14 bl[14] br[14] wl[186] vdd gnd cell_6t
Xbit_r187_c14 bl[14] br[14] wl[187] vdd gnd cell_6t
Xbit_r188_c14 bl[14] br[14] wl[188] vdd gnd cell_6t
Xbit_r189_c14 bl[14] br[14] wl[189] vdd gnd cell_6t
Xbit_r190_c14 bl[14] br[14] wl[190] vdd gnd cell_6t
Xbit_r191_c14 bl[14] br[14] wl[191] vdd gnd cell_6t
Xbit_r192_c14 bl[14] br[14] wl[192] vdd gnd cell_6t
Xbit_r193_c14 bl[14] br[14] wl[193] vdd gnd cell_6t
Xbit_r194_c14 bl[14] br[14] wl[194] vdd gnd cell_6t
Xbit_r195_c14 bl[14] br[14] wl[195] vdd gnd cell_6t
Xbit_r196_c14 bl[14] br[14] wl[196] vdd gnd cell_6t
Xbit_r197_c14 bl[14] br[14] wl[197] vdd gnd cell_6t
Xbit_r198_c14 bl[14] br[14] wl[198] vdd gnd cell_6t
Xbit_r199_c14 bl[14] br[14] wl[199] vdd gnd cell_6t
Xbit_r200_c14 bl[14] br[14] wl[200] vdd gnd cell_6t
Xbit_r201_c14 bl[14] br[14] wl[201] vdd gnd cell_6t
Xbit_r202_c14 bl[14] br[14] wl[202] vdd gnd cell_6t
Xbit_r203_c14 bl[14] br[14] wl[203] vdd gnd cell_6t
Xbit_r204_c14 bl[14] br[14] wl[204] vdd gnd cell_6t
Xbit_r205_c14 bl[14] br[14] wl[205] vdd gnd cell_6t
Xbit_r206_c14 bl[14] br[14] wl[206] vdd gnd cell_6t
Xbit_r207_c14 bl[14] br[14] wl[207] vdd gnd cell_6t
Xbit_r208_c14 bl[14] br[14] wl[208] vdd gnd cell_6t
Xbit_r209_c14 bl[14] br[14] wl[209] vdd gnd cell_6t
Xbit_r210_c14 bl[14] br[14] wl[210] vdd gnd cell_6t
Xbit_r211_c14 bl[14] br[14] wl[211] vdd gnd cell_6t
Xbit_r212_c14 bl[14] br[14] wl[212] vdd gnd cell_6t
Xbit_r213_c14 bl[14] br[14] wl[213] vdd gnd cell_6t
Xbit_r214_c14 bl[14] br[14] wl[214] vdd gnd cell_6t
Xbit_r215_c14 bl[14] br[14] wl[215] vdd gnd cell_6t
Xbit_r216_c14 bl[14] br[14] wl[216] vdd gnd cell_6t
Xbit_r217_c14 bl[14] br[14] wl[217] vdd gnd cell_6t
Xbit_r218_c14 bl[14] br[14] wl[218] vdd gnd cell_6t
Xbit_r219_c14 bl[14] br[14] wl[219] vdd gnd cell_6t
Xbit_r220_c14 bl[14] br[14] wl[220] vdd gnd cell_6t
Xbit_r221_c14 bl[14] br[14] wl[221] vdd gnd cell_6t
Xbit_r222_c14 bl[14] br[14] wl[222] vdd gnd cell_6t
Xbit_r223_c14 bl[14] br[14] wl[223] vdd gnd cell_6t
Xbit_r224_c14 bl[14] br[14] wl[224] vdd gnd cell_6t
Xbit_r225_c14 bl[14] br[14] wl[225] vdd gnd cell_6t
Xbit_r226_c14 bl[14] br[14] wl[226] vdd gnd cell_6t
Xbit_r227_c14 bl[14] br[14] wl[227] vdd gnd cell_6t
Xbit_r228_c14 bl[14] br[14] wl[228] vdd gnd cell_6t
Xbit_r229_c14 bl[14] br[14] wl[229] vdd gnd cell_6t
Xbit_r230_c14 bl[14] br[14] wl[230] vdd gnd cell_6t
Xbit_r231_c14 bl[14] br[14] wl[231] vdd gnd cell_6t
Xbit_r232_c14 bl[14] br[14] wl[232] vdd gnd cell_6t
Xbit_r233_c14 bl[14] br[14] wl[233] vdd gnd cell_6t
Xbit_r234_c14 bl[14] br[14] wl[234] vdd gnd cell_6t
Xbit_r235_c14 bl[14] br[14] wl[235] vdd gnd cell_6t
Xbit_r236_c14 bl[14] br[14] wl[236] vdd gnd cell_6t
Xbit_r237_c14 bl[14] br[14] wl[237] vdd gnd cell_6t
Xbit_r238_c14 bl[14] br[14] wl[238] vdd gnd cell_6t
Xbit_r239_c14 bl[14] br[14] wl[239] vdd gnd cell_6t
Xbit_r240_c14 bl[14] br[14] wl[240] vdd gnd cell_6t
Xbit_r241_c14 bl[14] br[14] wl[241] vdd gnd cell_6t
Xbit_r242_c14 bl[14] br[14] wl[242] vdd gnd cell_6t
Xbit_r243_c14 bl[14] br[14] wl[243] vdd gnd cell_6t
Xbit_r244_c14 bl[14] br[14] wl[244] vdd gnd cell_6t
Xbit_r245_c14 bl[14] br[14] wl[245] vdd gnd cell_6t
Xbit_r246_c14 bl[14] br[14] wl[246] vdd gnd cell_6t
Xbit_r247_c14 bl[14] br[14] wl[247] vdd gnd cell_6t
Xbit_r248_c14 bl[14] br[14] wl[248] vdd gnd cell_6t
Xbit_r249_c14 bl[14] br[14] wl[249] vdd gnd cell_6t
Xbit_r250_c14 bl[14] br[14] wl[250] vdd gnd cell_6t
Xbit_r251_c14 bl[14] br[14] wl[251] vdd gnd cell_6t
Xbit_r252_c14 bl[14] br[14] wl[252] vdd gnd cell_6t
Xbit_r253_c14 bl[14] br[14] wl[253] vdd gnd cell_6t
Xbit_r254_c14 bl[14] br[14] wl[254] vdd gnd cell_6t
Xbit_r255_c14 bl[14] br[14] wl[255] vdd gnd cell_6t
Xbit_r0_c15 bl[15] br[15] wl[0] vdd gnd cell_6t
Xbit_r1_c15 bl[15] br[15] wl[1] vdd gnd cell_6t
Xbit_r2_c15 bl[15] br[15] wl[2] vdd gnd cell_6t
Xbit_r3_c15 bl[15] br[15] wl[3] vdd gnd cell_6t
Xbit_r4_c15 bl[15] br[15] wl[4] vdd gnd cell_6t
Xbit_r5_c15 bl[15] br[15] wl[5] vdd gnd cell_6t
Xbit_r6_c15 bl[15] br[15] wl[6] vdd gnd cell_6t
Xbit_r7_c15 bl[15] br[15] wl[7] vdd gnd cell_6t
Xbit_r8_c15 bl[15] br[15] wl[8] vdd gnd cell_6t
Xbit_r9_c15 bl[15] br[15] wl[9] vdd gnd cell_6t
Xbit_r10_c15 bl[15] br[15] wl[10] vdd gnd cell_6t
Xbit_r11_c15 bl[15] br[15] wl[11] vdd gnd cell_6t
Xbit_r12_c15 bl[15] br[15] wl[12] vdd gnd cell_6t
Xbit_r13_c15 bl[15] br[15] wl[13] vdd gnd cell_6t
Xbit_r14_c15 bl[15] br[15] wl[14] vdd gnd cell_6t
Xbit_r15_c15 bl[15] br[15] wl[15] vdd gnd cell_6t
Xbit_r16_c15 bl[15] br[15] wl[16] vdd gnd cell_6t
Xbit_r17_c15 bl[15] br[15] wl[17] vdd gnd cell_6t
Xbit_r18_c15 bl[15] br[15] wl[18] vdd gnd cell_6t
Xbit_r19_c15 bl[15] br[15] wl[19] vdd gnd cell_6t
Xbit_r20_c15 bl[15] br[15] wl[20] vdd gnd cell_6t
Xbit_r21_c15 bl[15] br[15] wl[21] vdd gnd cell_6t
Xbit_r22_c15 bl[15] br[15] wl[22] vdd gnd cell_6t
Xbit_r23_c15 bl[15] br[15] wl[23] vdd gnd cell_6t
Xbit_r24_c15 bl[15] br[15] wl[24] vdd gnd cell_6t
Xbit_r25_c15 bl[15] br[15] wl[25] vdd gnd cell_6t
Xbit_r26_c15 bl[15] br[15] wl[26] vdd gnd cell_6t
Xbit_r27_c15 bl[15] br[15] wl[27] vdd gnd cell_6t
Xbit_r28_c15 bl[15] br[15] wl[28] vdd gnd cell_6t
Xbit_r29_c15 bl[15] br[15] wl[29] vdd gnd cell_6t
Xbit_r30_c15 bl[15] br[15] wl[30] vdd gnd cell_6t
Xbit_r31_c15 bl[15] br[15] wl[31] vdd gnd cell_6t
Xbit_r32_c15 bl[15] br[15] wl[32] vdd gnd cell_6t
Xbit_r33_c15 bl[15] br[15] wl[33] vdd gnd cell_6t
Xbit_r34_c15 bl[15] br[15] wl[34] vdd gnd cell_6t
Xbit_r35_c15 bl[15] br[15] wl[35] vdd gnd cell_6t
Xbit_r36_c15 bl[15] br[15] wl[36] vdd gnd cell_6t
Xbit_r37_c15 bl[15] br[15] wl[37] vdd gnd cell_6t
Xbit_r38_c15 bl[15] br[15] wl[38] vdd gnd cell_6t
Xbit_r39_c15 bl[15] br[15] wl[39] vdd gnd cell_6t
Xbit_r40_c15 bl[15] br[15] wl[40] vdd gnd cell_6t
Xbit_r41_c15 bl[15] br[15] wl[41] vdd gnd cell_6t
Xbit_r42_c15 bl[15] br[15] wl[42] vdd gnd cell_6t
Xbit_r43_c15 bl[15] br[15] wl[43] vdd gnd cell_6t
Xbit_r44_c15 bl[15] br[15] wl[44] vdd gnd cell_6t
Xbit_r45_c15 bl[15] br[15] wl[45] vdd gnd cell_6t
Xbit_r46_c15 bl[15] br[15] wl[46] vdd gnd cell_6t
Xbit_r47_c15 bl[15] br[15] wl[47] vdd gnd cell_6t
Xbit_r48_c15 bl[15] br[15] wl[48] vdd gnd cell_6t
Xbit_r49_c15 bl[15] br[15] wl[49] vdd gnd cell_6t
Xbit_r50_c15 bl[15] br[15] wl[50] vdd gnd cell_6t
Xbit_r51_c15 bl[15] br[15] wl[51] vdd gnd cell_6t
Xbit_r52_c15 bl[15] br[15] wl[52] vdd gnd cell_6t
Xbit_r53_c15 bl[15] br[15] wl[53] vdd gnd cell_6t
Xbit_r54_c15 bl[15] br[15] wl[54] vdd gnd cell_6t
Xbit_r55_c15 bl[15] br[15] wl[55] vdd gnd cell_6t
Xbit_r56_c15 bl[15] br[15] wl[56] vdd gnd cell_6t
Xbit_r57_c15 bl[15] br[15] wl[57] vdd gnd cell_6t
Xbit_r58_c15 bl[15] br[15] wl[58] vdd gnd cell_6t
Xbit_r59_c15 bl[15] br[15] wl[59] vdd gnd cell_6t
Xbit_r60_c15 bl[15] br[15] wl[60] vdd gnd cell_6t
Xbit_r61_c15 bl[15] br[15] wl[61] vdd gnd cell_6t
Xbit_r62_c15 bl[15] br[15] wl[62] vdd gnd cell_6t
Xbit_r63_c15 bl[15] br[15] wl[63] vdd gnd cell_6t
Xbit_r64_c15 bl[15] br[15] wl[64] vdd gnd cell_6t
Xbit_r65_c15 bl[15] br[15] wl[65] vdd gnd cell_6t
Xbit_r66_c15 bl[15] br[15] wl[66] vdd gnd cell_6t
Xbit_r67_c15 bl[15] br[15] wl[67] vdd gnd cell_6t
Xbit_r68_c15 bl[15] br[15] wl[68] vdd gnd cell_6t
Xbit_r69_c15 bl[15] br[15] wl[69] vdd gnd cell_6t
Xbit_r70_c15 bl[15] br[15] wl[70] vdd gnd cell_6t
Xbit_r71_c15 bl[15] br[15] wl[71] vdd gnd cell_6t
Xbit_r72_c15 bl[15] br[15] wl[72] vdd gnd cell_6t
Xbit_r73_c15 bl[15] br[15] wl[73] vdd gnd cell_6t
Xbit_r74_c15 bl[15] br[15] wl[74] vdd gnd cell_6t
Xbit_r75_c15 bl[15] br[15] wl[75] vdd gnd cell_6t
Xbit_r76_c15 bl[15] br[15] wl[76] vdd gnd cell_6t
Xbit_r77_c15 bl[15] br[15] wl[77] vdd gnd cell_6t
Xbit_r78_c15 bl[15] br[15] wl[78] vdd gnd cell_6t
Xbit_r79_c15 bl[15] br[15] wl[79] vdd gnd cell_6t
Xbit_r80_c15 bl[15] br[15] wl[80] vdd gnd cell_6t
Xbit_r81_c15 bl[15] br[15] wl[81] vdd gnd cell_6t
Xbit_r82_c15 bl[15] br[15] wl[82] vdd gnd cell_6t
Xbit_r83_c15 bl[15] br[15] wl[83] vdd gnd cell_6t
Xbit_r84_c15 bl[15] br[15] wl[84] vdd gnd cell_6t
Xbit_r85_c15 bl[15] br[15] wl[85] vdd gnd cell_6t
Xbit_r86_c15 bl[15] br[15] wl[86] vdd gnd cell_6t
Xbit_r87_c15 bl[15] br[15] wl[87] vdd gnd cell_6t
Xbit_r88_c15 bl[15] br[15] wl[88] vdd gnd cell_6t
Xbit_r89_c15 bl[15] br[15] wl[89] vdd gnd cell_6t
Xbit_r90_c15 bl[15] br[15] wl[90] vdd gnd cell_6t
Xbit_r91_c15 bl[15] br[15] wl[91] vdd gnd cell_6t
Xbit_r92_c15 bl[15] br[15] wl[92] vdd gnd cell_6t
Xbit_r93_c15 bl[15] br[15] wl[93] vdd gnd cell_6t
Xbit_r94_c15 bl[15] br[15] wl[94] vdd gnd cell_6t
Xbit_r95_c15 bl[15] br[15] wl[95] vdd gnd cell_6t
Xbit_r96_c15 bl[15] br[15] wl[96] vdd gnd cell_6t
Xbit_r97_c15 bl[15] br[15] wl[97] vdd gnd cell_6t
Xbit_r98_c15 bl[15] br[15] wl[98] vdd gnd cell_6t
Xbit_r99_c15 bl[15] br[15] wl[99] vdd gnd cell_6t
Xbit_r100_c15 bl[15] br[15] wl[100] vdd gnd cell_6t
Xbit_r101_c15 bl[15] br[15] wl[101] vdd gnd cell_6t
Xbit_r102_c15 bl[15] br[15] wl[102] vdd gnd cell_6t
Xbit_r103_c15 bl[15] br[15] wl[103] vdd gnd cell_6t
Xbit_r104_c15 bl[15] br[15] wl[104] vdd gnd cell_6t
Xbit_r105_c15 bl[15] br[15] wl[105] vdd gnd cell_6t
Xbit_r106_c15 bl[15] br[15] wl[106] vdd gnd cell_6t
Xbit_r107_c15 bl[15] br[15] wl[107] vdd gnd cell_6t
Xbit_r108_c15 bl[15] br[15] wl[108] vdd gnd cell_6t
Xbit_r109_c15 bl[15] br[15] wl[109] vdd gnd cell_6t
Xbit_r110_c15 bl[15] br[15] wl[110] vdd gnd cell_6t
Xbit_r111_c15 bl[15] br[15] wl[111] vdd gnd cell_6t
Xbit_r112_c15 bl[15] br[15] wl[112] vdd gnd cell_6t
Xbit_r113_c15 bl[15] br[15] wl[113] vdd gnd cell_6t
Xbit_r114_c15 bl[15] br[15] wl[114] vdd gnd cell_6t
Xbit_r115_c15 bl[15] br[15] wl[115] vdd gnd cell_6t
Xbit_r116_c15 bl[15] br[15] wl[116] vdd gnd cell_6t
Xbit_r117_c15 bl[15] br[15] wl[117] vdd gnd cell_6t
Xbit_r118_c15 bl[15] br[15] wl[118] vdd gnd cell_6t
Xbit_r119_c15 bl[15] br[15] wl[119] vdd gnd cell_6t
Xbit_r120_c15 bl[15] br[15] wl[120] vdd gnd cell_6t
Xbit_r121_c15 bl[15] br[15] wl[121] vdd gnd cell_6t
Xbit_r122_c15 bl[15] br[15] wl[122] vdd gnd cell_6t
Xbit_r123_c15 bl[15] br[15] wl[123] vdd gnd cell_6t
Xbit_r124_c15 bl[15] br[15] wl[124] vdd gnd cell_6t
Xbit_r125_c15 bl[15] br[15] wl[125] vdd gnd cell_6t
Xbit_r126_c15 bl[15] br[15] wl[126] vdd gnd cell_6t
Xbit_r127_c15 bl[15] br[15] wl[127] vdd gnd cell_6t
Xbit_r128_c15 bl[15] br[15] wl[128] vdd gnd cell_6t
Xbit_r129_c15 bl[15] br[15] wl[129] vdd gnd cell_6t
Xbit_r130_c15 bl[15] br[15] wl[130] vdd gnd cell_6t
Xbit_r131_c15 bl[15] br[15] wl[131] vdd gnd cell_6t
Xbit_r132_c15 bl[15] br[15] wl[132] vdd gnd cell_6t
Xbit_r133_c15 bl[15] br[15] wl[133] vdd gnd cell_6t
Xbit_r134_c15 bl[15] br[15] wl[134] vdd gnd cell_6t
Xbit_r135_c15 bl[15] br[15] wl[135] vdd gnd cell_6t
Xbit_r136_c15 bl[15] br[15] wl[136] vdd gnd cell_6t
Xbit_r137_c15 bl[15] br[15] wl[137] vdd gnd cell_6t
Xbit_r138_c15 bl[15] br[15] wl[138] vdd gnd cell_6t
Xbit_r139_c15 bl[15] br[15] wl[139] vdd gnd cell_6t
Xbit_r140_c15 bl[15] br[15] wl[140] vdd gnd cell_6t
Xbit_r141_c15 bl[15] br[15] wl[141] vdd gnd cell_6t
Xbit_r142_c15 bl[15] br[15] wl[142] vdd gnd cell_6t
Xbit_r143_c15 bl[15] br[15] wl[143] vdd gnd cell_6t
Xbit_r144_c15 bl[15] br[15] wl[144] vdd gnd cell_6t
Xbit_r145_c15 bl[15] br[15] wl[145] vdd gnd cell_6t
Xbit_r146_c15 bl[15] br[15] wl[146] vdd gnd cell_6t
Xbit_r147_c15 bl[15] br[15] wl[147] vdd gnd cell_6t
Xbit_r148_c15 bl[15] br[15] wl[148] vdd gnd cell_6t
Xbit_r149_c15 bl[15] br[15] wl[149] vdd gnd cell_6t
Xbit_r150_c15 bl[15] br[15] wl[150] vdd gnd cell_6t
Xbit_r151_c15 bl[15] br[15] wl[151] vdd gnd cell_6t
Xbit_r152_c15 bl[15] br[15] wl[152] vdd gnd cell_6t
Xbit_r153_c15 bl[15] br[15] wl[153] vdd gnd cell_6t
Xbit_r154_c15 bl[15] br[15] wl[154] vdd gnd cell_6t
Xbit_r155_c15 bl[15] br[15] wl[155] vdd gnd cell_6t
Xbit_r156_c15 bl[15] br[15] wl[156] vdd gnd cell_6t
Xbit_r157_c15 bl[15] br[15] wl[157] vdd gnd cell_6t
Xbit_r158_c15 bl[15] br[15] wl[158] vdd gnd cell_6t
Xbit_r159_c15 bl[15] br[15] wl[159] vdd gnd cell_6t
Xbit_r160_c15 bl[15] br[15] wl[160] vdd gnd cell_6t
Xbit_r161_c15 bl[15] br[15] wl[161] vdd gnd cell_6t
Xbit_r162_c15 bl[15] br[15] wl[162] vdd gnd cell_6t
Xbit_r163_c15 bl[15] br[15] wl[163] vdd gnd cell_6t
Xbit_r164_c15 bl[15] br[15] wl[164] vdd gnd cell_6t
Xbit_r165_c15 bl[15] br[15] wl[165] vdd gnd cell_6t
Xbit_r166_c15 bl[15] br[15] wl[166] vdd gnd cell_6t
Xbit_r167_c15 bl[15] br[15] wl[167] vdd gnd cell_6t
Xbit_r168_c15 bl[15] br[15] wl[168] vdd gnd cell_6t
Xbit_r169_c15 bl[15] br[15] wl[169] vdd gnd cell_6t
Xbit_r170_c15 bl[15] br[15] wl[170] vdd gnd cell_6t
Xbit_r171_c15 bl[15] br[15] wl[171] vdd gnd cell_6t
Xbit_r172_c15 bl[15] br[15] wl[172] vdd gnd cell_6t
Xbit_r173_c15 bl[15] br[15] wl[173] vdd gnd cell_6t
Xbit_r174_c15 bl[15] br[15] wl[174] vdd gnd cell_6t
Xbit_r175_c15 bl[15] br[15] wl[175] vdd gnd cell_6t
Xbit_r176_c15 bl[15] br[15] wl[176] vdd gnd cell_6t
Xbit_r177_c15 bl[15] br[15] wl[177] vdd gnd cell_6t
Xbit_r178_c15 bl[15] br[15] wl[178] vdd gnd cell_6t
Xbit_r179_c15 bl[15] br[15] wl[179] vdd gnd cell_6t
Xbit_r180_c15 bl[15] br[15] wl[180] vdd gnd cell_6t
Xbit_r181_c15 bl[15] br[15] wl[181] vdd gnd cell_6t
Xbit_r182_c15 bl[15] br[15] wl[182] vdd gnd cell_6t
Xbit_r183_c15 bl[15] br[15] wl[183] vdd gnd cell_6t
Xbit_r184_c15 bl[15] br[15] wl[184] vdd gnd cell_6t
Xbit_r185_c15 bl[15] br[15] wl[185] vdd gnd cell_6t
Xbit_r186_c15 bl[15] br[15] wl[186] vdd gnd cell_6t
Xbit_r187_c15 bl[15] br[15] wl[187] vdd gnd cell_6t
Xbit_r188_c15 bl[15] br[15] wl[188] vdd gnd cell_6t
Xbit_r189_c15 bl[15] br[15] wl[189] vdd gnd cell_6t
Xbit_r190_c15 bl[15] br[15] wl[190] vdd gnd cell_6t
Xbit_r191_c15 bl[15] br[15] wl[191] vdd gnd cell_6t
Xbit_r192_c15 bl[15] br[15] wl[192] vdd gnd cell_6t
Xbit_r193_c15 bl[15] br[15] wl[193] vdd gnd cell_6t
Xbit_r194_c15 bl[15] br[15] wl[194] vdd gnd cell_6t
Xbit_r195_c15 bl[15] br[15] wl[195] vdd gnd cell_6t
Xbit_r196_c15 bl[15] br[15] wl[196] vdd gnd cell_6t
Xbit_r197_c15 bl[15] br[15] wl[197] vdd gnd cell_6t
Xbit_r198_c15 bl[15] br[15] wl[198] vdd gnd cell_6t
Xbit_r199_c15 bl[15] br[15] wl[199] vdd gnd cell_6t
Xbit_r200_c15 bl[15] br[15] wl[200] vdd gnd cell_6t
Xbit_r201_c15 bl[15] br[15] wl[201] vdd gnd cell_6t
Xbit_r202_c15 bl[15] br[15] wl[202] vdd gnd cell_6t
Xbit_r203_c15 bl[15] br[15] wl[203] vdd gnd cell_6t
Xbit_r204_c15 bl[15] br[15] wl[204] vdd gnd cell_6t
Xbit_r205_c15 bl[15] br[15] wl[205] vdd gnd cell_6t
Xbit_r206_c15 bl[15] br[15] wl[206] vdd gnd cell_6t
Xbit_r207_c15 bl[15] br[15] wl[207] vdd gnd cell_6t
Xbit_r208_c15 bl[15] br[15] wl[208] vdd gnd cell_6t
Xbit_r209_c15 bl[15] br[15] wl[209] vdd gnd cell_6t
Xbit_r210_c15 bl[15] br[15] wl[210] vdd gnd cell_6t
Xbit_r211_c15 bl[15] br[15] wl[211] vdd gnd cell_6t
Xbit_r212_c15 bl[15] br[15] wl[212] vdd gnd cell_6t
Xbit_r213_c15 bl[15] br[15] wl[213] vdd gnd cell_6t
Xbit_r214_c15 bl[15] br[15] wl[214] vdd gnd cell_6t
Xbit_r215_c15 bl[15] br[15] wl[215] vdd gnd cell_6t
Xbit_r216_c15 bl[15] br[15] wl[216] vdd gnd cell_6t
Xbit_r217_c15 bl[15] br[15] wl[217] vdd gnd cell_6t
Xbit_r218_c15 bl[15] br[15] wl[218] vdd gnd cell_6t
Xbit_r219_c15 bl[15] br[15] wl[219] vdd gnd cell_6t
Xbit_r220_c15 bl[15] br[15] wl[220] vdd gnd cell_6t
Xbit_r221_c15 bl[15] br[15] wl[221] vdd gnd cell_6t
Xbit_r222_c15 bl[15] br[15] wl[222] vdd gnd cell_6t
Xbit_r223_c15 bl[15] br[15] wl[223] vdd gnd cell_6t
Xbit_r224_c15 bl[15] br[15] wl[224] vdd gnd cell_6t
Xbit_r225_c15 bl[15] br[15] wl[225] vdd gnd cell_6t
Xbit_r226_c15 bl[15] br[15] wl[226] vdd gnd cell_6t
Xbit_r227_c15 bl[15] br[15] wl[227] vdd gnd cell_6t
Xbit_r228_c15 bl[15] br[15] wl[228] vdd gnd cell_6t
Xbit_r229_c15 bl[15] br[15] wl[229] vdd gnd cell_6t
Xbit_r230_c15 bl[15] br[15] wl[230] vdd gnd cell_6t
Xbit_r231_c15 bl[15] br[15] wl[231] vdd gnd cell_6t
Xbit_r232_c15 bl[15] br[15] wl[232] vdd gnd cell_6t
Xbit_r233_c15 bl[15] br[15] wl[233] vdd gnd cell_6t
Xbit_r234_c15 bl[15] br[15] wl[234] vdd gnd cell_6t
Xbit_r235_c15 bl[15] br[15] wl[235] vdd gnd cell_6t
Xbit_r236_c15 bl[15] br[15] wl[236] vdd gnd cell_6t
Xbit_r237_c15 bl[15] br[15] wl[237] vdd gnd cell_6t
Xbit_r238_c15 bl[15] br[15] wl[238] vdd gnd cell_6t
Xbit_r239_c15 bl[15] br[15] wl[239] vdd gnd cell_6t
Xbit_r240_c15 bl[15] br[15] wl[240] vdd gnd cell_6t
Xbit_r241_c15 bl[15] br[15] wl[241] vdd gnd cell_6t
Xbit_r242_c15 bl[15] br[15] wl[242] vdd gnd cell_6t
Xbit_r243_c15 bl[15] br[15] wl[243] vdd gnd cell_6t
Xbit_r244_c15 bl[15] br[15] wl[244] vdd gnd cell_6t
Xbit_r245_c15 bl[15] br[15] wl[245] vdd gnd cell_6t
Xbit_r246_c15 bl[15] br[15] wl[246] vdd gnd cell_6t
Xbit_r247_c15 bl[15] br[15] wl[247] vdd gnd cell_6t
Xbit_r248_c15 bl[15] br[15] wl[248] vdd gnd cell_6t
Xbit_r249_c15 bl[15] br[15] wl[249] vdd gnd cell_6t
Xbit_r250_c15 bl[15] br[15] wl[250] vdd gnd cell_6t
Xbit_r251_c15 bl[15] br[15] wl[251] vdd gnd cell_6t
Xbit_r252_c15 bl[15] br[15] wl[252] vdd gnd cell_6t
Xbit_r253_c15 bl[15] br[15] wl[253] vdd gnd cell_6t
Xbit_r254_c15 bl[15] br[15] wl[254] vdd gnd cell_6t
Xbit_r255_c15 bl[15] br[15] wl[255] vdd gnd cell_6t
Xbit_r0_c16 bl[16] br[16] wl[0] vdd gnd cell_6t
Xbit_r1_c16 bl[16] br[16] wl[1] vdd gnd cell_6t
Xbit_r2_c16 bl[16] br[16] wl[2] vdd gnd cell_6t
Xbit_r3_c16 bl[16] br[16] wl[3] vdd gnd cell_6t
Xbit_r4_c16 bl[16] br[16] wl[4] vdd gnd cell_6t
Xbit_r5_c16 bl[16] br[16] wl[5] vdd gnd cell_6t
Xbit_r6_c16 bl[16] br[16] wl[6] vdd gnd cell_6t
Xbit_r7_c16 bl[16] br[16] wl[7] vdd gnd cell_6t
Xbit_r8_c16 bl[16] br[16] wl[8] vdd gnd cell_6t
Xbit_r9_c16 bl[16] br[16] wl[9] vdd gnd cell_6t
Xbit_r10_c16 bl[16] br[16] wl[10] vdd gnd cell_6t
Xbit_r11_c16 bl[16] br[16] wl[11] vdd gnd cell_6t
Xbit_r12_c16 bl[16] br[16] wl[12] vdd gnd cell_6t
Xbit_r13_c16 bl[16] br[16] wl[13] vdd gnd cell_6t
Xbit_r14_c16 bl[16] br[16] wl[14] vdd gnd cell_6t
Xbit_r15_c16 bl[16] br[16] wl[15] vdd gnd cell_6t
Xbit_r16_c16 bl[16] br[16] wl[16] vdd gnd cell_6t
Xbit_r17_c16 bl[16] br[16] wl[17] vdd gnd cell_6t
Xbit_r18_c16 bl[16] br[16] wl[18] vdd gnd cell_6t
Xbit_r19_c16 bl[16] br[16] wl[19] vdd gnd cell_6t
Xbit_r20_c16 bl[16] br[16] wl[20] vdd gnd cell_6t
Xbit_r21_c16 bl[16] br[16] wl[21] vdd gnd cell_6t
Xbit_r22_c16 bl[16] br[16] wl[22] vdd gnd cell_6t
Xbit_r23_c16 bl[16] br[16] wl[23] vdd gnd cell_6t
Xbit_r24_c16 bl[16] br[16] wl[24] vdd gnd cell_6t
Xbit_r25_c16 bl[16] br[16] wl[25] vdd gnd cell_6t
Xbit_r26_c16 bl[16] br[16] wl[26] vdd gnd cell_6t
Xbit_r27_c16 bl[16] br[16] wl[27] vdd gnd cell_6t
Xbit_r28_c16 bl[16] br[16] wl[28] vdd gnd cell_6t
Xbit_r29_c16 bl[16] br[16] wl[29] vdd gnd cell_6t
Xbit_r30_c16 bl[16] br[16] wl[30] vdd gnd cell_6t
Xbit_r31_c16 bl[16] br[16] wl[31] vdd gnd cell_6t
Xbit_r32_c16 bl[16] br[16] wl[32] vdd gnd cell_6t
Xbit_r33_c16 bl[16] br[16] wl[33] vdd gnd cell_6t
Xbit_r34_c16 bl[16] br[16] wl[34] vdd gnd cell_6t
Xbit_r35_c16 bl[16] br[16] wl[35] vdd gnd cell_6t
Xbit_r36_c16 bl[16] br[16] wl[36] vdd gnd cell_6t
Xbit_r37_c16 bl[16] br[16] wl[37] vdd gnd cell_6t
Xbit_r38_c16 bl[16] br[16] wl[38] vdd gnd cell_6t
Xbit_r39_c16 bl[16] br[16] wl[39] vdd gnd cell_6t
Xbit_r40_c16 bl[16] br[16] wl[40] vdd gnd cell_6t
Xbit_r41_c16 bl[16] br[16] wl[41] vdd gnd cell_6t
Xbit_r42_c16 bl[16] br[16] wl[42] vdd gnd cell_6t
Xbit_r43_c16 bl[16] br[16] wl[43] vdd gnd cell_6t
Xbit_r44_c16 bl[16] br[16] wl[44] vdd gnd cell_6t
Xbit_r45_c16 bl[16] br[16] wl[45] vdd gnd cell_6t
Xbit_r46_c16 bl[16] br[16] wl[46] vdd gnd cell_6t
Xbit_r47_c16 bl[16] br[16] wl[47] vdd gnd cell_6t
Xbit_r48_c16 bl[16] br[16] wl[48] vdd gnd cell_6t
Xbit_r49_c16 bl[16] br[16] wl[49] vdd gnd cell_6t
Xbit_r50_c16 bl[16] br[16] wl[50] vdd gnd cell_6t
Xbit_r51_c16 bl[16] br[16] wl[51] vdd gnd cell_6t
Xbit_r52_c16 bl[16] br[16] wl[52] vdd gnd cell_6t
Xbit_r53_c16 bl[16] br[16] wl[53] vdd gnd cell_6t
Xbit_r54_c16 bl[16] br[16] wl[54] vdd gnd cell_6t
Xbit_r55_c16 bl[16] br[16] wl[55] vdd gnd cell_6t
Xbit_r56_c16 bl[16] br[16] wl[56] vdd gnd cell_6t
Xbit_r57_c16 bl[16] br[16] wl[57] vdd gnd cell_6t
Xbit_r58_c16 bl[16] br[16] wl[58] vdd gnd cell_6t
Xbit_r59_c16 bl[16] br[16] wl[59] vdd gnd cell_6t
Xbit_r60_c16 bl[16] br[16] wl[60] vdd gnd cell_6t
Xbit_r61_c16 bl[16] br[16] wl[61] vdd gnd cell_6t
Xbit_r62_c16 bl[16] br[16] wl[62] vdd gnd cell_6t
Xbit_r63_c16 bl[16] br[16] wl[63] vdd gnd cell_6t
Xbit_r64_c16 bl[16] br[16] wl[64] vdd gnd cell_6t
Xbit_r65_c16 bl[16] br[16] wl[65] vdd gnd cell_6t
Xbit_r66_c16 bl[16] br[16] wl[66] vdd gnd cell_6t
Xbit_r67_c16 bl[16] br[16] wl[67] vdd gnd cell_6t
Xbit_r68_c16 bl[16] br[16] wl[68] vdd gnd cell_6t
Xbit_r69_c16 bl[16] br[16] wl[69] vdd gnd cell_6t
Xbit_r70_c16 bl[16] br[16] wl[70] vdd gnd cell_6t
Xbit_r71_c16 bl[16] br[16] wl[71] vdd gnd cell_6t
Xbit_r72_c16 bl[16] br[16] wl[72] vdd gnd cell_6t
Xbit_r73_c16 bl[16] br[16] wl[73] vdd gnd cell_6t
Xbit_r74_c16 bl[16] br[16] wl[74] vdd gnd cell_6t
Xbit_r75_c16 bl[16] br[16] wl[75] vdd gnd cell_6t
Xbit_r76_c16 bl[16] br[16] wl[76] vdd gnd cell_6t
Xbit_r77_c16 bl[16] br[16] wl[77] vdd gnd cell_6t
Xbit_r78_c16 bl[16] br[16] wl[78] vdd gnd cell_6t
Xbit_r79_c16 bl[16] br[16] wl[79] vdd gnd cell_6t
Xbit_r80_c16 bl[16] br[16] wl[80] vdd gnd cell_6t
Xbit_r81_c16 bl[16] br[16] wl[81] vdd gnd cell_6t
Xbit_r82_c16 bl[16] br[16] wl[82] vdd gnd cell_6t
Xbit_r83_c16 bl[16] br[16] wl[83] vdd gnd cell_6t
Xbit_r84_c16 bl[16] br[16] wl[84] vdd gnd cell_6t
Xbit_r85_c16 bl[16] br[16] wl[85] vdd gnd cell_6t
Xbit_r86_c16 bl[16] br[16] wl[86] vdd gnd cell_6t
Xbit_r87_c16 bl[16] br[16] wl[87] vdd gnd cell_6t
Xbit_r88_c16 bl[16] br[16] wl[88] vdd gnd cell_6t
Xbit_r89_c16 bl[16] br[16] wl[89] vdd gnd cell_6t
Xbit_r90_c16 bl[16] br[16] wl[90] vdd gnd cell_6t
Xbit_r91_c16 bl[16] br[16] wl[91] vdd gnd cell_6t
Xbit_r92_c16 bl[16] br[16] wl[92] vdd gnd cell_6t
Xbit_r93_c16 bl[16] br[16] wl[93] vdd gnd cell_6t
Xbit_r94_c16 bl[16] br[16] wl[94] vdd gnd cell_6t
Xbit_r95_c16 bl[16] br[16] wl[95] vdd gnd cell_6t
Xbit_r96_c16 bl[16] br[16] wl[96] vdd gnd cell_6t
Xbit_r97_c16 bl[16] br[16] wl[97] vdd gnd cell_6t
Xbit_r98_c16 bl[16] br[16] wl[98] vdd gnd cell_6t
Xbit_r99_c16 bl[16] br[16] wl[99] vdd gnd cell_6t
Xbit_r100_c16 bl[16] br[16] wl[100] vdd gnd cell_6t
Xbit_r101_c16 bl[16] br[16] wl[101] vdd gnd cell_6t
Xbit_r102_c16 bl[16] br[16] wl[102] vdd gnd cell_6t
Xbit_r103_c16 bl[16] br[16] wl[103] vdd gnd cell_6t
Xbit_r104_c16 bl[16] br[16] wl[104] vdd gnd cell_6t
Xbit_r105_c16 bl[16] br[16] wl[105] vdd gnd cell_6t
Xbit_r106_c16 bl[16] br[16] wl[106] vdd gnd cell_6t
Xbit_r107_c16 bl[16] br[16] wl[107] vdd gnd cell_6t
Xbit_r108_c16 bl[16] br[16] wl[108] vdd gnd cell_6t
Xbit_r109_c16 bl[16] br[16] wl[109] vdd gnd cell_6t
Xbit_r110_c16 bl[16] br[16] wl[110] vdd gnd cell_6t
Xbit_r111_c16 bl[16] br[16] wl[111] vdd gnd cell_6t
Xbit_r112_c16 bl[16] br[16] wl[112] vdd gnd cell_6t
Xbit_r113_c16 bl[16] br[16] wl[113] vdd gnd cell_6t
Xbit_r114_c16 bl[16] br[16] wl[114] vdd gnd cell_6t
Xbit_r115_c16 bl[16] br[16] wl[115] vdd gnd cell_6t
Xbit_r116_c16 bl[16] br[16] wl[116] vdd gnd cell_6t
Xbit_r117_c16 bl[16] br[16] wl[117] vdd gnd cell_6t
Xbit_r118_c16 bl[16] br[16] wl[118] vdd gnd cell_6t
Xbit_r119_c16 bl[16] br[16] wl[119] vdd gnd cell_6t
Xbit_r120_c16 bl[16] br[16] wl[120] vdd gnd cell_6t
Xbit_r121_c16 bl[16] br[16] wl[121] vdd gnd cell_6t
Xbit_r122_c16 bl[16] br[16] wl[122] vdd gnd cell_6t
Xbit_r123_c16 bl[16] br[16] wl[123] vdd gnd cell_6t
Xbit_r124_c16 bl[16] br[16] wl[124] vdd gnd cell_6t
Xbit_r125_c16 bl[16] br[16] wl[125] vdd gnd cell_6t
Xbit_r126_c16 bl[16] br[16] wl[126] vdd gnd cell_6t
Xbit_r127_c16 bl[16] br[16] wl[127] vdd gnd cell_6t
Xbit_r128_c16 bl[16] br[16] wl[128] vdd gnd cell_6t
Xbit_r129_c16 bl[16] br[16] wl[129] vdd gnd cell_6t
Xbit_r130_c16 bl[16] br[16] wl[130] vdd gnd cell_6t
Xbit_r131_c16 bl[16] br[16] wl[131] vdd gnd cell_6t
Xbit_r132_c16 bl[16] br[16] wl[132] vdd gnd cell_6t
Xbit_r133_c16 bl[16] br[16] wl[133] vdd gnd cell_6t
Xbit_r134_c16 bl[16] br[16] wl[134] vdd gnd cell_6t
Xbit_r135_c16 bl[16] br[16] wl[135] vdd gnd cell_6t
Xbit_r136_c16 bl[16] br[16] wl[136] vdd gnd cell_6t
Xbit_r137_c16 bl[16] br[16] wl[137] vdd gnd cell_6t
Xbit_r138_c16 bl[16] br[16] wl[138] vdd gnd cell_6t
Xbit_r139_c16 bl[16] br[16] wl[139] vdd gnd cell_6t
Xbit_r140_c16 bl[16] br[16] wl[140] vdd gnd cell_6t
Xbit_r141_c16 bl[16] br[16] wl[141] vdd gnd cell_6t
Xbit_r142_c16 bl[16] br[16] wl[142] vdd gnd cell_6t
Xbit_r143_c16 bl[16] br[16] wl[143] vdd gnd cell_6t
Xbit_r144_c16 bl[16] br[16] wl[144] vdd gnd cell_6t
Xbit_r145_c16 bl[16] br[16] wl[145] vdd gnd cell_6t
Xbit_r146_c16 bl[16] br[16] wl[146] vdd gnd cell_6t
Xbit_r147_c16 bl[16] br[16] wl[147] vdd gnd cell_6t
Xbit_r148_c16 bl[16] br[16] wl[148] vdd gnd cell_6t
Xbit_r149_c16 bl[16] br[16] wl[149] vdd gnd cell_6t
Xbit_r150_c16 bl[16] br[16] wl[150] vdd gnd cell_6t
Xbit_r151_c16 bl[16] br[16] wl[151] vdd gnd cell_6t
Xbit_r152_c16 bl[16] br[16] wl[152] vdd gnd cell_6t
Xbit_r153_c16 bl[16] br[16] wl[153] vdd gnd cell_6t
Xbit_r154_c16 bl[16] br[16] wl[154] vdd gnd cell_6t
Xbit_r155_c16 bl[16] br[16] wl[155] vdd gnd cell_6t
Xbit_r156_c16 bl[16] br[16] wl[156] vdd gnd cell_6t
Xbit_r157_c16 bl[16] br[16] wl[157] vdd gnd cell_6t
Xbit_r158_c16 bl[16] br[16] wl[158] vdd gnd cell_6t
Xbit_r159_c16 bl[16] br[16] wl[159] vdd gnd cell_6t
Xbit_r160_c16 bl[16] br[16] wl[160] vdd gnd cell_6t
Xbit_r161_c16 bl[16] br[16] wl[161] vdd gnd cell_6t
Xbit_r162_c16 bl[16] br[16] wl[162] vdd gnd cell_6t
Xbit_r163_c16 bl[16] br[16] wl[163] vdd gnd cell_6t
Xbit_r164_c16 bl[16] br[16] wl[164] vdd gnd cell_6t
Xbit_r165_c16 bl[16] br[16] wl[165] vdd gnd cell_6t
Xbit_r166_c16 bl[16] br[16] wl[166] vdd gnd cell_6t
Xbit_r167_c16 bl[16] br[16] wl[167] vdd gnd cell_6t
Xbit_r168_c16 bl[16] br[16] wl[168] vdd gnd cell_6t
Xbit_r169_c16 bl[16] br[16] wl[169] vdd gnd cell_6t
Xbit_r170_c16 bl[16] br[16] wl[170] vdd gnd cell_6t
Xbit_r171_c16 bl[16] br[16] wl[171] vdd gnd cell_6t
Xbit_r172_c16 bl[16] br[16] wl[172] vdd gnd cell_6t
Xbit_r173_c16 bl[16] br[16] wl[173] vdd gnd cell_6t
Xbit_r174_c16 bl[16] br[16] wl[174] vdd gnd cell_6t
Xbit_r175_c16 bl[16] br[16] wl[175] vdd gnd cell_6t
Xbit_r176_c16 bl[16] br[16] wl[176] vdd gnd cell_6t
Xbit_r177_c16 bl[16] br[16] wl[177] vdd gnd cell_6t
Xbit_r178_c16 bl[16] br[16] wl[178] vdd gnd cell_6t
Xbit_r179_c16 bl[16] br[16] wl[179] vdd gnd cell_6t
Xbit_r180_c16 bl[16] br[16] wl[180] vdd gnd cell_6t
Xbit_r181_c16 bl[16] br[16] wl[181] vdd gnd cell_6t
Xbit_r182_c16 bl[16] br[16] wl[182] vdd gnd cell_6t
Xbit_r183_c16 bl[16] br[16] wl[183] vdd gnd cell_6t
Xbit_r184_c16 bl[16] br[16] wl[184] vdd gnd cell_6t
Xbit_r185_c16 bl[16] br[16] wl[185] vdd gnd cell_6t
Xbit_r186_c16 bl[16] br[16] wl[186] vdd gnd cell_6t
Xbit_r187_c16 bl[16] br[16] wl[187] vdd gnd cell_6t
Xbit_r188_c16 bl[16] br[16] wl[188] vdd gnd cell_6t
Xbit_r189_c16 bl[16] br[16] wl[189] vdd gnd cell_6t
Xbit_r190_c16 bl[16] br[16] wl[190] vdd gnd cell_6t
Xbit_r191_c16 bl[16] br[16] wl[191] vdd gnd cell_6t
Xbit_r192_c16 bl[16] br[16] wl[192] vdd gnd cell_6t
Xbit_r193_c16 bl[16] br[16] wl[193] vdd gnd cell_6t
Xbit_r194_c16 bl[16] br[16] wl[194] vdd gnd cell_6t
Xbit_r195_c16 bl[16] br[16] wl[195] vdd gnd cell_6t
Xbit_r196_c16 bl[16] br[16] wl[196] vdd gnd cell_6t
Xbit_r197_c16 bl[16] br[16] wl[197] vdd gnd cell_6t
Xbit_r198_c16 bl[16] br[16] wl[198] vdd gnd cell_6t
Xbit_r199_c16 bl[16] br[16] wl[199] vdd gnd cell_6t
Xbit_r200_c16 bl[16] br[16] wl[200] vdd gnd cell_6t
Xbit_r201_c16 bl[16] br[16] wl[201] vdd gnd cell_6t
Xbit_r202_c16 bl[16] br[16] wl[202] vdd gnd cell_6t
Xbit_r203_c16 bl[16] br[16] wl[203] vdd gnd cell_6t
Xbit_r204_c16 bl[16] br[16] wl[204] vdd gnd cell_6t
Xbit_r205_c16 bl[16] br[16] wl[205] vdd gnd cell_6t
Xbit_r206_c16 bl[16] br[16] wl[206] vdd gnd cell_6t
Xbit_r207_c16 bl[16] br[16] wl[207] vdd gnd cell_6t
Xbit_r208_c16 bl[16] br[16] wl[208] vdd gnd cell_6t
Xbit_r209_c16 bl[16] br[16] wl[209] vdd gnd cell_6t
Xbit_r210_c16 bl[16] br[16] wl[210] vdd gnd cell_6t
Xbit_r211_c16 bl[16] br[16] wl[211] vdd gnd cell_6t
Xbit_r212_c16 bl[16] br[16] wl[212] vdd gnd cell_6t
Xbit_r213_c16 bl[16] br[16] wl[213] vdd gnd cell_6t
Xbit_r214_c16 bl[16] br[16] wl[214] vdd gnd cell_6t
Xbit_r215_c16 bl[16] br[16] wl[215] vdd gnd cell_6t
Xbit_r216_c16 bl[16] br[16] wl[216] vdd gnd cell_6t
Xbit_r217_c16 bl[16] br[16] wl[217] vdd gnd cell_6t
Xbit_r218_c16 bl[16] br[16] wl[218] vdd gnd cell_6t
Xbit_r219_c16 bl[16] br[16] wl[219] vdd gnd cell_6t
Xbit_r220_c16 bl[16] br[16] wl[220] vdd gnd cell_6t
Xbit_r221_c16 bl[16] br[16] wl[221] vdd gnd cell_6t
Xbit_r222_c16 bl[16] br[16] wl[222] vdd gnd cell_6t
Xbit_r223_c16 bl[16] br[16] wl[223] vdd gnd cell_6t
Xbit_r224_c16 bl[16] br[16] wl[224] vdd gnd cell_6t
Xbit_r225_c16 bl[16] br[16] wl[225] vdd gnd cell_6t
Xbit_r226_c16 bl[16] br[16] wl[226] vdd gnd cell_6t
Xbit_r227_c16 bl[16] br[16] wl[227] vdd gnd cell_6t
Xbit_r228_c16 bl[16] br[16] wl[228] vdd gnd cell_6t
Xbit_r229_c16 bl[16] br[16] wl[229] vdd gnd cell_6t
Xbit_r230_c16 bl[16] br[16] wl[230] vdd gnd cell_6t
Xbit_r231_c16 bl[16] br[16] wl[231] vdd gnd cell_6t
Xbit_r232_c16 bl[16] br[16] wl[232] vdd gnd cell_6t
Xbit_r233_c16 bl[16] br[16] wl[233] vdd gnd cell_6t
Xbit_r234_c16 bl[16] br[16] wl[234] vdd gnd cell_6t
Xbit_r235_c16 bl[16] br[16] wl[235] vdd gnd cell_6t
Xbit_r236_c16 bl[16] br[16] wl[236] vdd gnd cell_6t
Xbit_r237_c16 bl[16] br[16] wl[237] vdd gnd cell_6t
Xbit_r238_c16 bl[16] br[16] wl[238] vdd gnd cell_6t
Xbit_r239_c16 bl[16] br[16] wl[239] vdd gnd cell_6t
Xbit_r240_c16 bl[16] br[16] wl[240] vdd gnd cell_6t
Xbit_r241_c16 bl[16] br[16] wl[241] vdd gnd cell_6t
Xbit_r242_c16 bl[16] br[16] wl[242] vdd gnd cell_6t
Xbit_r243_c16 bl[16] br[16] wl[243] vdd gnd cell_6t
Xbit_r244_c16 bl[16] br[16] wl[244] vdd gnd cell_6t
Xbit_r245_c16 bl[16] br[16] wl[245] vdd gnd cell_6t
Xbit_r246_c16 bl[16] br[16] wl[246] vdd gnd cell_6t
Xbit_r247_c16 bl[16] br[16] wl[247] vdd gnd cell_6t
Xbit_r248_c16 bl[16] br[16] wl[248] vdd gnd cell_6t
Xbit_r249_c16 bl[16] br[16] wl[249] vdd gnd cell_6t
Xbit_r250_c16 bl[16] br[16] wl[250] vdd gnd cell_6t
Xbit_r251_c16 bl[16] br[16] wl[251] vdd gnd cell_6t
Xbit_r252_c16 bl[16] br[16] wl[252] vdd gnd cell_6t
Xbit_r253_c16 bl[16] br[16] wl[253] vdd gnd cell_6t
Xbit_r254_c16 bl[16] br[16] wl[254] vdd gnd cell_6t
Xbit_r255_c16 bl[16] br[16] wl[255] vdd gnd cell_6t
Xbit_r0_c17 bl[17] br[17] wl[0] vdd gnd cell_6t
Xbit_r1_c17 bl[17] br[17] wl[1] vdd gnd cell_6t
Xbit_r2_c17 bl[17] br[17] wl[2] vdd gnd cell_6t
Xbit_r3_c17 bl[17] br[17] wl[3] vdd gnd cell_6t
Xbit_r4_c17 bl[17] br[17] wl[4] vdd gnd cell_6t
Xbit_r5_c17 bl[17] br[17] wl[5] vdd gnd cell_6t
Xbit_r6_c17 bl[17] br[17] wl[6] vdd gnd cell_6t
Xbit_r7_c17 bl[17] br[17] wl[7] vdd gnd cell_6t
Xbit_r8_c17 bl[17] br[17] wl[8] vdd gnd cell_6t
Xbit_r9_c17 bl[17] br[17] wl[9] vdd gnd cell_6t
Xbit_r10_c17 bl[17] br[17] wl[10] vdd gnd cell_6t
Xbit_r11_c17 bl[17] br[17] wl[11] vdd gnd cell_6t
Xbit_r12_c17 bl[17] br[17] wl[12] vdd gnd cell_6t
Xbit_r13_c17 bl[17] br[17] wl[13] vdd gnd cell_6t
Xbit_r14_c17 bl[17] br[17] wl[14] vdd gnd cell_6t
Xbit_r15_c17 bl[17] br[17] wl[15] vdd gnd cell_6t
Xbit_r16_c17 bl[17] br[17] wl[16] vdd gnd cell_6t
Xbit_r17_c17 bl[17] br[17] wl[17] vdd gnd cell_6t
Xbit_r18_c17 bl[17] br[17] wl[18] vdd gnd cell_6t
Xbit_r19_c17 bl[17] br[17] wl[19] vdd gnd cell_6t
Xbit_r20_c17 bl[17] br[17] wl[20] vdd gnd cell_6t
Xbit_r21_c17 bl[17] br[17] wl[21] vdd gnd cell_6t
Xbit_r22_c17 bl[17] br[17] wl[22] vdd gnd cell_6t
Xbit_r23_c17 bl[17] br[17] wl[23] vdd gnd cell_6t
Xbit_r24_c17 bl[17] br[17] wl[24] vdd gnd cell_6t
Xbit_r25_c17 bl[17] br[17] wl[25] vdd gnd cell_6t
Xbit_r26_c17 bl[17] br[17] wl[26] vdd gnd cell_6t
Xbit_r27_c17 bl[17] br[17] wl[27] vdd gnd cell_6t
Xbit_r28_c17 bl[17] br[17] wl[28] vdd gnd cell_6t
Xbit_r29_c17 bl[17] br[17] wl[29] vdd gnd cell_6t
Xbit_r30_c17 bl[17] br[17] wl[30] vdd gnd cell_6t
Xbit_r31_c17 bl[17] br[17] wl[31] vdd gnd cell_6t
Xbit_r32_c17 bl[17] br[17] wl[32] vdd gnd cell_6t
Xbit_r33_c17 bl[17] br[17] wl[33] vdd gnd cell_6t
Xbit_r34_c17 bl[17] br[17] wl[34] vdd gnd cell_6t
Xbit_r35_c17 bl[17] br[17] wl[35] vdd gnd cell_6t
Xbit_r36_c17 bl[17] br[17] wl[36] vdd gnd cell_6t
Xbit_r37_c17 bl[17] br[17] wl[37] vdd gnd cell_6t
Xbit_r38_c17 bl[17] br[17] wl[38] vdd gnd cell_6t
Xbit_r39_c17 bl[17] br[17] wl[39] vdd gnd cell_6t
Xbit_r40_c17 bl[17] br[17] wl[40] vdd gnd cell_6t
Xbit_r41_c17 bl[17] br[17] wl[41] vdd gnd cell_6t
Xbit_r42_c17 bl[17] br[17] wl[42] vdd gnd cell_6t
Xbit_r43_c17 bl[17] br[17] wl[43] vdd gnd cell_6t
Xbit_r44_c17 bl[17] br[17] wl[44] vdd gnd cell_6t
Xbit_r45_c17 bl[17] br[17] wl[45] vdd gnd cell_6t
Xbit_r46_c17 bl[17] br[17] wl[46] vdd gnd cell_6t
Xbit_r47_c17 bl[17] br[17] wl[47] vdd gnd cell_6t
Xbit_r48_c17 bl[17] br[17] wl[48] vdd gnd cell_6t
Xbit_r49_c17 bl[17] br[17] wl[49] vdd gnd cell_6t
Xbit_r50_c17 bl[17] br[17] wl[50] vdd gnd cell_6t
Xbit_r51_c17 bl[17] br[17] wl[51] vdd gnd cell_6t
Xbit_r52_c17 bl[17] br[17] wl[52] vdd gnd cell_6t
Xbit_r53_c17 bl[17] br[17] wl[53] vdd gnd cell_6t
Xbit_r54_c17 bl[17] br[17] wl[54] vdd gnd cell_6t
Xbit_r55_c17 bl[17] br[17] wl[55] vdd gnd cell_6t
Xbit_r56_c17 bl[17] br[17] wl[56] vdd gnd cell_6t
Xbit_r57_c17 bl[17] br[17] wl[57] vdd gnd cell_6t
Xbit_r58_c17 bl[17] br[17] wl[58] vdd gnd cell_6t
Xbit_r59_c17 bl[17] br[17] wl[59] vdd gnd cell_6t
Xbit_r60_c17 bl[17] br[17] wl[60] vdd gnd cell_6t
Xbit_r61_c17 bl[17] br[17] wl[61] vdd gnd cell_6t
Xbit_r62_c17 bl[17] br[17] wl[62] vdd gnd cell_6t
Xbit_r63_c17 bl[17] br[17] wl[63] vdd gnd cell_6t
Xbit_r64_c17 bl[17] br[17] wl[64] vdd gnd cell_6t
Xbit_r65_c17 bl[17] br[17] wl[65] vdd gnd cell_6t
Xbit_r66_c17 bl[17] br[17] wl[66] vdd gnd cell_6t
Xbit_r67_c17 bl[17] br[17] wl[67] vdd gnd cell_6t
Xbit_r68_c17 bl[17] br[17] wl[68] vdd gnd cell_6t
Xbit_r69_c17 bl[17] br[17] wl[69] vdd gnd cell_6t
Xbit_r70_c17 bl[17] br[17] wl[70] vdd gnd cell_6t
Xbit_r71_c17 bl[17] br[17] wl[71] vdd gnd cell_6t
Xbit_r72_c17 bl[17] br[17] wl[72] vdd gnd cell_6t
Xbit_r73_c17 bl[17] br[17] wl[73] vdd gnd cell_6t
Xbit_r74_c17 bl[17] br[17] wl[74] vdd gnd cell_6t
Xbit_r75_c17 bl[17] br[17] wl[75] vdd gnd cell_6t
Xbit_r76_c17 bl[17] br[17] wl[76] vdd gnd cell_6t
Xbit_r77_c17 bl[17] br[17] wl[77] vdd gnd cell_6t
Xbit_r78_c17 bl[17] br[17] wl[78] vdd gnd cell_6t
Xbit_r79_c17 bl[17] br[17] wl[79] vdd gnd cell_6t
Xbit_r80_c17 bl[17] br[17] wl[80] vdd gnd cell_6t
Xbit_r81_c17 bl[17] br[17] wl[81] vdd gnd cell_6t
Xbit_r82_c17 bl[17] br[17] wl[82] vdd gnd cell_6t
Xbit_r83_c17 bl[17] br[17] wl[83] vdd gnd cell_6t
Xbit_r84_c17 bl[17] br[17] wl[84] vdd gnd cell_6t
Xbit_r85_c17 bl[17] br[17] wl[85] vdd gnd cell_6t
Xbit_r86_c17 bl[17] br[17] wl[86] vdd gnd cell_6t
Xbit_r87_c17 bl[17] br[17] wl[87] vdd gnd cell_6t
Xbit_r88_c17 bl[17] br[17] wl[88] vdd gnd cell_6t
Xbit_r89_c17 bl[17] br[17] wl[89] vdd gnd cell_6t
Xbit_r90_c17 bl[17] br[17] wl[90] vdd gnd cell_6t
Xbit_r91_c17 bl[17] br[17] wl[91] vdd gnd cell_6t
Xbit_r92_c17 bl[17] br[17] wl[92] vdd gnd cell_6t
Xbit_r93_c17 bl[17] br[17] wl[93] vdd gnd cell_6t
Xbit_r94_c17 bl[17] br[17] wl[94] vdd gnd cell_6t
Xbit_r95_c17 bl[17] br[17] wl[95] vdd gnd cell_6t
Xbit_r96_c17 bl[17] br[17] wl[96] vdd gnd cell_6t
Xbit_r97_c17 bl[17] br[17] wl[97] vdd gnd cell_6t
Xbit_r98_c17 bl[17] br[17] wl[98] vdd gnd cell_6t
Xbit_r99_c17 bl[17] br[17] wl[99] vdd gnd cell_6t
Xbit_r100_c17 bl[17] br[17] wl[100] vdd gnd cell_6t
Xbit_r101_c17 bl[17] br[17] wl[101] vdd gnd cell_6t
Xbit_r102_c17 bl[17] br[17] wl[102] vdd gnd cell_6t
Xbit_r103_c17 bl[17] br[17] wl[103] vdd gnd cell_6t
Xbit_r104_c17 bl[17] br[17] wl[104] vdd gnd cell_6t
Xbit_r105_c17 bl[17] br[17] wl[105] vdd gnd cell_6t
Xbit_r106_c17 bl[17] br[17] wl[106] vdd gnd cell_6t
Xbit_r107_c17 bl[17] br[17] wl[107] vdd gnd cell_6t
Xbit_r108_c17 bl[17] br[17] wl[108] vdd gnd cell_6t
Xbit_r109_c17 bl[17] br[17] wl[109] vdd gnd cell_6t
Xbit_r110_c17 bl[17] br[17] wl[110] vdd gnd cell_6t
Xbit_r111_c17 bl[17] br[17] wl[111] vdd gnd cell_6t
Xbit_r112_c17 bl[17] br[17] wl[112] vdd gnd cell_6t
Xbit_r113_c17 bl[17] br[17] wl[113] vdd gnd cell_6t
Xbit_r114_c17 bl[17] br[17] wl[114] vdd gnd cell_6t
Xbit_r115_c17 bl[17] br[17] wl[115] vdd gnd cell_6t
Xbit_r116_c17 bl[17] br[17] wl[116] vdd gnd cell_6t
Xbit_r117_c17 bl[17] br[17] wl[117] vdd gnd cell_6t
Xbit_r118_c17 bl[17] br[17] wl[118] vdd gnd cell_6t
Xbit_r119_c17 bl[17] br[17] wl[119] vdd gnd cell_6t
Xbit_r120_c17 bl[17] br[17] wl[120] vdd gnd cell_6t
Xbit_r121_c17 bl[17] br[17] wl[121] vdd gnd cell_6t
Xbit_r122_c17 bl[17] br[17] wl[122] vdd gnd cell_6t
Xbit_r123_c17 bl[17] br[17] wl[123] vdd gnd cell_6t
Xbit_r124_c17 bl[17] br[17] wl[124] vdd gnd cell_6t
Xbit_r125_c17 bl[17] br[17] wl[125] vdd gnd cell_6t
Xbit_r126_c17 bl[17] br[17] wl[126] vdd gnd cell_6t
Xbit_r127_c17 bl[17] br[17] wl[127] vdd gnd cell_6t
Xbit_r128_c17 bl[17] br[17] wl[128] vdd gnd cell_6t
Xbit_r129_c17 bl[17] br[17] wl[129] vdd gnd cell_6t
Xbit_r130_c17 bl[17] br[17] wl[130] vdd gnd cell_6t
Xbit_r131_c17 bl[17] br[17] wl[131] vdd gnd cell_6t
Xbit_r132_c17 bl[17] br[17] wl[132] vdd gnd cell_6t
Xbit_r133_c17 bl[17] br[17] wl[133] vdd gnd cell_6t
Xbit_r134_c17 bl[17] br[17] wl[134] vdd gnd cell_6t
Xbit_r135_c17 bl[17] br[17] wl[135] vdd gnd cell_6t
Xbit_r136_c17 bl[17] br[17] wl[136] vdd gnd cell_6t
Xbit_r137_c17 bl[17] br[17] wl[137] vdd gnd cell_6t
Xbit_r138_c17 bl[17] br[17] wl[138] vdd gnd cell_6t
Xbit_r139_c17 bl[17] br[17] wl[139] vdd gnd cell_6t
Xbit_r140_c17 bl[17] br[17] wl[140] vdd gnd cell_6t
Xbit_r141_c17 bl[17] br[17] wl[141] vdd gnd cell_6t
Xbit_r142_c17 bl[17] br[17] wl[142] vdd gnd cell_6t
Xbit_r143_c17 bl[17] br[17] wl[143] vdd gnd cell_6t
Xbit_r144_c17 bl[17] br[17] wl[144] vdd gnd cell_6t
Xbit_r145_c17 bl[17] br[17] wl[145] vdd gnd cell_6t
Xbit_r146_c17 bl[17] br[17] wl[146] vdd gnd cell_6t
Xbit_r147_c17 bl[17] br[17] wl[147] vdd gnd cell_6t
Xbit_r148_c17 bl[17] br[17] wl[148] vdd gnd cell_6t
Xbit_r149_c17 bl[17] br[17] wl[149] vdd gnd cell_6t
Xbit_r150_c17 bl[17] br[17] wl[150] vdd gnd cell_6t
Xbit_r151_c17 bl[17] br[17] wl[151] vdd gnd cell_6t
Xbit_r152_c17 bl[17] br[17] wl[152] vdd gnd cell_6t
Xbit_r153_c17 bl[17] br[17] wl[153] vdd gnd cell_6t
Xbit_r154_c17 bl[17] br[17] wl[154] vdd gnd cell_6t
Xbit_r155_c17 bl[17] br[17] wl[155] vdd gnd cell_6t
Xbit_r156_c17 bl[17] br[17] wl[156] vdd gnd cell_6t
Xbit_r157_c17 bl[17] br[17] wl[157] vdd gnd cell_6t
Xbit_r158_c17 bl[17] br[17] wl[158] vdd gnd cell_6t
Xbit_r159_c17 bl[17] br[17] wl[159] vdd gnd cell_6t
Xbit_r160_c17 bl[17] br[17] wl[160] vdd gnd cell_6t
Xbit_r161_c17 bl[17] br[17] wl[161] vdd gnd cell_6t
Xbit_r162_c17 bl[17] br[17] wl[162] vdd gnd cell_6t
Xbit_r163_c17 bl[17] br[17] wl[163] vdd gnd cell_6t
Xbit_r164_c17 bl[17] br[17] wl[164] vdd gnd cell_6t
Xbit_r165_c17 bl[17] br[17] wl[165] vdd gnd cell_6t
Xbit_r166_c17 bl[17] br[17] wl[166] vdd gnd cell_6t
Xbit_r167_c17 bl[17] br[17] wl[167] vdd gnd cell_6t
Xbit_r168_c17 bl[17] br[17] wl[168] vdd gnd cell_6t
Xbit_r169_c17 bl[17] br[17] wl[169] vdd gnd cell_6t
Xbit_r170_c17 bl[17] br[17] wl[170] vdd gnd cell_6t
Xbit_r171_c17 bl[17] br[17] wl[171] vdd gnd cell_6t
Xbit_r172_c17 bl[17] br[17] wl[172] vdd gnd cell_6t
Xbit_r173_c17 bl[17] br[17] wl[173] vdd gnd cell_6t
Xbit_r174_c17 bl[17] br[17] wl[174] vdd gnd cell_6t
Xbit_r175_c17 bl[17] br[17] wl[175] vdd gnd cell_6t
Xbit_r176_c17 bl[17] br[17] wl[176] vdd gnd cell_6t
Xbit_r177_c17 bl[17] br[17] wl[177] vdd gnd cell_6t
Xbit_r178_c17 bl[17] br[17] wl[178] vdd gnd cell_6t
Xbit_r179_c17 bl[17] br[17] wl[179] vdd gnd cell_6t
Xbit_r180_c17 bl[17] br[17] wl[180] vdd gnd cell_6t
Xbit_r181_c17 bl[17] br[17] wl[181] vdd gnd cell_6t
Xbit_r182_c17 bl[17] br[17] wl[182] vdd gnd cell_6t
Xbit_r183_c17 bl[17] br[17] wl[183] vdd gnd cell_6t
Xbit_r184_c17 bl[17] br[17] wl[184] vdd gnd cell_6t
Xbit_r185_c17 bl[17] br[17] wl[185] vdd gnd cell_6t
Xbit_r186_c17 bl[17] br[17] wl[186] vdd gnd cell_6t
Xbit_r187_c17 bl[17] br[17] wl[187] vdd gnd cell_6t
Xbit_r188_c17 bl[17] br[17] wl[188] vdd gnd cell_6t
Xbit_r189_c17 bl[17] br[17] wl[189] vdd gnd cell_6t
Xbit_r190_c17 bl[17] br[17] wl[190] vdd gnd cell_6t
Xbit_r191_c17 bl[17] br[17] wl[191] vdd gnd cell_6t
Xbit_r192_c17 bl[17] br[17] wl[192] vdd gnd cell_6t
Xbit_r193_c17 bl[17] br[17] wl[193] vdd gnd cell_6t
Xbit_r194_c17 bl[17] br[17] wl[194] vdd gnd cell_6t
Xbit_r195_c17 bl[17] br[17] wl[195] vdd gnd cell_6t
Xbit_r196_c17 bl[17] br[17] wl[196] vdd gnd cell_6t
Xbit_r197_c17 bl[17] br[17] wl[197] vdd gnd cell_6t
Xbit_r198_c17 bl[17] br[17] wl[198] vdd gnd cell_6t
Xbit_r199_c17 bl[17] br[17] wl[199] vdd gnd cell_6t
Xbit_r200_c17 bl[17] br[17] wl[200] vdd gnd cell_6t
Xbit_r201_c17 bl[17] br[17] wl[201] vdd gnd cell_6t
Xbit_r202_c17 bl[17] br[17] wl[202] vdd gnd cell_6t
Xbit_r203_c17 bl[17] br[17] wl[203] vdd gnd cell_6t
Xbit_r204_c17 bl[17] br[17] wl[204] vdd gnd cell_6t
Xbit_r205_c17 bl[17] br[17] wl[205] vdd gnd cell_6t
Xbit_r206_c17 bl[17] br[17] wl[206] vdd gnd cell_6t
Xbit_r207_c17 bl[17] br[17] wl[207] vdd gnd cell_6t
Xbit_r208_c17 bl[17] br[17] wl[208] vdd gnd cell_6t
Xbit_r209_c17 bl[17] br[17] wl[209] vdd gnd cell_6t
Xbit_r210_c17 bl[17] br[17] wl[210] vdd gnd cell_6t
Xbit_r211_c17 bl[17] br[17] wl[211] vdd gnd cell_6t
Xbit_r212_c17 bl[17] br[17] wl[212] vdd gnd cell_6t
Xbit_r213_c17 bl[17] br[17] wl[213] vdd gnd cell_6t
Xbit_r214_c17 bl[17] br[17] wl[214] vdd gnd cell_6t
Xbit_r215_c17 bl[17] br[17] wl[215] vdd gnd cell_6t
Xbit_r216_c17 bl[17] br[17] wl[216] vdd gnd cell_6t
Xbit_r217_c17 bl[17] br[17] wl[217] vdd gnd cell_6t
Xbit_r218_c17 bl[17] br[17] wl[218] vdd gnd cell_6t
Xbit_r219_c17 bl[17] br[17] wl[219] vdd gnd cell_6t
Xbit_r220_c17 bl[17] br[17] wl[220] vdd gnd cell_6t
Xbit_r221_c17 bl[17] br[17] wl[221] vdd gnd cell_6t
Xbit_r222_c17 bl[17] br[17] wl[222] vdd gnd cell_6t
Xbit_r223_c17 bl[17] br[17] wl[223] vdd gnd cell_6t
Xbit_r224_c17 bl[17] br[17] wl[224] vdd gnd cell_6t
Xbit_r225_c17 bl[17] br[17] wl[225] vdd gnd cell_6t
Xbit_r226_c17 bl[17] br[17] wl[226] vdd gnd cell_6t
Xbit_r227_c17 bl[17] br[17] wl[227] vdd gnd cell_6t
Xbit_r228_c17 bl[17] br[17] wl[228] vdd gnd cell_6t
Xbit_r229_c17 bl[17] br[17] wl[229] vdd gnd cell_6t
Xbit_r230_c17 bl[17] br[17] wl[230] vdd gnd cell_6t
Xbit_r231_c17 bl[17] br[17] wl[231] vdd gnd cell_6t
Xbit_r232_c17 bl[17] br[17] wl[232] vdd gnd cell_6t
Xbit_r233_c17 bl[17] br[17] wl[233] vdd gnd cell_6t
Xbit_r234_c17 bl[17] br[17] wl[234] vdd gnd cell_6t
Xbit_r235_c17 bl[17] br[17] wl[235] vdd gnd cell_6t
Xbit_r236_c17 bl[17] br[17] wl[236] vdd gnd cell_6t
Xbit_r237_c17 bl[17] br[17] wl[237] vdd gnd cell_6t
Xbit_r238_c17 bl[17] br[17] wl[238] vdd gnd cell_6t
Xbit_r239_c17 bl[17] br[17] wl[239] vdd gnd cell_6t
Xbit_r240_c17 bl[17] br[17] wl[240] vdd gnd cell_6t
Xbit_r241_c17 bl[17] br[17] wl[241] vdd gnd cell_6t
Xbit_r242_c17 bl[17] br[17] wl[242] vdd gnd cell_6t
Xbit_r243_c17 bl[17] br[17] wl[243] vdd gnd cell_6t
Xbit_r244_c17 bl[17] br[17] wl[244] vdd gnd cell_6t
Xbit_r245_c17 bl[17] br[17] wl[245] vdd gnd cell_6t
Xbit_r246_c17 bl[17] br[17] wl[246] vdd gnd cell_6t
Xbit_r247_c17 bl[17] br[17] wl[247] vdd gnd cell_6t
Xbit_r248_c17 bl[17] br[17] wl[248] vdd gnd cell_6t
Xbit_r249_c17 bl[17] br[17] wl[249] vdd gnd cell_6t
Xbit_r250_c17 bl[17] br[17] wl[250] vdd gnd cell_6t
Xbit_r251_c17 bl[17] br[17] wl[251] vdd gnd cell_6t
Xbit_r252_c17 bl[17] br[17] wl[252] vdd gnd cell_6t
Xbit_r253_c17 bl[17] br[17] wl[253] vdd gnd cell_6t
Xbit_r254_c17 bl[17] br[17] wl[254] vdd gnd cell_6t
Xbit_r255_c17 bl[17] br[17] wl[255] vdd gnd cell_6t
Xbit_r0_c18 bl[18] br[18] wl[0] vdd gnd cell_6t
Xbit_r1_c18 bl[18] br[18] wl[1] vdd gnd cell_6t
Xbit_r2_c18 bl[18] br[18] wl[2] vdd gnd cell_6t
Xbit_r3_c18 bl[18] br[18] wl[3] vdd gnd cell_6t
Xbit_r4_c18 bl[18] br[18] wl[4] vdd gnd cell_6t
Xbit_r5_c18 bl[18] br[18] wl[5] vdd gnd cell_6t
Xbit_r6_c18 bl[18] br[18] wl[6] vdd gnd cell_6t
Xbit_r7_c18 bl[18] br[18] wl[7] vdd gnd cell_6t
Xbit_r8_c18 bl[18] br[18] wl[8] vdd gnd cell_6t
Xbit_r9_c18 bl[18] br[18] wl[9] vdd gnd cell_6t
Xbit_r10_c18 bl[18] br[18] wl[10] vdd gnd cell_6t
Xbit_r11_c18 bl[18] br[18] wl[11] vdd gnd cell_6t
Xbit_r12_c18 bl[18] br[18] wl[12] vdd gnd cell_6t
Xbit_r13_c18 bl[18] br[18] wl[13] vdd gnd cell_6t
Xbit_r14_c18 bl[18] br[18] wl[14] vdd gnd cell_6t
Xbit_r15_c18 bl[18] br[18] wl[15] vdd gnd cell_6t
Xbit_r16_c18 bl[18] br[18] wl[16] vdd gnd cell_6t
Xbit_r17_c18 bl[18] br[18] wl[17] vdd gnd cell_6t
Xbit_r18_c18 bl[18] br[18] wl[18] vdd gnd cell_6t
Xbit_r19_c18 bl[18] br[18] wl[19] vdd gnd cell_6t
Xbit_r20_c18 bl[18] br[18] wl[20] vdd gnd cell_6t
Xbit_r21_c18 bl[18] br[18] wl[21] vdd gnd cell_6t
Xbit_r22_c18 bl[18] br[18] wl[22] vdd gnd cell_6t
Xbit_r23_c18 bl[18] br[18] wl[23] vdd gnd cell_6t
Xbit_r24_c18 bl[18] br[18] wl[24] vdd gnd cell_6t
Xbit_r25_c18 bl[18] br[18] wl[25] vdd gnd cell_6t
Xbit_r26_c18 bl[18] br[18] wl[26] vdd gnd cell_6t
Xbit_r27_c18 bl[18] br[18] wl[27] vdd gnd cell_6t
Xbit_r28_c18 bl[18] br[18] wl[28] vdd gnd cell_6t
Xbit_r29_c18 bl[18] br[18] wl[29] vdd gnd cell_6t
Xbit_r30_c18 bl[18] br[18] wl[30] vdd gnd cell_6t
Xbit_r31_c18 bl[18] br[18] wl[31] vdd gnd cell_6t
Xbit_r32_c18 bl[18] br[18] wl[32] vdd gnd cell_6t
Xbit_r33_c18 bl[18] br[18] wl[33] vdd gnd cell_6t
Xbit_r34_c18 bl[18] br[18] wl[34] vdd gnd cell_6t
Xbit_r35_c18 bl[18] br[18] wl[35] vdd gnd cell_6t
Xbit_r36_c18 bl[18] br[18] wl[36] vdd gnd cell_6t
Xbit_r37_c18 bl[18] br[18] wl[37] vdd gnd cell_6t
Xbit_r38_c18 bl[18] br[18] wl[38] vdd gnd cell_6t
Xbit_r39_c18 bl[18] br[18] wl[39] vdd gnd cell_6t
Xbit_r40_c18 bl[18] br[18] wl[40] vdd gnd cell_6t
Xbit_r41_c18 bl[18] br[18] wl[41] vdd gnd cell_6t
Xbit_r42_c18 bl[18] br[18] wl[42] vdd gnd cell_6t
Xbit_r43_c18 bl[18] br[18] wl[43] vdd gnd cell_6t
Xbit_r44_c18 bl[18] br[18] wl[44] vdd gnd cell_6t
Xbit_r45_c18 bl[18] br[18] wl[45] vdd gnd cell_6t
Xbit_r46_c18 bl[18] br[18] wl[46] vdd gnd cell_6t
Xbit_r47_c18 bl[18] br[18] wl[47] vdd gnd cell_6t
Xbit_r48_c18 bl[18] br[18] wl[48] vdd gnd cell_6t
Xbit_r49_c18 bl[18] br[18] wl[49] vdd gnd cell_6t
Xbit_r50_c18 bl[18] br[18] wl[50] vdd gnd cell_6t
Xbit_r51_c18 bl[18] br[18] wl[51] vdd gnd cell_6t
Xbit_r52_c18 bl[18] br[18] wl[52] vdd gnd cell_6t
Xbit_r53_c18 bl[18] br[18] wl[53] vdd gnd cell_6t
Xbit_r54_c18 bl[18] br[18] wl[54] vdd gnd cell_6t
Xbit_r55_c18 bl[18] br[18] wl[55] vdd gnd cell_6t
Xbit_r56_c18 bl[18] br[18] wl[56] vdd gnd cell_6t
Xbit_r57_c18 bl[18] br[18] wl[57] vdd gnd cell_6t
Xbit_r58_c18 bl[18] br[18] wl[58] vdd gnd cell_6t
Xbit_r59_c18 bl[18] br[18] wl[59] vdd gnd cell_6t
Xbit_r60_c18 bl[18] br[18] wl[60] vdd gnd cell_6t
Xbit_r61_c18 bl[18] br[18] wl[61] vdd gnd cell_6t
Xbit_r62_c18 bl[18] br[18] wl[62] vdd gnd cell_6t
Xbit_r63_c18 bl[18] br[18] wl[63] vdd gnd cell_6t
Xbit_r64_c18 bl[18] br[18] wl[64] vdd gnd cell_6t
Xbit_r65_c18 bl[18] br[18] wl[65] vdd gnd cell_6t
Xbit_r66_c18 bl[18] br[18] wl[66] vdd gnd cell_6t
Xbit_r67_c18 bl[18] br[18] wl[67] vdd gnd cell_6t
Xbit_r68_c18 bl[18] br[18] wl[68] vdd gnd cell_6t
Xbit_r69_c18 bl[18] br[18] wl[69] vdd gnd cell_6t
Xbit_r70_c18 bl[18] br[18] wl[70] vdd gnd cell_6t
Xbit_r71_c18 bl[18] br[18] wl[71] vdd gnd cell_6t
Xbit_r72_c18 bl[18] br[18] wl[72] vdd gnd cell_6t
Xbit_r73_c18 bl[18] br[18] wl[73] vdd gnd cell_6t
Xbit_r74_c18 bl[18] br[18] wl[74] vdd gnd cell_6t
Xbit_r75_c18 bl[18] br[18] wl[75] vdd gnd cell_6t
Xbit_r76_c18 bl[18] br[18] wl[76] vdd gnd cell_6t
Xbit_r77_c18 bl[18] br[18] wl[77] vdd gnd cell_6t
Xbit_r78_c18 bl[18] br[18] wl[78] vdd gnd cell_6t
Xbit_r79_c18 bl[18] br[18] wl[79] vdd gnd cell_6t
Xbit_r80_c18 bl[18] br[18] wl[80] vdd gnd cell_6t
Xbit_r81_c18 bl[18] br[18] wl[81] vdd gnd cell_6t
Xbit_r82_c18 bl[18] br[18] wl[82] vdd gnd cell_6t
Xbit_r83_c18 bl[18] br[18] wl[83] vdd gnd cell_6t
Xbit_r84_c18 bl[18] br[18] wl[84] vdd gnd cell_6t
Xbit_r85_c18 bl[18] br[18] wl[85] vdd gnd cell_6t
Xbit_r86_c18 bl[18] br[18] wl[86] vdd gnd cell_6t
Xbit_r87_c18 bl[18] br[18] wl[87] vdd gnd cell_6t
Xbit_r88_c18 bl[18] br[18] wl[88] vdd gnd cell_6t
Xbit_r89_c18 bl[18] br[18] wl[89] vdd gnd cell_6t
Xbit_r90_c18 bl[18] br[18] wl[90] vdd gnd cell_6t
Xbit_r91_c18 bl[18] br[18] wl[91] vdd gnd cell_6t
Xbit_r92_c18 bl[18] br[18] wl[92] vdd gnd cell_6t
Xbit_r93_c18 bl[18] br[18] wl[93] vdd gnd cell_6t
Xbit_r94_c18 bl[18] br[18] wl[94] vdd gnd cell_6t
Xbit_r95_c18 bl[18] br[18] wl[95] vdd gnd cell_6t
Xbit_r96_c18 bl[18] br[18] wl[96] vdd gnd cell_6t
Xbit_r97_c18 bl[18] br[18] wl[97] vdd gnd cell_6t
Xbit_r98_c18 bl[18] br[18] wl[98] vdd gnd cell_6t
Xbit_r99_c18 bl[18] br[18] wl[99] vdd gnd cell_6t
Xbit_r100_c18 bl[18] br[18] wl[100] vdd gnd cell_6t
Xbit_r101_c18 bl[18] br[18] wl[101] vdd gnd cell_6t
Xbit_r102_c18 bl[18] br[18] wl[102] vdd gnd cell_6t
Xbit_r103_c18 bl[18] br[18] wl[103] vdd gnd cell_6t
Xbit_r104_c18 bl[18] br[18] wl[104] vdd gnd cell_6t
Xbit_r105_c18 bl[18] br[18] wl[105] vdd gnd cell_6t
Xbit_r106_c18 bl[18] br[18] wl[106] vdd gnd cell_6t
Xbit_r107_c18 bl[18] br[18] wl[107] vdd gnd cell_6t
Xbit_r108_c18 bl[18] br[18] wl[108] vdd gnd cell_6t
Xbit_r109_c18 bl[18] br[18] wl[109] vdd gnd cell_6t
Xbit_r110_c18 bl[18] br[18] wl[110] vdd gnd cell_6t
Xbit_r111_c18 bl[18] br[18] wl[111] vdd gnd cell_6t
Xbit_r112_c18 bl[18] br[18] wl[112] vdd gnd cell_6t
Xbit_r113_c18 bl[18] br[18] wl[113] vdd gnd cell_6t
Xbit_r114_c18 bl[18] br[18] wl[114] vdd gnd cell_6t
Xbit_r115_c18 bl[18] br[18] wl[115] vdd gnd cell_6t
Xbit_r116_c18 bl[18] br[18] wl[116] vdd gnd cell_6t
Xbit_r117_c18 bl[18] br[18] wl[117] vdd gnd cell_6t
Xbit_r118_c18 bl[18] br[18] wl[118] vdd gnd cell_6t
Xbit_r119_c18 bl[18] br[18] wl[119] vdd gnd cell_6t
Xbit_r120_c18 bl[18] br[18] wl[120] vdd gnd cell_6t
Xbit_r121_c18 bl[18] br[18] wl[121] vdd gnd cell_6t
Xbit_r122_c18 bl[18] br[18] wl[122] vdd gnd cell_6t
Xbit_r123_c18 bl[18] br[18] wl[123] vdd gnd cell_6t
Xbit_r124_c18 bl[18] br[18] wl[124] vdd gnd cell_6t
Xbit_r125_c18 bl[18] br[18] wl[125] vdd gnd cell_6t
Xbit_r126_c18 bl[18] br[18] wl[126] vdd gnd cell_6t
Xbit_r127_c18 bl[18] br[18] wl[127] vdd gnd cell_6t
Xbit_r128_c18 bl[18] br[18] wl[128] vdd gnd cell_6t
Xbit_r129_c18 bl[18] br[18] wl[129] vdd gnd cell_6t
Xbit_r130_c18 bl[18] br[18] wl[130] vdd gnd cell_6t
Xbit_r131_c18 bl[18] br[18] wl[131] vdd gnd cell_6t
Xbit_r132_c18 bl[18] br[18] wl[132] vdd gnd cell_6t
Xbit_r133_c18 bl[18] br[18] wl[133] vdd gnd cell_6t
Xbit_r134_c18 bl[18] br[18] wl[134] vdd gnd cell_6t
Xbit_r135_c18 bl[18] br[18] wl[135] vdd gnd cell_6t
Xbit_r136_c18 bl[18] br[18] wl[136] vdd gnd cell_6t
Xbit_r137_c18 bl[18] br[18] wl[137] vdd gnd cell_6t
Xbit_r138_c18 bl[18] br[18] wl[138] vdd gnd cell_6t
Xbit_r139_c18 bl[18] br[18] wl[139] vdd gnd cell_6t
Xbit_r140_c18 bl[18] br[18] wl[140] vdd gnd cell_6t
Xbit_r141_c18 bl[18] br[18] wl[141] vdd gnd cell_6t
Xbit_r142_c18 bl[18] br[18] wl[142] vdd gnd cell_6t
Xbit_r143_c18 bl[18] br[18] wl[143] vdd gnd cell_6t
Xbit_r144_c18 bl[18] br[18] wl[144] vdd gnd cell_6t
Xbit_r145_c18 bl[18] br[18] wl[145] vdd gnd cell_6t
Xbit_r146_c18 bl[18] br[18] wl[146] vdd gnd cell_6t
Xbit_r147_c18 bl[18] br[18] wl[147] vdd gnd cell_6t
Xbit_r148_c18 bl[18] br[18] wl[148] vdd gnd cell_6t
Xbit_r149_c18 bl[18] br[18] wl[149] vdd gnd cell_6t
Xbit_r150_c18 bl[18] br[18] wl[150] vdd gnd cell_6t
Xbit_r151_c18 bl[18] br[18] wl[151] vdd gnd cell_6t
Xbit_r152_c18 bl[18] br[18] wl[152] vdd gnd cell_6t
Xbit_r153_c18 bl[18] br[18] wl[153] vdd gnd cell_6t
Xbit_r154_c18 bl[18] br[18] wl[154] vdd gnd cell_6t
Xbit_r155_c18 bl[18] br[18] wl[155] vdd gnd cell_6t
Xbit_r156_c18 bl[18] br[18] wl[156] vdd gnd cell_6t
Xbit_r157_c18 bl[18] br[18] wl[157] vdd gnd cell_6t
Xbit_r158_c18 bl[18] br[18] wl[158] vdd gnd cell_6t
Xbit_r159_c18 bl[18] br[18] wl[159] vdd gnd cell_6t
Xbit_r160_c18 bl[18] br[18] wl[160] vdd gnd cell_6t
Xbit_r161_c18 bl[18] br[18] wl[161] vdd gnd cell_6t
Xbit_r162_c18 bl[18] br[18] wl[162] vdd gnd cell_6t
Xbit_r163_c18 bl[18] br[18] wl[163] vdd gnd cell_6t
Xbit_r164_c18 bl[18] br[18] wl[164] vdd gnd cell_6t
Xbit_r165_c18 bl[18] br[18] wl[165] vdd gnd cell_6t
Xbit_r166_c18 bl[18] br[18] wl[166] vdd gnd cell_6t
Xbit_r167_c18 bl[18] br[18] wl[167] vdd gnd cell_6t
Xbit_r168_c18 bl[18] br[18] wl[168] vdd gnd cell_6t
Xbit_r169_c18 bl[18] br[18] wl[169] vdd gnd cell_6t
Xbit_r170_c18 bl[18] br[18] wl[170] vdd gnd cell_6t
Xbit_r171_c18 bl[18] br[18] wl[171] vdd gnd cell_6t
Xbit_r172_c18 bl[18] br[18] wl[172] vdd gnd cell_6t
Xbit_r173_c18 bl[18] br[18] wl[173] vdd gnd cell_6t
Xbit_r174_c18 bl[18] br[18] wl[174] vdd gnd cell_6t
Xbit_r175_c18 bl[18] br[18] wl[175] vdd gnd cell_6t
Xbit_r176_c18 bl[18] br[18] wl[176] vdd gnd cell_6t
Xbit_r177_c18 bl[18] br[18] wl[177] vdd gnd cell_6t
Xbit_r178_c18 bl[18] br[18] wl[178] vdd gnd cell_6t
Xbit_r179_c18 bl[18] br[18] wl[179] vdd gnd cell_6t
Xbit_r180_c18 bl[18] br[18] wl[180] vdd gnd cell_6t
Xbit_r181_c18 bl[18] br[18] wl[181] vdd gnd cell_6t
Xbit_r182_c18 bl[18] br[18] wl[182] vdd gnd cell_6t
Xbit_r183_c18 bl[18] br[18] wl[183] vdd gnd cell_6t
Xbit_r184_c18 bl[18] br[18] wl[184] vdd gnd cell_6t
Xbit_r185_c18 bl[18] br[18] wl[185] vdd gnd cell_6t
Xbit_r186_c18 bl[18] br[18] wl[186] vdd gnd cell_6t
Xbit_r187_c18 bl[18] br[18] wl[187] vdd gnd cell_6t
Xbit_r188_c18 bl[18] br[18] wl[188] vdd gnd cell_6t
Xbit_r189_c18 bl[18] br[18] wl[189] vdd gnd cell_6t
Xbit_r190_c18 bl[18] br[18] wl[190] vdd gnd cell_6t
Xbit_r191_c18 bl[18] br[18] wl[191] vdd gnd cell_6t
Xbit_r192_c18 bl[18] br[18] wl[192] vdd gnd cell_6t
Xbit_r193_c18 bl[18] br[18] wl[193] vdd gnd cell_6t
Xbit_r194_c18 bl[18] br[18] wl[194] vdd gnd cell_6t
Xbit_r195_c18 bl[18] br[18] wl[195] vdd gnd cell_6t
Xbit_r196_c18 bl[18] br[18] wl[196] vdd gnd cell_6t
Xbit_r197_c18 bl[18] br[18] wl[197] vdd gnd cell_6t
Xbit_r198_c18 bl[18] br[18] wl[198] vdd gnd cell_6t
Xbit_r199_c18 bl[18] br[18] wl[199] vdd gnd cell_6t
Xbit_r200_c18 bl[18] br[18] wl[200] vdd gnd cell_6t
Xbit_r201_c18 bl[18] br[18] wl[201] vdd gnd cell_6t
Xbit_r202_c18 bl[18] br[18] wl[202] vdd gnd cell_6t
Xbit_r203_c18 bl[18] br[18] wl[203] vdd gnd cell_6t
Xbit_r204_c18 bl[18] br[18] wl[204] vdd gnd cell_6t
Xbit_r205_c18 bl[18] br[18] wl[205] vdd gnd cell_6t
Xbit_r206_c18 bl[18] br[18] wl[206] vdd gnd cell_6t
Xbit_r207_c18 bl[18] br[18] wl[207] vdd gnd cell_6t
Xbit_r208_c18 bl[18] br[18] wl[208] vdd gnd cell_6t
Xbit_r209_c18 bl[18] br[18] wl[209] vdd gnd cell_6t
Xbit_r210_c18 bl[18] br[18] wl[210] vdd gnd cell_6t
Xbit_r211_c18 bl[18] br[18] wl[211] vdd gnd cell_6t
Xbit_r212_c18 bl[18] br[18] wl[212] vdd gnd cell_6t
Xbit_r213_c18 bl[18] br[18] wl[213] vdd gnd cell_6t
Xbit_r214_c18 bl[18] br[18] wl[214] vdd gnd cell_6t
Xbit_r215_c18 bl[18] br[18] wl[215] vdd gnd cell_6t
Xbit_r216_c18 bl[18] br[18] wl[216] vdd gnd cell_6t
Xbit_r217_c18 bl[18] br[18] wl[217] vdd gnd cell_6t
Xbit_r218_c18 bl[18] br[18] wl[218] vdd gnd cell_6t
Xbit_r219_c18 bl[18] br[18] wl[219] vdd gnd cell_6t
Xbit_r220_c18 bl[18] br[18] wl[220] vdd gnd cell_6t
Xbit_r221_c18 bl[18] br[18] wl[221] vdd gnd cell_6t
Xbit_r222_c18 bl[18] br[18] wl[222] vdd gnd cell_6t
Xbit_r223_c18 bl[18] br[18] wl[223] vdd gnd cell_6t
Xbit_r224_c18 bl[18] br[18] wl[224] vdd gnd cell_6t
Xbit_r225_c18 bl[18] br[18] wl[225] vdd gnd cell_6t
Xbit_r226_c18 bl[18] br[18] wl[226] vdd gnd cell_6t
Xbit_r227_c18 bl[18] br[18] wl[227] vdd gnd cell_6t
Xbit_r228_c18 bl[18] br[18] wl[228] vdd gnd cell_6t
Xbit_r229_c18 bl[18] br[18] wl[229] vdd gnd cell_6t
Xbit_r230_c18 bl[18] br[18] wl[230] vdd gnd cell_6t
Xbit_r231_c18 bl[18] br[18] wl[231] vdd gnd cell_6t
Xbit_r232_c18 bl[18] br[18] wl[232] vdd gnd cell_6t
Xbit_r233_c18 bl[18] br[18] wl[233] vdd gnd cell_6t
Xbit_r234_c18 bl[18] br[18] wl[234] vdd gnd cell_6t
Xbit_r235_c18 bl[18] br[18] wl[235] vdd gnd cell_6t
Xbit_r236_c18 bl[18] br[18] wl[236] vdd gnd cell_6t
Xbit_r237_c18 bl[18] br[18] wl[237] vdd gnd cell_6t
Xbit_r238_c18 bl[18] br[18] wl[238] vdd gnd cell_6t
Xbit_r239_c18 bl[18] br[18] wl[239] vdd gnd cell_6t
Xbit_r240_c18 bl[18] br[18] wl[240] vdd gnd cell_6t
Xbit_r241_c18 bl[18] br[18] wl[241] vdd gnd cell_6t
Xbit_r242_c18 bl[18] br[18] wl[242] vdd gnd cell_6t
Xbit_r243_c18 bl[18] br[18] wl[243] vdd gnd cell_6t
Xbit_r244_c18 bl[18] br[18] wl[244] vdd gnd cell_6t
Xbit_r245_c18 bl[18] br[18] wl[245] vdd gnd cell_6t
Xbit_r246_c18 bl[18] br[18] wl[246] vdd gnd cell_6t
Xbit_r247_c18 bl[18] br[18] wl[247] vdd gnd cell_6t
Xbit_r248_c18 bl[18] br[18] wl[248] vdd gnd cell_6t
Xbit_r249_c18 bl[18] br[18] wl[249] vdd gnd cell_6t
Xbit_r250_c18 bl[18] br[18] wl[250] vdd gnd cell_6t
Xbit_r251_c18 bl[18] br[18] wl[251] vdd gnd cell_6t
Xbit_r252_c18 bl[18] br[18] wl[252] vdd gnd cell_6t
Xbit_r253_c18 bl[18] br[18] wl[253] vdd gnd cell_6t
Xbit_r254_c18 bl[18] br[18] wl[254] vdd gnd cell_6t
Xbit_r255_c18 bl[18] br[18] wl[255] vdd gnd cell_6t
Xbit_r0_c19 bl[19] br[19] wl[0] vdd gnd cell_6t
Xbit_r1_c19 bl[19] br[19] wl[1] vdd gnd cell_6t
Xbit_r2_c19 bl[19] br[19] wl[2] vdd gnd cell_6t
Xbit_r3_c19 bl[19] br[19] wl[3] vdd gnd cell_6t
Xbit_r4_c19 bl[19] br[19] wl[4] vdd gnd cell_6t
Xbit_r5_c19 bl[19] br[19] wl[5] vdd gnd cell_6t
Xbit_r6_c19 bl[19] br[19] wl[6] vdd gnd cell_6t
Xbit_r7_c19 bl[19] br[19] wl[7] vdd gnd cell_6t
Xbit_r8_c19 bl[19] br[19] wl[8] vdd gnd cell_6t
Xbit_r9_c19 bl[19] br[19] wl[9] vdd gnd cell_6t
Xbit_r10_c19 bl[19] br[19] wl[10] vdd gnd cell_6t
Xbit_r11_c19 bl[19] br[19] wl[11] vdd gnd cell_6t
Xbit_r12_c19 bl[19] br[19] wl[12] vdd gnd cell_6t
Xbit_r13_c19 bl[19] br[19] wl[13] vdd gnd cell_6t
Xbit_r14_c19 bl[19] br[19] wl[14] vdd gnd cell_6t
Xbit_r15_c19 bl[19] br[19] wl[15] vdd gnd cell_6t
Xbit_r16_c19 bl[19] br[19] wl[16] vdd gnd cell_6t
Xbit_r17_c19 bl[19] br[19] wl[17] vdd gnd cell_6t
Xbit_r18_c19 bl[19] br[19] wl[18] vdd gnd cell_6t
Xbit_r19_c19 bl[19] br[19] wl[19] vdd gnd cell_6t
Xbit_r20_c19 bl[19] br[19] wl[20] vdd gnd cell_6t
Xbit_r21_c19 bl[19] br[19] wl[21] vdd gnd cell_6t
Xbit_r22_c19 bl[19] br[19] wl[22] vdd gnd cell_6t
Xbit_r23_c19 bl[19] br[19] wl[23] vdd gnd cell_6t
Xbit_r24_c19 bl[19] br[19] wl[24] vdd gnd cell_6t
Xbit_r25_c19 bl[19] br[19] wl[25] vdd gnd cell_6t
Xbit_r26_c19 bl[19] br[19] wl[26] vdd gnd cell_6t
Xbit_r27_c19 bl[19] br[19] wl[27] vdd gnd cell_6t
Xbit_r28_c19 bl[19] br[19] wl[28] vdd gnd cell_6t
Xbit_r29_c19 bl[19] br[19] wl[29] vdd gnd cell_6t
Xbit_r30_c19 bl[19] br[19] wl[30] vdd gnd cell_6t
Xbit_r31_c19 bl[19] br[19] wl[31] vdd gnd cell_6t
Xbit_r32_c19 bl[19] br[19] wl[32] vdd gnd cell_6t
Xbit_r33_c19 bl[19] br[19] wl[33] vdd gnd cell_6t
Xbit_r34_c19 bl[19] br[19] wl[34] vdd gnd cell_6t
Xbit_r35_c19 bl[19] br[19] wl[35] vdd gnd cell_6t
Xbit_r36_c19 bl[19] br[19] wl[36] vdd gnd cell_6t
Xbit_r37_c19 bl[19] br[19] wl[37] vdd gnd cell_6t
Xbit_r38_c19 bl[19] br[19] wl[38] vdd gnd cell_6t
Xbit_r39_c19 bl[19] br[19] wl[39] vdd gnd cell_6t
Xbit_r40_c19 bl[19] br[19] wl[40] vdd gnd cell_6t
Xbit_r41_c19 bl[19] br[19] wl[41] vdd gnd cell_6t
Xbit_r42_c19 bl[19] br[19] wl[42] vdd gnd cell_6t
Xbit_r43_c19 bl[19] br[19] wl[43] vdd gnd cell_6t
Xbit_r44_c19 bl[19] br[19] wl[44] vdd gnd cell_6t
Xbit_r45_c19 bl[19] br[19] wl[45] vdd gnd cell_6t
Xbit_r46_c19 bl[19] br[19] wl[46] vdd gnd cell_6t
Xbit_r47_c19 bl[19] br[19] wl[47] vdd gnd cell_6t
Xbit_r48_c19 bl[19] br[19] wl[48] vdd gnd cell_6t
Xbit_r49_c19 bl[19] br[19] wl[49] vdd gnd cell_6t
Xbit_r50_c19 bl[19] br[19] wl[50] vdd gnd cell_6t
Xbit_r51_c19 bl[19] br[19] wl[51] vdd gnd cell_6t
Xbit_r52_c19 bl[19] br[19] wl[52] vdd gnd cell_6t
Xbit_r53_c19 bl[19] br[19] wl[53] vdd gnd cell_6t
Xbit_r54_c19 bl[19] br[19] wl[54] vdd gnd cell_6t
Xbit_r55_c19 bl[19] br[19] wl[55] vdd gnd cell_6t
Xbit_r56_c19 bl[19] br[19] wl[56] vdd gnd cell_6t
Xbit_r57_c19 bl[19] br[19] wl[57] vdd gnd cell_6t
Xbit_r58_c19 bl[19] br[19] wl[58] vdd gnd cell_6t
Xbit_r59_c19 bl[19] br[19] wl[59] vdd gnd cell_6t
Xbit_r60_c19 bl[19] br[19] wl[60] vdd gnd cell_6t
Xbit_r61_c19 bl[19] br[19] wl[61] vdd gnd cell_6t
Xbit_r62_c19 bl[19] br[19] wl[62] vdd gnd cell_6t
Xbit_r63_c19 bl[19] br[19] wl[63] vdd gnd cell_6t
Xbit_r64_c19 bl[19] br[19] wl[64] vdd gnd cell_6t
Xbit_r65_c19 bl[19] br[19] wl[65] vdd gnd cell_6t
Xbit_r66_c19 bl[19] br[19] wl[66] vdd gnd cell_6t
Xbit_r67_c19 bl[19] br[19] wl[67] vdd gnd cell_6t
Xbit_r68_c19 bl[19] br[19] wl[68] vdd gnd cell_6t
Xbit_r69_c19 bl[19] br[19] wl[69] vdd gnd cell_6t
Xbit_r70_c19 bl[19] br[19] wl[70] vdd gnd cell_6t
Xbit_r71_c19 bl[19] br[19] wl[71] vdd gnd cell_6t
Xbit_r72_c19 bl[19] br[19] wl[72] vdd gnd cell_6t
Xbit_r73_c19 bl[19] br[19] wl[73] vdd gnd cell_6t
Xbit_r74_c19 bl[19] br[19] wl[74] vdd gnd cell_6t
Xbit_r75_c19 bl[19] br[19] wl[75] vdd gnd cell_6t
Xbit_r76_c19 bl[19] br[19] wl[76] vdd gnd cell_6t
Xbit_r77_c19 bl[19] br[19] wl[77] vdd gnd cell_6t
Xbit_r78_c19 bl[19] br[19] wl[78] vdd gnd cell_6t
Xbit_r79_c19 bl[19] br[19] wl[79] vdd gnd cell_6t
Xbit_r80_c19 bl[19] br[19] wl[80] vdd gnd cell_6t
Xbit_r81_c19 bl[19] br[19] wl[81] vdd gnd cell_6t
Xbit_r82_c19 bl[19] br[19] wl[82] vdd gnd cell_6t
Xbit_r83_c19 bl[19] br[19] wl[83] vdd gnd cell_6t
Xbit_r84_c19 bl[19] br[19] wl[84] vdd gnd cell_6t
Xbit_r85_c19 bl[19] br[19] wl[85] vdd gnd cell_6t
Xbit_r86_c19 bl[19] br[19] wl[86] vdd gnd cell_6t
Xbit_r87_c19 bl[19] br[19] wl[87] vdd gnd cell_6t
Xbit_r88_c19 bl[19] br[19] wl[88] vdd gnd cell_6t
Xbit_r89_c19 bl[19] br[19] wl[89] vdd gnd cell_6t
Xbit_r90_c19 bl[19] br[19] wl[90] vdd gnd cell_6t
Xbit_r91_c19 bl[19] br[19] wl[91] vdd gnd cell_6t
Xbit_r92_c19 bl[19] br[19] wl[92] vdd gnd cell_6t
Xbit_r93_c19 bl[19] br[19] wl[93] vdd gnd cell_6t
Xbit_r94_c19 bl[19] br[19] wl[94] vdd gnd cell_6t
Xbit_r95_c19 bl[19] br[19] wl[95] vdd gnd cell_6t
Xbit_r96_c19 bl[19] br[19] wl[96] vdd gnd cell_6t
Xbit_r97_c19 bl[19] br[19] wl[97] vdd gnd cell_6t
Xbit_r98_c19 bl[19] br[19] wl[98] vdd gnd cell_6t
Xbit_r99_c19 bl[19] br[19] wl[99] vdd gnd cell_6t
Xbit_r100_c19 bl[19] br[19] wl[100] vdd gnd cell_6t
Xbit_r101_c19 bl[19] br[19] wl[101] vdd gnd cell_6t
Xbit_r102_c19 bl[19] br[19] wl[102] vdd gnd cell_6t
Xbit_r103_c19 bl[19] br[19] wl[103] vdd gnd cell_6t
Xbit_r104_c19 bl[19] br[19] wl[104] vdd gnd cell_6t
Xbit_r105_c19 bl[19] br[19] wl[105] vdd gnd cell_6t
Xbit_r106_c19 bl[19] br[19] wl[106] vdd gnd cell_6t
Xbit_r107_c19 bl[19] br[19] wl[107] vdd gnd cell_6t
Xbit_r108_c19 bl[19] br[19] wl[108] vdd gnd cell_6t
Xbit_r109_c19 bl[19] br[19] wl[109] vdd gnd cell_6t
Xbit_r110_c19 bl[19] br[19] wl[110] vdd gnd cell_6t
Xbit_r111_c19 bl[19] br[19] wl[111] vdd gnd cell_6t
Xbit_r112_c19 bl[19] br[19] wl[112] vdd gnd cell_6t
Xbit_r113_c19 bl[19] br[19] wl[113] vdd gnd cell_6t
Xbit_r114_c19 bl[19] br[19] wl[114] vdd gnd cell_6t
Xbit_r115_c19 bl[19] br[19] wl[115] vdd gnd cell_6t
Xbit_r116_c19 bl[19] br[19] wl[116] vdd gnd cell_6t
Xbit_r117_c19 bl[19] br[19] wl[117] vdd gnd cell_6t
Xbit_r118_c19 bl[19] br[19] wl[118] vdd gnd cell_6t
Xbit_r119_c19 bl[19] br[19] wl[119] vdd gnd cell_6t
Xbit_r120_c19 bl[19] br[19] wl[120] vdd gnd cell_6t
Xbit_r121_c19 bl[19] br[19] wl[121] vdd gnd cell_6t
Xbit_r122_c19 bl[19] br[19] wl[122] vdd gnd cell_6t
Xbit_r123_c19 bl[19] br[19] wl[123] vdd gnd cell_6t
Xbit_r124_c19 bl[19] br[19] wl[124] vdd gnd cell_6t
Xbit_r125_c19 bl[19] br[19] wl[125] vdd gnd cell_6t
Xbit_r126_c19 bl[19] br[19] wl[126] vdd gnd cell_6t
Xbit_r127_c19 bl[19] br[19] wl[127] vdd gnd cell_6t
Xbit_r128_c19 bl[19] br[19] wl[128] vdd gnd cell_6t
Xbit_r129_c19 bl[19] br[19] wl[129] vdd gnd cell_6t
Xbit_r130_c19 bl[19] br[19] wl[130] vdd gnd cell_6t
Xbit_r131_c19 bl[19] br[19] wl[131] vdd gnd cell_6t
Xbit_r132_c19 bl[19] br[19] wl[132] vdd gnd cell_6t
Xbit_r133_c19 bl[19] br[19] wl[133] vdd gnd cell_6t
Xbit_r134_c19 bl[19] br[19] wl[134] vdd gnd cell_6t
Xbit_r135_c19 bl[19] br[19] wl[135] vdd gnd cell_6t
Xbit_r136_c19 bl[19] br[19] wl[136] vdd gnd cell_6t
Xbit_r137_c19 bl[19] br[19] wl[137] vdd gnd cell_6t
Xbit_r138_c19 bl[19] br[19] wl[138] vdd gnd cell_6t
Xbit_r139_c19 bl[19] br[19] wl[139] vdd gnd cell_6t
Xbit_r140_c19 bl[19] br[19] wl[140] vdd gnd cell_6t
Xbit_r141_c19 bl[19] br[19] wl[141] vdd gnd cell_6t
Xbit_r142_c19 bl[19] br[19] wl[142] vdd gnd cell_6t
Xbit_r143_c19 bl[19] br[19] wl[143] vdd gnd cell_6t
Xbit_r144_c19 bl[19] br[19] wl[144] vdd gnd cell_6t
Xbit_r145_c19 bl[19] br[19] wl[145] vdd gnd cell_6t
Xbit_r146_c19 bl[19] br[19] wl[146] vdd gnd cell_6t
Xbit_r147_c19 bl[19] br[19] wl[147] vdd gnd cell_6t
Xbit_r148_c19 bl[19] br[19] wl[148] vdd gnd cell_6t
Xbit_r149_c19 bl[19] br[19] wl[149] vdd gnd cell_6t
Xbit_r150_c19 bl[19] br[19] wl[150] vdd gnd cell_6t
Xbit_r151_c19 bl[19] br[19] wl[151] vdd gnd cell_6t
Xbit_r152_c19 bl[19] br[19] wl[152] vdd gnd cell_6t
Xbit_r153_c19 bl[19] br[19] wl[153] vdd gnd cell_6t
Xbit_r154_c19 bl[19] br[19] wl[154] vdd gnd cell_6t
Xbit_r155_c19 bl[19] br[19] wl[155] vdd gnd cell_6t
Xbit_r156_c19 bl[19] br[19] wl[156] vdd gnd cell_6t
Xbit_r157_c19 bl[19] br[19] wl[157] vdd gnd cell_6t
Xbit_r158_c19 bl[19] br[19] wl[158] vdd gnd cell_6t
Xbit_r159_c19 bl[19] br[19] wl[159] vdd gnd cell_6t
Xbit_r160_c19 bl[19] br[19] wl[160] vdd gnd cell_6t
Xbit_r161_c19 bl[19] br[19] wl[161] vdd gnd cell_6t
Xbit_r162_c19 bl[19] br[19] wl[162] vdd gnd cell_6t
Xbit_r163_c19 bl[19] br[19] wl[163] vdd gnd cell_6t
Xbit_r164_c19 bl[19] br[19] wl[164] vdd gnd cell_6t
Xbit_r165_c19 bl[19] br[19] wl[165] vdd gnd cell_6t
Xbit_r166_c19 bl[19] br[19] wl[166] vdd gnd cell_6t
Xbit_r167_c19 bl[19] br[19] wl[167] vdd gnd cell_6t
Xbit_r168_c19 bl[19] br[19] wl[168] vdd gnd cell_6t
Xbit_r169_c19 bl[19] br[19] wl[169] vdd gnd cell_6t
Xbit_r170_c19 bl[19] br[19] wl[170] vdd gnd cell_6t
Xbit_r171_c19 bl[19] br[19] wl[171] vdd gnd cell_6t
Xbit_r172_c19 bl[19] br[19] wl[172] vdd gnd cell_6t
Xbit_r173_c19 bl[19] br[19] wl[173] vdd gnd cell_6t
Xbit_r174_c19 bl[19] br[19] wl[174] vdd gnd cell_6t
Xbit_r175_c19 bl[19] br[19] wl[175] vdd gnd cell_6t
Xbit_r176_c19 bl[19] br[19] wl[176] vdd gnd cell_6t
Xbit_r177_c19 bl[19] br[19] wl[177] vdd gnd cell_6t
Xbit_r178_c19 bl[19] br[19] wl[178] vdd gnd cell_6t
Xbit_r179_c19 bl[19] br[19] wl[179] vdd gnd cell_6t
Xbit_r180_c19 bl[19] br[19] wl[180] vdd gnd cell_6t
Xbit_r181_c19 bl[19] br[19] wl[181] vdd gnd cell_6t
Xbit_r182_c19 bl[19] br[19] wl[182] vdd gnd cell_6t
Xbit_r183_c19 bl[19] br[19] wl[183] vdd gnd cell_6t
Xbit_r184_c19 bl[19] br[19] wl[184] vdd gnd cell_6t
Xbit_r185_c19 bl[19] br[19] wl[185] vdd gnd cell_6t
Xbit_r186_c19 bl[19] br[19] wl[186] vdd gnd cell_6t
Xbit_r187_c19 bl[19] br[19] wl[187] vdd gnd cell_6t
Xbit_r188_c19 bl[19] br[19] wl[188] vdd gnd cell_6t
Xbit_r189_c19 bl[19] br[19] wl[189] vdd gnd cell_6t
Xbit_r190_c19 bl[19] br[19] wl[190] vdd gnd cell_6t
Xbit_r191_c19 bl[19] br[19] wl[191] vdd gnd cell_6t
Xbit_r192_c19 bl[19] br[19] wl[192] vdd gnd cell_6t
Xbit_r193_c19 bl[19] br[19] wl[193] vdd gnd cell_6t
Xbit_r194_c19 bl[19] br[19] wl[194] vdd gnd cell_6t
Xbit_r195_c19 bl[19] br[19] wl[195] vdd gnd cell_6t
Xbit_r196_c19 bl[19] br[19] wl[196] vdd gnd cell_6t
Xbit_r197_c19 bl[19] br[19] wl[197] vdd gnd cell_6t
Xbit_r198_c19 bl[19] br[19] wl[198] vdd gnd cell_6t
Xbit_r199_c19 bl[19] br[19] wl[199] vdd gnd cell_6t
Xbit_r200_c19 bl[19] br[19] wl[200] vdd gnd cell_6t
Xbit_r201_c19 bl[19] br[19] wl[201] vdd gnd cell_6t
Xbit_r202_c19 bl[19] br[19] wl[202] vdd gnd cell_6t
Xbit_r203_c19 bl[19] br[19] wl[203] vdd gnd cell_6t
Xbit_r204_c19 bl[19] br[19] wl[204] vdd gnd cell_6t
Xbit_r205_c19 bl[19] br[19] wl[205] vdd gnd cell_6t
Xbit_r206_c19 bl[19] br[19] wl[206] vdd gnd cell_6t
Xbit_r207_c19 bl[19] br[19] wl[207] vdd gnd cell_6t
Xbit_r208_c19 bl[19] br[19] wl[208] vdd gnd cell_6t
Xbit_r209_c19 bl[19] br[19] wl[209] vdd gnd cell_6t
Xbit_r210_c19 bl[19] br[19] wl[210] vdd gnd cell_6t
Xbit_r211_c19 bl[19] br[19] wl[211] vdd gnd cell_6t
Xbit_r212_c19 bl[19] br[19] wl[212] vdd gnd cell_6t
Xbit_r213_c19 bl[19] br[19] wl[213] vdd gnd cell_6t
Xbit_r214_c19 bl[19] br[19] wl[214] vdd gnd cell_6t
Xbit_r215_c19 bl[19] br[19] wl[215] vdd gnd cell_6t
Xbit_r216_c19 bl[19] br[19] wl[216] vdd gnd cell_6t
Xbit_r217_c19 bl[19] br[19] wl[217] vdd gnd cell_6t
Xbit_r218_c19 bl[19] br[19] wl[218] vdd gnd cell_6t
Xbit_r219_c19 bl[19] br[19] wl[219] vdd gnd cell_6t
Xbit_r220_c19 bl[19] br[19] wl[220] vdd gnd cell_6t
Xbit_r221_c19 bl[19] br[19] wl[221] vdd gnd cell_6t
Xbit_r222_c19 bl[19] br[19] wl[222] vdd gnd cell_6t
Xbit_r223_c19 bl[19] br[19] wl[223] vdd gnd cell_6t
Xbit_r224_c19 bl[19] br[19] wl[224] vdd gnd cell_6t
Xbit_r225_c19 bl[19] br[19] wl[225] vdd gnd cell_6t
Xbit_r226_c19 bl[19] br[19] wl[226] vdd gnd cell_6t
Xbit_r227_c19 bl[19] br[19] wl[227] vdd gnd cell_6t
Xbit_r228_c19 bl[19] br[19] wl[228] vdd gnd cell_6t
Xbit_r229_c19 bl[19] br[19] wl[229] vdd gnd cell_6t
Xbit_r230_c19 bl[19] br[19] wl[230] vdd gnd cell_6t
Xbit_r231_c19 bl[19] br[19] wl[231] vdd gnd cell_6t
Xbit_r232_c19 bl[19] br[19] wl[232] vdd gnd cell_6t
Xbit_r233_c19 bl[19] br[19] wl[233] vdd gnd cell_6t
Xbit_r234_c19 bl[19] br[19] wl[234] vdd gnd cell_6t
Xbit_r235_c19 bl[19] br[19] wl[235] vdd gnd cell_6t
Xbit_r236_c19 bl[19] br[19] wl[236] vdd gnd cell_6t
Xbit_r237_c19 bl[19] br[19] wl[237] vdd gnd cell_6t
Xbit_r238_c19 bl[19] br[19] wl[238] vdd gnd cell_6t
Xbit_r239_c19 bl[19] br[19] wl[239] vdd gnd cell_6t
Xbit_r240_c19 bl[19] br[19] wl[240] vdd gnd cell_6t
Xbit_r241_c19 bl[19] br[19] wl[241] vdd gnd cell_6t
Xbit_r242_c19 bl[19] br[19] wl[242] vdd gnd cell_6t
Xbit_r243_c19 bl[19] br[19] wl[243] vdd gnd cell_6t
Xbit_r244_c19 bl[19] br[19] wl[244] vdd gnd cell_6t
Xbit_r245_c19 bl[19] br[19] wl[245] vdd gnd cell_6t
Xbit_r246_c19 bl[19] br[19] wl[246] vdd gnd cell_6t
Xbit_r247_c19 bl[19] br[19] wl[247] vdd gnd cell_6t
Xbit_r248_c19 bl[19] br[19] wl[248] vdd gnd cell_6t
Xbit_r249_c19 bl[19] br[19] wl[249] vdd gnd cell_6t
Xbit_r250_c19 bl[19] br[19] wl[250] vdd gnd cell_6t
Xbit_r251_c19 bl[19] br[19] wl[251] vdd gnd cell_6t
Xbit_r252_c19 bl[19] br[19] wl[252] vdd gnd cell_6t
Xbit_r253_c19 bl[19] br[19] wl[253] vdd gnd cell_6t
Xbit_r254_c19 bl[19] br[19] wl[254] vdd gnd cell_6t
Xbit_r255_c19 bl[19] br[19] wl[255] vdd gnd cell_6t
Xbit_r0_c20 bl[20] br[20] wl[0] vdd gnd cell_6t
Xbit_r1_c20 bl[20] br[20] wl[1] vdd gnd cell_6t
Xbit_r2_c20 bl[20] br[20] wl[2] vdd gnd cell_6t
Xbit_r3_c20 bl[20] br[20] wl[3] vdd gnd cell_6t
Xbit_r4_c20 bl[20] br[20] wl[4] vdd gnd cell_6t
Xbit_r5_c20 bl[20] br[20] wl[5] vdd gnd cell_6t
Xbit_r6_c20 bl[20] br[20] wl[6] vdd gnd cell_6t
Xbit_r7_c20 bl[20] br[20] wl[7] vdd gnd cell_6t
Xbit_r8_c20 bl[20] br[20] wl[8] vdd gnd cell_6t
Xbit_r9_c20 bl[20] br[20] wl[9] vdd gnd cell_6t
Xbit_r10_c20 bl[20] br[20] wl[10] vdd gnd cell_6t
Xbit_r11_c20 bl[20] br[20] wl[11] vdd gnd cell_6t
Xbit_r12_c20 bl[20] br[20] wl[12] vdd gnd cell_6t
Xbit_r13_c20 bl[20] br[20] wl[13] vdd gnd cell_6t
Xbit_r14_c20 bl[20] br[20] wl[14] vdd gnd cell_6t
Xbit_r15_c20 bl[20] br[20] wl[15] vdd gnd cell_6t
Xbit_r16_c20 bl[20] br[20] wl[16] vdd gnd cell_6t
Xbit_r17_c20 bl[20] br[20] wl[17] vdd gnd cell_6t
Xbit_r18_c20 bl[20] br[20] wl[18] vdd gnd cell_6t
Xbit_r19_c20 bl[20] br[20] wl[19] vdd gnd cell_6t
Xbit_r20_c20 bl[20] br[20] wl[20] vdd gnd cell_6t
Xbit_r21_c20 bl[20] br[20] wl[21] vdd gnd cell_6t
Xbit_r22_c20 bl[20] br[20] wl[22] vdd gnd cell_6t
Xbit_r23_c20 bl[20] br[20] wl[23] vdd gnd cell_6t
Xbit_r24_c20 bl[20] br[20] wl[24] vdd gnd cell_6t
Xbit_r25_c20 bl[20] br[20] wl[25] vdd gnd cell_6t
Xbit_r26_c20 bl[20] br[20] wl[26] vdd gnd cell_6t
Xbit_r27_c20 bl[20] br[20] wl[27] vdd gnd cell_6t
Xbit_r28_c20 bl[20] br[20] wl[28] vdd gnd cell_6t
Xbit_r29_c20 bl[20] br[20] wl[29] vdd gnd cell_6t
Xbit_r30_c20 bl[20] br[20] wl[30] vdd gnd cell_6t
Xbit_r31_c20 bl[20] br[20] wl[31] vdd gnd cell_6t
Xbit_r32_c20 bl[20] br[20] wl[32] vdd gnd cell_6t
Xbit_r33_c20 bl[20] br[20] wl[33] vdd gnd cell_6t
Xbit_r34_c20 bl[20] br[20] wl[34] vdd gnd cell_6t
Xbit_r35_c20 bl[20] br[20] wl[35] vdd gnd cell_6t
Xbit_r36_c20 bl[20] br[20] wl[36] vdd gnd cell_6t
Xbit_r37_c20 bl[20] br[20] wl[37] vdd gnd cell_6t
Xbit_r38_c20 bl[20] br[20] wl[38] vdd gnd cell_6t
Xbit_r39_c20 bl[20] br[20] wl[39] vdd gnd cell_6t
Xbit_r40_c20 bl[20] br[20] wl[40] vdd gnd cell_6t
Xbit_r41_c20 bl[20] br[20] wl[41] vdd gnd cell_6t
Xbit_r42_c20 bl[20] br[20] wl[42] vdd gnd cell_6t
Xbit_r43_c20 bl[20] br[20] wl[43] vdd gnd cell_6t
Xbit_r44_c20 bl[20] br[20] wl[44] vdd gnd cell_6t
Xbit_r45_c20 bl[20] br[20] wl[45] vdd gnd cell_6t
Xbit_r46_c20 bl[20] br[20] wl[46] vdd gnd cell_6t
Xbit_r47_c20 bl[20] br[20] wl[47] vdd gnd cell_6t
Xbit_r48_c20 bl[20] br[20] wl[48] vdd gnd cell_6t
Xbit_r49_c20 bl[20] br[20] wl[49] vdd gnd cell_6t
Xbit_r50_c20 bl[20] br[20] wl[50] vdd gnd cell_6t
Xbit_r51_c20 bl[20] br[20] wl[51] vdd gnd cell_6t
Xbit_r52_c20 bl[20] br[20] wl[52] vdd gnd cell_6t
Xbit_r53_c20 bl[20] br[20] wl[53] vdd gnd cell_6t
Xbit_r54_c20 bl[20] br[20] wl[54] vdd gnd cell_6t
Xbit_r55_c20 bl[20] br[20] wl[55] vdd gnd cell_6t
Xbit_r56_c20 bl[20] br[20] wl[56] vdd gnd cell_6t
Xbit_r57_c20 bl[20] br[20] wl[57] vdd gnd cell_6t
Xbit_r58_c20 bl[20] br[20] wl[58] vdd gnd cell_6t
Xbit_r59_c20 bl[20] br[20] wl[59] vdd gnd cell_6t
Xbit_r60_c20 bl[20] br[20] wl[60] vdd gnd cell_6t
Xbit_r61_c20 bl[20] br[20] wl[61] vdd gnd cell_6t
Xbit_r62_c20 bl[20] br[20] wl[62] vdd gnd cell_6t
Xbit_r63_c20 bl[20] br[20] wl[63] vdd gnd cell_6t
Xbit_r64_c20 bl[20] br[20] wl[64] vdd gnd cell_6t
Xbit_r65_c20 bl[20] br[20] wl[65] vdd gnd cell_6t
Xbit_r66_c20 bl[20] br[20] wl[66] vdd gnd cell_6t
Xbit_r67_c20 bl[20] br[20] wl[67] vdd gnd cell_6t
Xbit_r68_c20 bl[20] br[20] wl[68] vdd gnd cell_6t
Xbit_r69_c20 bl[20] br[20] wl[69] vdd gnd cell_6t
Xbit_r70_c20 bl[20] br[20] wl[70] vdd gnd cell_6t
Xbit_r71_c20 bl[20] br[20] wl[71] vdd gnd cell_6t
Xbit_r72_c20 bl[20] br[20] wl[72] vdd gnd cell_6t
Xbit_r73_c20 bl[20] br[20] wl[73] vdd gnd cell_6t
Xbit_r74_c20 bl[20] br[20] wl[74] vdd gnd cell_6t
Xbit_r75_c20 bl[20] br[20] wl[75] vdd gnd cell_6t
Xbit_r76_c20 bl[20] br[20] wl[76] vdd gnd cell_6t
Xbit_r77_c20 bl[20] br[20] wl[77] vdd gnd cell_6t
Xbit_r78_c20 bl[20] br[20] wl[78] vdd gnd cell_6t
Xbit_r79_c20 bl[20] br[20] wl[79] vdd gnd cell_6t
Xbit_r80_c20 bl[20] br[20] wl[80] vdd gnd cell_6t
Xbit_r81_c20 bl[20] br[20] wl[81] vdd gnd cell_6t
Xbit_r82_c20 bl[20] br[20] wl[82] vdd gnd cell_6t
Xbit_r83_c20 bl[20] br[20] wl[83] vdd gnd cell_6t
Xbit_r84_c20 bl[20] br[20] wl[84] vdd gnd cell_6t
Xbit_r85_c20 bl[20] br[20] wl[85] vdd gnd cell_6t
Xbit_r86_c20 bl[20] br[20] wl[86] vdd gnd cell_6t
Xbit_r87_c20 bl[20] br[20] wl[87] vdd gnd cell_6t
Xbit_r88_c20 bl[20] br[20] wl[88] vdd gnd cell_6t
Xbit_r89_c20 bl[20] br[20] wl[89] vdd gnd cell_6t
Xbit_r90_c20 bl[20] br[20] wl[90] vdd gnd cell_6t
Xbit_r91_c20 bl[20] br[20] wl[91] vdd gnd cell_6t
Xbit_r92_c20 bl[20] br[20] wl[92] vdd gnd cell_6t
Xbit_r93_c20 bl[20] br[20] wl[93] vdd gnd cell_6t
Xbit_r94_c20 bl[20] br[20] wl[94] vdd gnd cell_6t
Xbit_r95_c20 bl[20] br[20] wl[95] vdd gnd cell_6t
Xbit_r96_c20 bl[20] br[20] wl[96] vdd gnd cell_6t
Xbit_r97_c20 bl[20] br[20] wl[97] vdd gnd cell_6t
Xbit_r98_c20 bl[20] br[20] wl[98] vdd gnd cell_6t
Xbit_r99_c20 bl[20] br[20] wl[99] vdd gnd cell_6t
Xbit_r100_c20 bl[20] br[20] wl[100] vdd gnd cell_6t
Xbit_r101_c20 bl[20] br[20] wl[101] vdd gnd cell_6t
Xbit_r102_c20 bl[20] br[20] wl[102] vdd gnd cell_6t
Xbit_r103_c20 bl[20] br[20] wl[103] vdd gnd cell_6t
Xbit_r104_c20 bl[20] br[20] wl[104] vdd gnd cell_6t
Xbit_r105_c20 bl[20] br[20] wl[105] vdd gnd cell_6t
Xbit_r106_c20 bl[20] br[20] wl[106] vdd gnd cell_6t
Xbit_r107_c20 bl[20] br[20] wl[107] vdd gnd cell_6t
Xbit_r108_c20 bl[20] br[20] wl[108] vdd gnd cell_6t
Xbit_r109_c20 bl[20] br[20] wl[109] vdd gnd cell_6t
Xbit_r110_c20 bl[20] br[20] wl[110] vdd gnd cell_6t
Xbit_r111_c20 bl[20] br[20] wl[111] vdd gnd cell_6t
Xbit_r112_c20 bl[20] br[20] wl[112] vdd gnd cell_6t
Xbit_r113_c20 bl[20] br[20] wl[113] vdd gnd cell_6t
Xbit_r114_c20 bl[20] br[20] wl[114] vdd gnd cell_6t
Xbit_r115_c20 bl[20] br[20] wl[115] vdd gnd cell_6t
Xbit_r116_c20 bl[20] br[20] wl[116] vdd gnd cell_6t
Xbit_r117_c20 bl[20] br[20] wl[117] vdd gnd cell_6t
Xbit_r118_c20 bl[20] br[20] wl[118] vdd gnd cell_6t
Xbit_r119_c20 bl[20] br[20] wl[119] vdd gnd cell_6t
Xbit_r120_c20 bl[20] br[20] wl[120] vdd gnd cell_6t
Xbit_r121_c20 bl[20] br[20] wl[121] vdd gnd cell_6t
Xbit_r122_c20 bl[20] br[20] wl[122] vdd gnd cell_6t
Xbit_r123_c20 bl[20] br[20] wl[123] vdd gnd cell_6t
Xbit_r124_c20 bl[20] br[20] wl[124] vdd gnd cell_6t
Xbit_r125_c20 bl[20] br[20] wl[125] vdd gnd cell_6t
Xbit_r126_c20 bl[20] br[20] wl[126] vdd gnd cell_6t
Xbit_r127_c20 bl[20] br[20] wl[127] vdd gnd cell_6t
Xbit_r128_c20 bl[20] br[20] wl[128] vdd gnd cell_6t
Xbit_r129_c20 bl[20] br[20] wl[129] vdd gnd cell_6t
Xbit_r130_c20 bl[20] br[20] wl[130] vdd gnd cell_6t
Xbit_r131_c20 bl[20] br[20] wl[131] vdd gnd cell_6t
Xbit_r132_c20 bl[20] br[20] wl[132] vdd gnd cell_6t
Xbit_r133_c20 bl[20] br[20] wl[133] vdd gnd cell_6t
Xbit_r134_c20 bl[20] br[20] wl[134] vdd gnd cell_6t
Xbit_r135_c20 bl[20] br[20] wl[135] vdd gnd cell_6t
Xbit_r136_c20 bl[20] br[20] wl[136] vdd gnd cell_6t
Xbit_r137_c20 bl[20] br[20] wl[137] vdd gnd cell_6t
Xbit_r138_c20 bl[20] br[20] wl[138] vdd gnd cell_6t
Xbit_r139_c20 bl[20] br[20] wl[139] vdd gnd cell_6t
Xbit_r140_c20 bl[20] br[20] wl[140] vdd gnd cell_6t
Xbit_r141_c20 bl[20] br[20] wl[141] vdd gnd cell_6t
Xbit_r142_c20 bl[20] br[20] wl[142] vdd gnd cell_6t
Xbit_r143_c20 bl[20] br[20] wl[143] vdd gnd cell_6t
Xbit_r144_c20 bl[20] br[20] wl[144] vdd gnd cell_6t
Xbit_r145_c20 bl[20] br[20] wl[145] vdd gnd cell_6t
Xbit_r146_c20 bl[20] br[20] wl[146] vdd gnd cell_6t
Xbit_r147_c20 bl[20] br[20] wl[147] vdd gnd cell_6t
Xbit_r148_c20 bl[20] br[20] wl[148] vdd gnd cell_6t
Xbit_r149_c20 bl[20] br[20] wl[149] vdd gnd cell_6t
Xbit_r150_c20 bl[20] br[20] wl[150] vdd gnd cell_6t
Xbit_r151_c20 bl[20] br[20] wl[151] vdd gnd cell_6t
Xbit_r152_c20 bl[20] br[20] wl[152] vdd gnd cell_6t
Xbit_r153_c20 bl[20] br[20] wl[153] vdd gnd cell_6t
Xbit_r154_c20 bl[20] br[20] wl[154] vdd gnd cell_6t
Xbit_r155_c20 bl[20] br[20] wl[155] vdd gnd cell_6t
Xbit_r156_c20 bl[20] br[20] wl[156] vdd gnd cell_6t
Xbit_r157_c20 bl[20] br[20] wl[157] vdd gnd cell_6t
Xbit_r158_c20 bl[20] br[20] wl[158] vdd gnd cell_6t
Xbit_r159_c20 bl[20] br[20] wl[159] vdd gnd cell_6t
Xbit_r160_c20 bl[20] br[20] wl[160] vdd gnd cell_6t
Xbit_r161_c20 bl[20] br[20] wl[161] vdd gnd cell_6t
Xbit_r162_c20 bl[20] br[20] wl[162] vdd gnd cell_6t
Xbit_r163_c20 bl[20] br[20] wl[163] vdd gnd cell_6t
Xbit_r164_c20 bl[20] br[20] wl[164] vdd gnd cell_6t
Xbit_r165_c20 bl[20] br[20] wl[165] vdd gnd cell_6t
Xbit_r166_c20 bl[20] br[20] wl[166] vdd gnd cell_6t
Xbit_r167_c20 bl[20] br[20] wl[167] vdd gnd cell_6t
Xbit_r168_c20 bl[20] br[20] wl[168] vdd gnd cell_6t
Xbit_r169_c20 bl[20] br[20] wl[169] vdd gnd cell_6t
Xbit_r170_c20 bl[20] br[20] wl[170] vdd gnd cell_6t
Xbit_r171_c20 bl[20] br[20] wl[171] vdd gnd cell_6t
Xbit_r172_c20 bl[20] br[20] wl[172] vdd gnd cell_6t
Xbit_r173_c20 bl[20] br[20] wl[173] vdd gnd cell_6t
Xbit_r174_c20 bl[20] br[20] wl[174] vdd gnd cell_6t
Xbit_r175_c20 bl[20] br[20] wl[175] vdd gnd cell_6t
Xbit_r176_c20 bl[20] br[20] wl[176] vdd gnd cell_6t
Xbit_r177_c20 bl[20] br[20] wl[177] vdd gnd cell_6t
Xbit_r178_c20 bl[20] br[20] wl[178] vdd gnd cell_6t
Xbit_r179_c20 bl[20] br[20] wl[179] vdd gnd cell_6t
Xbit_r180_c20 bl[20] br[20] wl[180] vdd gnd cell_6t
Xbit_r181_c20 bl[20] br[20] wl[181] vdd gnd cell_6t
Xbit_r182_c20 bl[20] br[20] wl[182] vdd gnd cell_6t
Xbit_r183_c20 bl[20] br[20] wl[183] vdd gnd cell_6t
Xbit_r184_c20 bl[20] br[20] wl[184] vdd gnd cell_6t
Xbit_r185_c20 bl[20] br[20] wl[185] vdd gnd cell_6t
Xbit_r186_c20 bl[20] br[20] wl[186] vdd gnd cell_6t
Xbit_r187_c20 bl[20] br[20] wl[187] vdd gnd cell_6t
Xbit_r188_c20 bl[20] br[20] wl[188] vdd gnd cell_6t
Xbit_r189_c20 bl[20] br[20] wl[189] vdd gnd cell_6t
Xbit_r190_c20 bl[20] br[20] wl[190] vdd gnd cell_6t
Xbit_r191_c20 bl[20] br[20] wl[191] vdd gnd cell_6t
Xbit_r192_c20 bl[20] br[20] wl[192] vdd gnd cell_6t
Xbit_r193_c20 bl[20] br[20] wl[193] vdd gnd cell_6t
Xbit_r194_c20 bl[20] br[20] wl[194] vdd gnd cell_6t
Xbit_r195_c20 bl[20] br[20] wl[195] vdd gnd cell_6t
Xbit_r196_c20 bl[20] br[20] wl[196] vdd gnd cell_6t
Xbit_r197_c20 bl[20] br[20] wl[197] vdd gnd cell_6t
Xbit_r198_c20 bl[20] br[20] wl[198] vdd gnd cell_6t
Xbit_r199_c20 bl[20] br[20] wl[199] vdd gnd cell_6t
Xbit_r200_c20 bl[20] br[20] wl[200] vdd gnd cell_6t
Xbit_r201_c20 bl[20] br[20] wl[201] vdd gnd cell_6t
Xbit_r202_c20 bl[20] br[20] wl[202] vdd gnd cell_6t
Xbit_r203_c20 bl[20] br[20] wl[203] vdd gnd cell_6t
Xbit_r204_c20 bl[20] br[20] wl[204] vdd gnd cell_6t
Xbit_r205_c20 bl[20] br[20] wl[205] vdd gnd cell_6t
Xbit_r206_c20 bl[20] br[20] wl[206] vdd gnd cell_6t
Xbit_r207_c20 bl[20] br[20] wl[207] vdd gnd cell_6t
Xbit_r208_c20 bl[20] br[20] wl[208] vdd gnd cell_6t
Xbit_r209_c20 bl[20] br[20] wl[209] vdd gnd cell_6t
Xbit_r210_c20 bl[20] br[20] wl[210] vdd gnd cell_6t
Xbit_r211_c20 bl[20] br[20] wl[211] vdd gnd cell_6t
Xbit_r212_c20 bl[20] br[20] wl[212] vdd gnd cell_6t
Xbit_r213_c20 bl[20] br[20] wl[213] vdd gnd cell_6t
Xbit_r214_c20 bl[20] br[20] wl[214] vdd gnd cell_6t
Xbit_r215_c20 bl[20] br[20] wl[215] vdd gnd cell_6t
Xbit_r216_c20 bl[20] br[20] wl[216] vdd gnd cell_6t
Xbit_r217_c20 bl[20] br[20] wl[217] vdd gnd cell_6t
Xbit_r218_c20 bl[20] br[20] wl[218] vdd gnd cell_6t
Xbit_r219_c20 bl[20] br[20] wl[219] vdd gnd cell_6t
Xbit_r220_c20 bl[20] br[20] wl[220] vdd gnd cell_6t
Xbit_r221_c20 bl[20] br[20] wl[221] vdd gnd cell_6t
Xbit_r222_c20 bl[20] br[20] wl[222] vdd gnd cell_6t
Xbit_r223_c20 bl[20] br[20] wl[223] vdd gnd cell_6t
Xbit_r224_c20 bl[20] br[20] wl[224] vdd gnd cell_6t
Xbit_r225_c20 bl[20] br[20] wl[225] vdd gnd cell_6t
Xbit_r226_c20 bl[20] br[20] wl[226] vdd gnd cell_6t
Xbit_r227_c20 bl[20] br[20] wl[227] vdd gnd cell_6t
Xbit_r228_c20 bl[20] br[20] wl[228] vdd gnd cell_6t
Xbit_r229_c20 bl[20] br[20] wl[229] vdd gnd cell_6t
Xbit_r230_c20 bl[20] br[20] wl[230] vdd gnd cell_6t
Xbit_r231_c20 bl[20] br[20] wl[231] vdd gnd cell_6t
Xbit_r232_c20 bl[20] br[20] wl[232] vdd gnd cell_6t
Xbit_r233_c20 bl[20] br[20] wl[233] vdd gnd cell_6t
Xbit_r234_c20 bl[20] br[20] wl[234] vdd gnd cell_6t
Xbit_r235_c20 bl[20] br[20] wl[235] vdd gnd cell_6t
Xbit_r236_c20 bl[20] br[20] wl[236] vdd gnd cell_6t
Xbit_r237_c20 bl[20] br[20] wl[237] vdd gnd cell_6t
Xbit_r238_c20 bl[20] br[20] wl[238] vdd gnd cell_6t
Xbit_r239_c20 bl[20] br[20] wl[239] vdd gnd cell_6t
Xbit_r240_c20 bl[20] br[20] wl[240] vdd gnd cell_6t
Xbit_r241_c20 bl[20] br[20] wl[241] vdd gnd cell_6t
Xbit_r242_c20 bl[20] br[20] wl[242] vdd gnd cell_6t
Xbit_r243_c20 bl[20] br[20] wl[243] vdd gnd cell_6t
Xbit_r244_c20 bl[20] br[20] wl[244] vdd gnd cell_6t
Xbit_r245_c20 bl[20] br[20] wl[245] vdd gnd cell_6t
Xbit_r246_c20 bl[20] br[20] wl[246] vdd gnd cell_6t
Xbit_r247_c20 bl[20] br[20] wl[247] vdd gnd cell_6t
Xbit_r248_c20 bl[20] br[20] wl[248] vdd gnd cell_6t
Xbit_r249_c20 bl[20] br[20] wl[249] vdd gnd cell_6t
Xbit_r250_c20 bl[20] br[20] wl[250] vdd gnd cell_6t
Xbit_r251_c20 bl[20] br[20] wl[251] vdd gnd cell_6t
Xbit_r252_c20 bl[20] br[20] wl[252] vdd gnd cell_6t
Xbit_r253_c20 bl[20] br[20] wl[253] vdd gnd cell_6t
Xbit_r254_c20 bl[20] br[20] wl[254] vdd gnd cell_6t
Xbit_r255_c20 bl[20] br[20] wl[255] vdd gnd cell_6t
Xbit_r0_c21 bl[21] br[21] wl[0] vdd gnd cell_6t
Xbit_r1_c21 bl[21] br[21] wl[1] vdd gnd cell_6t
Xbit_r2_c21 bl[21] br[21] wl[2] vdd gnd cell_6t
Xbit_r3_c21 bl[21] br[21] wl[3] vdd gnd cell_6t
Xbit_r4_c21 bl[21] br[21] wl[4] vdd gnd cell_6t
Xbit_r5_c21 bl[21] br[21] wl[5] vdd gnd cell_6t
Xbit_r6_c21 bl[21] br[21] wl[6] vdd gnd cell_6t
Xbit_r7_c21 bl[21] br[21] wl[7] vdd gnd cell_6t
Xbit_r8_c21 bl[21] br[21] wl[8] vdd gnd cell_6t
Xbit_r9_c21 bl[21] br[21] wl[9] vdd gnd cell_6t
Xbit_r10_c21 bl[21] br[21] wl[10] vdd gnd cell_6t
Xbit_r11_c21 bl[21] br[21] wl[11] vdd gnd cell_6t
Xbit_r12_c21 bl[21] br[21] wl[12] vdd gnd cell_6t
Xbit_r13_c21 bl[21] br[21] wl[13] vdd gnd cell_6t
Xbit_r14_c21 bl[21] br[21] wl[14] vdd gnd cell_6t
Xbit_r15_c21 bl[21] br[21] wl[15] vdd gnd cell_6t
Xbit_r16_c21 bl[21] br[21] wl[16] vdd gnd cell_6t
Xbit_r17_c21 bl[21] br[21] wl[17] vdd gnd cell_6t
Xbit_r18_c21 bl[21] br[21] wl[18] vdd gnd cell_6t
Xbit_r19_c21 bl[21] br[21] wl[19] vdd gnd cell_6t
Xbit_r20_c21 bl[21] br[21] wl[20] vdd gnd cell_6t
Xbit_r21_c21 bl[21] br[21] wl[21] vdd gnd cell_6t
Xbit_r22_c21 bl[21] br[21] wl[22] vdd gnd cell_6t
Xbit_r23_c21 bl[21] br[21] wl[23] vdd gnd cell_6t
Xbit_r24_c21 bl[21] br[21] wl[24] vdd gnd cell_6t
Xbit_r25_c21 bl[21] br[21] wl[25] vdd gnd cell_6t
Xbit_r26_c21 bl[21] br[21] wl[26] vdd gnd cell_6t
Xbit_r27_c21 bl[21] br[21] wl[27] vdd gnd cell_6t
Xbit_r28_c21 bl[21] br[21] wl[28] vdd gnd cell_6t
Xbit_r29_c21 bl[21] br[21] wl[29] vdd gnd cell_6t
Xbit_r30_c21 bl[21] br[21] wl[30] vdd gnd cell_6t
Xbit_r31_c21 bl[21] br[21] wl[31] vdd gnd cell_6t
Xbit_r32_c21 bl[21] br[21] wl[32] vdd gnd cell_6t
Xbit_r33_c21 bl[21] br[21] wl[33] vdd gnd cell_6t
Xbit_r34_c21 bl[21] br[21] wl[34] vdd gnd cell_6t
Xbit_r35_c21 bl[21] br[21] wl[35] vdd gnd cell_6t
Xbit_r36_c21 bl[21] br[21] wl[36] vdd gnd cell_6t
Xbit_r37_c21 bl[21] br[21] wl[37] vdd gnd cell_6t
Xbit_r38_c21 bl[21] br[21] wl[38] vdd gnd cell_6t
Xbit_r39_c21 bl[21] br[21] wl[39] vdd gnd cell_6t
Xbit_r40_c21 bl[21] br[21] wl[40] vdd gnd cell_6t
Xbit_r41_c21 bl[21] br[21] wl[41] vdd gnd cell_6t
Xbit_r42_c21 bl[21] br[21] wl[42] vdd gnd cell_6t
Xbit_r43_c21 bl[21] br[21] wl[43] vdd gnd cell_6t
Xbit_r44_c21 bl[21] br[21] wl[44] vdd gnd cell_6t
Xbit_r45_c21 bl[21] br[21] wl[45] vdd gnd cell_6t
Xbit_r46_c21 bl[21] br[21] wl[46] vdd gnd cell_6t
Xbit_r47_c21 bl[21] br[21] wl[47] vdd gnd cell_6t
Xbit_r48_c21 bl[21] br[21] wl[48] vdd gnd cell_6t
Xbit_r49_c21 bl[21] br[21] wl[49] vdd gnd cell_6t
Xbit_r50_c21 bl[21] br[21] wl[50] vdd gnd cell_6t
Xbit_r51_c21 bl[21] br[21] wl[51] vdd gnd cell_6t
Xbit_r52_c21 bl[21] br[21] wl[52] vdd gnd cell_6t
Xbit_r53_c21 bl[21] br[21] wl[53] vdd gnd cell_6t
Xbit_r54_c21 bl[21] br[21] wl[54] vdd gnd cell_6t
Xbit_r55_c21 bl[21] br[21] wl[55] vdd gnd cell_6t
Xbit_r56_c21 bl[21] br[21] wl[56] vdd gnd cell_6t
Xbit_r57_c21 bl[21] br[21] wl[57] vdd gnd cell_6t
Xbit_r58_c21 bl[21] br[21] wl[58] vdd gnd cell_6t
Xbit_r59_c21 bl[21] br[21] wl[59] vdd gnd cell_6t
Xbit_r60_c21 bl[21] br[21] wl[60] vdd gnd cell_6t
Xbit_r61_c21 bl[21] br[21] wl[61] vdd gnd cell_6t
Xbit_r62_c21 bl[21] br[21] wl[62] vdd gnd cell_6t
Xbit_r63_c21 bl[21] br[21] wl[63] vdd gnd cell_6t
Xbit_r64_c21 bl[21] br[21] wl[64] vdd gnd cell_6t
Xbit_r65_c21 bl[21] br[21] wl[65] vdd gnd cell_6t
Xbit_r66_c21 bl[21] br[21] wl[66] vdd gnd cell_6t
Xbit_r67_c21 bl[21] br[21] wl[67] vdd gnd cell_6t
Xbit_r68_c21 bl[21] br[21] wl[68] vdd gnd cell_6t
Xbit_r69_c21 bl[21] br[21] wl[69] vdd gnd cell_6t
Xbit_r70_c21 bl[21] br[21] wl[70] vdd gnd cell_6t
Xbit_r71_c21 bl[21] br[21] wl[71] vdd gnd cell_6t
Xbit_r72_c21 bl[21] br[21] wl[72] vdd gnd cell_6t
Xbit_r73_c21 bl[21] br[21] wl[73] vdd gnd cell_6t
Xbit_r74_c21 bl[21] br[21] wl[74] vdd gnd cell_6t
Xbit_r75_c21 bl[21] br[21] wl[75] vdd gnd cell_6t
Xbit_r76_c21 bl[21] br[21] wl[76] vdd gnd cell_6t
Xbit_r77_c21 bl[21] br[21] wl[77] vdd gnd cell_6t
Xbit_r78_c21 bl[21] br[21] wl[78] vdd gnd cell_6t
Xbit_r79_c21 bl[21] br[21] wl[79] vdd gnd cell_6t
Xbit_r80_c21 bl[21] br[21] wl[80] vdd gnd cell_6t
Xbit_r81_c21 bl[21] br[21] wl[81] vdd gnd cell_6t
Xbit_r82_c21 bl[21] br[21] wl[82] vdd gnd cell_6t
Xbit_r83_c21 bl[21] br[21] wl[83] vdd gnd cell_6t
Xbit_r84_c21 bl[21] br[21] wl[84] vdd gnd cell_6t
Xbit_r85_c21 bl[21] br[21] wl[85] vdd gnd cell_6t
Xbit_r86_c21 bl[21] br[21] wl[86] vdd gnd cell_6t
Xbit_r87_c21 bl[21] br[21] wl[87] vdd gnd cell_6t
Xbit_r88_c21 bl[21] br[21] wl[88] vdd gnd cell_6t
Xbit_r89_c21 bl[21] br[21] wl[89] vdd gnd cell_6t
Xbit_r90_c21 bl[21] br[21] wl[90] vdd gnd cell_6t
Xbit_r91_c21 bl[21] br[21] wl[91] vdd gnd cell_6t
Xbit_r92_c21 bl[21] br[21] wl[92] vdd gnd cell_6t
Xbit_r93_c21 bl[21] br[21] wl[93] vdd gnd cell_6t
Xbit_r94_c21 bl[21] br[21] wl[94] vdd gnd cell_6t
Xbit_r95_c21 bl[21] br[21] wl[95] vdd gnd cell_6t
Xbit_r96_c21 bl[21] br[21] wl[96] vdd gnd cell_6t
Xbit_r97_c21 bl[21] br[21] wl[97] vdd gnd cell_6t
Xbit_r98_c21 bl[21] br[21] wl[98] vdd gnd cell_6t
Xbit_r99_c21 bl[21] br[21] wl[99] vdd gnd cell_6t
Xbit_r100_c21 bl[21] br[21] wl[100] vdd gnd cell_6t
Xbit_r101_c21 bl[21] br[21] wl[101] vdd gnd cell_6t
Xbit_r102_c21 bl[21] br[21] wl[102] vdd gnd cell_6t
Xbit_r103_c21 bl[21] br[21] wl[103] vdd gnd cell_6t
Xbit_r104_c21 bl[21] br[21] wl[104] vdd gnd cell_6t
Xbit_r105_c21 bl[21] br[21] wl[105] vdd gnd cell_6t
Xbit_r106_c21 bl[21] br[21] wl[106] vdd gnd cell_6t
Xbit_r107_c21 bl[21] br[21] wl[107] vdd gnd cell_6t
Xbit_r108_c21 bl[21] br[21] wl[108] vdd gnd cell_6t
Xbit_r109_c21 bl[21] br[21] wl[109] vdd gnd cell_6t
Xbit_r110_c21 bl[21] br[21] wl[110] vdd gnd cell_6t
Xbit_r111_c21 bl[21] br[21] wl[111] vdd gnd cell_6t
Xbit_r112_c21 bl[21] br[21] wl[112] vdd gnd cell_6t
Xbit_r113_c21 bl[21] br[21] wl[113] vdd gnd cell_6t
Xbit_r114_c21 bl[21] br[21] wl[114] vdd gnd cell_6t
Xbit_r115_c21 bl[21] br[21] wl[115] vdd gnd cell_6t
Xbit_r116_c21 bl[21] br[21] wl[116] vdd gnd cell_6t
Xbit_r117_c21 bl[21] br[21] wl[117] vdd gnd cell_6t
Xbit_r118_c21 bl[21] br[21] wl[118] vdd gnd cell_6t
Xbit_r119_c21 bl[21] br[21] wl[119] vdd gnd cell_6t
Xbit_r120_c21 bl[21] br[21] wl[120] vdd gnd cell_6t
Xbit_r121_c21 bl[21] br[21] wl[121] vdd gnd cell_6t
Xbit_r122_c21 bl[21] br[21] wl[122] vdd gnd cell_6t
Xbit_r123_c21 bl[21] br[21] wl[123] vdd gnd cell_6t
Xbit_r124_c21 bl[21] br[21] wl[124] vdd gnd cell_6t
Xbit_r125_c21 bl[21] br[21] wl[125] vdd gnd cell_6t
Xbit_r126_c21 bl[21] br[21] wl[126] vdd gnd cell_6t
Xbit_r127_c21 bl[21] br[21] wl[127] vdd gnd cell_6t
Xbit_r128_c21 bl[21] br[21] wl[128] vdd gnd cell_6t
Xbit_r129_c21 bl[21] br[21] wl[129] vdd gnd cell_6t
Xbit_r130_c21 bl[21] br[21] wl[130] vdd gnd cell_6t
Xbit_r131_c21 bl[21] br[21] wl[131] vdd gnd cell_6t
Xbit_r132_c21 bl[21] br[21] wl[132] vdd gnd cell_6t
Xbit_r133_c21 bl[21] br[21] wl[133] vdd gnd cell_6t
Xbit_r134_c21 bl[21] br[21] wl[134] vdd gnd cell_6t
Xbit_r135_c21 bl[21] br[21] wl[135] vdd gnd cell_6t
Xbit_r136_c21 bl[21] br[21] wl[136] vdd gnd cell_6t
Xbit_r137_c21 bl[21] br[21] wl[137] vdd gnd cell_6t
Xbit_r138_c21 bl[21] br[21] wl[138] vdd gnd cell_6t
Xbit_r139_c21 bl[21] br[21] wl[139] vdd gnd cell_6t
Xbit_r140_c21 bl[21] br[21] wl[140] vdd gnd cell_6t
Xbit_r141_c21 bl[21] br[21] wl[141] vdd gnd cell_6t
Xbit_r142_c21 bl[21] br[21] wl[142] vdd gnd cell_6t
Xbit_r143_c21 bl[21] br[21] wl[143] vdd gnd cell_6t
Xbit_r144_c21 bl[21] br[21] wl[144] vdd gnd cell_6t
Xbit_r145_c21 bl[21] br[21] wl[145] vdd gnd cell_6t
Xbit_r146_c21 bl[21] br[21] wl[146] vdd gnd cell_6t
Xbit_r147_c21 bl[21] br[21] wl[147] vdd gnd cell_6t
Xbit_r148_c21 bl[21] br[21] wl[148] vdd gnd cell_6t
Xbit_r149_c21 bl[21] br[21] wl[149] vdd gnd cell_6t
Xbit_r150_c21 bl[21] br[21] wl[150] vdd gnd cell_6t
Xbit_r151_c21 bl[21] br[21] wl[151] vdd gnd cell_6t
Xbit_r152_c21 bl[21] br[21] wl[152] vdd gnd cell_6t
Xbit_r153_c21 bl[21] br[21] wl[153] vdd gnd cell_6t
Xbit_r154_c21 bl[21] br[21] wl[154] vdd gnd cell_6t
Xbit_r155_c21 bl[21] br[21] wl[155] vdd gnd cell_6t
Xbit_r156_c21 bl[21] br[21] wl[156] vdd gnd cell_6t
Xbit_r157_c21 bl[21] br[21] wl[157] vdd gnd cell_6t
Xbit_r158_c21 bl[21] br[21] wl[158] vdd gnd cell_6t
Xbit_r159_c21 bl[21] br[21] wl[159] vdd gnd cell_6t
Xbit_r160_c21 bl[21] br[21] wl[160] vdd gnd cell_6t
Xbit_r161_c21 bl[21] br[21] wl[161] vdd gnd cell_6t
Xbit_r162_c21 bl[21] br[21] wl[162] vdd gnd cell_6t
Xbit_r163_c21 bl[21] br[21] wl[163] vdd gnd cell_6t
Xbit_r164_c21 bl[21] br[21] wl[164] vdd gnd cell_6t
Xbit_r165_c21 bl[21] br[21] wl[165] vdd gnd cell_6t
Xbit_r166_c21 bl[21] br[21] wl[166] vdd gnd cell_6t
Xbit_r167_c21 bl[21] br[21] wl[167] vdd gnd cell_6t
Xbit_r168_c21 bl[21] br[21] wl[168] vdd gnd cell_6t
Xbit_r169_c21 bl[21] br[21] wl[169] vdd gnd cell_6t
Xbit_r170_c21 bl[21] br[21] wl[170] vdd gnd cell_6t
Xbit_r171_c21 bl[21] br[21] wl[171] vdd gnd cell_6t
Xbit_r172_c21 bl[21] br[21] wl[172] vdd gnd cell_6t
Xbit_r173_c21 bl[21] br[21] wl[173] vdd gnd cell_6t
Xbit_r174_c21 bl[21] br[21] wl[174] vdd gnd cell_6t
Xbit_r175_c21 bl[21] br[21] wl[175] vdd gnd cell_6t
Xbit_r176_c21 bl[21] br[21] wl[176] vdd gnd cell_6t
Xbit_r177_c21 bl[21] br[21] wl[177] vdd gnd cell_6t
Xbit_r178_c21 bl[21] br[21] wl[178] vdd gnd cell_6t
Xbit_r179_c21 bl[21] br[21] wl[179] vdd gnd cell_6t
Xbit_r180_c21 bl[21] br[21] wl[180] vdd gnd cell_6t
Xbit_r181_c21 bl[21] br[21] wl[181] vdd gnd cell_6t
Xbit_r182_c21 bl[21] br[21] wl[182] vdd gnd cell_6t
Xbit_r183_c21 bl[21] br[21] wl[183] vdd gnd cell_6t
Xbit_r184_c21 bl[21] br[21] wl[184] vdd gnd cell_6t
Xbit_r185_c21 bl[21] br[21] wl[185] vdd gnd cell_6t
Xbit_r186_c21 bl[21] br[21] wl[186] vdd gnd cell_6t
Xbit_r187_c21 bl[21] br[21] wl[187] vdd gnd cell_6t
Xbit_r188_c21 bl[21] br[21] wl[188] vdd gnd cell_6t
Xbit_r189_c21 bl[21] br[21] wl[189] vdd gnd cell_6t
Xbit_r190_c21 bl[21] br[21] wl[190] vdd gnd cell_6t
Xbit_r191_c21 bl[21] br[21] wl[191] vdd gnd cell_6t
Xbit_r192_c21 bl[21] br[21] wl[192] vdd gnd cell_6t
Xbit_r193_c21 bl[21] br[21] wl[193] vdd gnd cell_6t
Xbit_r194_c21 bl[21] br[21] wl[194] vdd gnd cell_6t
Xbit_r195_c21 bl[21] br[21] wl[195] vdd gnd cell_6t
Xbit_r196_c21 bl[21] br[21] wl[196] vdd gnd cell_6t
Xbit_r197_c21 bl[21] br[21] wl[197] vdd gnd cell_6t
Xbit_r198_c21 bl[21] br[21] wl[198] vdd gnd cell_6t
Xbit_r199_c21 bl[21] br[21] wl[199] vdd gnd cell_6t
Xbit_r200_c21 bl[21] br[21] wl[200] vdd gnd cell_6t
Xbit_r201_c21 bl[21] br[21] wl[201] vdd gnd cell_6t
Xbit_r202_c21 bl[21] br[21] wl[202] vdd gnd cell_6t
Xbit_r203_c21 bl[21] br[21] wl[203] vdd gnd cell_6t
Xbit_r204_c21 bl[21] br[21] wl[204] vdd gnd cell_6t
Xbit_r205_c21 bl[21] br[21] wl[205] vdd gnd cell_6t
Xbit_r206_c21 bl[21] br[21] wl[206] vdd gnd cell_6t
Xbit_r207_c21 bl[21] br[21] wl[207] vdd gnd cell_6t
Xbit_r208_c21 bl[21] br[21] wl[208] vdd gnd cell_6t
Xbit_r209_c21 bl[21] br[21] wl[209] vdd gnd cell_6t
Xbit_r210_c21 bl[21] br[21] wl[210] vdd gnd cell_6t
Xbit_r211_c21 bl[21] br[21] wl[211] vdd gnd cell_6t
Xbit_r212_c21 bl[21] br[21] wl[212] vdd gnd cell_6t
Xbit_r213_c21 bl[21] br[21] wl[213] vdd gnd cell_6t
Xbit_r214_c21 bl[21] br[21] wl[214] vdd gnd cell_6t
Xbit_r215_c21 bl[21] br[21] wl[215] vdd gnd cell_6t
Xbit_r216_c21 bl[21] br[21] wl[216] vdd gnd cell_6t
Xbit_r217_c21 bl[21] br[21] wl[217] vdd gnd cell_6t
Xbit_r218_c21 bl[21] br[21] wl[218] vdd gnd cell_6t
Xbit_r219_c21 bl[21] br[21] wl[219] vdd gnd cell_6t
Xbit_r220_c21 bl[21] br[21] wl[220] vdd gnd cell_6t
Xbit_r221_c21 bl[21] br[21] wl[221] vdd gnd cell_6t
Xbit_r222_c21 bl[21] br[21] wl[222] vdd gnd cell_6t
Xbit_r223_c21 bl[21] br[21] wl[223] vdd gnd cell_6t
Xbit_r224_c21 bl[21] br[21] wl[224] vdd gnd cell_6t
Xbit_r225_c21 bl[21] br[21] wl[225] vdd gnd cell_6t
Xbit_r226_c21 bl[21] br[21] wl[226] vdd gnd cell_6t
Xbit_r227_c21 bl[21] br[21] wl[227] vdd gnd cell_6t
Xbit_r228_c21 bl[21] br[21] wl[228] vdd gnd cell_6t
Xbit_r229_c21 bl[21] br[21] wl[229] vdd gnd cell_6t
Xbit_r230_c21 bl[21] br[21] wl[230] vdd gnd cell_6t
Xbit_r231_c21 bl[21] br[21] wl[231] vdd gnd cell_6t
Xbit_r232_c21 bl[21] br[21] wl[232] vdd gnd cell_6t
Xbit_r233_c21 bl[21] br[21] wl[233] vdd gnd cell_6t
Xbit_r234_c21 bl[21] br[21] wl[234] vdd gnd cell_6t
Xbit_r235_c21 bl[21] br[21] wl[235] vdd gnd cell_6t
Xbit_r236_c21 bl[21] br[21] wl[236] vdd gnd cell_6t
Xbit_r237_c21 bl[21] br[21] wl[237] vdd gnd cell_6t
Xbit_r238_c21 bl[21] br[21] wl[238] vdd gnd cell_6t
Xbit_r239_c21 bl[21] br[21] wl[239] vdd gnd cell_6t
Xbit_r240_c21 bl[21] br[21] wl[240] vdd gnd cell_6t
Xbit_r241_c21 bl[21] br[21] wl[241] vdd gnd cell_6t
Xbit_r242_c21 bl[21] br[21] wl[242] vdd gnd cell_6t
Xbit_r243_c21 bl[21] br[21] wl[243] vdd gnd cell_6t
Xbit_r244_c21 bl[21] br[21] wl[244] vdd gnd cell_6t
Xbit_r245_c21 bl[21] br[21] wl[245] vdd gnd cell_6t
Xbit_r246_c21 bl[21] br[21] wl[246] vdd gnd cell_6t
Xbit_r247_c21 bl[21] br[21] wl[247] vdd gnd cell_6t
Xbit_r248_c21 bl[21] br[21] wl[248] vdd gnd cell_6t
Xbit_r249_c21 bl[21] br[21] wl[249] vdd gnd cell_6t
Xbit_r250_c21 bl[21] br[21] wl[250] vdd gnd cell_6t
Xbit_r251_c21 bl[21] br[21] wl[251] vdd gnd cell_6t
Xbit_r252_c21 bl[21] br[21] wl[252] vdd gnd cell_6t
Xbit_r253_c21 bl[21] br[21] wl[253] vdd gnd cell_6t
Xbit_r254_c21 bl[21] br[21] wl[254] vdd gnd cell_6t
Xbit_r255_c21 bl[21] br[21] wl[255] vdd gnd cell_6t
Xbit_r0_c22 bl[22] br[22] wl[0] vdd gnd cell_6t
Xbit_r1_c22 bl[22] br[22] wl[1] vdd gnd cell_6t
Xbit_r2_c22 bl[22] br[22] wl[2] vdd gnd cell_6t
Xbit_r3_c22 bl[22] br[22] wl[3] vdd gnd cell_6t
Xbit_r4_c22 bl[22] br[22] wl[4] vdd gnd cell_6t
Xbit_r5_c22 bl[22] br[22] wl[5] vdd gnd cell_6t
Xbit_r6_c22 bl[22] br[22] wl[6] vdd gnd cell_6t
Xbit_r7_c22 bl[22] br[22] wl[7] vdd gnd cell_6t
Xbit_r8_c22 bl[22] br[22] wl[8] vdd gnd cell_6t
Xbit_r9_c22 bl[22] br[22] wl[9] vdd gnd cell_6t
Xbit_r10_c22 bl[22] br[22] wl[10] vdd gnd cell_6t
Xbit_r11_c22 bl[22] br[22] wl[11] vdd gnd cell_6t
Xbit_r12_c22 bl[22] br[22] wl[12] vdd gnd cell_6t
Xbit_r13_c22 bl[22] br[22] wl[13] vdd gnd cell_6t
Xbit_r14_c22 bl[22] br[22] wl[14] vdd gnd cell_6t
Xbit_r15_c22 bl[22] br[22] wl[15] vdd gnd cell_6t
Xbit_r16_c22 bl[22] br[22] wl[16] vdd gnd cell_6t
Xbit_r17_c22 bl[22] br[22] wl[17] vdd gnd cell_6t
Xbit_r18_c22 bl[22] br[22] wl[18] vdd gnd cell_6t
Xbit_r19_c22 bl[22] br[22] wl[19] vdd gnd cell_6t
Xbit_r20_c22 bl[22] br[22] wl[20] vdd gnd cell_6t
Xbit_r21_c22 bl[22] br[22] wl[21] vdd gnd cell_6t
Xbit_r22_c22 bl[22] br[22] wl[22] vdd gnd cell_6t
Xbit_r23_c22 bl[22] br[22] wl[23] vdd gnd cell_6t
Xbit_r24_c22 bl[22] br[22] wl[24] vdd gnd cell_6t
Xbit_r25_c22 bl[22] br[22] wl[25] vdd gnd cell_6t
Xbit_r26_c22 bl[22] br[22] wl[26] vdd gnd cell_6t
Xbit_r27_c22 bl[22] br[22] wl[27] vdd gnd cell_6t
Xbit_r28_c22 bl[22] br[22] wl[28] vdd gnd cell_6t
Xbit_r29_c22 bl[22] br[22] wl[29] vdd gnd cell_6t
Xbit_r30_c22 bl[22] br[22] wl[30] vdd gnd cell_6t
Xbit_r31_c22 bl[22] br[22] wl[31] vdd gnd cell_6t
Xbit_r32_c22 bl[22] br[22] wl[32] vdd gnd cell_6t
Xbit_r33_c22 bl[22] br[22] wl[33] vdd gnd cell_6t
Xbit_r34_c22 bl[22] br[22] wl[34] vdd gnd cell_6t
Xbit_r35_c22 bl[22] br[22] wl[35] vdd gnd cell_6t
Xbit_r36_c22 bl[22] br[22] wl[36] vdd gnd cell_6t
Xbit_r37_c22 bl[22] br[22] wl[37] vdd gnd cell_6t
Xbit_r38_c22 bl[22] br[22] wl[38] vdd gnd cell_6t
Xbit_r39_c22 bl[22] br[22] wl[39] vdd gnd cell_6t
Xbit_r40_c22 bl[22] br[22] wl[40] vdd gnd cell_6t
Xbit_r41_c22 bl[22] br[22] wl[41] vdd gnd cell_6t
Xbit_r42_c22 bl[22] br[22] wl[42] vdd gnd cell_6t
Xbit_r43_c22 bl[22] br[22] wl[43] vdd gnd cell_6t
Xbit_r44_c22 bl[22] br[22] wl[44] vdd gnd cell_6t
Xbit_r45_c22 bl[22] br[22] wl[45] vdd gnd cell_6t
Xbit_r46_c22 bl[22] br[22] wl[46] vdd gnd cell_6t
Xbit_r47_c22 bl[22] br[22] wl[47] vdd gnd cell_6t
Xbit_r48_c22 bl[22] br[22] wl[48] vdd gnd cell_6t
Xbit_r49_c22 bl[22] br[22] wl[49] vdd gnd cell_6t
Xbit_r50_c22 bl[22] br[22] wl[50] vdd gnd cell_6t
Xbit_r51_c22 bl[22] br[22] wl[51] vdd gnd cell_6t
Xbit_r52_c22 bl[22] br[22] wl[52] vdd gnd cell_6t
Xbit_r53_c22 bl[22] br[22] wl[53] vdd gnd cell_6t
Xbit_r54_c22 bl[22] br[22] wl[54] vdd gnd cell_6t
Xbit_r55_c22 bl[22] br[22] wl[55] vdd gnd cell_6t
Xbit_r56_c22 bl[22] br[22] wl[56] vdd gnd cell_6t
Xbit_r57_c22 bl[22] br[22] wl[57] vdd gnd cell_6t
Xbit_r58_c22 bl[22] br[22] wl[58] vdd gnd cell_6t
Xbit_r59_c22 bl[22] br[22] wl[59] vdd gnd cell_6t
Xbit_r60_c22 bl[22] br[22] wl[60] vdd gnd cell_6t
Xbit_r61_c22 bl[22] br[22] wl[61] vdd gnd cell_6t
Xbit_r62_c22 bl[22] br[22] wl[62] vdd gnd cell_6t
Xbit_r63_c22 bl[22] br[22] wl[63] vdd gnd cell_6t
Xbit_r64_c22 bl[22] br[22] wl[64] vdd gnd cell_6t
Xbit_r65_c22 bl[22] br[22] wl[65] vdd gnd cell_6t
Xbit_r66_c22 bl[22] br[22] wl[66] vdd gnd cell_6t
Xbit_r67_c22 bl[22] br[22] wl[67] vdd gnd cell_6t
Xbit_r68_c22 bl[22] br[22] wl[68] vdd gnd cell_6t
Xbit_r69_c22 bl[22] br[22] wl[69] vdd gnd cell_6t
Xbit_r70_c22 bl[22] br[22] wl[70] vdd gnd cell_6t
Xbit_r71_c22 bl[22] br[22] wl[71] vdd gnd cell_6t
Xbit_r72_c22 bl[22] br[22] wl[72] vdd gnd cell_6t
Xbit_r73_c22 bl[22] br[22] wl[73] vdd gnd cell_6t
Xbit_r74_c22 bl[22] br[22] wl[74] vdd gnd cell_6t
Xbit_r75_c22 bl[22] br[22] wl[75] vdd gnd cell_6t
Xbit_r76_c22 bl[22] br[22] wl[76] vdd gnd cell_6t
Xbit_r77_c22 bl[22] br[22] wl[77] vdd gnd cell_6t
Xbit_r78_c22 bl[22] br[22] wl[78] vdd gnd cell_6t
Xbit_r79_c22 bl[22] br[22] wl[79] vdd gnd cell_6t
Xbit_r80_c22 bl[22] br[22] wl[80] vdd gnd cell_6t
Xbit_r81_c22 bl[22] br[22] wl[81] vdd gnd cell_6t
Xbit_r82_c22 bl[22] br[22] wl[82] vdd gnd cell_6t
Xbit_r83_c22 bl[22] br[22] wl[83] vdd gnd cell_6t
Xbit_r84_c22 bl[22] br[22] wl[84] vdd gnd cell_6t
Xbit_r85_c22 bl[22] br[22] wl[85] vdd gnd cell_6t
Xbit_r86_c22 bl[22] br[22] wl[86] vdd gnd cell_6t
Xbit_r87_c22 bl[22] br[22] wl[87] vdd gnd cell_6t
Xbit_r88_c22 bl[22] br[22] wl[88] vdd gnd cell_6t
Xbit_r89_c22 bl[22] br[22] wl[89] vdd gnd cell_6t
Xbit_r90_c22 bl[22] br[22] wl[90] vdd gnd cell_6t
Xbit_r91_c22 bl[22] br[22] wl[91] vdd gnd cell_6t
Xbit_r92_c22 bl[22] br[22] wl[92] vdd gnd cell_6t
Xbit_r93_c22 bl[22] br[22] wl[93] vdd gnd cell_6t
Xbit_r94_c22 bl[22] br[22] wl[94] vdd gnd cell_6t
Xbit_r95_c22 bl[22] br[22] wl[95] vdd gnd cell_6t
Xbit_r96_c22 bl[22] br[22] wl[96] vdd gnd cell_6t
Xbit_r97_c22 bl[22] br[22] wl[97] vdd gnd cell_6t
Xbit_r98_c22 bl[22] br[22] wl[98] vdd gnd cell_6t
Xbit_r99_c22 bl[22] br[22] wl[99] vdd gnd cell_6t
Xbit_r100_c22 bl[22] br[22] wl[100] vdd gnd cell_6t
Xbit_r101_c22 bl[22] br[22] wl[101] vdd gnd cell_6t
Xbit_r102_c22 bl[22] br[22] wl[102] vdd gnd cell_6t
Xbit_r103_c22 bl[22] br[22] wl[103] vdd gnd cell_6t
Xbit_r104_c22 bl[22] br[22] wl[104] vdd gnd cell_6t
Xbit_r105_c22 bl[22] br[22] wl[105] vdd gnd cell_6t
Xbit_r106_c22 bl[22] br[22] wl[106] vdd gnd cell_6t
Xbit_r107_c22 bl[22] br[22] wl[107] vdd gnd cell_6t
Xbit_r108_c22 bl[22] br[22] wl[108] vdd gnd cell_6t
Xbit_r109_c22 bl[22] br[22] wl[109] vdd gnd cell_6t
Xbit_r110_c22 bl[22] br[22] wl[110] vdd gnd cell_6t
Xbit_r111_c22 bl[22] br[22] wl[111] vdd gnd cell_6t
Xbit_r112_c22 bl[22] br[22] wl[112] vdd gnd cell_6t
Xbit_r113_c22 bl[22] br[22] wl[113] vdd gnd cell_6t
Xbit_r114_c22 bl[22] br[22] wl[114] vdd gnd cell_6t
Xbit_r115_c22 bl[22] br[22] wl[115] vdd gnd cell_6t
Xbit_r116_c22 bl[22] br[22] wl[116] vdd gnd cell_6t
Xbit_r117_c22 bl[22] br[22] wl[117] vdd gnd cell_6t
Xbit_r118_c22 bl[22] br[22] wl[118] vdd gnd cell_6t
Xbit_r119_c22 bl[22] br[22] wl[119] vdd gnd cell_6t
Xbit_r120_c22 bl[22] br[22] wl[120] vdd gnd cell_6t
Xbit_r121_c22 bl[22] br[22] wl[121] vdd gnd cell_6t
Xbit_r122_c22 bl[22] br[22] wl[122] vdd gnd cell_6t
Xbit_r123_c22 bl[22] br[22] wl[123] vdd gnd cell_6t
Xbit_r124_c22 bl[22] br[22] wl[124] vdd gnd cell_6t
Xbit_r125_c22 bl[22] br[22] wl[125] vdd gnd cell_6t
Xbit_r126_c22 bl[22] br[22] wl[126] vdd gnd cell_6t
Xbit_r127_c22 bl[22] br[22] wl[127] vdd gnd cell_6t
Xbit_r128_c22 bl[22] br[22] wl[128] vdd gnd cell_6t
Xbit_r129_c22 bl[22] br[22] wl[129] vdd gnd cell_6t
Xbit_r130_c22 bl[22] br[22] wl[130] vdd gnd cell_6t
Xbit_r131_c22 bl[22] br[22] wl[131] vdd gnd cell_6t
Xbit_r132_c22 bl[22] br[22] wl[132] vdd gnd cell_6t
Xbit_r133_c22 bl[22] br[22] wl[133] vdd gnd cell_6t
Xbit_r134_c22 bl[22] br[22] wl[134] vdd gnd cell_6t
Xbit_r135_c22 bl[22] br[22] wl[135] vdd gnd cell_6t
Xbit_r136_c22 bl[22] br[22] wl[136] vdd gnd cell_6t
Xbit_r137_c22 bl[22] br[22] wl[137] vdd gnd cell_6t
Xbit_r138_c22 bl[22] br[22] wl[138] vdd gnd cell_6t
Xbit_r139_c22 bl[22] br[22] wl[139] vdd gnd cell_6t
Xbit_r140_c22 bl[22] br[22] wl[140] vdd gnd cell_6t
Xbit_r141_c22 bl[22] br[22] wl[141] vdd gnd cell_6t
Xbit_r142_c22 bl[22] br[22] wl[142] vdd gnd cell_6t
Xbit_r143_c22 bl[22] br[22] wl[143] vdd gnd cell_6t
Xbit_r144_c22 bl[22] br[22] wl[144] vdd gnd cell_6t
Xbit_r145_c22 bl[22] br[22] wl[145] vdd gnd cell_6t
Xbit_r146_c22 bl[22] br[22] wl[146] vdd gnd cell_6t
Xbit_r147_c22 bl[22] br[22] wl[147] vdd gnd cell_6t
Xbit_r148_c22 bl[22] br[22] wl[148] vdd gnd cell_6t
Xbit_r149_c22 bl[22] br[22] wl[149] vdd gnd cell_6t
Xbit_r150_c22 bl[22] br[22] wl[150] vdd gnd cell_6t
Xbit_r151_c22 bl[22] br[22] wl[151] vdd gnd cell_6t
Xbit_r152_c22 bl[22] br[22] wl[152] vdd gnd cell_6t
Xbit_r153_c22 bl[22] br[22] wl[153] vdd gnd cell_6t
Xbit_r154_c22 bl[22] br[22] wl[154] vdd gnd cell_6t
Xbit_r155_c22 bl[22] br[22] wl[155] vdd gnd cell_6t
Xbit_r156_c22 bl[22] br[22] wl[156] vdd gnd cell_6t
Xbit_r157_c22 bl[22] br[22] wl[157] vdd gnd cell_6t
Xbit_r158_c22 bl[22] br[22] wl[158] vdd gnd cell_6t
Xbit_r159_c22 bl[22] br[22] wl[159] vdd gnd cell_6t
Xbit_r160_c22 bl[22] br[22] wl[160] vdd gnd cell_6t
Xbit_r161_c22 bl[22] br[22] wl[161] vdd gnd cell_6t
Xbit_r162_c22 bl[22] br[22] wl[162] vdd gnd cell_6t
Xbit_r163_c22 bl[22] br[22] wl[163] vdd gnd cell_6t
Xbit_r164_c22 bl[22] br[22] wl[164] vdd gnd cell_6t
Xbit_r165_c22 bl[22] br[22] wl[165] vdd gnd cell_6t
Xbit_r166_c22 bl[22] br[22] wl[166] vdd gnd cell_6t
Xbit_r167_c22 bl[22] br[22] wl[167] vdd gnd cell_6t
Xbit_r168_c22 bl[22] br[22] wl[168] vdd gnd cell_6t
Xbit_r169_c22 bl[22] br[22] wl[169] vdd gnd cell_6t
Xbit_r170_c22 bl[22] br[22] wl[170] vdd gnd cell_6t
Xbit_r171_c22 bl[22] br[22] wl[171] vdd gnd cell_6t
Xbit_r172_c22 bl[22] br[22] wl[172] vdd gnd cell_6t
Xbit_r173_c22 bl[22] br[22] wl[173] vdd gnd cell_6t
Xbit_r174_c22 bl[22] br[22] wl[174] vdd gnd cell_6t
Xbit_r175_c22 bl[22] br[22] wl[175] vdd gnd cell_6t
Xbit_r176_c22 bl[22] br[22] wl[176] vdd gnd cell_6t
Xbit_r177_c22 bl[22] br[22] wl[177] vdd gnd cell_6t
Xbit_r178_c22 bl[22] br[22] wl[178] vdd gnd cell_6t
Xbit_r179_c22 bl[22] br[22] wl[179] vdd gnd cell_6t
Xbit_r180_c22 bl[22] br[22] wl[180] vdd gnd cell_6t
Xbit_r181_c22 bl[22] br[22] wl[181] vdd gnd cell_6t
Xbit_r182_c22 bl[22] br[22] wl[182] vdd gnd cell_6t
Xbit_r183_c22 bl[22] br[22] wl[183] vdd gnd cell_6t
Xbit_r184_c22 bl[22] br[22] wl[184] vdd gnd cell_6t
Xbit_r185_c22 bl[22] br[22] wl[185] vdd gnd cell_6t
Xbit_r186_c22 bl[22] br[22] wl[186] vdd gnd cell_6t
Xbit_r187_c22 bl[22] br[22] wl[187] vdd gnd cell_6t
Xbit_r188_c22 bl[22] br[22] wl[188] vdd gnd cell_6t
Xbit_r189_c22 bl[22] br[22] wl[189] vdd gnd cell_6t
Xbit_r190_c22 bl[22] br[22] wl[190] vdd gnd cell_6t
Xbit_r191_c22 bl[22] br[22] wl[191] vdd gnd cell_6t
Xbit_r192_c22 bl[22] br[22] wl[192] vdd gnd cell_6t
Xbit_r193_c22 bl[22] br[22] wl[193] vdd gnd cell_6t
Xbit_r194_c22 bl[22] br[22] wl[194] vdd gnd cell_6t
Xbit_r195_c22 bl[22] br[22] wl[195] vdd gnd cell_6t
Xbit_r196_c22 bl[22] br[22] wl[196] vdd gnd cell_6t
Xbit_r197_c22 bl[22] br[22] wl[197] vdd gnd cell_6t
Xbit_r198_c22 bl[22] br[22] wl[198] vdd gnd cell_6t
Xbit_r199_c22 bl[22] br[22] wl[199] vdd gnd cell_6t
Xbit_r200_c22 bl[22] br[22] wl[200] vdd gnd cell_6t
Xbit_r201_c22 bl[22] br[22] wl[201] vdd gnd cell_6t
Xbit_r202_c22 bl[22] br[22] wl[202] vdd gnd cell_6t
Xbit_r203_c22 bl[22] br[22] wl[203] vdd gnd cell_6t
Xbit_r204_c22 bl[22] br[22] wl[204] vdd gnd cell_6t
Xbit_r205_c22 bl[22] br[22] wl[205] vdd gnd cell_6t
Xbit_r206_c22 bl[22] br[22] wl[206] vdd gnd cell_6t
Xbit_r207_c22 bl[22] br[22] wl[207] vdd gnd cell_6t
Xbit_r208_c22 bl[22] br[22] wl[208] vdd gnd cell_6t
Xbit_r209_c22 bl[22] br[22] wl[209] vdd gnd cell_6t
Xbit_r210_c22 bl[22] br[22] wl[210] vdd gnd cell_6t
Xbit_r211_c22 bl[22] br[22] wl[211] vdd gnd cell_6t
Xbit_r212_c22 bl[22] br[22] wl[212] vdd gnd cell_6t
Xbit_r213_c22 bl[22] br[22] wl[213] vdd gnd cell_6t
Xbit_r214_c22 bl[22] br[22] wl[214] vdd gnd cell_6t
Xbit_r215_c22 bl[22] br[22] wl[215] vdd gnd cell_6t
Xbit_r216_c22 bl[22] br[22] wl[216] vdd gnd cell_6t
Xbit_r217_c22 bl[22] br[22] wl[217] vdd gnd cell_6t
Xbit_r218_c22 bl[22] br[22] wl[218] vdd gnd cell_6t
Xbit_r219_c22 bl[22] br[22] wl[219] vdd gnd cell_6t
Xbit_r220_c22 bl[22] br[22] wl[220] vdd gnd cell_6t
Xbit_r221_c22 bl[22] br[22] wl[221] vdd gnd cell_6t
Xbit_r222_c22 bl[22] br[22] wl[222] vdd gnd cell_6t
Xbit_r223_c22 bl[22] br[22] wl[223] vdd gnd cell_6t
Xbit_r224_c22 bl[22] br[22] wl[224] vdd gnd cell_6t
Xbit_r225_c22 bl[22] br[22] wl[225] vdd gnd cell_6t
Xbit_r226_c22 bl[22] br[22] wl[226] vdd gnd cell_6t
Xbit_r227_c22 bl[22] br[22] wl[227] vdd gnd cell_6t
Xbit_r228_c22 bl[22] br[22] wl[228] vdd gnd cell_6t
Xbit_r229_c22 bl[22] br[22] wl[229] vdd gnd cell_6t
Xbit_r230_c22 bl[22] br[22] wl[230] vdd gnd cell_6t
Xbit_r231_c22 bl[22] br[22] wl[231] vdd gnd cell_6t
Xbit_r232_c22 bl[22] br[22] wl[232] vdd gnd cell_6t
Xbit_r233_c22 bl[22] br[22] wl[233] vdd gnd cell_6t
Xbit_r234_c22 bl[22] br[22] wl[234] vdd gnd cell_6t
Xbit_r235_c22 bl[22] br[22] wl[235] vdd gnd cell_6t
Xbit_r236_c22 bl[22] br[22] wl[236] vdd gnd cell_6t
Xbit_r237_c22 bl[22] br[22] wl[237] vdd gnd cell_6t
Xbit_r238_c22 bl[22] br[22] wl[238] vdd gnd cell_6t
Xbit_r239_c22 bl[22] br[22] wl[239] vdd gnd cell_6t
Xbit_r240_c22 bl[22] br[22] wl[240] vdd gnd cell_6t
Xbit_r241_c22 bl[22] br[22] wl[241] vdd gnd cell_6t
Xbit_r242_c22 bl[22] br[22] wl[242] vdd gnd cell_6t
Xbit_r243_c22 bl[22] br[22] wl[243] vdd gnd cell_6t
Xbit_r244_c22 bl[22] br[22] wl[244] vdd gnd cell_6t
Xbit_r245_c22 bl[22] br[22] wl[245] vdd gnd cell_6t
Xbit_r246_c22 bl[22] br[22] wl[246] vdd gnd cell_6t
Xbit_r247_c22 bl[22] br[22] wl[247] vdd gnd cell_6t
Xbit_r248_c22 bl[22] br[22] wl[248] vdd gnd cell_6t
Xbit_r249_c22 bl[22] br[22] wl[249] vdd gnd cell_6t
Xbit_r250_c22 bl[22] br[22] wl[250] vdd gnd cell_6t
Xbit_r251_c22 bl[22] br[22] wl[251] vdd gnd cell_6t
Xbit_r252_c22 bl[22] br[22] wl[252] vdd gnd cell_6t
Xbit_r253_c22 bl[22] br[22] wl[253] vdd gnd cell_6t
Xbit_r254_c22 bl[22] br[22] wl[254] vdd gnd cell_6t
Xbit_r255_c22 bl[22] br[22] wl[255] vdd gnd cell_6t
Xbit_r0_c23 bl[23] br[23] wl[0] vdd gnd cell_6t
Xbit_r1_c23 bl[23] br[23] wl[1] vdd gnd cell_6t
Xbit_r2_c23 bl[23] br[23] wl[2] vdd gnd cell_6t
Xbit_r3_c23 bl[23] br[23] wl[3] vdd gnd cell_6t
Xbit_r4_c23 bl[23] br[23] wl[4] vdd gnd cell_6t
Xbit_r5_c23 bl[23] br[23] wl[5] vdd gnd cell_6t
Xbit_r6_c23 bl[23] br[23] wl[6] vdd gnd cell_6t
Xbit_r7_c23 bl[23] br[23] wl[7] vdd gnd cell_6t
Xbit_r8_c23 bl[23] br[23] wl[8] vdd gnd cell_6t
Xbit_r9_c23 bl[23] br[23] wl[9] vdd gnd cell_6t
Xbit_r10_c23 bl[23] br[23] wl[10] vdd gnd cell_6t
Xbit_r11_c23 bl[23] br[23] wl[11] vdd gnd cell_6t
Xbit_r12_c23 bl[23] br[23] wl[12] vdd gnd cell_6t
Xbit_r13_c23 bl[23] br[23] wl[13] vdd gnd cell_6t
Xbit_r14_c23 bl[23] br[23] wl[14] vdd gnd cell_6t
Xbit_r15_c23 bl[23] br[23] wl[15] vdd gnd cell_6t
Xbit_r16_c23 bl[23] br[23] wl[16] vdd gnd cell_6t
Xbit_r17_c23 bl[23] br[23] wl[17] vdd gnd cell_6t
Xbit_r18_c23 bl[23] br[23] wl[18] vdd gnd cell_6t
Xbit_r19_c23 bl[23] br[23] wl[19] vdd gnd cell_6t
Xbit_r20_c23 bl[23] br[23] wl[20] vdd gnd cell_6t
Xbit_r21_c23 bl[23] br[23] wl[21] vdd gnd cell_6t
Xbit_r22_c23 bl[23] br[23] wl[22] vdd gnd cell_6t
Xbit_r23_c23 bl[23] br[23] wl[23] vdd gnd cell_6t
Xbit_r24_c23 bl[23] br[23] wl[24] vdd gnd cell_6t
Xbit_r25_c23 bl[23] br[23] wl[25] vdd gnd cell_6t
Xbit_r26_c23 bl[23] br[23] wl[26] vdd gnd cell_6t
Xbit_r27_c23 bl[23] br[23] wl[27] vdd gnd cell_6t
Xbit_r28_c23 bl[23] br[23] wl[28] vdd gnd cell_6t
Xbit_r29_c23 bl[23] br[23] wl[29] vdd gnd cell_6t
Xbit_r30_c23 bl[23] br[23] wl[30] vdd gnd cell_6t
Xbit_r31_c23 bl[23] br[23] wl[31] vdd gnd cell_6t
Xbit_r32_c23 bl[23] br[23] wl[32] vdd gnd cell_6t
Xbit_r33_c23 bl[23] br[23] wl[33] vdd gnd cell_6t
Xbit_r34_c23 bl[23] br[23] wl[34] vdd gnd cell_6t
Xbit_r35_c23 bl[23] br[23] wl[35] vdd gnd cell_6t
Xbit_r36_c23 bl[23] br[23] wl[36] vdd gnd cell_6t
Xbit_r37_c23 bl[23] br[23] wl[37] vdd gnd cell_6t
Xbit_r38_c23 bl[23] br[23] wl[38] vdd gnd cell_6t
Xbit_r39_c23 bl[23] br[23] wl[39] vdd gnd cell_6t
Xbit_r40_c23 bl[23] br[23] wl[40] vdd gnd cell_6t
Xbit_r41_c23 bl[23] br[23] wl[41] vdd gnd cell_6t
Xbit_r42_c23 bl[23] br[23] wl[42] vdd gnd cell_6t
Xbit_r43_c23 bl[23] br[23] wl[43] vdd gnd cell_6t
Xbit_r44_c23 bl[23] br[23] wl[44] vdd gnd cell_6t
Xbit_r45_c23 bl[23] br[23] wl[45] vdd gnd cell_6t
Xbit_r46_c23 bl[23] br[23] wl[46] vdd gnd cell_6t
Xbit_r47_c23 bl[23] br[23] wl[47] vdd gnd cell_6t
Xbit_r48_c23 bl[23] br[23] wl[48] vdd gnd cell_6t
Xbit_r49_c23 bl[23] br[23] wl[49] vdd gnd cell_6t
Xbit_r50_c23 bl[23] br[23] wl[50] vdd gnd cell_6t
Xbit_r51_c23 bl[23] br[23] wl[51] vdd gnd cell_6t
Xbit_r52_c23 bl[23] br[23] wl[52] vdd gnd cell_6t
Xbit_r53_c23 bl[23] br[23] wl[53] vdd gnd cell_6t
Xbit_r54_c23 bl[23] br[23] wl[54] vdd gnd cell_6t
Xbit_r55_c23 bl[23] br[23] wl[55] vdd gnd cell_6t
Xbit_r56_c23 bl[23] br[23] wl[56] vdd gnd cell_6t
Xbit_r57_c23 bl[23] br[23] wl[57] vdd gnd cell_6t
Xbit_r58_c23 bl[23] br[23] wl[58] vdd gnd cell_6t
Xbit_r59_c23 bl[23] br[23] wl[59] vdd gnd cell_6t
Xbit_r60_c23 bl[23] br[23] wl[60] vdd gnd cell_6t
Xbit_r61_c23 bl[23] br[23] wl[61] vdd gnd cell_6t
Xbit_r62_c23 bl[23] br[23] wl[62] vdd gnd cell_6t
Xbit_r63_c23 bl[23] br[23] wl[63] vdd gnd cell_6t
Xbit_r64_c23 bl[23] br[23] wl[64] vdd gnd cell_6t
Xbit_r65_c23 bl[23] br[23] wl[65] vdd gnd cell_6t
Xbit_r66_c23 bl[23] br[23] wl[66] vdd gnd cell_6t
Xbit_r67_c23 bl[23] br[23] wl[67] vdd gnd cell_6t
Xbit_r68_c23 bl[23] br[23] wl[68] vdd gnd cell_6t
Xbit_r69_c23 bl[23] br[23] wl[69] vdd gnd cell_6t
Xbit_r70_c23 bl[23] br[23] wl[70] vdd gnd cell_6t
Xbit_r71_c23 bl[23] br[23] wl[71] vdd gnd cell_6t
Xbit_r72_c23 bl[23] br[23] wl[72] vdd gnd cell_6t
Xbit_r73_c23 bl[23] br[23] wl[73] vdd gnd cell_6t
Xbit_r74_c23 bl[23] br[23] wl[74] vdd gnd cell_6t
Xbit_r75_c23 bl[23] br[23] wl[75] vdd gnd cell_6t
Xbit_r76_c23 bl[23] br[23] wl[76] vdd gnd cell_6t
Xbit_r77_c23 bl[23] br[23] wl[77] vdd gnd cell_6t
Xbit_r78_c23 bl[23] br[23] wl[78] vdd gnd cell_6t
Xbit_r79_c23 bl[23] br[23] wl[79] vdd gnd cell_6t
Xbit_r80_c23 bl[23] br[23] wl[80] vdd gnd cell_6t
Xbit_r81_c23 bl[23] br[23] wl[81] vdd gnd cell_6t
Xbit_r82_c23 bl[23] br[23] wl[82] vdd gnd cell_6t
Xbit_r83_c23 bl[23] br[23] wl[83] vdd gnd cell_6t
Xbit_r84_c23 bl[23] br[23] wl[84] vdd gnd cell_6t
Xbit_r85_c23 bl[23] br[23] wl[85] vdd gnd cell_6t
Xbit_r86_c23 bl[23] br[23] wl[86] vdd gnd cell_6t
Xbit_r87_c23 bl[23] br[23] wl[87] vdd gnd cell_6t
Xbit_r88_c23 bl[23] br[23] wl[88] vdd gnd cell_6t
Xbit_r89_c23 bl[23] br[23] wl[89] vdd gnd cell_6t
Xbit_r90_c23 bl[23] br[23] wl[90] vdd gnd cell_6t
Xbit_r91_c23 bl[23] br[23] wl[91] vdd gnd cell_6t
Xbit_r92_c23 bl[23] br[23] wl[92] vdd gnd cell_6t
Xbit_r93_c23 bl[23] br[23] wl[93] vdd gnd cell_6t
Xbit_r94_c23 bl[23] br[23] wl[94] vdd gnd cell_6t
Xbit_r95_c23 bl[23] br[23] wl[95] vdd gnd cell_6t
Xbit_r96_c23 bl[23] br[23] wl[96] vdd gnd cell_6t
Xbit_r97_c23 bl[23] br[23] wl[97] vdd gnd cell_6t
Xbit_r98_c23 bl[23] br[23] wl[98] vdd gnd cell_6t
Xbit_r99_c23 bl[23] br[23] wl[99] vdd gnd cell_6t
Xbit_r100_c23 bl[23] br[23] wl[100] vdd gnd cell_6t
Xbit_r101_c23 bl[23] br[23] wl[101] vdd gnd cell_6t
Xbit_r102_c23 bl[23] br[23] wl[102] vdd gnd cell_6t
Xbit_r103_c23 bl[23] br[23] wl[103] vdd gnd cell_6t
Xbit_r104_c23 bl[23] br[23] wl[104] vdd gnd cell_6t
Xbit_r105_c23 bl[23] br[23] wl[105] vdd gnd cell_6t
Xbit_r106_c23 bl[23] br[23] wl[106] vdd gnd cell_6t
Xbit_r107_c23 bl[23] br[23] wl[107] vdd gnd cell_6t
Xbit_r108_c23 bl[23] br[23] wl[108] vdd gnd cell_6t
Xbit_r109_c23 bl[23] br[23] wl[109] vdd gnd cell_6t
Xbit_r110_c23 bl[23] br[23] wl[110] vdd gnd cell_6t
Xbit_r111_c23 bl[23] br[23] wl[111] vdd gnd cell_6t
Xbit_r112_c23 bl[23] br[23] wl[112] vdd gnd cell_6t
Xbit_r113_c23 bl[23] br[23] wl[113] vdd gnd cell_6t
Xbit_r114_c23 bl[23] br[23] wl[114] vdd gnd cell_6t
Xbit_r115_c23 bl[23] br[23] wl[115] vdd gnd cell_6t
Xbit_r116_c23 bl[23] br[23] wl[116] vdd gnd cell_6t
Xbit_r117_c23 bl[23] br[23] wl[117] vdd gnd cell_6t
Xbit_r118_c23 bl[23] br[23] wl[118] vdd gnd cell_6t
Xbit_r119_c23 bl[23] br[23] wl[119] vdd gnd cell_6t
Xbit_r120_c23 bl[23] br[23] wl[120] vdd gnd cell_6t
Xbit_r121_c23 bl[23] br[23] wl[121] vdd gnd cell_6t
Xbit_r122_c23 bl[23] br[23] wl[122] vdd gnd cell_6t
Xbit_r123_c23 bl[23] br[23] wl[123] vdd gnd cell_6t
Xbit_r124_c23 bl[23] br[23] wl[124] vdd gnd cell_6t
Xbit_r125_c23 bl[23] br[23] wl[125] vdd gnd cell_6t
Xbit_r126_c23 bl[23] br[23] wl[126] vdd gnd cell_6t
Xbit_r127_c23 bl[23] br[23] wl[127] vdd gnd cell_6t
Xbit_r128_c23 bl[23] br[23] wl[128] vdd gnd cell_6t
Xbit_r129_c23 bl[23] br[23] wl[129] vdd gnd cell_6t
Xbit_r130_c23 bl[23] br[23] wl[130] vdd gnd cell_6t
Xbit_r131_c23 bl[23] br[23] wl[131] vdd gnd cell_6t
Xbit_r132_c23 bl[23] br[23] wl[132] vdd gnd cell_6t
Xbit_r133_c23 bl[23] br[23] wl[133] vdd gnd cell_6t
Xbit_r134_c23 bl[23] br[23] wl[134] vdd gnd cell_6t
Xbit_r135_c23 bl[23] br[23] wl[135] vdd gnd cell_6t
Xbit_r136_c23 bl[23] br[23] wl[136] vdd gnd cell_6t
Xbit_r137_c23 bl[23] br[23] wl[137] vdd gnd cell_6t
Xbit_r138_c23 bl[23] br[23] wl[138] vdd gnd cell_6t
Xbit_r139_c23 bl[23] br[23] wl[139] vdd gnd cell_6t
Xbit_r140_c23 bl[23] br[23] wl[140] vdd gnd cell_6t
Xbit_r141_c23 bl[23] br[23] wl[141] vdd gnd cell_6t
Xbit_r142_c23 bl[23] br[23] wl[142] vdd gnd cell_6t
Xbit_r143_c23 bl[23] br[23] wl[143] vdd gnd cell_6t
Xbit_r144_c23 bl[23] br[23] wl[144] vdd gnd cell_6t
Xbit_r145_c23 bl[23] br[23] wl[145] vdd gnd cell_6t
Xbit_r146_c23 bl[23] br[23] wl[146] vdd gnd cell_6t
Xbit_r147_c23 bl[23] br[23] wl[147] vdd gnd cell_6t
Xbit_r148_c23 bl[23] br[23] wl[148] vdd gnd cell_6t
Xbit_r149_c23 bl[23] br[23] wl[149] vdd gnd cell_6t
Xbit_r150_c23 bl[23] br[23] wl[150] vdd gnd cell_6t
Xbit_r151_c23 bl[23] br[23] wl[151] vdd gnd cell_6t
Xbit_r152_c23 bl[23] br[23] wl[152] vdd gnd cell_6t
Xbit_r153_c23 bl[23] br[23] wl[153] vdd gnd cell_6t
Xbit_r154_c23 bl[23] br[23] wl[154] vdd gnd cell_6t
Xbit_r155_c23 bl[23] br[23] wl[155] vdd gnd cell_6t
Xbit_r156_c23 bl[23] br[23] wl[156] vdd gnd cell_6t
Xbit_r157_c23 bl[23] br[23] wl[157] vdd gnd cell_6t
Xbit_r158_c23 bl[23] br[23] wl[158] vdd gnd cell_6t
Xbit_r159_c23 bl[23] br[23] wl[159] vdd gnd cell_6t
Xbit_r160_c23 bl[23] br[23] wl[160] vdd gnd cell_6t
Xbit_r161_c23 bl[23] br[23] wl[161] vdd gnd cell_6t
Xbit_r162_c23 bl[23] br[23] wl[162] vdd gnd cell_6t
Xbit_r163_c23 bl[23] br[23] wl[163] vdd gnd cell_6t
Xbit_r164_c23 bl[23] br[23] wl[164] vdd gnd cell_6t
Xbit_r165_c23 bl[23] br[23] wl[165] vdd gnd cell_6t
Xbit_r166_c23 bl[23] br[23] wl[166] vdd gnd cell_6t
Xbit_r167_c23 bl[23] br[23] wl[167] vdd gnd cell_6t
Xbit_r168_c23 bl[23] br[23] wl[168] vdd gnd cell_6t
Xbit_r169_c23 bl[23] br[23] wl[169] vdd gnd cell_6t
Xbit_r170_c23 bl[23] br[23] wl[170] vdd gnd cell_6t
Xbit_r171_c23 bl[23] br[23] wl[171] vdd gnd cell_6t
Xbit_r172_c23 bl[23] br[23] wl[172] vdd gnd cell_6t
Xbit_r173_c23 bl[23] br[23] wl[173] vdd gnd cell_6t
Xbit_r174_c23 bl[23] br[23] wl[174] vdd gnd cell_6t
Xbit_r175_c23 bl[23] br[23] wl[175] vdd gnd cell_6t
Xbit_r176_c23 bl[23] br[23] wl[176] vdd gnd cell_6t
Xbit_r177_c23 bl[23] br[23] wl[177] vdd gnd cell_6t
Xbit_r178_c23 bl[23] br[23] wl[178] vdd gnd cell_6t
Xbit_r179_c23 bl[23] br[23] wl[179] vdd gnd cell_6t
Xbit_r180_c23 bl[23] br[23] wl[180] vdd gnd cell_6t
Xbit_r181_c23 bl[23] br[23] wl[181] vdd gnd cell_6t
Xbit_r182_c23 bl[23] br[23] wl[182] vdd gnd cell_6t
Xbit_r183_c23 bl[23] br[23] wl[183] vdd gnd cell_6t
Xbit_r184_c23 bl[23] br[23] wl[184] vdd gnd cell_6t
Xbit_r185_c23 bl[23] br[23] wl[185] vdd gnd cell_6t
Xbit_r186_c23 bl[23] br[23] wl[186] vdd gnd cell_6t
Xbit_r187_c23 bl[23] br[23] wl[187] vdd gnd cell_6t
Xbit_r188_c23 bl[23] br[23] wl[188] vdd gnd cell_6t
Xbit_r189_c23 bl[23] br[23] wl[189] vdd gnd cell_6t
Xbit_r190_c23 bl[23] br[23] wl[190] vdd gnd cell_6t
Xbit_r191_c23 bl[23] br[23] wl[191] vdd gnd cell_6t
Xbit_r192_c23 bl[23] br[23] wl[192] vdd gnd cell_6t
Xbit_r193_c23 bl[23] br[23] wl[193] vdd gnd cell_6t
Xbit_r194_c23 bl[23] br[23] wl[194] vdd gnd cell_6t
Xbit_r195_c23 bl[23] br[23] wl[195] vdd gnd cell_6t
Xbit_r196_c23 bl[23] br[23] wl[196] vdd gnd cell_6t
Xbit_r197_c23 bl[23] br[23] wl[197] vdd gnd cell_6t
Xbit_r198_c23 bl[23] br[23] wl[198] vdd gnd cell_6t
Xbit_r199_c23 bl[23] br[23] wl[199] vdd gnd cell_6t
Xbit_r200_c23 bl[23] br[23] wl[200] vdd gnd cell_6t
Xbit_r201_c23 bl[23] br[23] wl[201] vdd gnd cell_6t
Xbit_r202_c23 bl[23] br[23] wl[202] vdd gnd cell_6t
Xbit_r203_c23 bl[23] br[23] wl[203] vdd gnd cell_6t
Xbit_r204_c23 bl[23] br[23] wl[204] vdd gnd cell_6t
Xbit_r205_c23 bl[23] br[23] wl[205] vdd gnd cell_6t
Xbit_r206_c23 bl[23] br[23] wl[206] vdd gnd cell_6t
Xbit_r207_c23 bl[23] br[23] wl[207] vdd gnd cell_6t
Xbit_r208_c23 bl[23] br[23] wl[208] vdd gnd cell_6t
Xbit_r209_c23 bl[23] br[23] wl[209] vdd gnd cell_6t
Xbit_r210_c23 bl[23] br[23] wl[210] vdd gnd cell_6t
Xbit_r211_c23 bl[23] br[23] wl[211] vdd gnd cell_6t
Xbit_r212_c23 bl[23] br[23] wl[212] vdd gnd cell_6t
Xbit_r213_c23 bl[23] br[23] wl[213] vdd gnd cell_6t
Xbit_r214_c23 bl[23] br[23] wl[214] vdd gnd cell_6t
Xbit_r215_c23 bl[23] br[23] wl[215] vdd gnd cell_6t
Xbit_r216_c23 bl[23] br[23] wl[216] vdd gnd cell_6t
Xbit_r217_c23 bl[23] br[23] wl[217] vdd gnd cell_6t
Xbit_r218_c23 bl[23] br[23] wl[218] vdd gnd cell_6t
Xbit_r219_c23 bl[23] br[23] wl[219] vdd gnd cell_6t
Xbit_r220_c23 bl[23] br[23] wl[220] vdd gnd cell_6t
Xbit_r221_c23 bl[23] br[23] wl[221] vdd gnd cell_6t
Xbit_r222_c23 bl[23] br[23] wl[222] vdd gnd cell_6t
Xbit_r223_c23 bl[23] br[23] wl[223] vdd gnd cell_6t
Xbit_r224_c23 bl[23] br[23] wl[224] vdd gnd cell_6t
Xbit_r225_c23 bl[23] br[23] wl[225] vdd gnd cell_6t
Xbit_r226_c23 bl[23] br[23] wl[226] vdd gnd cell_6t
Xbit_r227_c23 bl[23] br[23] wl[227] vdd gnd cell_6t
Xbit_r228_c23 bl[23] br[23] wl[228] vdd gnd cell_6t
Xbit_r229_c23 bl[23] br[23] wl[229] vdd gnd cell_6t
Xbit_r230_c23 bl[23] br[23] wl[230] vdd gnd cell_6t
Xbit_r231_c23 bl[23] br[23] wl[231] vdd gnd cell_6t
Xbit_r232_c23 bl[23] br[23] wl[232] vdd gnd cell_6t
Xbit_r233_c23 bl[23] br[23] wl[233] vdd gnd cell_6t
Xbit_r234_c23 bl[23] br[23] wl[234] vdd gnd cell_6t
Xbit_r235_c23 bl[23] br[23] wl[235] vdd gnd cell_6t
Xbit_r236_c23 bl[23] br[23] wl[236] vdd gnd cell_6t
Xbit_r237_c23 bl[23] br[23] wl[237] vdd gnd cell_6t
Xbit_r238_c23 bl[23] br[23] wl[238] vdd gnd cell_6t
Xbit_r239_c23 bl[23] br[23] wl[239] vdd gnd cell_6t
Xbit_r240_c23 bl[23] br[23] wl[240] vdd gnd cell_6t
Xbit_r241_c23 bl[23] br[23] wl[241] vdd gnd cell_6t
Xbit_r242_c23 bl[23] br[23] wl[242] vdd gnd cell_6t
Xbit_r243_c23 bl[23] br[23] wl[243] vdd gnd cell_6t
Xbit_r244_c23 bl[23] br[23] wl[244] vdd gnd cell_6t
Xbit_r245_c23 bl[23] br[23] wl[245] vdd gnd cell_6t
Xbit_r246_c23 bl[23] br[23] wl[246] vdd gnd cell_6t
Xbit_r247_c23 bl[23] br[23] wl[247] vdd gnd cell_6t
Xbit_r248_c23 bl[23] br[23] wl[248] vdd gnd cell_6t
Xbit_r249_c23 bl[23] br[23] wl[249] vdd gnd cell_6t
Xbit_r250_c23 bl[23] br[23] wl[250] vdd gnd cell_6t
Xbit_r251_c23 bl[23] br[23] wl[251] vdd gnd cell_6t
Xbit_r252_c23 bl[23] br[23] wl[252] vdd gnd cell_6t
Xbit_r253_c23 bl[23] br[23] wl[253] vdd gnd cell_6t
Xbit_r254_c23 bl[23] br[23] wl[254] vdd gnd cell_6t
Xbit_r255_c23 bl[23] br[23] wl[255] vdd gnd cell_6t
Xbit_r0_c24 bl[24] br[24] wl[0] vdd gnd cell_6t
Xbit_r1_c24 bl[24] br[24] wl[1] vdd gnd cell_6t
Xbit_r2_c24 bl[24] br[24] wl[2] vdd gnd cell_6t
Xbit_r3_c24 bl[24] br[24] wl[3] vdd gnd cell_6t
Xbit_r4_c24 bl[24] br[24] wl[4] vdd gnd cell_6t
Xbit_r5_c24 bl[24] br[24] wl[5] vdd gnd cell_6t
Xbit_r6_c24 bl[24] br[24] wl[6] vdd gnd cell_6t
Xbit_r7_c24 bl[24] br[24] wl[7] vdd gnd cell_6t
Xbit_r8_c24 bl[24] br[24] wl[8] vdd gnd cell_6t
Xbit_r9_c24 bl[24] br[24] wl[9] vdd gnd cell_6t
Xbit_r10_c24 bl[24] br[24] wl[10] vdd gnd cell_6t
Xbit_r11_c24 bl[24] br[24] wl[11] vdd gnd cell_6t
Xbit_r12_c24 bl[24] br[24] wl[12] vdd gnd cell_6t
Xbit_r13_c24 bl[24] br[24] wl[13] vdd gnd cell_6t
Xbit_r14_c24 bl[24] br[24] wl[14] vdd gnd cell_6t
Xbit_r15_c24 bl[24] br[24] wl[15] vdd gnd cell_6t
Xbit_r16_c24 bl[24] br[24] wl[16] vdd gnd cell_6t
Xbit_r17_c24 bl[24] br[24] wl[17] vdd gnd cell_6t
Xbit_r18_c24 bl[24] br[24] wl[18] vdd gnd cell_6t
Xbit_r19_c24 bl[24] br[24] wl[19] vdd gnd cell_6t
Xbit_r20_c24 bl[24] br[24] wl[20] vdd gnd cell_6t
Xbit_r21_c24 bl[24] br[24] wl[21] vdd gnd cell_6t
Xbit_r22_c24 bl[24] br[24] wl[22] vdd gnd cell_6t
Xbit_r23_c24 bl[24] br[24] wl[23] vdd gnd cell_6t
Xbit_r24_c24 bl[24] br[24] wl[24] vdd gnd cell_6t
Xbit_r25_c24 bl[24] br[24] wl[25] vdd gnd cell_6t
Xbit_r26_c24 bl[24] br[24] wl[26] vdd gnd cell_6t
Xbit_r27_c24 bl[24] br[24] wl[27] vdd gnd cell_6t
Xbit_r28_c24 bl[24] br[24] wl[28] vdd gnd cell_6t
Xbit_r29_c24 bl[24] br[24] wl[29] vdd gnd cell_6t
Xbit_r30_c24 bl[24] br[24] wl[30] vdd gnd cell_6t
Xbit_r31_c24 bl[24] br[24] wl[31] vdd gnd cell_6t
Xbit_r32_c24 bl[24] br[24] wl[32] vdd gnd cell_6t
Xbit_r33_c24 bl[24] br[24] wl[33] vdd gnd cell_6t
Xbit_r34_c24 bl[24] br[24] wl[34] vdd gnd cell_6t
Xbit_r35_c24 bl[24] br[24] wl[35] vdd gnd cell_6t
Xbit_r36_c24 bl[24] br[24] wl[36] vdd gnd cell_6t
Xbit_r37_c24 bl[24] br[24] wl[37] vdd gnd cell_6t
Xbit_r38_c24 bl[24] br[24] wl[38] vdd gnd cell_6t
Xbit_r39_c24 bl[24] br[24] wl[39] vdd gnd cell_6t
Xbit_r40_c24 bl[24] br[24] wl[40] vdd gnd cell_6t
Xbit_r41_c24 bl[24] br[24] wl[41] vdd gnd cell_6t
Xbit_r42_c24 bl[24] br[24] wl[42] vdd gnd cell_6t
Xbit_r43_c24 bl[24] br[24] wl[43] vdd gnd cell_6t
Xbit_r44_c24 bl[24] br[24] wl[44] vdd gnd cell_6t
Xbit_r45_c24 bl[24] br[24] wl[45] vdd gnd cell_6t
Xbit_r46_c24 bl[24] br[24] wl[46] vdd gnd cell_6t
Xbit_r47_c24 bl[24] br[24] wl[47] vdd gnd cell_6t
Xbit_r48_c24 bl[24] br[24] wl[48] vdd gnd cell_6t
Xbit_r49_c24 bl[24] br[24] wl[49] vdd gnd cell_6t
Xbit_r50_c24 bl[24] br[24] wl[50] vdd gnd cell_6t
Xbit_r51_c24 bl[24] br[24] wl[51] vdd gnd cell_6t
Xbit_r52_c24 bl[24] br[24] wl[52] vdd gnd cell_6t
Xbit_r53_c24 bl[24] br[24] wl[53] vdd gnd cell_6t
Xbit_r54_c24 bl[24] br[24] wl[54] vdd gnd cell_6t
Xbit_r55_c24 bl[24] br[24] wl[55] vdd gnd cell_6t
Xbit_r56_c24 bl[24] br[24] wl[56] vdd gnd cell_6t
Xbit_r57_c24 bl[24] br[24] wl[57] vdd gnd cell_6t
Xbit_r58_c24 bl[24] br[24] wl[58] vdd gnd cell_6t
Xbit_r59_c24 bl[24] br[24] wl[59] vdd gnd cell_6t
Xbit_r60_c24 bl[24] br[24] wl[60] vdd gnd cell_6t
Xbit_r61_c24 bl[24] br[24] wl[61] vdd gnd cell_6t
Xbit_r62_c24 bl[24] br[24] wl[62] vdd gnd cell_6t
Xbit_r63_c24 bl[24] br[24] wl[63] vdd gnd cell_6t
Xbit_r64_c24 bl[24] br[24] wl[64] vdd gnd cell_6t
Xbit_r65_c24 bl[24] br[24] wl[65] vdd gnd cell_6t
Xbit_r66_c24 bl[24] br[24] wl[66] vdd gnd cell_6t
Xbit_r67_c24 bl[24] br[24] wl[67] vdd gnd cell_6t
Xbit_r68_c24 bl[24] br[24] wl[68] vdd gnd cell_6t
Xbit_r69_c24 bl[24] br[24] wl[69] vdd gnd cell_6t
Xbit_r70_c24 bl[24] br[24] wl[70] vdd gnd cell_6t
Xbit_r71_c24 bl[24] br[24] wl[71] vdd gnd cell_6t
Xbit_r72_c24 bl[24] br[24] wl[72] vdd gnd cell_6t
Xbit_r73_c24 bl[24] br[24] wl[73] vdd gnd cell_6t
Xbit_r74_c24 bl[24] br[24] wl[74] vdd gnd cell_6t
Xbit_r75_c24 bl[24] br[24] wl[75] vdd gnd cell_6t
Xbit_r76_c24 bl[24] br[24] wl[76] vdd gnd cell_6t
Xbit_r77_c24 bl[24] br[24] wl[77] vdd gnd cell_6t
Xbit_r78_c24 bl[24] br[24] wl[78] vdd gnd cell_6t
Xbit_r79_c24 bl[24] br[24] wl[79] vdd gnd cell_6t
Xbit_r80_c24 bl[24] br[24] wl[80] vdd gnd cell_6t
Xbit_r81_c24 bl[24] br[24] wl[81] vdd gnd cell_6t
Xbit_r82_c24 bl[24] br[24] wl[82] vdd gnd cell_6t
Xbit_r83_c24 bl[24] br[24] wl[83] vdd gnd cell_6t
Xbit_r84_c24 bl[24] br[24] wl[84] vdd gnd cell_6t
Xbit_r85_c24 bl[24] br[24] wl[85] vdd gnd cell_6t
Xbit_r86_c24 bl[24] br[24] wl[86] vdd gnd cell_6t
Xbit_r87_c24 bl[24] br[24] wl[87] vdd gnd cell_6t
Xbit_r88_c24 bl[24] br[24] wl[88] vdd gnd cell_6t
Xbit_r89_c24 bl[24] br[24] wl[89] vdd gnd cell_6t
Xbit_r90_c24 bl[24] br[24] wl[90] vdd gnd cell_6t
Xbit_r91_c24 bl[24] br[24] wl[91] vdd gnd cell_6t
Xbit_r92_c24 bl[24] br[24] wl[92] vdd gnd cell_6t
Xbit_r93_c24 bl[24] br[24] wl[93] vdd gnd cell_6t
Xbit_r94_c24 bl[24] br[24] wl[94] vdd gnd cell_6t
Xbit_r95_c24 bl[24] br[24] wl[95] vdd gnd cell_6t
Xbit_r96_c24 bl[24] br[24] wl[96] vdd gnd cell_6t
Xbit_r97_c24 bl[24] br[24] wl[97] vdd gnd cell_6t
Xbit_r98_c24 bl[24] br[24] wl[98] vdd gnd cell_6t
Xbit_r99_c24 bl[24] br[24] wl[99] vdd gnd cell_6t
Xbit_r100_c24 bl[24] br[24] wl[100] vdd gnd cell_6t
Xbit_r101_c24 bl[24] br[24] wl[101] vdd gnd cell_6t
Xbit_r102_c24 bl[24] br[24] wl[102] vdd gnd cell_6t
Xbit_r103_c24 bl[24] br[24] wl[103] vdd gnd cell_6t
Xbit_r104_c24 bl[24] br[24] wl[104] vdd gnd cell_6t
Xbit_r105_c24 bl[24] br[24] wl[105] vdd gnd cell_6t
Xbit_r106_c24 bl[24] br[24] wl[106] vdd gnd cell_6t
Xbit_r107_c24 bl[24] br[24] wl[107] vdd gnd cell_6t
Xbit_r108_c24 bl[24] br[24] wl[108] vdd gnd cell_6t
Xbit_r109_c24 bl[24] br[24] wl[109] vdd gnd cell_6t
Xbit_r110_c24 bl[24] br[24] wl[110] vdd gnd cell_6t
Xbit_r111_c24 bl[24] br[24] wl[111] vdd gnd cell_6t
Xbit_r112_c24 bl[24] br[24] wl[112] vdd gnd cell_6t
Xbit_r113_c24 bl[24] br[24] wl[113] vdd gnd cell_6t
Xbit_r114_c24 bl[24] br[24] wl[114] vdd gnd cell_6t
Xbit_r115_c24 bl[24] br[24] wl[115] vdd gnd cell_6t
Xbit_r116_c24 bl[24] br[24] wl[116] vdd gnd cell_6t
Xbit_r117_c24 bl[24] br[24] wl[117] vdd gnd cell_6t
Xbit_r118_c24 bl[24] br[24] wl[118] vdd gnd cell_6t
Xbit_r119_c24 bl[24] br[24] wl[119] vdd gnd cell_6t
Xbit_r120_c24 bl[24] br[24] wl[120] vdd gnd cell_6t
Xbit_r121_c24 bl[24] br[24] wl[121] vdd gnd cell_6t
Xbit_r122_c24 bl[24] br[24] wl[122] vdd gnd cell_6t
Xbit_r123_c24 bl[24] br[24] wl[123] vdd gnd cell_6t
Xbit_r124_c24 bl[24] br[24] wl[124] vdd gnd cell_6t
Xbit_r125_c24 bl[24] br[24] wl[125] vdd gnd cell_6t
Xbit_r126_c24 bl[24] br[24] wl[126] vdd gnd cell_6t
Xbit_r127_c24 bl[24] br[24] wl[127] vdd gnd cell_6t
Xbit_r128_c24 bl[24] br[24] wl[128] vdd gnd cell_6t
Xbit_r129_c24 bl[24] br[24] wl[129] vdd gnd cell_6t
Xbit_r130_c24 bl[24] br[24] wl[130] vdd gnd cell_6t
Xbit_r131_c24 bl[24] br[24] wl[131] vdd gnd cell_6t
Xbit_r132_c24 bl[24] br[24] wl[132] vdd gnd cell_6t
Xbit_r133_c24 bl[24] br[24] wl[133] vdd gnd cell_6t
Xbit_r134_c24 bl[24] br[24] wl[134] vdd gnd cell_6t
Xbit_r135_c24 bl[24] br[24] wl[135] vdd gnd cell_6t
Xbit_r136_c24 bl[24] br[24] wl[136] vdd gnd cell_6t
Xbit_r137_c24 bl[24] br[24] wl[137] vdd gnd cell_6t
Xbit_r138_c24 bl[24] br[24] wl[138] vdd gnd cell_6t
Xbit_r139_c24 bl[24] br[24] wl[139] vdd gnd cell_6t
Xbit_r140_c24 bl[24] br[24] wl[140] vdd gnd cell_6t
Xbit_r141_c24 bl[24] br[24] wl[141] vdd gnd cell_6t
Xbit_r142_c24 bl[24] br[24] wl[142] vdd gnd cell_6t
Xbit_r143_c24 bl[24] br[24] wl[143] vdd gnd cell_6t
Xbit_r144_c24 bl[24] br[24] wl[144] vdd gnd cell_6t
Xbit_r145_c24 bl[24] br[24] wl[145] vdd gnd cell_6t
Xbit_r146_c24 bl[24] br[24] wl[146] vdd gnd cell_6t
Xbit_r147_c24 bl[24] br[24] wl[147] vdd gnd cell_6t
Xbit_r148_c24 bl[24] br[24] wl[148] vdd gnd cell_6t
Xbit_r149_c24 bl[24] br[24] wl[149] vdd gnd cell_6t
Xbit_r150_c24 bl[24] br[24] wl[150] vdd gnd cell_6t
Xbit_r151_c24 bl[24] br[24] wl[151] vdd gnd cell_6t
Xbit_r152_c24 bl[24] br[24] wl[152] vdd gnd cell_6t
Xbit_r153_c24 bl[24] br[24] wl[153] vdd gnd cell_6t
Xbit_r154_c24 bl[24] br[24] wl[154] vdd gnd cell_6t
Xbit_r155_c24 bl[24] br[24] wl[155] vdd gnd cell_6t
Xbit_r156_c24 bl[24] br[24] wl[156] vdd gnd cell_6t
Xbit_r157_c24 bl[24] br[24] wl[157] vdd gnd cell_6t
Xbit_r158_c24 bl[24] br[24] wl[158] vdd gnd cell_6t
Xbit_r159_c24 bl[24] br[24] wl[159] vdd gnd cell_6t
Xbit_r160_c24 bl[24] br[24] wl[160] vdd gnd cell_6t
Xbit_r161_c24 bl[24] br[24] wl[161] vdd gnd cell_6t
Xbit_r162_c24 bl[24] br[24] wl[162] vdd gnd cell_6t
Xbit_r163_c24 bl[24] br[24] wl[163] vdd gnd cell_6t
Xbit_r164_c24 bl[24] br[24] wl[164] vdd gnd cell_6t
Xbit_r165_c24 bl[24] br[24] wl[165] vdd gnd cell_6t
Xbit_r166_c24 bl[24] br[24] wl[166] vdd gnd cell_6t
Xbit_r167_c24 bl[24] br[24] wl[167] vdd gnd cell_6t
Xbit_r168_c24 bl[24] br[24] wl[168] vdd gnd cell_6t
Xbit_r169_c24 bl[24] br[24] wl[169] vdd gnd cell_6t
Xbit_r170_c24 bl[24] br[24] wl[170] vdd gnd cell_6t
Xbit_r171_c24 bl[24] br[24] wl[171] vdd gnd cell_6t
Xbit_r172_c24 bl[24] br[24] wl[172] vdd gnd cell_6t
Xbit_r173_c24 bl[24] br[24] wl[173] vdd gnd cell_6t
Xbit_r174_c24 bl[24] br[24] wl[174] vdd gnd cell_6t
Xbit_r175_c24 bl[24] br[24] wl[175] vdd gnd cell_6t
Xbit_r176_c24 bl[24] br[24] wl[176] vdd gnd cell_6t
Xbit_r177_c24 bl[24] br[24] wl[177] vdd gnd cell_6t
Xbit_r178_c24 bl[24] br[24] wl[178] vdd gnd cell_6t
Xbit_r179_c24 bl[24] br[24] wl[179] vdd gnd cell_6t
Xbit_r180_c24 bl[24] br[24] wl[180] vdd gnd cell_6t
Xbit_r181_c24 bl[24] br[24] wl[181] vdd gnd cell_6t
Xbit_r182_c24 bl[24] br[24] wl[182] vdd gnd cell_6t
Xbit_r183_c24 bl[24] br[24] wl[183] vdd gnd cell_6t
Xbit_r184_c24 bl[24] br[24] wl[184] vdd gnd cell_6t
Xbit_r185_c24 bl[24] br[24] wl[185] vdd gnd cell_6t
Xbit_r186_c24 bl[24] br[24] wl[186] vdd gnd cell_6t
Xbit_r187_c24 bl[24] br[24] wl[187] vdd gnd cell_6t
Xbit_r188_c24 bl[24] br[24] wl[188] vdd gnd cell_6t
Xbit_r189_c24 bl[24] br[24] wl[189] vdd gnd cell_6t
Xbit_r190_c24 bl[24] br[24] wl[190] vdd gnd cell_6t
Xbit_r191_c24 bl[24] br[24] wl[191] vdd gnd cell_6t
Xbit_r192_c24 bl[24] br[24] wl[192] vdd gnd cell_6t
Xbit_r193_c24 bl[24] br[24] wl[193] vdd gnd cell_6t
Xbit_r194_c24 bl[24] br[24] wl[194] vdd gnd cell_6t
Xbit_r195_c24 bl[24] br[24] wl[195] vdd gnd cell_6t
Xbit_r196_c24 bl[24] br[24] wl[196] vdd gnd cell_6t
Xbit_r197_c24 bl[24] br[24] wl[197] vdd gnd cell_6t
Xbit_r198_c24 bl[24] br[24] wl[198] vdd gnd cell_6t
Xbit_r199_c24 bl[24] br[24] wl[199] vdd gnd cell_6t
Xbit_r200_c24 bl[24] br[24] wl[200] vdd gnd cell_6t
Xbit_r201_c24 bl[24] br[24] wl[201] vdd gnd cell_6t
Xbit_r202_c24 bl[24] br[24] wl[202] vdd gnd cell_6t
Xbit_r203_c24 bl[24] br[24] wl[203] vdd gnd cell_6t
Xbit_r204_c24 bl[24] br[24] wl[204] vdd gnd cell_6t
Xbit_r205_c24 bl[24] br[24] wl[205] vdd gnd cell_6t
Xbit_r206_c24 bl[24] br[24] wl[206] vdd gnd cell_6t
Xbit_r207_c24 bl[24] br[24] wl[207] vdd gnd cell_6t
Xbit_r208_c24 bl[24] br[24] wl[208] vdd gnd cell_6t
Xbit_r209_c24 bl[24] br[24] wl[209] vdd gnd cell_6t
Xbit_r210_c24 bl[24] br[24] wl[210] vdd gnd cell_6t
Xbit_r211_c24 bl[24] br[24] wl[211] vdd gnd cell_6t
Xbit_r212_c24 bl[24] br[24] wl[212] vdd gnd cell_6t
Xbit_r213_c24 bl[24] br[24] wl[213] vdd gnd cell_6t
Xbit_r214_c24 bl[24] br[24] wl[214] vdd gnd cell_6t
Xbit_r215_c24 bl[24] br[24] wl[215] vdd gnd cell_6t
Xbit_r216_c24 bl[24] br[24] wl[216] vdd gnd cell_6t
Xbit_r217_c24 bl[24] br[24] wl[217] vdd gnd cell_6t
Xbit_r218_c24 bl[24] br[24] wl[218] vdd gnd cell_6t
Xbit_r219_c24 bl[24] br[24] wl[219] vdd gnd cell_6t
Xbit_r220_c24 bl[24] br[24] wl[220] vdd gnd cell_6t
Xbit_r221_c24 bl[24] br[24] wl[221] vdd gnd cell_6t
Xbit_r222_c24 bl[24] br[24] wl[222] vdd gnd cell_6t
Xbit_r223_c24 bl[24] br[24] wl[223] vdd gnd cell_6t
Xbit_r224_c24 bl[24] br[24] wl[224] vdd gnd cell_6t
Xbit_r225_c24 bl[24] br[24] wl[225] vdd gnd cell_6t
Xbit_r226_c24 bl[24] br[24] wl[226] vdd gnd cell_6t
Xbit_r227_c24 bl[24] br[24] wl[227] vdd gnd cell_6t
Xbit_r228_c24 bl[24] br[24] wl[228] vdd gnd cell_6t
Xbit_r229_c24 bl[24] br[24] wl[229] vdd gnd cell_6t
Xbit_r230_c24 bl[24] br[24] wl[230] vdd gnd cell_6t
Xbit_r231_c24 bl[24] br[24] wl[231] vdd gnd cell_6t
Xbit_r232_c24 bl[24] br[24] wl[232] vdd gnd cell_6t
Xbit_r233_c24 bl[24] br[24] wl[233] vdd gnd cell_6t
Xbit_r234_c24 bl[24] br[24] wl[234] vdd gnd cell_6t
Xbit_r235_c24 bl[24] br[24] wl[235] vdd gnd cell_6t
Xbit_r236_c24 bl[24] br[24] wl[236] vdd gnd cell_6t
Xbit_r237_c24 bl[24] br[24] wl[237] vdd gnd cell_6t
Xbit_r238_c24 bl[24] br[24] wl[238] vdd gnd cell_6t
Xbit_r239_c24 bl[24] br[24] wl[239] vdd gnd cell_6t
Xbit_r240_c24 bl[24] br[24] wl[240] vdd gnd cell_6t
Xbit_r241_c24 bl[24] br[24] wl[241] vdd gnd cell_6t
Xbit_r242_c24 bl[24] br[24] wl[242] vdd gnd cell_6t
Xbit_r243_c24 bl[24] br[24] wl[243] vdd gnd cell_6t
Xbit_r244_c24 bl[24] br[24] wl[244] vdd gnd cell_6t
Xbit_r245_c24 bl[24] br[24] wl[245] vdd gnd cell_6t
Xbit_r246_c24 bl[24] br[24] wl[246] vdd gnd cell_6t
Xbit_r247_c24 bl[24] br[24] wl[247] vdd gnd cell_6t
Xbit_r248_c24 bl[24] br[24] wl[248] vdd gnd cell_6t
Xbit_r249_c24 bl[24] br[24] wl[249] vdd gnd cell_6t
Xbit_r250_c24 bl[24] br[24] wl[250] vdd gnd cell_6t
Xbit_r251_c24 bl[24] br[24] wl[251] vdd gnd cell_6t
Xbit_r252_c24 bl[24] br[24] wl[252] vdd gnd cell_6t
Xbit_r253_c24 bl[24] br[24] wl[253] vdd gnd cell_6t
Xbit_r254_c24 bl[24] br[24] wl[254] vdd gnd cell_6t
Xbit_r255_c24 bl[24] br[24] wl[255] vdd gnd cell_6t
Xbit_r0_c25 bl[25] br[25] wl[0] vdd gnd cell_6t
Xbit_r1_c25 bl[25] br[25] wl[1] vdd gnd cell_6t
Xbit_r2_c25 bl[25] br[25] wl[2] vdd gnd cell_6t
Xbit_r3_c25 bl[25] br[25] wl[3] vdd gnd cell_6t
Xbit_r4_c25 bl[25] br[25] wl[4] vdd gnd cell_6t
Xbit_r5_c25 bl[25] br[25] wl[5] vdd gnd cell_6t
Xbit_r6_c25 bl[25] br[25] wl[6] vdd gnd cell_6t
Xbit_r7_c25 bl[25] br[25] wl[7] vdd gnd cell_6t
Xbit_r8_c25 bl[25] br[25] wl[8] vdd gnd cell_6t
Xbit_r9_c25 bl[25] br[25] wl[9] vdd gnd cell_6t
Xbit_r10_c25 bl[25] br[25] wl[10] vdd gnd cell_6t
Xbit_r11_c25 bl[25] br[25] wl[11] vdd gnd cell_6t
Xbit_r12_c25 bl[25] br[25] wl[12] vdd gnd cell_6t
Xbit_r13_c25 bl[25] br[25] wl[13] vdd gnd cell_6t
Xbit_r14_c25 bl[25] br[25] wl[14] vdd gnd cell_6t
Xbit_r15_c25 bl[25] br[25] wl[15] vdd gnd cell_6t
Xbit_r16_c25 bl[25] br[25] wl[16] vdd gnd cell_6t
Xbit_r17_c25 bl[25] br[25] wl[17] vdd gnd cell_6t
Xbit_r18_c25 bl[25] br[25] wl[18] vdd gnd cell_6t
Xbit_r19_c25 bl[25] br[25] wl[19] vdd gnd cell_6t
Xbit_r20_c25 bl[25] br[25] wl[20] vdd gnd cell_6t
Xbit_r21_c25 bl[25] br[25] wl[21] vdd gnd cell_6t
Xbit_r22_c25 bl[25] br[25] wl[22] vdd gnd cell_6t
Xbit_r23_c25 bl[25] br[25] wl[23] vdd gnd cell_6t
Xbit_r24_c25 bl[25] br[25] wl[24] vdd gnd cell_6t
Xbit_r25_c25 bl[25] br[25] wl[25] vdd gnd cell_6t
Xbit_r26_c25 bl[25] br[25] wl[26] vdd gnd cell_6t
Xbit_r27_c25 bl[25] br[25] wl[27] vdd gnd cell_6t
Xbit_r28_c25 bl[25] br[25] wl[28] vdd gnd cell_6t
Xbit_r29_c25 bl[25] br[25] wl[29] vdd gnd cell_6t
Xbit_r30_c25 bl[25] br[25] wl[30] vdd gnd cell_6t
Xbit_r31_c25 bl[25] br[25] wl[31] vdd gnd cell_6t
Xbit_r32_c25 bl[25] br[25] wl[32] vdd gnd cell_6t
Xbit_r33_c25 bl[25] br[25] wl[33] vdd gnd cell_6t
Xbit_r34_c25 bl[25] br[25] wl[34] vdd gnd cell_6t
Xbit_r35_c25 bl[25] br[25] wl[35] vdd gnd cell_6t
Xbit_r36_c25 bl[25] br[25] wl[36] vdd gnd cell_6t
Xbit_r37_c25 bl[25] br[25] wl[37] vdd gnd cell_6t
Xbit_r38_c25 bl[25] br[25] wl[38] vdd gnd cell_6t
Xbit_r39_c25 bl[25] br[25] wl[39] vdd gnd cell_6t
Xbit_r40_c25 bl[25] br[25] wl[40] vdd gnd cell_6t
Xbit_r41_c25 bl[25] br[25] wl[41] vdd gnd cell_6t
Xbit_r42_c25 bl[25] br[25] wl[42] vdd gnd cell_6t
Xbit_r43_c25 bl[25] br[25] wl[43] vdd gnd cell_6t
Xbit_r44_c25 bl[25] br[25] wl[44] vdd gnd cell_6t
Xbit_r45_c25 bl[25] br[25] wl[45] vdd gnd cell_6t
Xbit_r46_c25 bl[25] br[25] wl[46] vdd gnd cell_6t
Xbit_r47_c25 bl[25] br[25] wl[47] vdd gnd cell_6t
Xbit_r48_c25 bl[25] br[25] wl[48] vdd gnd cell_6t
Xbit_r49_c25 bl[25] br[25] wl[49] vdd gnd cell_6t
Xbit_r50_c25 bl[25] br[25] wl[50] vdd gnd cell_6t
Xbit_r51_c25 bl[25] br[25] wl[51] vdd gnd cell_6t
Xbit_r52_c25 bl[25] br[25] wl[52] vdd gnd cell_6t
Xbit_r53_c25 bl[25] br[25] wl[53] vdd gnd cell_6t
Xbit_r54_c25 bl[25] br[25] wl[54] vdd gnd cell_6t
Xbit_r55_c25 bl[25] br[25] wl[55] vdd gnd cell_6t
Xbit_r56_c25 bl[25] br[25] wl[56] vdd gnd cell_6t
Xbit_r57_c25 bl[25] br[25] wl[57] vdd gnd cell_6t
Xbit_r58_c25 bl[25] br[25] wl[58] vdd gnd cell_6t
Xbit_r59_c25 bl[25] br[25] wl[59] vdd gnd cell_6t
Xbit_r60_c25 bl[25] br[25] wl[60] vdd gnd cell_6t
Xbit_r61_c25 bl[25] br[25] wl[61] vdd gnd cell_6t
Xbit_r62_c25 bl[25] br[25] wl[62] vdd gnd cell_6t
Xbit_r63_c25 bl[25] br[25] wl[63] vdd gnd cell_6t
Xbit_r64_c25 bl[25] br[25] wl[64] vdd gnd cell_6t
Xbit_r65_c25 bl[25] br[25] wl[65] vdd gnd cell_6t
Xbit_r66_c25 bl[25] br[25] wl[66] vdd gnd cell_6t
Xbit_r67_c25 bl[25] br[25] wl[67] vdd gnd cell_6t
Xbit_r68_c25 bl[25] br[25] wl[68] vdd gnd cell_6t
Xbit_r69_c25 bl[25] br[25] wl[69] vdd gnd cell_6t
Xbit_r70_c25 bl[25] br[25] wl[70] vdd gnd cell_6t
Xbit_r71_c25 bl[25] br[25] wl[71] vdd gnd cell_6t
Xbit_r72_c25 bl[25] br[25] wl[72] vdd gnd cell_6t
Xbit_r73_c25 bl[25] br[25] wl[73] vdd gnd cell_6t
Xbit_r74_c25 bl[25] br[25] wl[74] vdd gnd cell_6t
Xbit_r75_c25 bl[25] br[25] wl[75] vdd gnd cell_6t
Xbit_r76_c25 bl[25] br[25] wl[76] vdd gnd cell_6t
Xbit_r77_c25 bl[25] br[25] wl[77] vdd gnd cell_6t
Xbit_r78_c25 bl[25] br[25] wl[78] vdd gnd cell_6t
Xbit_r79_c25 bl[25] br[25] wl[79] vdd gnd cell_6t
Xbit_r80_c25 bl[25] br[25] wl[80] vdd gnd cell_6t
Xbit_r81_c25 bl[25] br[25] wl[81] vdd gnd cell_6t
Xbit_r82_c25 bl[25] br[25] wl[82] vdd gnd cell_6t
Xbit_r83_c25 bl[25] br[25] wl[83] vdd gnd cell_6t
Xbit_r84_c25 bl[25] br[25] wl[84] vdd gnd cell_6t
Xbit_r85_c25 bl[25] br[25] wl[85] vdd gnd cell_6t
Xbit_r86_c25 bl[25] br[25] wl[86] vdd gnd cell_6t
Xbit_r87_c25 bl[25] br[25] wl[87] vdd gnd cell_6t
Xbit_r88_c25 bl[25] br[25] wl[88] vdd gnd cell_6t
Xbit_r89_c25 bl[25] br[25] wl[89] vdd gnd cell_6t
Xbit_r90_c25 bl[25] br[25] wl[90] vdd gnd cell_6t
Xbit_r91_c25 bl[25] br[25] wl[91] vdd gnd cell_6t
Xbit_r92_c25 bl[25] br[25] wl[92] vdd gnd cell_6t
Xbit_r93_c25 bl[25] br[25] wl[93] vdd gnd cell_6t
Xbit_r94_c25 bl[25] br[25] wl[94] vdd gnd cell_6t
Xbit_r95_c25 bl[25] br[25] wl[95] vdd gnd cell_6t
Xbit_r96_c25 bl[25] br[25] wl[96] vdd gnd cell_6t
Xbit_r97_c25 bl[25] br[25] wl[97] vdd gnd cell_6t
Xbit_r98_c25 bl[25] br[25] wl[98] vdd gnd cell_6t
Xbit_r99_c25 bl[25] br[25] wl[99] vdd gnd cell_6t
Xbit_r100_c25 bl[25] br[25] wl[100] vdd gnd cell_6t
Xbit_r101_c25 bl[25] br[25] wl[101] vdd gnd cell_6t
Xbit_r102_c25 bl[25] br[25] wl[102] vdd gnd cell_6t
Xbit_r103_c25 bl[25] br[25] wl[103] vdd gnd cell_6t
Xbit_r104_c25 bl[25] br[25] wl[104] vdd gnd cell_6t
Xbit_r105_c25 bl[25] br[25] wl[105] vdd gnd cell_6t
Xbit_r106_c25 bl[25] br[25] wl[106] vdd gnd cell_6t
Xbit_r107_c25 bl[25] br[25] wl[107] vdd gnd cell_6t
Xbit_r108_c25 bl[25] br[25] wl[108] vdd gnd cell_6t
Xbit_r109_c25 bl[25] br[25] wl[109] vdd gnd cell_6t
Xbit_r110_c25 bl[25] br[25] wl[110] vdd gnd cell_6t
Xbit_r111_c25 bl[25] br[25] wl[111] vdd gnd cell_6t
Xbit_r112_c25 bl[25] br[25] wl[112] vdd gnd cell_6t
Xbit_r113_c25 bl[25] br[25] wl[113] vdd gnd cell_6t
Xbit_r114_c25 bl[25] br[25] wl[114] vdd gnd cell_6t
Xbit_r115_c25 bl[25] br[25] wl[115] vdd gnd cell_6t
Xbit_r116_c25 bl[25] br[25] wl[116] vdd gnd cell_6t
Xbit_r117_c25 bl[25] br[25] wl[117] vdd gnd cell_6t
Xbit_r118_c25 bl[25] br[25] wl[118] vdd gnd cell_6t
Xbit_r119_c25 bl[25] br[25] wl[119] vdd gnd cell_6t
Xbit_r120_c25 bl[25] br[25] wl[120] vdd gnd cell_6t
Xbit_r121_c25 bl[25] br[25] wl[121] vdd gnd cell_6t
Xbit_r122_c25 bl[25] br[25] wl[122] vdd gnd cell_6t
Xbit_r123_c25 bl[25] br[25] wl[123] vdd gnd cell_6t
Xbit_r124_c25 bl[25] br[25] wl[124] vdd gnd cell_6t
Xbit_r125_c25 bl[25] br[25] wl[125] vdd gnd cell_6t
Xbit_r126_c25 bl[25] br[25] wl[126] vdd gnd cell_6t
Xbit_r127_c25 bl[25] br[25] wl[127] vdd gnd cell_6t
Xbit_r128_c25 bl[25] br[25] wl[128] vdd gnd cell_6t
Xbit_r129_c25 bl[25] br[25] wl[129] vdd gnd cell_6t
Xbit_r130_c25 bl[25] br[25] wl[130] vdd gnd cell_6t
Xbit_r131_c25 bl[25] br[25] wl[131] vdd gnd cell_6t
Xbit_r132_c25 bl[25] br[25] wl[132] vdd gnd cell_6t
Xbit_r133_c25 bl[25] br[25] wl[133] vdd gnd cell_6t
Xbit_r134_c25 bl[25] br[25] wl[134] vdd gnd cell_6t
Xbit_r135_c25 bl[25] br[25] wl[135] vdd gnd cell_6t
Xbit_r136_c25 bl[25] br[25] wl[136] vdd gnd cell_6t
Xbit_r137_c25 bl[25] br[25] wl[137] vdd gnd cell_6t
Xbit_r138_c25 bl[25] br[25] wl[138] vdd gnd cell_6t
Xbit_r139_c25 bl[25] br[25] wl[139] vdd gnd cell_6t
Xbit_r140_c25 bl[25] br[25] wl[140] vdd gnd cell_6t
Xbit_r141_c25 bl[25] br[25] wl[141] vdd gnd cell_6t
Xbit_r142_c25 bl[25] br[25] wl[142] vdd gnd cell_6t
Xbit_r143_c25 bl[25] br[25] wl[143] vdd gnd cell_6t
Xbit_r144_c25 bl[25] br[25] wl[144] vdd gnd cell_6t
Xbit_r145_c25 bl[25] br[25] wl[145] vdd gnd cell_6t
Xbit_r146_c25 bl[25] br[25] wl[146] vdd gnd cell_6t
Xbit_r147_c25 bl[25] br[25] wl[147] vdd gnd cell_6t
Xbit_r148_c25 bl[25] br[25] wl[148] vdd gnd cell_6t
Xbit_r149_c25 bl[25] br[25] wl[149] vdd gnd cell_6t
Xbit_r150_c25 bl[25] br[25] wl[150] vdd gnd cell_6t
Xbit_r151_c25 bl[25] br[25] wl[151] vdd gnd cell_6t
Xbit_r152_c25 bl[25] br[25] wl[152] vdd gnd cell_6t
Xbit_r153_c25 bl[25] br[25] wl[153] vdd gnd cell_6t
Xbit_r154_c25 bl[25] br[25] wl[154] vdd gnd cell_6t
Xbit_r155_c25 bl[25] br[25] wl[155] vdd gnd cell_6t
Xbit_r156_c25 bl[25] br[25] wl[156] vdd gnd cell_6t
Xbit_r157_c25 bl[25] br[25] wl[157] vdd gnd cell_6t
Xbit_r158_c25 bl[25] br[25] wl[158] vdd gnd cell_6t
Xbit_r159_c25 bl[25] br[25] wl[159] vdd gnd cell_6t
Xbit_r160_c25 bl[25] br[25] wl[160] vdd gnd cell_6t
Xbit_r161_c25 bl[25] br[25] wl[161] vdd gnd cell_6t
Xbit_r162_c25 bl[25] br[25] wl[162] vdd gnd cell_6t
Xbit_r163_c25 bl[25] br[25] wl[163] vdd gnd cell_6t
Xbit_r164_c25 bl[25] br[25] wl[164] vdd gnd cell_6t
Xbit_r165_c25 bl[25] br[25] wl[165] vdd gnd cell_6t
Xbit_r166_c25 bl[25] br[25] wl[166] vdd gnd cell_6t
Xbit_r167_c25 bl[25] br[25] wl[167] vdd gnd cell_6t
Xbit_r168_c25 bl[25] br[25] wl[168] vdd gnd cell_6t
Xbit_r169_c25 bl[25] br[25] wl[169] vdd gnd cell_6t
Xbit_r170_c25 bl[25] br[25] wl[170] vdd gnd cell_6t
Xbit_r171_c25 bl[25] br[25] wl[171] vdd gnd cell_6t
Xbit_r172_c25 bl[25] br[25] wl[172] vdd gnd cell_6t
Xbit_r173_c25 bl[25] br[25] wl[173] vdd gnd cell_6t
Xbit_r174_c25 bl[25] br[25] wl[174] vdd gnd cell_6t
Xbit_r175_c25 bl[25] br[25] wl[175] vdd gnd cell_6t
Xbit_r176_c25 bl[25] br[25] wl[176] vdd gnd cell_6t
Xbit_r177_c25 bl[25] br[25] wl[177] vdd gnd cell_6t
Xbit_r178_c25 bl[25] br[25] wl[178] vdd gnd cell_6t
Xbit_r179_c25 bl[25] br[25] wl[179] vdd gnd cell_6t
Xbit_r180_c25 bl[25] br[25] wl[180] vdd gnd cell_6t
Xbit_r181_c25 bl[25] br[25] wl[181] vdd gnd cell_6t
Xbit_r182_c25 bl[25] br[25] wl[182] vdd gnd cell_6t
Xbit_r183_c25 bl[25] br[25] wl[183] vdd gnd cell_6t
Xbit_r184_c25 bl[25] br[25] wl[184] vdd gnd cell_6t
Xbit_r185_c25 bl[25] br[25] wl[185] vdd gnd cell_6t
Xbit_r186_c25 bl[25] br[25] wl[186] vdd gnd cell_6t
Xbit_r187_c25 bl[25] br[25] wl[187] vdd gnd cell_6t
Xbit_r188_c25 bl[25] br[25] wl[188] vdd gnd cell_6t
Xbit_r189_c25 bl[25] br[25] wl[189] vdd gnd cell_6t
Xbit_r190_c25 bl[25] br[25] wl[190] vdd gnd cell_6t
Xbit_r191_c25 bl[25] br[25] wl[191] vdd gnd cell_6t
Xbit_r192_c25 bl[25] br[25] wl[192] vdd gnd cell_6t
Xbit_r193_c25 bl[25] br[25] wl[193] vdd gnd cell_6t
Xbit_r194_c25 bl[25] br[25] wl[194] vdd gnd cell_6t
Xbit_r195_c25 bl[25] br[25] wl[195] vdd gnd cell_6t
Xbit_r196_c25 bl[25] br[25] wl[196] vdd gnd cell_6t
Xbit_r197_c25 bl[25] br[25] wl[197] vdd gnd cell_6t
Xbit_r198_c25 bl[25] br[25] wl[198] vdd gnd cell_6t
Xbit_r199_c25 bl[25] br[25] wl[199] vdd gnd cell_6t
Xbit_r200_c25 bl[25] br[25] wl[200] vdd gnd cell_6t
Xbit_r201_c25 bl[25] br[25] wl[201] vdd gnd cell_6t
Xbit_r202_c25 bl[25] br[25] wl[202] vdd gnd cell_6t
Xbit_r203_c25 bl[25] br[25] wl[203] vdd gnd cell_6t
Xbit_r204_c25 bl[25] br[25] wl[204] vdd gnd cell_6t
Xbit_r205_c25 bl[25] br[25] wl[205] vdd gnd cell_6t
Xbit_r206_c25 bl[25] br[25] wl[206] vdd gnd cell_6t
Xbit_r207_c25 bl[25] br[25] wl[207] vdd gnd cell_6t
Xbit_r208_c25 bl[25] br[25] wl[208] vdd gnd cell_6t
Xbit_r209_c25 bl[25] br[25] wl[209] vdd gnd cell_6t
Xbit_r210_c25 bl[25] br[25] wl[210] vdd gnd cell_6t
Xbit_r211_c25 bl[25] br[25] wl[211] vdd gnd cell_6t
Xbit_r212_c25 bl[25] br[25] wl[212] vdd gnd cell_6t
Xbit_r213_c25 bl[25] br[25] wl[213] vdd gnd cell_6t
Xbit_r214_c25 bl[25] br[25] wl[214] vdd gnd cell_6t
Xbit_r215_c25 bl[25] br[25] wl[215] vdd gnd cell_6t
Xbit_r216_c25 bl[25] br[25] wl[216] vdd gnd cell_6t
Xbit_r217_c25 bl[25] br[25] wl[217] vdd gnd cell_6t
Xbit_r218_c25 bl[25] br[25] wl[218] vdd gnd cell_6t
Xbit_r219_c25 bl[25] br[25] wl[219] vdd gnd cell_6t
Xbit_r220_c25 bl[25] br[25] wl[220] vdd gnd cell_6t
Xbit_r221_c25 bl[25] br[25] wl[221] vdd gnd cell_6t
Xbit_r222_c25 bl[25] br[25] wl[222] vdd gnd cell_6t
Xbit_r223_c25 bl[25] br[25] wl[223] vdd gnd cell_6t
Xbit_r224_c25 bl[25] br[25] wl[224] vdd gnd cell_6t
Xbit_r225_c25 bl[25] br[25] wl[225] vdd gnd cell_6t
Xbit_r226_c25 bl[25] br[25] wl[226] vdd gnd cell_6t
Xbit_r227_c25 bl[25] br[25] wl[227] vdd gnd cell_6t
Xbit_r228_c25 bl[25] br[25] wl[228] vdd gnd cell_6t
Xbit_r229_c25 bl[25] br[25] wl[229] vdd gnd cell_6t
Xbit_r230_c25 bl[25] br[25] wl[230] vdd gnd cell_6t
Xbit_r231_c25 bl[25] br[25] wl[231] vdd gnd cell_6t
Xbit_r232_c25 bl[25] br[25] wl[232] vdd gnd cell_6t
Xbit_r233_c25 bl[25] br[25] wl[233] vdd gnd cell_6t
Xbit_r234_c25 bl[25] br[25] wl[234] vdd gnd cell_6t
Xbit_r235_c25 bl[25] br[25] wl[235] vdd gnd cell_6t
Xbit_r236_c25 bl[25] br[25] wl[236] vdd gnd cell_6t
Xbit_r237_c25 bl[25] br[25] wl[237] vdd gnd cell_6t
Xbit_r238_c25 bl[25] br[25] wl[238] vdd gnd cell_6t
Xbit_r239_c25 bl[25] br[25] wl[239] vdd gnd cell_6t
Xbit_r240_c25 bl[25] br[25] wl[240] vdd gnd cell_6t
Xbit_r241_c25 bl[25] br[25] wl[241] vdd gnd cell_6t
Xbit_r242_c25 bl[25] br[25] wl[242] vdd gnd cell_6t
Xbit_r243_c25 bl[25] br[25] wl[243] vdd gnd cell_6t
Xbit_r244_c25 bl[25] br[25] wl[244] vdd gnd cell_6t
Xbit_r245_c25 bl[25] br[25] wl[245] vdd gnd cell_6t
Xbit_r246_c25 bl[25] br[25] wl[246] vdd gnd cell_6t
Xbit_r247_c25 bl[25] br[25] wl[247] vdd gnd cell_6t
Xbit_r248_c25 bl[25] br[25] wl[248] vdd gnd cell_6t
Xbit_r249_c25 bl[25] br[25] wl[249] vdd gnd cell_6t
Xbit_r250_c25 bl[25] br[25] wl[250] vdd gnd cell_6t
Xbit_r251_c25 bl[25] br[25] wl[251] vdd gnd cell_6t
Xbit_r252_c25 bl[25] br[25] wl[252] vdd gnd cell_6t
Xbit_r253_c25 bl[25] br[25] wl[253] vdd gnd cell_6t
Xbit_r254_c25 bl[25] br[25] wl[254] vdd gnd cell_6t
Xbit_r255_c25 bl[25] br[25] wl[255] vdd gnd cell_6t
Xbit_r0_c26 bl[26] br[26] wl[0] vdd gnd cell_6t
Xbit_r1_c26 bl[26] br[26] wl[1] vdd gnd cell_6t
Xbit_r2_c26 bl[26] br[26] wl[2] vdd gnd cell_6t
Xbit_r3_c26 bl[26] br[26] wl[3] vdd gnd cell_6t
Xbit_r4_c26 bl[26] br[26] wl[4] vdd gnd cell_6t
Xbit_r5_c26 bl[26] br[26] wl[5] vdd gnd cell_6t
Xbit_r6_c26 bl[26] br[26] wl[6] vdd gnd cell_6t
Xbit_r7_c26 bl[26] br[26] wl[7] vdd gnd cell_6t
Xbit_r8_c26 bl[26] br[26] wl[8] vdd gnd cell_6t
Xbit_r9_c26 bl[26] br[26] wl[9] vdd gnd cell_6t
Xbit_r10_c26 bl[26] br[26] wl[10] vdd gnd cell_6t
Xbit_r11_c26 bl[26] br[26] wl[11] vdd gnd cell_6t
Xbit_r12_c26 bl[26] br[26] wl[12] vdd gnd cell_6t
Xbit_r13_c26 bl[26] br[26] wl[13] vdd gnd cell_6t
Xbit_r14_c26 bl[26] br[26] wl[14] vdd gnd cell_6t
Xbit_r15_c26 bl[26] br[26] wl[15] vdd gnd cell_6t
Xbit_r16_c26 bl[26] br[26] wl[16] vdd gnd cell_6t
Xbit_r17_c26 bl[26] br[26] wl[17] vdd gnd cell_6t
Xbit_r18_c26 bl[26] br[26] wl[18] vdd gnd cell_6t
Xbit_r19_c26 bl[26] br[26] wl[19] vdd gnd cell_6t
Xbit_r20_c26 bl[26] br[26] wl[20] vdd gnd cell_6t
Xbit_r21_c26 bl[26] br[26] wl[21] vdd gnd cell_6t
Xbit_r22_c26 bl[26] br[26] wl[22] vdd gnd cell_6t
Xbit_r23_c26 bl[26] br[26] wl[23] vdd gnd cell_6t
Xbit_r24_c26 bl[26] br[26] wl[24] vdd gnd cell_6t
Xbit_r25_c26 bl[26] br[26] wl[25] vdd gnd cell_6t
Xbit_r26_c26 bl[26] br[26] wl[26] vdd gnd cell_6t
Xbit_r27_c26 bl[26] br[26] wl[27] vdd gnd cell_6t
Xbit_r28_c26 bl[26] br[26] wl[28] vdd gnd cell_6t
Xbit_r29_c26 bl[26] br[26] wl[29] vdd gnd cell_6t
Xbit_r30_c26 bl[26] br[26] wl[30] vdd gnd cell_6t
Xbit_r31_c26 bl[26] br[26] wl[31] vdd gnd cell_6t
Xbit_r32_c26 bl[26] br[26] wl[32] vdd gnd cell_6t
Xbit_r33_c26 bl[26] br[26] wl[33] vdd gnd cell_6t
Xbit_r34_c26 bl[26] br[26] wl[34] vdd gnd cell_6t
Xbit_r35_c26 bl[26] br[26] wl[35] vdd gnd cell_6t
Xbit_r36_c26 bl[26] br[26] wl[36] vdd gnd cell_6t
Xbit_r37_c26 bl[26] br[26] wl[37] vdd gnd cell_6t
Xbit_r38_c26 bl[26] br[26] wl[38] vdd gnd cell_6t
Xbit_r39_c26 bl[26] br[26] wl[39] vdd gnd cell_6t
Xbit_r40_c26 bl[26] br[26] wl[40] vdd gnd cell_6t
Xbit_r41_c26 bl[26] br[26] wl[41] vdd gnd cell_6t
Xbit_r42_c26 bl[26] br[26] wl[42] vdd gnd cell_6t
Xbit_r43_c26 bl[26] br[26] wl[43] vdd gnd cell_6t
Xbit_r44_c26 bl[26] br[26] wl[44] vdd gnd cell_6t
Xbit_r45_c26 bl[26] br[26] wl[45] vdd gnd cell_6t
Xbit_r46_c26 bl[26] br[26] wl[46] vdd gnd cell_6t
Xbit_r47_c26 bl[26] br[26] wl[47] vdd gnd cell_6t
Xbit_r48_c26 bl[26] br[26] wl[48] vdd gnd cell_6t
Xbit_r49_c26 bl[26] br[26] wl[49] vdd gnd cell_6t
Xbit_r50_c26 bl[26] br[26] wl[50] vdd gnd cell_6t
Xbit_r51_c26 bl[26] br[26] wl[51] vdd gnd cell_6t
Xbit_r52_c26 bl[26] br[26] wl[52] vdd gnd cell_6t
Xbit_r53_c26 bl[26] br[26] wl[53] vdd gnd cell_6t
Xbit_r54_c26 bl[26] br[26] wl[54] vdd gnd cell_6t
Xbit_r55_c26 bl[26] br[26] wl[55] vdd gnd cell_6t
Xbit_r56_c26 bl[26] br[26] wl[56] vdd gnd cell_6t
Xbit_r57_c26 bl[26] br[26] wl[57] vdd gnd cell_6t
Xbit_r58_c26 bl[26] br[26] wl[58] vdd gnd cell_6t
Xbit_r59_c26 bl[26] br[26] wl[59] vdd gnd cell_6t
Xbit_r60_c26 bl[26] br[26] wl[60] vdd gnd cell_6t
Xbit_r61_c26 bl[26] br[26] wl[61] vdd gnd cell_6t
Xbit_r62_c26 bl[26] br[26] wl[62] vdd gnd cell_6t
Xbit_r63_c26 bl[26] br[26] wl[63] vdd gnd cell_6t
Xbit_r64_c26 bl[26] br[26] wl[64] vdd gnd cell_6t
Xbit_r65_c26 bl[26] br[26] wl[65] vdd gnd cell_6t
Xbit_r66_c26 bl[26] br[26] wl[66] vdd gnd cell_6t
Xbit_r67_c26 bl[26] br[26] wl[67] vdd gnd cell_6t
Xbit_r68_c26 bl[26] br[26] wl[68] vdd gnd cell_6t
Xbit_r69_c26 bl[26] br[26] wl[69] vdd gnd cell_6t
Xbit_r70_c26 bl[26] br[26] wl[70] vdd gnd cell_6t
Xbit_r71_c26 bl[26] br[26] wl[71] vdd gnd cell_6t
Xbit_r72_c26 bl[26] br[26] wl[72] vdd gnd cell_6t
Xbit_r73_c26 bl[26] br[26] wl[73] vdd gnd cell_6t
Xbit_r74_c26 bl[26] br[26] wl[74] vdd gnd cell_6t
Xbit_r75_c26 bl[26] br[26] wl[75] vdd gnd cell_6t
Xbit_r76_c26 bl[26] br[26] wl[76] vdd gnd cell_6t
Xbit_r77_c26 bl[26] br[26] wl[77] vdd gnd cell_6t
Xbit_r78_c26 bl[26] br[26] wl[78] vdd gnd cell_6t
Xbit_r79_c26 bl[26] br[26] wl[79] vdd gnd cell_6t
Xbit_r80_c26 bl[26] br[26] wl[80] vdd gnd cell_6t
Xbit_r81_c26 bl[26] br[26] wl[81] vdd gnd cell_6t
Xbit_r82_c26 bl[26] br[26] wl[82] vdd gnd cell_6t
Xbit_r83_c26 bl[26] br[26] wl[83] vdd gnd cell_6t
Xbit_r84_c26 bl[26] br[26] wl[84] vdd gnd cell_6t
Xbit_r85_c26 bl[26] br[26] wl[85] vdd gnd cell_6t
Xbit_r86_c26 bl[26] br[26] wl[86] vdd gnd cell_6t
Xbit_r87_c26 bl[26] br[26] wl[87] vdd gnd cell_6t
Xbit_r88_c26 bl[26] br[26] wl[88] vdd gnd cell_6t
Xbit_r89_c26 bl[26] br[26] wl[89] vdd gnd cell_6t
Xbit_r90_c26 bl[26] br[26] wl[90] vdd gnd cell_6t
Xbit_r91_c26 bl[26] br[26] wl[91] vdd gnd cell_6t
Xbit_r92_c26 bl[26] br[26] wl[92] vdd gnd cell_6t
Xbit_r93_c26 bl[26] br[26] wl[93] vdd gnd cell_6t
Xbit_r94_c26 bl[26] br[26] wl[94] vdd gnd cell_6t
Xbit_r95_c26 bl[26] br[26] wl[95] vdd gnd cell_6t
Xbit_r96_c26 bl[26] br[26] wl[96] vdd gnd cell_6t
Xbit_r97_c26 bl[26] br[26] wl[97] vdd gnd cell_6t
Xbit_r98_c26 bl[26] br[26] wl[98] vdd gnd cell_6t
Xbit_r99_c26 bl[26] br[26] wl[99] vdd gnd cell_6t
Xbit_r100_c26 bl[26] br[26] wl[100] vdd gnd cell_6t
Xbit_r101_c26 bl[26] br[26] wl[101] vdd gnd cell_6t
Xbit_r102_c26 bl[26] br[26] wl[102] vdd gnd cell_6t
Xbit_r103_c26 bl[26] br[26] wl[103] vdd gnd cell_6t
Xbit_r104_c26 bl[26] br[26] wl[104] vdd gnd cell_6t
Xbit_r105_c26 bl[26] br[26] wl[105] vdd gnd cell_6t
Xbit_r106_c26 bl[26] br[26] wl[106] vdd gnd cell_6t
Xbit_r107_c26 bl[26] br[26] wl[107] vdd gnd cell_6t
Xbit_r108_c26 bl[26] br[26] wl[108] vdd gnd cell_6t
Xbit_r109_c26 bl[26] br[26] wl[109] vdd gnd cell_6t
Xbit_r110_c26 bl[26] br[26] wl[110] vdd gnd cell_6t
Xbit_r111_c26 bl[26] br[26] wl[111] vdd gnd cell_6t
Xbit_r112_c26 bl[26] br[26] wl[112] vdd gnd cell_6t
Xbit_r113_c26 bl[26] br[26] wl[113] vdd gnd cell_6t
Xbit_r114_c26 bl[26] br[26] wl[114] vdd gnd cell_6t
Xbit_r115_c26 bl[26] br[26] wl[115] vdd gnd cell_6t
Xbit_r116_c26 bl[26] br[26] wl[116] vdd gnd cell_6t
Xbit_r117_c26 bl[26] br[26] wl[117] vdd gnd cell_6t
Xbit_r118_c26 bl[26] br[26] wl[118] vdd gnd cell_6t
Xbit_r119_c26 bl[26] br[26] wl[119] vdd gnd cell_6t
Xbit_r120_c26 bl[26] br[26] wl[120] vdd gnd cell_6t
Xbit_r121_c26 bl[26] br[26] wl[121] vdd gnd cell_6t
Xbit_r122_c26 bl[26] br[26] wl[122] vdd gnd cell_6t
Xbit_r123_c26 bl[26] br[26] wl[123] vdd gnd cell_6t
Xbit_r124_c26 bl[26] br[26] wl[124] vdd gnd cell_6t
Xbit_r125_c26 bl[26] br[26] wl[125] vdd gnd cell_6t
Xbit_r126_c26 bl[26] br[26] wl[126] vdd gnd cell_6t
Xbit_r127_c26 bl[26] br[26] wl[127] vdd gnd cell_6t
Xbit_r128_c26 bl[26] br[26] wl[128] vdd gnd cell_6t
Xbit_r129_c26 bl[26] br[26] wl[129] vdd gnd cell_6t
Xbit_r130_c26 bl[26] br[26] wl[130] vdd gnd cell_6t
Xbit_r131_c26 bl[26] br[26] wl[131] vdd gnd cell_6t
Xbit_r132_c26 bl[26] br[26] wl[132] vdd gnd cell_6t
Xbit_r133_c26 bl[26] br[26] wl[133] vdd gnd cell_6t
Xbit_r134_c26 bl[26] br[26] wl[134] vdd gnd cell_6t
Xbit_r135_c26 bl[26] br[26] wl[135] vdd gnd cell_6t
Xbit_r136_c26 bl[26] br[26] wl[136] vdd gnd cell_6t
Xbit_r137_c26 bl[26] br[26] wl[137] vdd gnd cell_6t
Xbit_r138_c26 bl[26] br[26] wl[138] vdd gnd cell_6t
Xbit_r139_c26 bl[26] br[26] wl[139] vdd gnd cell_6t
Xbit_r140_c26 bl[26] br[26] wl[140] vdd gnd cell_6t
Xbit_r141_c26 bl[26] br[26] wl[141] vdd gnd cell_6t
Xbit_r142_c26 bl[26] br[26] wl[142] vdd gnd cell_6t
Xbit_r143_c26 bl[26] br[26] wl[143] vdd gnd cell_6t
Xbit_r144_c26 bl[26] br[26] wl[144] vdd gnd cell_6t
Xbit_r145_c26 bl[26] br[26] wl[145] vdd gnd cell_6t
Xbit_r146_c26 bl[26] br[26] wl[146] vdd gnd cell_6t
Xbit_r147_c26 bl[26] br[26] wl[147] vdd gnd cell_6t
Xbit_r148_c26 bl[26] br[26] wl[148] vdd gnd cell_6t
Xbit_r149_c26 bl[26] br[26] wl[149] vdd gnd cell_6t
Xbit_r150_c26 bl[26] br[26] wl[150] vdd gnd cell_6t
Xbit_r151_c26 bl[26] br[26] wl[151] vdd gnd cell_6t
Xbit_r152_c26 bl[26] br[26] wl[152] vdd gnd cell_6t
Xbit_r153_c26 bl[26] br[26] wl[153] vdd gnd cell_6t
Xbit_r154_c26 bl[26] br[26] wl[154] vdd gnd cell_6t
Xbit_r155_c26 bl[26] br[26] wl[155] vdd gnd cell_6t
Xbit_r156_c26 bl[26] br[26] wl[156] vdd gnd cell_6t
Xbit_r157_c26 bl[26] br[26] wl[157] vdd gnd cell_6t
Xbit_r158_c26 bl[26] br[26] wl[158] vdd gnd cell_6t
Xbit_r159_c26 bl[26] br[26] wl[159] vdd gnd cell_6t
Xbit_r160_c26 bl[26] br[26] wl[160] vdd gnd cell_6t
Xbit_r161_c26 bl[26] br[26] wl[161] vdd gnd cell_6t
Xbit_r162_c26 bl[26] br[26] wl[162] vdd gnd cell_6t
Xbit_r163_c26 bl[26] br[26] wl[163] vdd gnd cell_6t
Xbit_r164_c26 bl[26] br[26] wl[164] vdd gnd cell_6t
Xbit_r165_c26 bl[26] br[26] wl[165] vdd gnd cell_6t
Xbit_r166_c26 bl[26] br[26] wl[166] vdd gnd cell_6t
Xbit_r167_c26 bl[26] br[26] wl[167] vdd gnd cell_6t
Xbit_r168_c26 bl[26] br[26] wl[168] vdd gnd cell_6t
Xbit_r169_c26 bl[26] br[26] wl[169] vdd gnd cell_6t
Xbit_r170_c26 bl[26] br[26] wl[170] vdd gnd cell_6t
Xbit_r171_c26 bl[26] br[26] wl[171] vdd gnd cell_6t
Xbit_r172_c26 bl[26] br[26] wl[172] vdd gnd cell_6t
Xbit_r173_c26 bl[26] br[26] wl[173] vdd gnd cell_6t
Xbit_r174_c26 bl[26] br[26] wl[174] vdd gnd cell_6t
Xbit_r175_c26 bl[26] br[26] wl[175] vdd gnd cell_6t
Xbit_r176_c26 bl[26] br[26] wl[176] vdd gnd cell_6t
Xbit_r177_c26 bl[26] br[26] wl[177] vdd gnd cell_6t
Xbit_r178_c26 bl[26] br[26] wl[178] vdd gnd cell_6t
Xbit_r179_c26 bl[26] br[26] wl[179] vdd gnd cell_6t
Xbit_r180_c26 bl[26] br[26] wl[180] vdd gnd cell_6t
Xbit_r181_c26 bl[26] br[26] wl[181] vdd gnd cell_6t
Xbit_r182_c26 bl[26] br[26] wl[182] vdd gnd cell_6t
Xbit_r183_c26 bl[26] br[26] wl[183] vdd gnd cell_6t
Xbit_r184_c26 bl[26] br[26] wl[184] vdd gnd cell_6t
Xbit_r185_c26 bl[26] br[26] wl[185] vdd gnd cell_6t
Xbit_r186_c26 bl[26] br[26] wl[186] vdd gnd cell_6t
Xbit_r187_c26 bl[26] br[26] wl[187] vdd gnd cell_6t
Xbit_r188_c26 bl[26] br[26] wl[188] vdd gnd cell_6t
Xbit_r189_c26 bl[26] br[26] wl[189] vdd gnd cell_6t
Xbit_r190_c26 bl[26] br[26] wl[190] vdd gnd cell_6t
Xbit_r191_c26 bl[26] br[26] wl[191] vdd gnd cell_6t
Xbit_r192_c26 bl[26] br[26] wl[192] vdd gnd cell_6t
Xbit_r193_c26 bl[26] br[26] wl[193] vdd gnd cell_6t
Xbit_r194_c26 bl[26] br[26] wl[194] vdd gnd cell_6t
Xbit_r195_c26 bl[26] br[26] wl[195] vdd gnd cell_6t
Xbit_r196_c26 bl[26] br[26] wl[196] vdd gnd cell_6t
Xbit_r197_c26 bl[26] br[26] wl[197] vdd gnd cell_6t
Xbit_r198_c26 bl[26] br[26] wl[198] vdd gnd cell_6t
Xbit_r199_c26 bl[26] br[26] wl[199] vdd gnd cell_6t
Xbit_r200_c26 bl[26] br[26] wl[200] vdd gnd cell_6t
Xbit_r201_c26 bl[26] br[26] wl[201] vdd gnd cell_6t
Xbit_r202_c26 bl[26] br[26] wl[202] vdd gnd cell_6t
Xbit_r203_c26 bl[26] br[26] wl[203] vdd gnd cell_6t
Xbit_r204_c26 bl[26] br[26] wl[204] vdd gnd cell_6t
Xbit_r205_c26 bl[26] br[26] wl[205] vdd gnd cell_6t
Xbit_r206_c26 bl[26] br[26] wl[206] vdd gnd cell_6t
Xbit_r207_c26 bl[26] br[26] wl[207] vdd gnd cell_6t
Xbit_r208_c26 bl[26] br[26] wl[208] vdd gnd cell_6t
Xbit_r209_c26 bl[26] br[26] wl[209] vdd gnd cell_6t
Xbit_r210_c26 bl[26] br[26] wl[210] vdd gnd cell_6t
Xbit_r211_c26 bl[26] br[26] wl[211] vdd gnd cell_6t
Xbit_r212_c26 bl[26] br[26] wl[212] vdd gnd cell_6t
Xbit_r213_c26 bl[26] br[26] wl[213] vdd gnd cell_6t
Xbit_r214_c26 bl[26] br[26] wl[214] vdd gnd cell_6t
Xbit_r215_c26 bl[26] br[26] wl[215] vdd gnd cell_6t
Xbit_r216_c26 bl[26] br[26] wl[216] vdd gnd cell_6t
Xbit_r217_c26 bl[26] br[26] wl[217] vdd gnd cell_6t
Xbit_r218_c26 bl[26] br[26] wl[218] vdd gnd cell_6t
Xbit_r219_c26 bl[26] br[26] wl[219] vdd gnd cell_6t
Xbit_r220_c26 bl[26] br[26] wl[220] vdd gnd cell_6t
Xbit_r221_c26 bl[26] br[26] wl[221] vdd gnd cell_6t
Xbit_r222_c26 bl[26] br[26] wl[222] vdd gnd cell_6t
Xbit_r223_c26 bl[26] br[26] wl[223] vdd gnd cell_6t
Xbit_r224_c26 bl[26] br[26] wl[224] vdd gnd cell_6t
Xbit_r225_c26 bl[26] br[26] wl[225] vdd gnd cell_6t
Xbit_r226_c26 bl[26] br[26] wl[226] vdd gnd cell_6t
Xbit_r227_c26 bl[26] br[26] wl[227] vdd gnd cell_6t
Xbit_r228_c26 bl[26] br[26] wl[228] vdd gnd cell_6t
Xbit_r229_c26 bl[26] br[26] wl[229] vdd gnd cell_6t
Xbit_r230_c26 bl[26] br[26] wl[230] vdd gnd cell_6t
Xbit_r231_c26 bl[26] br[26] wl[231] vdd gnd cell_6t
Xbit_r232_c26 bl[26] br[26] wl[232] vdd gnd cell_6t
Xbit_r233_c26 bl[26] br[26] wl[233] vdd gnd cell_6t
Xbit_r234_c26 bl[26] br[26] wl[234] vdd gnd cell_6t
Xbit_r235_c26 bl[26] br[26] wl[235] vdd gnd cell_6t
Xbit_r236_c26 bl[26] br[26] wl[236] vdd gnd cell_6t
Xbit_r237_c26 bl[26] br[26] wl[237] vdd gnd cell_6t
Xbit_r238_c26 bl[26] br[26] wl[238] vdd gnd cell_6t
Xbit_r239_c26 bl[26] br[26] wl[239] vdd gnd cell_6t
Xbit_r240_c26 bl[26] br[26] wl[240] vdd gnd cell_6t
Xbit_r241_c26 bl[26] br[26] wl[241] vdd gnd cell_6t
Xbit_r242_c26 bl[26] br[26] wl[242] vdd gnd cell_6t
Xbit_r243_c26 bl[26] br[26] wl[243] vdd gnd cell_6t
Xbit_r244_c26 bl[26] br[26] wl[244] vdd gnd cell_6t
Xbit_r245_c26 bl[26] br[26] wl[245] vdd gnd cell_6t
Xbit_r246_c26 bl[26] br[26] wl[246] vdd gnd cell_6t
Xbit_r247_c26 bl[26] br[26] wl[247] vdd gnd cell_6t
Xbit_r248_c26 bl[26] br[26] wl[248] vdd gnd cell_6t
Xbit_r249_c26 bl[26] br[26] wl[249] vdd gnd cell_6t
Xbit_r250_c26 bl[26] br[26] wl[250] vdd gnd cell_6t
Xbit_r251_c26 bl[26] br[26] wl[251] vdd gnd cell_6t
Xbit_r252_c26 bl[26] br[26] wl[252] vdd gnd cell_6t
Xbit_r253_c26 bl[26] br[26] wl[253] vdd gnd cell_6t
Xbit_r254_c26 bl[26] br[26] wl[254] vdd gnd cell_6t
Xbit_r255_c26 bl[26] br[26] wl[255] vdd gnd cell_6t
Xbit_r0_c27 bl[27] br[27] wl[0] vdd gnd cell_6t
Xbit_r1_c27 bl[27] br[27] wl[1] vdd gnd cell_6t
Xbit_r2_c27 bl[27] br[27] wl[2] vdd gnd cell_6t
Xbit_r3_c27 bl[27] br[27] wl[3] vdd gnd cell_6t
Xbit_r4_c27 bl[27] br[27] wl[4] vdd gnd cell_6t
Xbit_r5_c27 bl[27] br[27] wl[5] vdd gnd cell_6t
Xbit_r6_c27 bl[27] br[27] wl[6] vdd gnd cell_6t
Xbit_r7_c27 bl[27] br[27] wl[7] vdd gnd cell_6t
Xbit_r8_c27 bl[27] br[27] wl[8] vdd gnd cell_6t
Xbit_r9_c27 bl[27] br[27] wl[9] vdd gnd cell_6t
Xbit_r10_c27 bl[27] br[27] wl[10] vdd gnd cell_6t
Xbit_r11_c27 bl[27] br[27] wl[11] vdd gnd cell_6t
Xbit_r12_c27 bl[27] br[27] wl[12] vdd gnd cell_6t
Xbit_r13_c27 bl[27] br[27] wl[13] vdd gnd cell_6t
Xbit_r14_c27 bl[27] br[27] wl[14] vdd gnd cell_6t
Xbit_r15_c27 bl[27] br[27] wl[15] vdd gnd cell_6t
Xbit_r16_c27 bl[27] br[27] wl[16] vdd gnd cell_6t
Xbit_r17_c27 bl[27] br[27] wl[17] vdd gnd cell_6t
Xbit_r18_c27 bl[27] br[27] wl[18] vdd gnd cell_6t
Xbit_r19_c27 bl[27] br[27] wl[19] vdd gnd cell_6t
Xbit_r20_c27 bl[27] br[27] wl[20] vdd gnd cell_6t
Xbit_r21_c27 bl[27] br[27] wl[21] vdd gnd cell_6t
Xbit_r22_c27 bl[27] br[27] wl[22] vdd gnd cell_6t
Xbit_r23_c27 bl[27] br[27] wl[23] vdd gnd cell_6t
Xbit_r24_c27 bl[27] br[27] wl[24] vdd gnd cell_6t
Xbit_r25_c27 bl[27] br[27] wl[25] vdd gnd cell_6t
Xbit_r26_c27 bl[27] br[27] wl[26] vdd gnd cell_6t
Xbit_r27_c27 bl[27] br[27] wl[27] vdd gnd cell_6t
Xbit_r28_c27 bl[27] br[27] wl[28] vdd gnd cell_6t
Xbit_r29_c27 bl[27] br[27] wl[29] vdd gnd cell_6t
Xbit_r30_c27 bl[27] br[27] wl[30] vdd gnd cell_6t
Xbit_r31_c27 bl[27] br[27] wl[31] vdd gnd cell_6t
Xbit_r32_c27 bl[27] br[27] wl[32] vdd gnd cell_6t
Xbit_r33_c27 bl[27] br[27] wl[33] vdd gnd cell_6t
Xbit_r34_c27 bl[27] br[27] wl[34] vdd gnd cell_6t
Xbit_r35_c27 bl[27] br[27] wl[35] vdd gnd cell_6t
Xbit_r36_c27 bl[27] br[27] wl[36] vdd gnd cell_6t
Xbit_r37_c27 bl[27] br[27] wl[37] vdd gnd cell_6t
Xbit_r38_c27 bl[27] br[27] wl[38] vdd gnd cell_6t
Xbit_r39_c27 bl[27] br[27] wl[39] vdd gnd cell_6t
Xbit_r40_c27 bl[27] br[27] wl[40] vdd gnd cell_6t
Xbit_r41_c27 bl[27] br[27] wl[41] vdd gnd cell_6t
Xbit_r42_c27 bl[27] br[27] wl[42] vdd gnd cell_6t
Xbit_r43_c27 bl[27] br[27] wl[43] vdd gnd cell_6t
Xbit_r44_c27 bl[27] br[27] wl[44] vdd gnd cell_6t
Xbit_r45_c27 bl[27] br[27] wl[45] vdd gnd cell_6t
Xbit_r46_c27 bl[27] br[27] wl[46] vdd gnd cell_6t
Xbit_r47_c27 bl[27] br[27] wl[47] vdd gnd cell_6t
Xbit_r48_c27 bl[27] br[27] wl[48] vdd gnd cell_6t
Xbit_r49_c27 bl[27] br[27] wl[49] vdd gnd cell_6t
Xbit_r50_c27 bl[27] br[27] wl[50] vdd gnd cell_6t
Xbit_r51_c27 bl[27] br[27] wl[51] vdd gnd cell_6t
Xbit_r52_c27 bl[27] br[27] wl[52] vdd gnd cell_6t
Xbit_r53_c27 bl[27] br[27] wl[53] vdd gnd cell_6t
Xbit_r54_c27 bl[27] br[27] wl[54] vdd gnd cell_6t
Xbit_r55_c27 bl[27] br[27] wl[55] vdd gnd cell_6t
Xbit_r56_c27 bl[27] br[27] wl[56] vdd gnd cell_6t
Xbit_r57_c27 bl[27] br[27] wl[57] vdd gnd cell_6t
Xbit_r58_c27 bl[27] br[27] wl[58] vdd gnd cell_6t
Xbit_r59_c27 bl[27] br[27] wl[59] vdd gnd cell_6t
Xbit_r60_c27 bl[27] br[27] wl[60] vdd gnd cell_6t
Xbit_r61_c27 bl[27] br[27] wl[61] vdd gnd cell_6t
Xbit_r62_c27 bl[27] br[27] wl[62] vdd gnd cell_6t
Xbit_r63_c27 bl[27] br[27] wl[63] vdd gnd cell_6t
Xbit_r64_c27 bl[27] br[27] wl[64] vdd gnd cell_6t
Xbit_r65_c27 bl[27] br[27] wl[65] vdd gnd cell_6t
Xbit_r66_c27 bl[27] br[27] wl[66] vdd gnd cell_6t
Xbit_r67_c27 bl[27] br[27] wl[67] vdd gnd cell_6t
Xbit_r68_c27 bl[27] br[27] wl[68] vdd gnd cell_6t
Xbit_r69_c27 bl[27] br[27] wl[69] vdd gnd cell_6t
Xbit_r70_c27 bl[27] br[27] wl[70] vdd gnd cell_6t
Xbit_r71_c27 bl[27] br[27] wl[71] vdd gnd cell_6t
Xbit_r72_c27 bl[27] br[27] wl[72] vdd gnd cell_6t
Xbit_r73_c27 bl[27] br[27] wl[73] vdd gnd cell_6t
Xbit_r74_c27 bl[27] br[27] wl[74] vdd gnd cell_6t
Xbit_r75_c27 bl[27] br[27] wl[75] vdd gnd cell_6t
Xbit_r76_c27 bl[27] br[27] wl[76] vdd gnd cell_6t
Xbit_r77_c27 bl[27] br[27] wl[77] vdd gnd cell_6t
Xbit_r78_c27 bl[27] br[27] wl[78] vdd gnd cell_6t
Xbit_r79_c27 bl[27] br[27] wl[79] vdd gnd cell_6t
Xbit_r80_c27 bl[27] br[27] wl[80] vdd gnd cell_6t
Xbit_r81_c27 bl[27] br[27] wl[81] vdd gnd cell_6t
Xbit_r82_c27 bl[27] br[27] wl[82] vdd gnd cell_6t
Xbit_r83_c27 bl[27] br[27] wl[83] vdd gnd cell_6t
Xbit_r84_c27 bl[27] br[27] wl[84] vdd gnd cell_6t
Xbit_r85_c27 bl[27] br[27] wl[85] vdd gnd cell_6t
Xbit_r86_c27 bl[27] br[27] wl[86] vdd gnd cell_6t
Xbit_r87_c27 bl[27] br[27] wl[87] vdd gnd cell_6t
Xbit_r88_c27 bl[27] br[27] wl[88] vdd gnd cell_6t
Xbit_r89_c27 bl[27] br[27] wl[89] vdd gnd cell_6t
Xbit_r90_c27 bl[27] br[27] wl[90] vdd gnd cell_6t
Xbit_r91_c27 bl[27] br[27] wl[91] vdd gnd cell_6t
Xbit_r92_c27 bl[27] br[27] wl[92] vdd gnd cell_6t
Xbit_r93_c27 bl[27] br[27] wl[93] vdd gnd cell_6t
Xbit_r94_c27 bl[27] br[27] wl[94] vdd gnd cell_6t
Xbit_r95_c27 bl[27] br[27] wl[95] vdd gnd cell_6t
Xbit_r96_c27 bl[27] br[27] wl[96] vdd gnd cell_6t
Xbit_r97_c27 bl[27] br[27] wl[97] vdd gnd cell_6t
Xbit_r98_c27 bl[27] br[27] wl[98] vdd gnd cell_6t
Xbit_r99_c27 bl[27] br[27] wl[99] vdd gnd cell_6t
Xbit_r100_c27 bl[27] br[27] wl[100] vdd gnd cell_6t
Xbit_r101_c27 bl[27] br[27] wl[101] vdd gnd cell_6t
Xbit_r102_c27 bl[27] br[27] wl[102] vdd gnd cell_6t
Xbit_r103_c27 bl[27] br[27] wl[103] vdd gnd cell_6t
Xbit_r104_c27 bl[27] br[27] wl[104] vdd gnd cell_6t
Xbit_r105_c27 bl[27] br[27] wl[105] vdd gnd cell_6t
Xbit_r106_c27 bl[27] br[27] wl[106] vdd gnd cell_6t
Xbit_r107_c27 bl[27] br[27] wl[107] vdd gnd cell_6t
Xbit_r108_c27 bl[27] br[27] wl[108] vdd gnd cell_6t
Xbit_r109_c27 bl[27] br[27] wl[109] vdd gnd cell_6t
Xbit_r110_c27 bl[27] br[27] wl[110] vdd gnd cell_6t
Xbit_r111_c27 bl[27] br[27] wl[111] vdd gnd cell_6t
Xbit_r112_c27 bl[27] br[27] wl[112] vdd gnd cell_6t
Xbit_r113_c27 bl[27] br[27] wl[113] vdd gnd cell_6t
Xbit_r114_c27 bl[27] br[27] wl[114] vdd gnd cell_6t
Xbit_r115_c27 bl[27] br[27] wl[115] vdd gnd cell_6t
Xbit_r116_c27 bl[27] br[27] wl[116] vdd gnd cell_6t
Xbit_r117_c27 bl[27] br[27] wl[117] vdd gnd cell_6t
Xbit_r118_c27 bl[27] br[27] wl[118] vdd gnd cell_6t
Xbit_r119_c27 bl[27] br[27] wl[119] vdd gnd cell_6t
Xbit_r120_c27 bl[27] br[27] wl[120] vdd gnd cell_6t
Xbit_r121_c27 bl[27] br[27] wl[121] vdd gnd cell_6t
Xbit_r122_c27 bl[27] br[27] wl[122] vdd gnd cell_6t
Xbit_r123_c27 bl[27] br[27] wl[123] vdd gnd cell_6t
Xbit_r124_c27 bl[27] br[27] wl[124] vdd gnd cell_6t
Xbit_r125_c27 bl[27] br[27] wl[125] vdd gnd cell_6t
Xbit_r126_c27 bl[27] br[27] wl[126] vdd gnd cell_6t
Xbit_r127_c27 bl[27] br[27] wl[127] vdd gnd cell_6t
Xbit_r128_c27 bl[27] br[27] wl[128] vdd gnd cell_6t
Xbit_r129_c27 bl[27] br[27] wl[129] vdd gnd cell_6t
Xbit_r130_c27 bl[27] br[27] wl[130] vdd gnd cell_6t
Xbit_r131_c27 bl[27] br[27] wl[131] vdd gnd cell_6t
Xbit_r132_c27 bl[27] br[27] wl[132] vdd gnd cell_6t
Xbit_r133_c27 bl[27] br[27] wl[133] vdd gnd cell_6t
Xbit_r134_c27 bl[27] br[27] wl[134] vdd gnd cell_6t
Xbit_r135_c27 bl[27] br[27] wl[135] vdd gnd cell_6t
Xbit_r136_c27 bl[27] br[27] wl[136] vdd gnd cell_6t
Xbit_r137_c27 bl[27] br[27] wl[137] vdd gnd cell_6t
Xbit_r138_c27 bl[27] br[27] wl[138] vdd gnd cell_6t
Xbit_r139_c27 bl[27] br[27] wl[139] vdd gnd cell_6t
Xbit_r140_c27 bl[27] br[27] wl[140] vdd gnd cell_6t
Xbit_r141_c27 bl[27] br[27] wl[141] vdd gnd cell_6t
Xbit_r142_c27 bl[27] br[27] wl[142] vdd gnd cell_6t
Xbit_r143_c27 bl[27] br[27] wl[143] vdd gnd cell_6t
Xbit_r144_c27 bl[27] br[27] wl[144] vdd gnd cell_6t
Xbit_r145_c27 bl[27] br[27] wl[145] vdd gnd cell_6t
Xbit_r146_c27 bl[27] br[27] wl[146] vdd gnd cell_6t
Xbit_r147_c27 bl[27] br[27] wl[147] vdd gnd cell_6t
Xbit_r148_c27 bl[27] br[27] wl[148] vdd gnd cell_6t
Xbit_r149_c27 bl[27] br[27] wl[149] vdd gnd cell_6t
Xbit_r150_c27 bl[27] br[27] wl[150] vdd gnd cell_6t
Xbit_r151_c27 bl[27] br[27] wl[151] vdd gnd cell_6t
Xbit_r152_c27 bl[27] br[27] wl[152] vdd gnd cell_6t
Xbit_r153_c27 bl[27] br[27] wl[153] vdd gnd cell_6t
Xbit_r154_c27 bl[27] br[27] wl[154] vdd gnd cell_6t
Xbit_r155_c27 bl[27] br[27] wl[155] vdd gnd cell_6t
Xbit_r156_c27 bl[27] br[27] wl[156] vdd gnd cell_6t
Xbit_r157_c27 bl[27] br[27] wl[157] vdd gnd cell_6t
Xbit_r158_c27 bl[27] br[27] wl[158] vdd gnd cell_6t
Xbit_r159_c27 bl[27] br[27] wl[159] vdd gnd cell_6t
Xbit_r160_c27 bl[27] br[27] wl[160] vdd gnd cell_6t
Xbit_r161_c27 bl[27] br[27] wl[161] vdd gnd cell_6t
Xbit_r162_c27 bl[27] br[27] wl[162] vdd gnd cell_6t
Xbit_r163_c27 bl[27] br[27] wl[163] vdd gnd cell_6t
Xbit_r164_c27 bl[27] br[27] wl[164] vdd gnd cell_6t
Xbit_r165_c27 bl[27] br[27] wl[165] vdd gnd cell_6t
Xbit_r166_c27 bl[27] br[27] wl[166] vdd gnd cell_6t
Xbit_r167_c27 bl[27] br[27] wl[167] vdd gnd cell_6t
Xbit_r168_c27 bl[27] br[27] wl[168] vdd gnd cell_6t
Xbit_r169_c27 bl[27] br[27] wl[169] vdd gnd cell_6t
Xbit_r170_c27 bl[27] br[27] wl[170] vdd gnd cell_6t
Xbit_r171_c27 bl[27] br[27] wl[171] vdd gnd cell_6t
Xbit_r172_c27 bl[27] br[27] wl[172] vdd gnd cell_6t
Xbit_r173_c27 bl[27] br[27] wl[173] vdd gnd cell_6t
Xbit_r174_c27 bl[27] br[27] wl[174] vdd gnd cell_6t
Xbit_r175_c27 bl[27] br[27] wl[175] vdd gnd cell_6t
Xbit_r176_c27 bl[27] br[27] wl[176] vdd gnd cell_6t
Xbit_r177_c27 bl[27] br[27] wl[177] vdd gnd cell_6t
Xbit_r178_c27 bl[27] br[27] wl[178] vdd gnd cell_6t
Xbit_r179_c27 bl[27] br[27] wl[179] vdd gnd cell_6t
Xbit_r180_c27 bl[27] br[27] wl[180] vdd gnd cell_6t
Xbit_r181_c27 bl[27] br[27] wl[181] vdd gnd cell_6t
Xbit_r182_c27 bl[27] br[27] wl[182] vdd gnd cell_6t
Xbit_r183_c27 bl[27] br[27] wl[183] vdd gnd cell_6t
Xbit_r184_c27 bl[27] br[27] wl[184] vdd gnd cell_6t
Xbit_r185_c27 bl[27] br[27] wl[185] vdd gnd cell_6t
Xbit_r186_c27 bl[27] br[27] wl[186] vdd gnd cell_6t
Xbit_r187_c27 bl[27] br[27] wl[187] vdd gnd cell_6t
Xbit_r188_c27 bl[27] br[27] wl[188] vdd gnd cell_6t
Xbit_r189_c27 bl[27] br[27] wl[189] vdd gnd cell_6t
Xbit_r190_c27 bl[27] br[27] wl[190] vdd gnd cell_6t
Xbit_r191_c27 bl[27] br[27] wl[191] vdd gnd cell_6t
Xbit_r192_c27 bl[27] br[27] wl[192] vdd gnd cell_6t
Xbit_r193_c27 bl[27] br[27] wl[193] vdd gnd cell_6t
Xbit_r194_c27 bl[27] br[27] wl[194] vdd gnd cell_6t
Xbit_r195_c27 bl[27] br[27] wl[195] vdd gnd cell_6t
Xbit_r196_c27 bl[27] br[27] wl[196] vdd gnd cell_6t
Xbit_r197_c27 bl[27] br[27] wl[197] vdd gnd cell_6t
Xbit_r198_c27 bl[27] br[27] wl[198] vdd gnd cell_6t
Xbit_r199_c27 bl[27] br[27] wl[199] vdd gnd cell_6t
Xbit_r200_c27 bl[27] br[27] wl[200] vdd gnd cell_6t
Xbit_r201_c27 bl[27] br[27] wl[201] vdd gnd cell_6t
Xbit_r202_c27 bl[27] br[27] wl[202] vdd gnd cell_6t
Xbit_r203_c27 bl[27] br[27] wl[203] vdd gnd cell_6t
Xbit_r204_c27 bl[27] br[27] wl[204] vdd gnd cell_6t
Xbit_r205_c27 bl[27] br[27] wl[205] vdd gnd cell_6t
Xbit_r206_c27 bl[27] br[27] wl[206] vdd gnd cell_6t
Xbit_r207_c27 bl[27] br[27] wl[207] vdd gnd cell_6t
Xbit_r208_c27 bl[27] br[27] wl[208] vdd gnd cell_6t
Xbit_r209_c27 bl[27] br[27] wl[209] vdd gnd cell_6t
Xbit_r210_c27 bl[27] br[27] wl[210] vdd gnd cell_6t
Xbit_r211_c27 bl[27] br[27] wl[211] vdd gnd cell_6t
Xbit_r212_c27 bl[27] br[27] wl[212] vdd gnd cell_6t
Xbit_r213_c27 bl[27] br[27] wl[213] vdd gnd cell_6t
Xbit_r214_c27 bl[27] br[27] wl[214] vdd gnd cell_6t
Xbit_r215_c27 bl[27] br[27] wl[215] vdd gnd cell_6t
Xbit_r216_c27 bl[27] br[27] wl[216] vdd gnd cell_6t
Xbit_r217_c27 bl[27] br[27] wl[217] vdd gnd cell_6t
Xbit_r218_c27 bl[27] br[27] wl[218] vdd gnd cell_6t
Xbit_r219_c27 bl[27] br[27] wl[219] vdd gnd cell_6t
Xbit_r220_c27 bl[27] br[27] wl[220] vdd gnd cell_6t
Xbit_r221_c27 bl[27] br[27] wl[221] vdd gnd cell_6t
Xbit_r222_c27 bl[27] br[27] wl[222] vdd gnd cell_6t
Xbit_r223_c27 bl[27] br[27] wl[223] vdd gnd cell_6t
Xbit_r224_c27 bl[27] br[27] wl[224] vdd gnd cell_6t
Xbit_r225_c27 bl[27] br[27] wl[225] vdd gnd cell_6t
Xbit_r226_c27 bl[27] br[27] wl[226] vdd gnd cell_6t
Xbit_r227_c27 bl[27] br[27] wl[227] vdd gnd cell_6t
Xbit_r228_c27 bl[27] br[27] wl[228] vdd gnd cell_6t
Xbit_r229_c27 bl[27] br[27] wl[229] vdd gnd cell_6t
Xbit_r230_c27 bl[27] br[27] wl[230] vdd gnd cell_6t
Xbit_r231_c27 bl[27] br[27] wl[231] vdd gnd cell_6t
Xbit_r232_c27 bl[27] br[27] wl[232] vdd gnd cell_6t
Xbit_r233_c27 bl[27] br[27] wl[233] vdd gnd cell_6t
Xbit_r234_c27 bl[27] br[27] wl[234] vdd gnd cell_6t
Xbit_r235_c27 bl[27] br[27] wl[235] vdd gnd cell_6t
Xbit_r236_c27 bl[27] br[27] wl[236] vdd gnd cell_6t
Xbit_r237_c27 bl[27] br[27] wl[237] vdd gnd cell_6t
Xbit_r238_c27 bl[27] br[27] wl[238] vdd gnd cell_6t
Xbit_r239_c27 bl[27] br[27] wl[239] vdd gnd cell_6t
Xbit_r240_c27 bl[27] br[27] wl[240] vdd gnd cell_6t
Xbit_r241_c27 bl[27] br[27] wl[241] vdd gnd cell_6t
Xbit_r242_c27 bl[27] br[27] wl[242] vdd gnd cell_6t
Xbit_r243_c27 bl[27] br[27] wl[243] vdd gnd cell_6t
Xbit_r244_c27 bl[27] br[27] wl[244] vdd gnd cell_6t
Xbit_r245_c27 bl[27] br[27] wl[245] vdd gnd cell_6t
Xbit_r246_c27 bl[27] br[27] wl[246] vdd gnd cell_6t
Xbit_r247_c27 bl[27] br[27] wl[247] vdd gnd cell_6t
Xbit_r248_c27 bl[27] br[27] wl[248] vdd gnd cell_6t
Xbit_r249_c27 bl[27] br[27] wl[249] vdd gnd cell_6t
Xbit_r250_c27 bl[27] br[27] wl[250] vdd gnd cell_6t
Xbit_r251_c27 bl[27] br[27] wl[251] vdd gnd cell_6t
Xbit_r252_c27 bl[27] br[27] wl[252] vdd gnd cell_6t
Xbit_r253_c27 bl[27] br[27] wl[253] vdd gnd cell_6t
Xbit_r254_c27 bl[27] br[27] wl[254] vdd gnd cell_6t
Xbit_r255_c27 bl[27] br[27] wl[255] vdd gnd cell_6t
Xbit_r0_c28 bl[28] br[28] wl[0] vdd gnd cell_6t
Xbit_r1_c28 bl[28] br[28] wl[1] vdd gnd cell_6t
Xbit_r2_c28 bl[28] br[28] wl[2] vdd gnd cell_6t
Xbit_r3_c28 bl[28] br[28] wl[3] vdd gnd cell_6t
Xbit_r4_c28 bl[28] br[28] wl[4] vdd gnd cell_6t
Xbit_r5_c28 bl[28] br[28] wl[5] vdd gnd cell_6t
Xbit_r6_c28 bl[28] br[28] wl[6] vdd gnd cell_6t
Xbit_r7_c28 bl[28] br[28] wl[7] vdd gnd cell_6t
Xbit_r8_c28 bl[28] br[28] wl[8] vdd gnd cell_6t
Xbit_r9_c28 bl[28] br[28] wl[9] vdd gnd cell_6t
Xbit_r10_c28 bl[28] br[28] wl[10] vdd gnd cell_6t
Xbit_r11_c28 bl[28] br[28] wl[11] vdd gnd cell_6t
Xbit_r12_c28 bl[28] br[28] wl[12] vdd gnd cell_6t
Xbit_r13_c28 bl[28] br[28] wl[13] vdd gnd cell_6t
Xbit_r14_c28 bl[28] br[28] wl[14] vdd gnd cell_6t
Xbit_r15_c28 bl[28] br[28] wl[15] vdd gnd cell_6t
Xbit_r16_c28 bl[28] br[28] wl[16] vdd gnd cell_6t
Xbit_r17_c28 bl[28] br[28] wl[17] vdd gnd cell_6t
Xbit_r18_c28 bl[28] br[28] wl[18] vdd gnd cell_6t
Xbit_r19_c28 bl[28] br[28] wl[19] vdd gnd cell_6t
Xbit_r20_c28 bl[28] br[28] wl[20] vdd gnd cell_6t
Xbit_r21_c28 bl[28] br[28] wl[21] vdd gnd cell_6t
Xbit_r22_c28 bl[28] br[28] wl[22] vdd gnd cell_6t
Xbit_r23_c28 bl[28] br[28] wl[23] vdd gnd cell_6t
Xbit_r24_c28 bl[28] br[28] wl[24] vdd gnd cell_6t
Xbit_r25_c28 bl[28] br[28] wl[25] vdd gnd cell_6t
Xbit_r26_c28 bl[28] br[28] wl[26] vdd gnd cell_6t
Xbit_r27_c28 bl[28] br[28] wl[27] vdd gnd cell_6t
Xbit_r28_c28 bl[28] br[28] wl[28] vdd gnd cell_6t
Xbit_r29_c28 bl[28] br[28] wl[29] vdd gnd cell_6t
Xbit_r30_c28 bl[28] br[28] wl[30] vdd gnd cell_6t
Xbit_r31_c28 bl[28] br[28] wl[31] vdd gnd cell_6t
Xbit_r32_c28 bl[28] br[28] wl[32] vdd gnd cell_6t
Xbit_r33_c28 bl[28] br[28] wl[33] vdd gnd cell_6t
Xbit_r34_c28 bl[28] br[28] wl[34] vdd gnd cell_6t
Xbit_r35_c28 bl[28] br[28] wl[35] vdd gnd cell_6t
Xbit_r36_c28 bl[28] br[28] wl[36] vdd gnd cell_6t
Xbit_r37_c28 bl[28] br[28] wl[37] vdd gnd cell_6t
Xbit_r38_c28 bl[28] br[28] wl[38] vdd gnd cell_6t
Xbit_r39_c28 bl[28] br[28] wl[39] vdd gnd cell_6t
Xbit_r40_c28 bl[28] br[28] wl[40] vdd gnd cell_6t
Xbit_r41_c28 bl[28] br[28] wl[41] vdd gnd cell_6t
Xbit_r42_c28 bl[28] br[28] wl[42] vdd gnd cell_6t
Xbit_r43_c28 bl[28] br[28] wl[43] vdd gnd cell_6t
Xbit_r44_c28 bl[28] br[28] wl[44] vdd gnd cell_6t
Xbit_r45_c28 bl[28] br[28] wl[45] vdd gnd cell_6t
Xbit_r46_c28 bl[28] br[28] wl[46] vdd gnd cell_6t
Xbit_r47_c28 bl[28] br[28] wl[47] vdd gnd cell_6t
Xbit_r48_c28 bl[28] br[28] wl[48] vdd gnd cell_6t
Xbit_r49_c28 bl[28] br[28] wl[49] vdd gnd cell_6t
Xbit_r50_c28 bl[28] br[28] wl[50] vdd gnd cell_6t
Xbit_r51_c28 bl[28] br[28] wl[51] vdd gnd cell_6t
Xbit_r52_c28 bl[28] br[28] wl[52] vdd gnd cell_6t
Xbit_r53_c28 bl[28] br[28] wl[53] vdd gnd cell_6t
Xbit_r54_c28 bl[28] br[28] wl[54] vdd gnd cell_6t
Xbit_r55_c28 bl[28] br[28] wl[55] vdd gnd cell_6t
Xbit_r56_c28 bl[28] br[28] wl[56] vdd gnd cell_6t
Xbit_r57_c28 bl[28] br[28] wl[57] vdd gnd cell_6t
Xbit_r58_c28 bl[28] br[28] wl[58] vdd gnd cell_6t
Xbit_r59_c28 bl[28] br[28] wl[59] vdd gnd cell_6t
Xbit_r60_c28 bl[28] br[28] wl[60] vdd gnd cell_6t
Xbit_r61_c28 bl[28] br[28] wl[61] vdd gnd cell_6t
Xbit_r62_c28 bl[28] br[28] wl[62] vdd gnd cell_6t
Xbit_r63_c28 bl[28] br[28] wl[63] vdd gnd cell_6t
Xbit_r64_c28 bl[28] br[28] wl[64] vdd gnd cell_6t
Xbit_r65_c28 bl[28] br[28] wl[65] vdd gnd cell_6t
Xbit_r66_c28 bl[28] br[28] wl[66] vdd gnd cell_6t
Xbit_r67_c28 bl[28] br[28] wl[67] vdd gnd cell_6t
Xbit_r68_c28 bl[28] br[28] wl[68] vdd gnd cell_6t
Xbit_r69_c28 bl[28] br[28] wl[69] vdd gnd cell_6t
Xbit_r70_c28 bl[28] br[28] wl[70] vdd gnd cell_6t
Xbit_r71_c28 bl[28] br[28] wl[71] vdd gnd cell_6t
Xbit_r72_c28 bl[28] br[28] wl[72] vdd gnd cell_6t
Xbit_r73_c28 bl[28] br[28] wl[73] vdd gnd cell_6t
Xbit_r74_c28 bl[28] br[28] wl[74] vdd gnd cell_6t
Xbit_r75_c28 bl[28] br[28] wl[75] vdd gnd cell_6t
Xbit_r76_c28 bl[28] br[28] wl[76] vdd gnd cell_6t
Xbit_r77_c28 bl[28] br[28] wl[77] vdd gnd cell_6t
Xbit_r78_c28 bl[28] br[28] wl[78] vdd gnd cell_6t
Xbit_r79_c28 bl[28] br[28] wl[79] vdd gnd cell_6t
Xbit_r80_c28 bl[28] br[28] wl[80] vdd gnd cell_6t
Xbit_r81_c28 bl[28] br[28] wl[81] vdd gnd cell_6t
Xbit_r82_c28 bl[28] br[28] wl[82] vdd gnd cell_6t
Xbit_r83_c28 bl[28] br[28] wl[83] vdd gnd cell_6t
Xbit_r84_c28 bl[28] br[28] wl[84] vdd gnd cell_6t
Xbit_r85_c28 bl[28] br[28] wl[85] vdd gnd cell_6t
Xbit_r86_c28 bl[28] br[28] wl[86] vdd gnd cell_6t
Xbit_r87_c28 bl[28] br[28] wl[87] vdd gnd cell_6t
Xbit_r88_c28 bl[28] br[28] wl[88] vdd gnd cell_6t
Xbit_r89_c28 bl[28] br[28] wl[89] vdd gnd cell_6t
Xbit_r90_c28 bl[28] br[28] wl[90] vdd gnd cell_6t
Xbit_r91_c28 bl[28] br[28] wl[91] vdd gnd cell_6t
Xbit_r92_c28 bl[28] br[28] wl[92] vdd gnd cell_6t
Xbit_r93_c28 bl[28] br[28] wl[93] vdd gnd cell_6t
Xbit_r94_c28 bl[28] br[28] wl[94] vdd gnd cell_6t
Xbit_r95_c28 bl[28] br[28] wl[95] vdd gnd cell_6t
Xbit_r96_c28 bl[28] br[28] wl[96] vdd gnd cell_6t
Xbit_r97_c28 bl[28] br[28] wl[97] vdd gnd cell_6t
Xbit_r98_c28 bl[28] br[28] wl[98] vdd gnd cell_6t
Xbit_r99_c28 bl[28] br[28] wl[99] vdd gnd cell_6t
Xbit_r100_c28 bl[28] br[28] wl[100] vdd gnd cell_6t
Xbit_r101_c28 bl[28] br[28] wl[101] vdd gnd cell_6t
Xbit_r102_c28 bl[28] br[28] wl[102] vdd gnd cell_6t
Xbit_r103_c28 bl[28] br[28] wl[103] vdd gnd cell_6t
Xbit_r104_c28 bl[28] br[28] wl[104] vdd gnd cell_6t
Xbit_r105_c28 bl[28] br[28] wl[105] vdd gnd cell_6t
Xbit_r106_c28 bl[28] br[28] wl[106] vdd gnd cell_6t
Xbit_r107_c28 bl[28] br[28] wl[107] vdd gnd cell_6t
Xbit_r108_c28 bl[28] br[28] wl[108] vdd gnd cell_6t
Xbit_r109_c28 bl[28] br[28] wl[109] vdd gnd cell_6t
Xbit_r110_c28 bl[28] br[28] wl[110] vdd gnd cell_6t
Xbit_r111_c28 bl[28] br[28] wl[111] vdd gnd cell_6t
Xbit_r112_c28 bl[28] br[28] wl[112] vdd gnd cell_6t
Xbit_r113_c28 bl[28] br[28] wl[113] vdd gnd cell_6t
Xbit_r114_c28 bl[28] br[28] wl[114] vdd gnd cell_6t
Xbit_r115_c28 bl[28] br[28] wl[115] vdd gnd cell_6t
Xbit_r116_c28 bl[28] br[28] wl[116] vdd gnd cell_6t
Xbit_r117_c28 bl[28] br[28] wl[117] vdd gnd cell_6t
Xbit_r118_c28 bl[28] br[28] wl[118] vdd gnd cell_6t
Xbit_r119_c28 bl[28] br[28] wl[119] vdd gnd cell_6t
Xbit_r120_c28 bl[28] br[28] wl[120] vdd gnd cell_6t
Xbit_r121_c28 bl[28] br[28] wl[121] vdd gnd cell_6t
Xbit_r122_c28 bl[28] br[28] wl[122] vdd gnd cell_6t
Xbit_r123_c28 bl[28] br[28] wl[123] vdd gnd cell_6t
Xbit_r124_c28 bl[28] br[28] wl[124] vdd gnd cell_6t
Xbit_r125_c28 bl[28] br[28] wl[125] vdd gnd cell_6t
Xbit_r126_c28 bl[28] br[28] wl[126] vdd gnd cell_6t
Xbit_r127_c28 bl[28] br[28] wl[127] vdd gnd cell_6t
Xbit_r128_c28 bl[28] br[28] wl[128] vdd gnd cell_6t
Xbit_r129_c28 bl[28] br[28] wl[129] vdd gnd cell_6t
Xbit_r130_c28 bl[28] br[28] wl[130] vdd gnd cell_6t
Xbit_r131_c28 bl[28] br[28] wl[131] vdd gnd cell_6t
Xbit_r132_c28 bl[28] br[28] wl[132] vdd gnd cell_6t
Xbit_r133_c28 bl[28] br[28] wl[133] vdd gnd cell_6t
Xbit_r134_c28 bl[28] br[28] wl[134] vdd gnd cell_6t
Xbit_r135_c28 bl[28] br[28] wl[135] vdd gnd cell_6t
Xbit_r136_c28 bl[28] br[28] wl[136] vdd gnd cell_6t
Xbit_r137_c28 bl[28] br[28] wl[137] vdd gnd cell_6t
Xbit_r138_c28 bl[28] br[28] wl[138] vdd gnd cell_6t
Xbit_r139_c28 bl[28] br[28] wl[139] vdd gnd cell_6t
Xbit_r140_c28 bl[28] br[28] wl[140] vdd gnd cell_6t
Xbit_r141_c28 bl[28] br[28] wl[141] vdd gnd cell_6t
Xbit_r142_c28 bl[28] br[28] wl[142] vdd gnd cell_6t
Xbit_r143_c28 bl[28] br[28] wl[143] vdd gnd cell_6t
Xbit_r144_c28 bl[28] br[28] wl[144] vdd gnd cell_6t
Xbit_r145_c28 bl[28] br[28] wl[145] vdd gnd cell_6t
Xbit_r146_c28 bl[28] br[28] wl[146] vdd gnd cell_6t
Xbit_r147_c28 bl[28] br[28] wl[147] vdd gnd cell_6t
Xbit_r148_c28 bl[28] br[28] wl[148] vdd gnd cell_6t
Xbit_r149_c28 bl[28] br[28] wl[149] vdd gnd cell_6t
Xbit_r150_c28 bl[28] br[28] wl[150] vdd gnd cell_6t
Xbit_r151_c28 bl[28] br[28] wl[151] vdd gnd cell_6t
Xbit_r152_c28 bl[28] br[28] wl[152] vdd gnd cell_6t
Xbit_r153_c28 bl[28] br[28] wl[153] vdd gnd cell_6t
Xbit_r154_c28 bl[28] br[28] wl[154] vdd gnd cell_6t
Xbit_r155_c28 bl[28] br[28] wl[155] vdd gnd cell_6t
Xbit_r156_c28 bl[28] br[28] wl[156] vdd gnd cell_6t
Xbit_r157_c28 bl[28] br[28] wl[157] vdd gnd cell_6t
Xbit_r158_c28 bl[28] br[28] wl[158] vdd gnd cell_6t
Xbit_r159_c28 bl[28] br[28] wl[159] vdd gnd cell_6t
Xbit_r160_c28 bl[28] br[28] wl[160] vdd gnd cell_6t
Xbit_r161_c28 bl[28] br[28] wl[161] vdd gnd cell_6t
Xbit_r162_c28 bl[28] br[28] wl[162] vdd gnd cell_6t
Xbit_r163_c28 bl[28] br[28] wl[163] vdd gnd cell_6t
Xbit_r164_c28 bl[28] br[28] wl[164] vdd gnd cell_6t
Xbit_r165_c28 bl[28] br[28] wl[165] vdd gnd cell_6t
Xbit_r166_c28 bl[28] br[28] wl[166] vdd gnd cell_6t
Xbit_r167_c28 bl[28] br[28] wl[167] vdd gnd cell_6t
Xbit_r168_c28 bl[28] br[28] wl[168] vdd gnd cell_6t
Xbit_r169_c28 bl[28] br[28] wl[169] vdd gnd cell_6t
Xbit_r170_c28 bl[28] br[28] wl[170] vdd gnd cell_6t
Xbit_r171_c28 bl[28] br[28] wl[171] vdd gnd cell_6t
Xbit_r172_c28 bl[28] br[28] wl[172] vdd gnd cell_6t
Xbit_r173_c28 bl[28] br[28] wl[173] vdd gnd cell_6t
Xbit_r174_c28 bl[28] br[28] wl[174] vdd gnd cell_6t
Xbit_r175_c28 bl[28] br[28] wl[175] vdd gnd cell_6t
Xbit_r176_c28 bl[28] br[28] wl[176] vdd gnd cell_6t
Xbit_r177_c28 bl[28] br[28] wl[177] vdd gnd cell_6t
Xbit_r178_c28 bl[28] br[28] wl[178] vdd gnd cell_6t
Xbit_r179_c28 bl[28] br[28] wl[179] vdd gnd cell_6t
Xbit_r180_c28 bl[28] br[28] wl[180] vdd gnd cell_6t
Xbit_r181_c28 bl[28] br[28] wl[181] vdd gnd cell_6t
Xbit_r182_c28 bl[28] br[28] wl[182] vdd gnd cell_6t
Xbit_r183_c28 bl[28] br[28] wl[183] vdd gnd cell_6t
Xbit_r184_c28 bl[28] br[28] wl[184] vdd gnd cell_6t
Xbit_r185_c28 bl[28] br[28] wl[185] vdd gnd cell_6t
Xbit_r186_c28 bl[28] br[28] wl[186] vdd gnd cell_6t
Xbit_r187_c28 bl[28] br[28] wl[187] vdd gnd cell_6t
Xbit_r188_c28 bl[28] br[28] wl[188] vdd gnd cell_6t
Xbit_r189_c28 bl[28] br[28] wl[189] vdd gnd cell_6t
Xbit_r190_c28 bl[28] br[28] wl[190] vdd gnd cell_6t
Xbit_r191_c28 bl[28] br[28] wl[191] vdd gnd cell_6t
Xbit_r192_c28 bl[28] br[28] wl[192] vdd gnd cell_6t
Xbit_r193_c28 bl[28] br[28] wl[193] vdd gnd cell_6t
Xbit_r194_c28 bl[28] br[28] wl[194] vdd gnd cell_6t
Xbit_r195_c28 bl[28] br[28] wl[195] vdd gnd cell_6t
Xbit_r196_c28 bl[28] br[28] wl[196] vdd gnd cell_6t
Xbit_r197_c28 bl[28] br[28] wl[197] vdd gnd cell_6t
Xbit_r198_c28 bl[28] br[28] wl[198] vdd gnd cell_6t
Xbit_r199_c28 bl[28] br[28] wl[199] vdd gnd cell_6t
Xbit_r200_c28 bl[28] br[28] wl[200] vdd gnd cell_6t
Xbit_r201_c28 bl[28] br[28] wl[201] vdd gnd cell_6t
Xbit_r202_c28 bl[28] br[28] wl[202] vdd gnd cell_6t
Xbit_r203_c28 bl[28] br[28] wl[203] vdd gnd cell_6t
Xbit_r204_c28 bl[28] br[28] wl[204] vdd gnd cell_6t
Xbit_r205_c28 bl[28] br[28] wl[205] vdd gnd cell_6t
Xbit_r206_c28 bl[28] br[28] wl[206] vdd gnd cell_6t
Xbit_r207_c28 bl[28] br[28] wl[207] vdd gnd cell_6t
Xbit_r208_c28 bl[28] br[28] wl[208] vdd gnd cell_6t
Xbit_r209_c28 bl[28] br[28] wl[209] vdd gnd cell_6t
Xbit_r210_c28 bl[28] br[28] wl[210] vdd gnd cell_6t
Xbit_r211_c28 bl[28] br[28] wl[211] vdd gnd cell_6t
Xbit_r212_c28 bl[28] br[28] wl[212] vdd gnd cell_6t
Xbit_r213_c28 bl[28] br[28] wl[213] vdd gnd cell_6t
Xbit_r214_c28 bl[28] br[28] wl[214] vdd gnd cell_6t
Xbit_r215_c28 bl[28] br[28] wl[215] vdd gnd cell_6t
Xbit_r216_c28 bl[28] br[28] wl[216] vdd gnd cell_6t
Xbit_r217_c28 bl[28] br[28] wl[217] vdd gnd cell_6t
Xbit_r218_c28 bl[28] br[28] wl[218] vdd gnd cell_6t
Xbit_r219_c28 bl[28] br[28] wl[219] vdd gnd cell_6t
Xbit_r220_c28 bl[28] br[28] wl[220] vdd gnd cell_6t
Xbit_r221_c28 bl[28] br[28] wl[221] vdd gnd cell_6t
Xbit_r222_c28 bl[28] br[28] wl[222] vdd gnd cell_6t
Xbit_r223_c28 bl[28] br[28] wl[223] vdd gnd cell_6t
Xbit_r224_c28 bl[28] br[28] wl[224] vdd gnd cell_6t
Xbit_r225_c28 bl[28] br[28] wl[225] vdd gnd cell_6t
Xbit_r226_c28 bl[28] br[28] wl[226] vdd gnd cell_6t
Xbit_r227_c28 bl[28] br[28] wl[227] vdd gnd cell_6t
Xbit_r228_c28 bl[28] br[28] wl[228] vdd gnd cell_6t
Xbit_r229_c28 bl[28] br[28] wl[229] vdd gnd cell_6t
Xbit_r230_c28 bl[28] br[28] wl[230] vdd gnd cell_6t
Xbit_r231_c28 bl[28] br[28] wl[231] vdd gnd cell_6t
Xbit_r232_c28 bl[28] br[28] wl[232] vdd gnd cell_6t
Xbit_r233_c28 bl[28] br[28] wl[233] vdd gnd cell_6t
Xbit_r234_c28 bl[28] br[28] wl[234] vdd gnd cell_6t
Xbit_r235_c28 bl[28] br[28] wl[235] vdd gnd cell_6t
Xbit_r236_c28 bl[28] br[28] wl[236] vdd gnd cell_6t
Xbit_r237_c28 bl[28] br[28] wl[237] vdd gnd cell_6t
Xbit_r238_c28 bl[28] br[28] wl[238] vdd gnd cell_6t
Xbit_r239_c28 bl[28] br[28] wl[239] vdd gnd cell_6t
Xbit_r240_c28 bl[28] br[28] wl[240] vdd gnd cell_6t
Xbit_r241_c28 bl[28] br[28] wl[241] vdd gnd cell_6t
Xbit_r242_c28 bl[28] br[28] wl[242] vdd gnd cell_6t
Xbit_r243_c28 bl[28] br[28] wl[243] vdd gnd cell_6t
Xbit_r244_c28 bl[28] br[28] wl[244] vdd gnd cell_6t
Xbit_r245_c28 bl[28] br[28] wl[245] vdd gnd cell_6t
Xbit_r246_c28 bl[28] br[28] wl[246] vdd gnd cell_6t
Xbit_r247_c28 bl[28] br[28] wl[247] vdd gnd cell_6t
Xbit_r248_c28 bl[28] br[28] wl[248] vdd gnd cell_6t
Xbit_r249_c28 bl[28] br[28] wl[249] vdd gnd cell_6t
Xbit_r250_c28 bl[28] br[28] wl[250] vdd gnd cell_6t
Xbit_r251_c28 bl[28] br[28] wl[251] vdd gnd cell_6t
Xbit_r252_c28 bl[28] br[28] wl[252] vdd gnd cell_6t
Xbit_r253_c28 bl[28] br[28] wl[253] vdd gnd cell_6t
Xbit_r254_c28 bl[28] br[28] wl[254] vdd gnd cell_6t
Xbit_r255_c28 bl[28] br[28] wl[255] vdd gnd cell_6t
Xbit_r0_c29 bl[29] br[29] wl[0] vdd gnd cell_6t
Xbit_r1_c29 bl[29] br[29] wl[1] vdd gnd cell_6t
Xbit_r2_c29 bl[29] br[29] wl[2] vdd gnd cell_6t
Xbit_r3_c29 bl[29] br[29] wl[3] vdd gnd cell_6t
Xbit_r4_c29 bl[29] br[29] wl[4] vdd gnd cell_6t
Xbit_r5_c29 bl[29] br[29] wl[5] vdd gnd cell_6t
Xbit_r6_c29 bl[29] br[29] wl[6] vdd gnd cell_6t
Xbit_r7_c29 bl[29] br[29] wl[7] vdd gnd cell_6t
Xbit_r8_c29 bl[29] br[29] wl[8] vdd gnd cell_6t
Xbit_r9_c29 bl[29] br[29] wl[9] vdd gnd cell_6t
Xbit_r10_c29 bl[29] br[29] wl[10] vdd gnd cell_6t
Xbit_r11_c29 bl[29] br[29] wl[11] vdd gnd cell_6t
Xbit_r12_c29 bl[29] br[29] wl[12] vdd gnd cell_6t
Xbit_r13_c29 bl[29] br[29] wl[13] vdd gnd cell_6t
Xbit_r14_c29 bl[29] br[29] wl[14] vdd gnd cell_6t
Xbit_r15_c29 bl[29] br[29] wl[15] vdd gnd cell_6t
Xbit_r16_c29 bl[29] br[29] wl[16] vdd gnd cell_6t
Xbit_r17_c29 bl[29] br[29] wl[17] vdd gnd cell_6t
Xbit_r18_c29 bl[29] br[29] wl[18] vdd gnd cell_6t
Xbit_r19_c29 bl[29] br[29] wl[19] vdd gnd cell_6t
Xbit_r20_c29 bl[29] br[29] wl[20] vdd gnd cell_6t
Xbit_r21_c29 bl[29] br[29] wl[21] vdd gnd cell_6t
Xbit_r22_c29 bl[29] br[29] wl[22] vdd gnd cell_6t
Xbit_r23_c29 bl[29] br[29] wl[23] vdd gnd cell_6t
Xbit_r24_c29 bl[29] br[29] wl[24] vdd gnd cell_6t
Xbit_r25_c29 bl[29] br[29] wl[25] vdd gnd cell_6t
Xbit_r26_c29 bl[29] br[29] wl[26] vdd gnd cell_6t
Xbit_r27_c29 bl[29] br[29] wl[27] vdd gnd cell_6t
Xbit_r28_c29 bl[29] br[29] wl[28] vdd gnd cell_6t
Xbit_r29_c29 bl[29] br[29] wl[29] vdd gnd cell_6t
Xbit_r30_c29 bl[29] br[29] wl[30] vdd gnd cell_6t
Xbit_r31_c29 bl[29] br[29] wl[31] vdd gnd cell_6t
Xbit_r32_c29 bl[29] br[29] wl[32] vdd gnd cell_6t
Xbit_r33_c29 bl[29] br[29] wl[33] vdd gnd cell_6t
Xbit_r34_c29 bl[29] br[29] wl[34] vdd gnd cell_6t
Xbit_r35_c29 bl[29] br[29] wl[35] vdd gnd cell_6t
Xbit_r36_c29 bl[29] br[29] wl[36] vdd gnd cell_6t
Xbit_r37_c29 bl[29] br[29] wl[37] vdd gnd cell_6t
Xbit_r38_c29 bl[29] br[29] wl[38] vdd gnd cell_6t
Xbit_r39_c29 bl[29] br[29] wl[39] vdd gnd cell_6t
Xbit_r40_c29 bl[29] br[29] wl[40] vdd gnd cell_6t
Xbit_r41_c29 bl[29] br[29] wl[41] vdd gnd cell_6t
Xbit_r42_c29 bl[29] br[29] wl[42] vdd gnd cell_6t
Xbit_r43_c29 bl[29] br[29] wl[43] vdd gnd cell_6t
Xbit_r44_c29 bl[29] br[29] wl[44] vdd gnd cell_6t
Xbit_r45_c29 bl[29] br[29] wl[45] vdd gnd cell_6t
Xbit_r46_c29 bl[29] br[29] wl[46] vdd gnd cell_6t
Xbit_r47_c29 bl[29] br[29] wl[47] vdd gnd cell_6t
Xbit_r48_c29 bl[29] br[29] wl[48] vdd gnd cell_6t
Xbit_r49_c29 bl[29] br[29] wl[49] vdd gnd cell_6t
Xbit_r50_c29 bl[29] br[29] wl[50] vdd gnd cell_6t
Xbit_r51_c29 bl[29] br[29] wl[51] vdd gnd cell_6t
Xbit_r52_c29 bl[29] br[29] wl[52] vdd gnd cell_6t
Xbit_r53_c29 bl[29] br[29] wl[53] vdd gnd cell_6t
Xbit_r54_c29 bl[29] br[29] wl[54] vdd gnd cell_6t
Xbit_r55_c29 bl[29] br[29] wl[55] vdd gnd cell_6t
Xbit_r56_c29 bl[29] br[29] wl[56] vdd gnd cell_6t
Xbit_r57_c29 bl[29] br[29] wl[57] vdd gnd cell_6t
Xbit_r58_c29 bl[29] br[29] wl[58] vdd gnd cell_6t
Xbit_r59_c29 bl[29] br[29] wl[59] vdd gnd cell_6t
Xbit_r60_c29 bl[29] br[29] wl[60] vdd gnd cell_6t
Xbit_r61_c29 bl[29] br[29] wl[61] vdd gnd cell_6t
Xbit_r62_c29 bl[29] br[29] wl[62] vdd gnd cell_6t
Xbit_r63_c29 bl[29] br[29] wl[63] vdd gnd cell_6t
Xbit_r64_c29 bl[29] br[29] wl[64] vdd gnd cell_6t
Xbit_r65_c29 bl[29] br[29] wl[65] vdd gnd cell_6t
Xbit_r66_c29 bl[29] br[29] wl[66] vdd gnd cell_6t
Xbit_r67_c29 bl[29] br[29] wl[67] vdd gnd cell_6t
Xbit_r68_c29 bl[29] br[29] wl[68] vdd gnd cell_6t
Xbit_r69_c29 bl[29] br[29] wl[69] vdd gnd cell_6t
Xbit_r70_c29 bl[29] br[29] wl[70] vdd gnd cell_6t
Xbit_r71_c29 bl[29] br[29] wl[71] vdd gnd cell_6t
Xbit_r72_c29 bl[29] br[29] wl[72] vdd gnd cell_6t
Xbit_r73_c29 bl[29] br[29] wl[73] vdd gnd cell_6t
Xbit_r74_c29 bl[29] br[29] wl[74] vdd gnd cell_6t
Xbit_r75_c29 bl[29] br[29] wl[75] vdd gnd cell_6t
Xbit_r76_c29 bl[29] br[29] wl[76] vdd gnd cell_6t
Xbit_r77_c29 bl[29] br[29] wl[77] vdd gnd cell_6t
Xbit_r78_c29 bl[29] br[29] wl[78] vdd gnd cell_6t
Xbit_r79_c29 bl[29] br[29] wl[79] vdd gnd cell_6t
Xbit_r80_c29 bl[29] br[29] wl[80] vdd gnd cell_6t
Xbit_r81_c29 bl[29] br[29] wl[81] vdd gnd cell_6t
Xbit_r82_c29 bl[29] br[29] wl[82] vdd gnd cell_6t
Xbit_r83_c29 bl[29] br[29] wl[83] vdd gnd cell_6t
Xbit_r84_c29 bl[29] br[29] wl[84] vdd gnd cell_6t
Xbit_r85_c29 bl[29] br[29] wl[85] vdd gnd cell_6t
Xbit_r86_c29 bl[29] br[29] wl[86] vdd gnd cell_6t
Xbit_r87_c29 bl[29] br[29] wl[87] vdd gnd cell_6t
Xbit_r88_c29 bl[29] br[29] wl[88] vdd gnd cell_6t
Xbit_r89_c29 bl[29] br[29] wl[89] vdd gnd cell_6t
Xbit_r90_c29 bl[29] br[29] wl[90] vdd gnd cell_6t
Xbit_r91_c29 bl[29] br[29] wl[91] vdd gnd cell_6t
Xbit_r92_c29 bl[29] br[29] wl[92] vdd gnd cell_6t
Xbit_r93_c29 bl[29] br[29] wl[93] vdd gnd cell_6t
Xbit_r94_c29 bl[29] br[29] wl[94] vdd gnd cell_6t
Xbit_r95_c29 bl[29] br[29] wl[95] vdd gnd cell_6t
Xbit_r96_c29 bl[29] br[29] wl[96] vdd gnd cell_6t
Xbit_r97_c29 bl[29] br[29] wl[97] vdd gnd cell_6t
Xbit_r98_c29 bl[29] br[29] wl[98] vdd gnd cell_6t
Xbit_r99_c29 bl[29] br[29] wl[99] vdd gnd cell_6t
Xbit_r100_c29 bl[29] br[29] wl[100] vdd gnd cell_6t
Xbit_r101_c29 bl[29] br[29] wl[101] vdd gnd cell_6t
Xbit_r102_c29 bl[29] br[29] wl[102] vdd gnd cell_6t
Xbit_r103_c29 bl[29] br[29] wl[103] vdd gnd cell_6t
Xbit_r104_c29 bl[29] br[29] wl[104] vdd gnd cell_6t
Xbit_r105_c29 bl[29] br[29] wl[105] vdd gnd cell_6t
Xbit_r106_c29 bl[29] br[29] wl[106] vdd gnd cell_6t
Xbit_r107_c29 bl[29] br[29] wl[107] vdd gnd cell_6t
Xbit_r108_c29 bl[29] br[29] wl[108] vdd gnd cell_6t
Xbit_r109_c29 bl[29] br[29] wl[109] vdd gnd cell_6t
Xbit_r110_c29 bl[29] br[29] wl[110] vdd gnd cell_6t
Xbit_r111_c29 bl[29] br[29] wl[111] vdd gnd cell_6t
Xbit_r112_c29 bl[29] br[29] wl[112] vdd gnd cell_6t
Xbit_r113_c29 bl[29] br[29] wl[113] vdd gnd cell_6t
Xbit_r114_c29 bl[29] br[29] wl[114] vdd gnd cell_6t
Xbit_r115_c29 bl[29] br[29] wl[115] vdd gnd cell_6t
Xbit_r116_c29 bl[29] br[29] wl[116] vdd gnd cell_6t
Xbit_r117_c29 bl[29] br[29] wl[117] vdd gnd cell_6t
Xbit_r118_c29 bl[29] br[29] wl[118] vdd gnd cell_6t
Xbit_r119_c29 bl[29] br[29] wl[119] vdd gnd cell_6t
Xbit_r120_c29 bl[29] br[29] wl[120] vdd gnd cell_6t
Xbit_r121_c29 bl[29] br[29] wl[121] vdd gnd cell_6t
Xbit_r122_c29 bl[29] br[29] wl[122] vdd gnd cell_6t
Xbit_r123_c29 bl[29] br[29] wl[123] vdd gnd cell_6t
Xbit_r124_c29 bl[29] br[29] wl[124] vdd gnd cell_6t
Xbit_r125_c29 bl[29] br[29] wl[125] vdd gnd cell_6t
Xbit_r126_c29 bl[29] br[29] wl[126] vdd gnd cell_6t
Xbit_r127_c29 bl[29] br[29] wl[127] vdd gnd cell_6t
Xbit_r128_c29 bl[29] br[29] wl[128] vdd gnd cell_6t
Xbit_r129_c29 bl[29] br[29] wl[129] vdd gnd cell_6t
Xbit_r130_c29 bl[29] br[29] wl[130] vdd gnd cell_6t
Xbit_r131_c29 bl[29] br[29] wl[131] vdd gnd cell_6t
Xbit_r132_c29 bl[29] br[29] wl[132] vdd gnd cell_6t
Xbit_r133_c29 bl[29] br[29] wl[133] vdd gnd cell_6t
Xbit_r134_c29 bl[29] br[29] wl[134] vdd gnd cell_6t
Xbit_r135_c29 bl[29] br[29] wl[135] vdd gnd cell_6t
Xbit_r136_c29 bl[29] br[29] wl[136] vdd gnd cell_6t
Xbit_r137_c29 bl[29] br[29] wl[137] vdd gnd cell_6t
Xbit_r138_c29 bl[29] br[29] wl[138] vdd gnd cell_6t
Xbit_r139_c29 bl[29] br[29] wl[139] vdd gnd cell_6t
Xbit_r140_c29 bl[29] br[29] wl[140] vdd gnd cell_6t
Xbit_r141_c29 bl[29] br[29] wl[141] vdd gnd cell_6t
Xbit_r142_c29 bl[29] br[29] wl[142] vdd gnd cell_6t
Xbit_r143_c29 bl[29] br[29] wl[143] vdd gnd cell_6t
Xbit_r144_c29 bl[29] br[29] wl[144] vdd gnd cell_6t
Xbit_r145_c29 bl[29] br[29] wl[145] vdd gnd cell_6t
Xbit_r146_c29 bl[29] br[29] wl[146] vdd gnd cell_6t
Xbit_r147_c29 bl[29] br[29] wl[147] vdd gnd cell_6t
Xbit_r148_c29 bl[29] br[29] wl[148] vdd gnd cell_6t
Xbit_r149_c29 bl[29] br[29] wl[149] vdd gnd cell_6t
Xbit_r150_c29 bl[29] br[29] wl[150] vdd gnd cell_6t
Xbit_r151_c29 bl[29] br[29] wl[151] vdd gnd cell_6t
Xbit_r152_c29 bl[29] br[29] wl[152] vdd gnd cell_6t
Xbit_r153_c29 bl[29] br[29] wl[153] vdd gnd cell_6t
Xbit_r154_c29 bl[29] br[29] wl[154] vdd gnd cell_6t
Xbit_r155_c29 bl[29] br[29] wl[155] vdd gnd cell_6t
Xbit_r156_c29 bl[29] br[29] wl[156] vdd gnd cell_6t
Xbit_r157_c29 bl[29] br[29] wl[157] vdd gnd cell_6t
Xbit_r158_c29 bl[29] br[29] wl[158] vdd gnd cell_6t
Xbit_r159_c29 bl[29] br[29] wl[159] vdd gnd cell_6t
Xbit_r160_c29 bl[29] br[29] wl[160] vdd gnd cell_6t
Xbit_r161_c29 bl[29] br[29] wl[161] vdd gnd cell_6t
Xbit_r162_c29 bl[29] br[29] wl[162] vdd gnd cell_6t
Xbit_r163_c29 bl[29] br[29] wl[163] vdd gnd cell_6t
Xbit_r164_c29 bl[29] br[29] wl[164] vdd gnd cell_6t
Xbit_r165_c29 bl[29] br[29] wl[165] vdd gnd cell_6t
Xbit_r166_c29 bl[29] br[29] wl[166] vdd gnd cell_6t
Xbit_r167_c29 bl[29] br[29] wl[167] vdd gnd cell_6t
Xbit_r168_c29 bl[29] br[29] wl[168] vdd gnd cell_6t
Xbit_r169_c29 bl[29] br[29] wl[169] vdd gnd cell_6t
Xbit_r170_c29 bl[29] br[29] wl[170] vdd gnd cell_6t
Xbit_r171_c29 bl[29] br[29] wl[171] vdd gnd cell_6t
Xbit_r172_c29 bl[29] br[29] wl[172] vdd gnd cell_6t
Xbit_r173_c29 bl[29] br[29] wl[173] vdd gnd cell_6t
Xbit_r174_c29 bl[29] br[29] wl[174] vdd gnd cell_6t
Xbit_r175_c29 bl[29] br[29] wl[175] vdd gnd cell_6t
Xbit_r176_c29 bl[29] br[29] wl[176] vdd gnd cell_6t
Xbit_r177_c29 bl[29] br[29] wl[177] vdd gnd cell_6t
Xbit_r178_c29 bl[29] br[29] wl[178] vdd gnd cell_6t
Xbit_r179_c29 bl[29] br[29] wl[179] vdd gnd cell_6t
Xbit_r180_c29 bl[29] br[29] wl[180] vdd gnd cell_6t
Xbit_r181_c29 bl[29] br[29] wl[181] vdd gnd cell_6t
Xbit_r182_c29 bl[29] br[29] wl[182] vdd gnd cell_6t
Xbit_r183_c29 bl[29] br[29] wl[183] vdd gnd cell_6t
Xbit_r184_c29 bl[29] br[29] wl[184] vdd gnd cell_6t
Xbit_r185_c29 bl[29] br[29] wl[185] vdd gnd cell_6t
Xbit_r186_c29 bl[29] br[29] wl[186] vdd gnd cell_6t
Xbit_r187_c29 bl[29] br[29] wl[187] vdd gnd cell_6t
Xbit_r188_c29 bl[29] br[29] wl[188] vdd gnd cell_6t
Xbit_r189_c29 bl[29] br[29] wl[189] vdd gnd cell_6t
Xbit_r190_c29 bl[29] br[29] wl[190] vdd gnd cell_6t
Xbit_r191_c29 bl[29] br[29] wl[191] vdd gnd cell_6t
Xbit_r192_c29 bl[29] br[29] wl[192] vdd gnd cell_6t
Xbit_r193_c29 bl[29] br[29] wl[193] vdd gnd cell_6t
Xbit_r194_c29 bl[29] br[29] wl[194] vdd gnd cell_6t
Xbit_r195_c29 bl[29] br[29] wl[195] vdd gnd cell_6t
Xbit_r196_c29 bl[29] br[29] wl[196] vdd gnd cell_6t
Xbit_r197_c29 bl[29] br[29] wl[197] vdd gnd cell_6t
Xbit_r198_c29 bl[29] br[29] wl[198] vdd gnd cell_6t
Xbit_r199_c29 bl[29] br[29] wl[199] vdd gnd cell_6t
Xbit_r200_c29 bl[29] br[29] wl[200] vdd gnd cell_6t
Xbit_r201_c29 bl[29] br[29] wl[201] vdd gnd cell_6t
Xbit_r202_c29 bl[29] br[29] wl[202] vdd gnd cell_6t
Xbit_r203_c29 bl[29] br[29] wl[203] vdd gnd cell_6t
Xbit_r204_c29 bl[29] br[29] wl[204] vdd gnd cell_6t
Xbit_r205_c29 bl[29] br[29] wl[205] vdd gnd cell_6t
Xbit_r206_c29 bl[29] br[29] wl[206] vdd gnd cell_6t
Xbit_r207_c29 bl[29] br[29] wl[207] vdd gnd cell_6t
Xbit_r208_c29 bl[29] br[29] wl[208] vdd gnd cell_6t
Xbit_r209_c29 bl[29] br[29] wl[209] vdd gnd cell_6t
Xbit_r210_c29 bl[29] br[29] wl[210] vdd gnd cell_6t
Xbit_r211_c29 bl[29] br[29] wl[211] vdd gnd cell_6t
Xbit_r212_c29 bl[29] br[29] wl[212] vdd gnd cell_6t
Xbit_r213_c29 bl[29] br[29] wl[213] vdd gnd cell_6t
Xbit_r214_c29 bl[29] br[29] wl[214] vdd gnd cell_6t
Xbit_r215_c29 bl[29] br[29] wl[215] vdd gnd cell_6t
Xbit_r216_c29 bl[29] br[29] wl[216] vdd gnd cell_6t
Xbit_r217_c29 bl[29] br[29] wl[217] vdd gnd cell_6t
Xbit_r218_c29 bl[29] br[29] wl[218] vdd gnd cell_6t
Xbit_r219_c29 bl[29] br[29] wl[219] vdd gnd cell_6t
Xbit_r220_c29 bl[29] br[29] wl[220] vdd gnd cell_6t
Xbit_r221_c29 bl[29] br[29] wl[221] vdd gnd cell_6t
Xbit_r222_c29 bl[29] br[29] wl[222] vdd gnd cell_6t
Xbit_r223_c29 bl[29] br[29] wl[223] vdd gnd cell_6t
Xbit_r224_c29 bl[29] br[29] wl[224] vdd gnd cell_6t
Xbit_r225_c29 bl[29] br[29] wl[225] vdd gnd cell_6t
Xbit_r226_c29 bl[29] br[29] wl[226] vdd gnd cell_6t
Xbit_r227_c29 bl[29] br[29] wl[227] vdd gnd cell_6t
Xbit_r228_c29 bl[29] br[29] wl[228] vdd gnd cell_6t
Xbit_r229_c29 bl[29] br[29] wl[229] vdd gnd cell_6t
Xbit_r230_c29 bl[29] br[29] wl[230] vdd gnd cell_6t
Xbit_r231_c29 bl[29] br[29] wl[231] vdd gnd cell_6t
Xbit_r232_c29 bl[29] br[29] wl[232] vdd gnd cell_6t
Xbit_r233_c29 bl[29] br[29] wl[233] vdd gnd cell_6t
Xbit_r234_c29 bl[29] br[29] wl[234] vdd gnd cell_6t
Xbit_r235_c29 bl[29] br[29] wl[235] vdd gnd cell_6t
Xbit_r236_c29 bl[29] br[29] wl[236] vdd gnd cell_6t
Xbit_r237_c29 bl[29] br[29] wl[237] vdd gnd cell_6t
Xbit_r238_c29 bl[29] br[29] wl[238] vdd gnd cell_6t
Xbit_r239_c29 bl[29] br[29] wl[239] vdd gnd cell_6t
Xbit_r240_c29 bl[29] br[29] wl[240] vdd gnd cell_6t
Xbit_r241_c29 bl[29] br[29] wl[241] vdd gnd cell_6t
Xbit_r242_c29 bl[29] br[29] wl[242] vdd gnd cell_6t
Xbit_r243_c29 bl[29] br[29] wl[243] vdd gnd cell_6t
Xbit_r244_c29 bl[29] br[29] wl[244] vdd gnd cell_6t
Xbit_r245_c29 bl[29] br[29] wl[245] vdd gnd cell_6t
Xbit_r246_c29 bl[29] br[29] wl[246] vdd gnd cell_6t
Xbit_r247_c29 bl[29] br[29] wl[247] vdd gnd cell_6t
Xbit_r248_c29 bl[29] br[29] wl[248] vdd gnd cell_6t
Xbit_r249_c29 bl[29] br[29] wl[249] vdd gnd cell_6t
Xbit_r250_c29 bl[29] br[29] wl[250] vdd gnd cell_6t
Xbit_r251_c29 bl[29] br[29] wl[251] vdd gnd cell_6t
Xbit_r252_c29 bl[29] br[29] wl[252] vdd gnd cell_6t
Xbit_r253_c29 bl[29] br[29] wl[253] vdd gnd cell_6t
Xbit_r254_c29 bl[29] br[29] wl[254] vdd gnd cell_6t
Xbit_r255_c29 bl[29] br[29] wl[255] vdd gnd cell_6t
Xbit_r0_c30 bl[30] br[30] wl[0] vdd gnd cell_6t
Xbit_r1_c30 bl[30] br[30] wl[1] vdd gnd cell_6t
Xbit_r2_c30 bl[30] br[30] wl[2] vdd gnd cell_6t
Xbit_r3_c30 bl[30] br[30] wl[3] vdd gnd cell_6t
Xbit_r4_c30 bl[30] br[30] wl[4] vdd gnd cell_6t
Xbit_r5_c30 bl[30] br[30] wl[5] vdd gnd cell_6t
Xbit_r6_c30 bl[30] br[30] wl[6] vdd gnd cell_6t
Xbit_r7_c30 bl[30] br[30] wl[7] vdd gnd cell_6t
Xbit_r8_c30 bl[30] br[30] wl[8] vdd gnd cell_6t
Xbit_r9_c30 bl[30] br[30] wl[9] vdd gnd cell_6t
Xbit_r10_c30 bl[30] br[30] wl[10] vdd gnd cell_6t
Xbit_r11_c30 bl[30] br[30] wl[11] vdd gnd cell_6t
Xbit_r12_c30 bl[30] br[30] wl[12] vdd gnd cell_6t
Xbit_r13_c30 bl[30] br[30] wl[13] vdd gnd cell_6t
Xbit_r14_c30 bl[30] br[30] wl[14] vdd gnd cell_6t
Xbit_r15_c30 bl[30] br[30] wl[15] vdd gnd cell_6t
Xbit_r16_c30 bl[30] br[30] wl[16] vdd gnd cell_6t
Xbit_r17_c30 bl[30] br[30] wl[17] vdd gnd cell_6t
Xbit_r18_c30 bl[30] br[30] wl[18] vdd gnd cell_6t
Xbit_r19_c30 bl[30] br[30] wl[19] vdd gnd cell_6t
Xbit_r20_c30 bl[30] br[30] wl[20] vdd gnd cell_6t
Xbit_r21_c30 bl[30] br[30] wl[21] vdd gnd cell_6t
Xbit_r22_c30 bl[30] br[30] wl[22] vdd gnd cell_6t
Xbit_r23_c30 bl[30] br[30] wl[23] vdd gnd cell_6t
Xbit_r24_c30 bl[30] br[30] wl[24] vdd gnd cell_6t
Xbit_r25_c30 bl[30] br[30] wl[25] vdd gnd cell_6t
Xbit_r26_c30 bl[30] br[30] wl[26] vdd gnd cell_6t
Xbit_r27_c30 bl[30] br[30] wl[27] vdd gnd cell_6t
Xbit_r28_c30 bl[30] br[30] wl[28] vdd gnd cell_6t
Xbit_r29_c30 bl[30] br[30] wl[29] vdd gnd cell_6t
Xbit_r30_c30 bl[30] br[30] wl[30] vdd gnd cell_6t
Xbit_r31_c30 bl[30] br[30] wl[31] vdd gnd cell_6t
Xbit_r32_c30 bl[30] br[30] wl[32] vdd gnd cell_6t
Xbit_r33_c30 bl[30] br[30] wl[33] vdd gnd cell_6t
Xbit_r34_c30 bl[30] br[30] wl[34] vdd gnd cell_6t
Xbit_r35_c30 bl[30] br[30] wl[35] vdd gnd cell_6t
Xbit_r36_c30 bl[30] br[30] wl[36] vdd gnd cell_6t
Xbit_r37_c30 bl[30] br[30] wl[37] vdd gnd cell_6t
Xbit_r38_c30 bl[30] br[30] wl[38] vdd gnd cell_6t
Xbit_r39_c30 bl[30] br[30] wl[39] vdd gnd cell_6t
Xbit_r40_c30 bl[30] br[30] wl[40] vdd gnd cell_6t
Xbit_r41_c30 bl[30] br[30] wl[41] vdd gnd cell_6t
Xbit_r42_c30 bl[30] br[30] wl[42] vdd gnd cell_6t
Xbit_r43_c30 bl[30] br[30] wl[43] vdd gnd cell_6t
Xbit_r44_c30 bl[30] br[30] wl[44] vdd gnd cell_6t
Xbit_r45_c30 bl[30] br[30] wl[45] vdd gnd cell_6t
Xbit_r46_c30 bl[30] br[30] wl[46] vdd gnd cell_6t
Xbit_r47_c30 bl[30] br[30] wl[47] vdd gnd cell_6t
Xbit_r48_c30 bl[30] br[30] wl[48] vdd gnd cell_6t
Xbit_r49_c30 bl[30] br[30] wl[49] vdd gnd cell_6t
Xbit_r50_c30 bl[30] br[30] wl[50] vdd gnd cell_6t
Xbit_r51_c30 bl[30] br[30] wl[51] vdd gnd cell_6t
Xbit_r52_c30 bl[30] br[30] wl[52] vdd gnd cell_6t
Xbit_r53_c30 bl[30] br[30] wl[53] vdd gnd cell_6t
Xbit_r54_c30 bl[30] br[30] wl[54] vdd gnd cell_6t
Xbit_r55_c30 bl[30] br[30] wl[55] vdd gnd cell_6t
Xbit_r56_c30 bl[30] br[30] wl[56] vdd gnd cell_6t
Xbit_r57_c30 bl[30] br[30] wl[57] vdd gnd cell_6t
Xbit_r58_c30 bl[30] br[30] wl[58] vdd gnd cell_6t
Xbit_r59_c30 bl[30] br[30] wl[59] vdd gnd cell_6t
Xbit_r60_c30 bl[30] br[30] wl[60] vdd gnd cell_6t
Xbit_r61_c30 bl[30] br[30] wl[61] vdd gnd cell_6t
Xbit_r62_c30 bl[30] br[30] wl[62] vdd gnd cell_6t
Xbit_r63_c30 bl[30] br[30] wl[63] vdd gnd cell_6t
Xbit_r64_c30 bl[30] br[30] wl[64] vdd gnd cell_6t
Xbit_r65_c30 bl[30] br[30] wl[65] vdd gnd cell_6t
Xbit_r66_c30 bl[30] br[30] wl[66] vdd gnd cell_6t
Xbit_r67_c30 bl[30] br[30] wl[67] vdd gnd cell_6t
Xbit_r68_c30 bl[30] br[30] wl[68] vdd gnd cell_6t
Xbit_r69_c30 bl[30] br[30] wl[69] vdd gnd cell_6t
Xbit_r70_c30 bl[30] br[30] wl[70] vdd gnd cell_6t
Xbit_r71_c30 bl[30] br[30] wl[71] vdd gnd cell_6t
Xbit_r72_c30 bl[30] br[30] wl[72] vdd gnd cell_6t
Xbit_r73_c30 bl[30] br[30] wl[73] vdd gnd cell_6t
Xbit_r74_c30 bl[30] br[30] wl[74] vdd gnd cell_6t
Xbit_r75_c30 bl[30] br[30] wl[75] vdd gnd cell_6t
Xbit_r76_c30 bl[30] br[30] wl[76] vdd gnd cell_6t
Xbit_r77_c30 bl[30] br[30] wl[77] vdd gnd cell_6t
Xbit_r78_c30 bl[30] br[30] wl[78] vdd gnd cell_6t
Xbit_r79_c30 bl[30] br[30] wl[79] vdd gnd cell_6t
Xbit_r80_c30 bl[30] br[30] wl[80] vdd gnd cell_6t
Xbit_r81_c30 bl[30] br[30] wl[81] vdd gnd cell_6t
Xbit_r82_c30 bl[30] br[30] wl[82] vdd gnd cell_6t
Xbit_r83_c30 bl[30] br[30] wl[83] vdd gnd cell_6t
Xbit_r84_c30 bl[30] br[30] wl[84] vdd gnd cell_6t
Xbit_r85_c30 bl[30] br[30] wl[85] vdd gnd cell_6t
Xbit_r86_c30 bl[30] br[30] wl[86] vdd gnd cell_6t
Xbit_r87_c30 bl[30] br[30] wl[87] vdd gnd cell_6t
Xbit_r88_c30 bl[30] br[30] wl[88] vdd gnd cell_6t
Xbit_r89_c30 bl[30] br[30] wl[89] vdd gnd cell_6t
Xbit_r90_c30 bl[30] br[30] wl[90] vdd gnd cell_6t
Xbit_r91_c30 bl[30] br[30] wl[91] vdd gnd cell_6t
Xbit_r92_c30 bl[30] br[30] wl[92] vdd gnd cell_6t
Xbit_r93_c30 bl[30] br[30] wl[93] vdd gnd cell_6t
Xbit_r94_c30 bl[30] br[30] wl[94] vdd gnd cell_6t
Xbit_r95_c30 bl[30] br[30] wl[95] vdd gnd cell_6t
Xbit_r96_c30 bl[30] br[30] wl[96] vdd gnd cell_6t
Xbit_r97_c30 bl[30] br[30] wl[97] vdd gnd cell_6t
Xbit_r98_c30 bl[30] br[30] wl[98] vdd gnd cell_6t
Xbit_r99_c30 bl[30] br[30] wl[99] vdd gnd cell_6t
Xbit_r100_c30 bl[30] br[30] wl[100] vdd gnd cell_6t
Xbit_r101_c30 bl[30] br[30] wl[101] vdd gnd cell_6t
Xbit_r102_c30 bl[30] br[30] wl[102] vdd gnd cell_6t
Xbit_r103_c30 bl[30] br[30] wl[103] vdd gnd cell_6t
Xbit_r104_c30 bl[30] br[30] wl[104] vdd gnd cell_6t
Xbit_r105_c30 bl[30] br[30] wl[105] vdd gnd cell_6t
Xbit_r106_c30 bl[30] br[30] wl[106] vdd gnd cell_6t
Xbit_r107_c30 bl[30] br[30] wl[107] vdd gnd cell_6t
Xbit_r108_c30 bl[30] br[30] wl[108] vdd gnd cell_6t
Xbit_r109_c30 bl[30] br[30] wl[109] vdd gnd cell_6t
Xbit_r110_c30 bl[30] br[30] wl[110] vdd gnd cell_6t
Xbit_r111_c30 bl[30] br[30] wl[111] vdd gnd cell_6t
Xbit_r112_c30 bl[30] br[30] wl[112] vdd gnd cell_6t
Xbit_r113_c30 bl[30] br[30] wl[113] vdd gnd cell_6t
Xbit_r114_c30 bl[30] br[30] wl[114] vdd gnd cell_6t
Xbit_r115_c30 bl[30] br[30] wl[115] vdd gnd cell_6t
Xbit_r116_c30 bl[30] br[30] wl[116] vdd gnd cell_6t
Xbit_r117_c30 bl[30] br[30] wl[117] vdd gnd cell_6t
Xbit_r118_c30 bl[30] br[30] wl[118] vdd gnd cell_6t
Xbit_r119_c30 bl[30] br[30] wl[119] vdd gnd cell_6t
Xbit_r120_c30 bl[30] br[30] wl[120] vdd gnd cell_6t
Xbit_r121_c30 bl[30] br[30] wl[121] vdd gnd cell_6t
Xbit_r122_c30 bl[30] br[30] wl[122] vdd gnd cell_6t
Xbit_r123_c30 bl[30] br[30] wl[123] vdd gnd cell_6t
Xbit_r124_c30 bl[30] br[30] wl[124] vdd gnd cell_6t
Xbit_r125_c30 bl[30] br[30] wl[125] vdd gnd cell_6t
Xbit_r126_c30 bl[30] br[30] wl[126] vdd gnd cell_6t
Xbit_r127_c30 bl[30] br[30] wl[127] vdd gnd cell_6t
Xbit_r128_c30 bl[30] br[30] wl[128] vdd gnd cell_6t
Xbit_r129_c30 bl[30] br[30] wl[129] vdd gnd cell_6t
Xbit_r130_c30 bl[30] br[30] wl[130] vdd gnd cell_6t
Xbit_r131_c30 bl[30] br[30] wl[131] vdd gnd cell_6t
Xbit_r132_c30 bl[30] br[30] wl[132] vdd gnd cell_6t
Xbit_r133_c30 bl[30] br[30] wl[133] vdd gnd cell_6t
Xbit_r134_c30 bl[30] br[30] wl[134] vdd gnd cell_6t
Xbit_r135_c30 bl[30] br[30] wl[135] vdd gnd cell_6t
Xbit_r136_c30 bl[30] br[30] wl[136] vdd gnd cell_6t
Xbit_r137_c30 bl[30] br[30] wl[137] vdd gnd cell_6t
Xbit_r138_c30 bl[30] br[30] wl[138] vdd gnd cell_6t
Xbit_r139_c30 bl[30] br[30] wl[139] vdd gnd cell_6t
Xbit_r140_c30 bl[30] br[30] wl[140] vdd gnd cell_6t
Xbit_r141_c30 bl[30] br[30] wl[141] vdd gnd cell_6t
Xbit_r142_c30 bl[30] br[30] wl[142] vdd gnd cell_6t
Xbit_r143_c30 bl[30] br[30] wl[143] vdd gnd cell_6t
Xbit_r144_c30 bl[30] br[30] wl[144] vdd gnd cell_6t
Xbit_r145_c30 bl[30] br[30] wl[145] vdd gnd cell_6t
Xbit_r146_c30 bl[30] br[30] wl[146] vdd gnd cell_6t
Xbit_r147_c30 bl[30] br[30] wl[147] vdd gnd cell_6t
Xbit_r148_c30 bl[30] br[30] wl[148] vdd gnd cell_6t
Xbit_r149_c30 bl[30] br[30] wl[149] vdd gnd cell_6t
Xbit_r150_c30 bl[30] br[30] wl[150] vdd gnd cell_6t
Xbit_r151_c30 bl[30] br[30] wl[151] vdd gnd cell_6t
Xbit_r152_c30 bl[30] br[30] wl[152] vdd gnd cell_6t
Xbit_r153_c30 bl[30] br[30] wl[153] vdd gnd cell_6t
Xbit_r154_c30 bl[30] br[30] wl[154] vdd gnd cell_6t
Xbit_r155_c30 bl[30] br[30] wl[155] vdd gnd cell_6t
Xbit_r156_c30 bl[30] br[30] wl[156] vdd gnd cell_6t
Xbit_r157_c30 bl[30] br[30] wl[157] vdd gnd cell_6t
Xbit_r158_c30 bl[30] br[30] wl[158] vdd gnd cell_6t
Xbit_r159_c30 bl[30] br[30] wl[159] vdd gnd cell_6t
Xbit_r160_c30 bl[30] br[30] wl[160] vdd gnd cell_6t
Xbit_r161_c30 bl[30] br[30] wl[161] vdd gnd cell_6t
Xbit_r162_c30 bl[30] br[30] wl[162] vdd gnd cell_6t
Xbit_r163_c30 bl[30] br[30] wl[163] vdd gnd cell_6t
Xbit_r164_c30 bl[30] br[30] wl[164] vdd gnd cell_6t
Xbit_r165_c30 bl[30] br[30] wl[165] vdd gnd cell_6t
Xbit_r166_c30 bl[30] br[30] wl[166] vdd gnd cell_6t
Xbit_r167_c30 bl[30] br[30] wl[167] vdd gnd cell_6t
Xbit_r168_c30 bl[30] br[30] wl[168] vdd gnd cell_6t
Xbit_r169_c30 bl[30] br[30] wl[169] vdd gnd cell_6t
Xbit_r170_c30 bl[30] br[30] wl[170] vdd gnd cell_6t
Xbit_r171_c30 bl[30] br[30] wl[171] vdd gnd cell_6t
Xbit_r172_c30 bl[30] br[30] wl[172] vdd gnd cell_6t
Xbit_r173_c30 bl[30] br[30] wl[173] vdd gnd cell_6t
Xbit_r174_c30 bl[30] br[30] wl[174] vdd gnd cell_6t
Xbit_r175_c30 bl[30] br[30] wl[175] vdd gnd cell_6t
Xbit_r176_c30 bl[30] br[30] wl[176] vdd gnd cell_6t
Xbit_r177_c30 bl[30] br[30] wl[177] vdd gnd cell_6t
Xbit_r178_c30 bl[30] br[30] wl[178] vdd gnd cell_6t
Xbit_r179_c30 bl[30] br[30] wl[179] vdd gnd cell_6t
Xbit_r180_c30 bl[30] br[30] wl[180] vdd gnd cell_6t
Xbit_r181_c30 bl[30] br[30] wl[181] vdd gnd cell_6t
Xbit_r182_c30 bl[30] br[30] wl[182] vdd gnd cell_6t
Xbit_r183_c30 bl[30] br[30] wl[183] vdd gnd cell_6t
Xbit_r184_c30 bl[30] br[30] wl[184] vdd gnd cell_6t
Xbit_r185_c30 bl[30] br[30] wl[185] vdd gnd cell_6t
Xbit_r186_c30 bl[30] br[30] wl[186] vdd gnd cell_6t
Xbit_r187_c30 bl[30] br[30] wl[187] vdd gnd cell_6t
Xbit_r188_c30 bl[30] br[30] wl[188] vdd gnd cell_6t
Xbit_r189_c30 bl[30] br[30] wl[189] vdd gnd cell_6t
Xbit_r190_c30 bl[30] br[30] wl[190] vdd gnd cell_6t
Xbit_r191_c30 bl[30] br[30] wl[191] vdd gnd cell_6t
Xbit_r192_c30 bl[30] br[30] wl[192] vdd gnd cell_6t
Xbit_r193_c30 bl[30] br[30] wl[193] vdd gnd cell_6t
Xbit_r194_c30 bl[30] br[30] wl[194] vdd gnd cell_6t
Xbit_r195_c30 bl[30] br[30] wl[195] vdd gnd cell_6t
Xbit_r196_c30 bl[30] br[30] wl[196] vdd gnd cell_6t
Xbit_r197_c30 bl[30] br[30] wl[197] vdd gnd cell_6t
Xbit_r198_c30 bl[30] br[30] wl[198] vdd gnd cell_6t
Xbit_r199_c30 bl[30] br[30] wl[199] vdd gnd cell_6t
Xbit_r200_c30 bl[30] br[30] wl[200] vdd gnd cell_6t
Xbit_r201_c30 bl[30] br[30] wl[201] vdd gnd cell_6t
Xbit_r202_c30 bl[30] br[30] wl[202] vdd gnd cell_6t
Xbit_r203_c30 bl[30] br[30] wl[203] vdd gnd cell_6t
Xbit_r204_c30 bl[30] br[30] wl[204] vdd gnd cell_6t
Xbit_r205_c30 bl[30] br[30] wl[205] vdd gnd cell_6t
Xbit_r206_c30 bl[30] br[30] wl[206] vdd gnd cell_6t
Xbit_r207_c30 bl[30] br[30] wl[207] vdd gnd cell_6t
Xbit_r208_c30 bl[30] br[30] wl[208] vdd gnd cell_6t
Xbit_r209_c30 bl[30] br[30] wl[209] vdd gnd cell_6t
Xbit_r210_c30 bl[30] br[30] wl[210] vdd gnd cell_6t
Xbit_r211_c30 bl[30] br[30] wl[211] vdd gnd cell_6t
Xbit_r212_c30 bl[30] br[30] wl[212] vdd gnd cell_6t
Xbit_r213_c30 bl[30] br[30] wl[213] vdd gnd cell_6t
Xbit_r214_c30 bl[30] br[30] wl[214] vdd gnd cell_6t
Xbit_r215_c30 bl[30] br[30] wl[215] vdd gnd cell_6t
Xbit_r216_c30 bl[30] br[30] wl[216] vdd gnd cell_6t
Xbit_r217_c30 bl[30] br[30] wl[217] vdd gnd cell_6t
Xbit_r218_c30 bl[30] br[30] wl[218] vdd gnd cell_6t
Xbit_r219_c30 bl[30] br[30] wl[219] vdd gnd cell_6t
Xbit_r220_c30 bl[30] br[30] wl[220] vdd gnd cell_6t
Xbit_r221_c30 bl[30] br[30] wl[221] vdd gnd cell_6t
Xbit_r222_c30 bl[30] br[30] wl[222] vdd gnd cell_6t
Xbit_r223_c30 bl[30] br[30] wl[223] vdd gnd cell_6t
Xbit_r224_c30 bl[30] br[30] wl[224] vdd gnd cell_6t
Xbit_r225_c30 bl[30] br[30] wl[225] vdd gnd cell_6t
Xbit_r226_c30 bl[30] br[30] wl[226] vdd gnd cell_6t
Xbit_r227_c30 bl[30] br[30] wl[227] vdd gnd cell_6t
Xbit_r228_c30 bl[30] br[30] wl[228] vdd gnd cell_6t
Xbit_r229_c30 bl[30] br[30] wl[229] vdd gnd cell_6t
Xbit_r230_c30 bl[30] br[30] wl[230] vdd gnd cell_6t
Xbit_r231_c30 bl[30] br[30] wl[231] vdd gnd cell_6t
Xbit_r232_c30 bl[30] br[30] wl[232] vdd gnd cell_6t
Xbit_r233_c30 bl[30] br[30] wl[233] vdd gnd cell_6t
Xbit_r234_c30 bl[30] br[30] wl[234] vdd gnd cell_6t
Xbit_r235_c30 bl[30] br[30] wl[235] vdd gnd cell_6t
Xbit_r236_c30 bl[30] br[30] wl[236] vdd gnd cell_6t
Xbit_r237_c30 bl[30] br[30] wl[237] vdd gnd cell_6t
Xbit_r238_c30 bl[30] br[30] wl[238] vdd gnd cell_6t
Xbit_r239_c30 bl[30] br[30] wl[239] vdd gnd cell_6t
Xbit_r240_c30 bl[30] br[30] wl[240] vdd gnd cell_6t
Xbit_r241_c30 bl[30] br[30] wl[241] vdd gnd cell_6t
Xbit_r242_c30 bl[30] br[30] wl[242] vdd gnd cell_6t
Xbit_r243_c30 bl[30] br[30] wl[243] vdd gnd cell_6t
Xbit_r244_c30 bl[30] br[30] wl[244] vdd gnd cell_6t
Xbit_r245_c30 bl[30] br[30] wl[245] vdd gnd cell_6t
Xbit_r246_c30 bl[30] br[30] wl[246] vdd gnd cell_6t
Xbit_r247_c30 bl[30] br[30] wl[247] vdd gnd cell_6t
Xbit_r248_c30 bl[30] br[30] wl[248] vdd gnd cell_6t
Xbit_r249_c30 bl[30] br[30] wl[249] vdd gnd cell_6t
Xbit_r250_c30 bl[30] br[30] wl[250] vdd gnd cell_6t
Xbit_r251_c30 bl[30] br[30] wl[251] vdd gnd cell_6t
Xbit_r252_c30 bl[30] br[30] wl[252] vdd gnd cell_6t
Xbit_r253_c30 bl[30] br[30] wl[253] vdd gnd cell_6t
Xbit_r254_c30 bl[30] br[30] wl[254] vdd gnd cell_6t
Xbit_r255_c30 bl[30] br[30] wl[255] vdd gnd cell_6t
Xbit_r0_c31 bl[31] br[31] wl[0] vdd gnd cell_6t
Xbit_r1_c31 bl[31] br[31] wl[1] vdd gnd cell_6t
Xbit_r2_c31 bl[31] br[31] wl[2] vdd gnd cell_6t
Xbit_r3_c31 bl[31] br[31] wl[3] vdd gnd cell_6t
Xbit_r4_c31 bl[31] br[31] wl[4] vdd gnd cell_6t
Xbit_r5_c31 bl[31] br[31] wl[5] vdd gnd cell_6t
Xbit_r6_c31 bl[31] br[31] wl[6] vdd gnd cell_6t
Xbit_r7_c31 bl[31] br[31] wl[7] vdd gnd cell_6t
Xbit_r8_c31 bl[31] br[31] wl[8] vdd gnd cell_6t
Xbit_r9_c31 bl[31] br[31] wl[9] vdd gnd cell_6t
Xbit_r10_c31 bl[31] br[31] wl[10] vdd gnd cell_6t
Xbit_r11_c31 bl[31] br[31] wl[11] vdd gnd cell_6t
Xbit_r12_c31 bl[31] br[31] wl[12] vdd gnd cell_6t
Xbit_r13_c31 bl[31] br[31] wl[13] vdd gnd cell_6t
Xbit_r14_c31 bl[31] br[31] wl[14] vdd gnd cell_6t
Xbit_r15_c31 bl[31] br[31] wl[15] vdd gnd cell_6t
Xbit_r16_c31 bl[31] br[31] wl[16] vdd gnd cell_6t
Xbit_r17_c31 bl[31] br[31] wl[17] vdd gnd cell_6t
Xbit_r18_c31 bl[31] br[31] wl[18] vdd gnd cell_6t
Xbit_r19_c31 bl[31] br[31] wl[19] vdd gnd cell_6t
Xbit_r20_c31 bl[31] br[31] wl[20] vdd gnd cell_6t
Xbit_r21_c31 bl[31] br[31] wl[21] vdd gnd cell_6t
Xbit_r22_c31 bl[31] br[31] wl[22] vdd gnd cell_6t
Xbit_r23_c31 bl[31] br[31] wl[23] vdd gnd cell_6t
Xbit_r24_c31 bl[31] br[31] wl[24] vdd gnd cell_6t
Xbit_r25_c31 bl[31] br[31] wl[25] vdd gnd cell_6t
Xbit_r26_c31 bl[31] br[31] wl[26] vdd gnd cell_6t
Xbit_r27_c31 bl[31] br[31] wl[27] vdd gnd cell_6t
Xbit_r28_c31 bl[31] br[31] wl[28] vdd gnd cell_6t
Xbit_r29_c31 bl[31] br[31] wl[29] vdd gnd cell_6t
Xbit_r30_c31 bl[31] br[31] wl[30] vdd gnd cell_6t
Xbit_r31_c31 bl[31] br[31] wl[31] vdd gnd cell_6t
Xbit_r32_c31 bl[31] br[31] wl[32] vdd gnd cell_6t
Xbit_r33_c31 bl[31] br[31] wl[33] vdd gnd cell_6t
Xbit_r34_c31 bl[31] br[31] wl[34] vdd gnd cell_6t
Xbit_r35_c31 bl[31] br[31] wl[35] vdd gnd cell_6t
Xbit_r36_c31 bl[31] br[31] wl[36] vdd gnd cell_6t
Xbit_r37_c31 bl[31] br[31] wl[37] vdd gnd cell_6t
Xbit_r38_c31 bl[31] br[31] wl[38] vdd gnd cell_6t
Xbit_r39_c31 bl[31] br[31] wl[39] vdd gnd cell_6t
Xbit_r40_c31 bl[31] br[31] wl[40] vdd gnd cell_6t
Xbit_r41_c31 bl[31] br[31] wl[41] vdd gnd cell_6t
Xbit_r42_c31 bl[31] br[31] wl[42] vdd gnd cell_6t
Xbit_r43_c31 bl[31] br[31] wl[43] vdd gnd cell_6t
Xbit_r44_c31 bl[31] br[31] wl[44] vdd gnd cell_6t
Xbit_r45_c31 bl[31] br[31] wl[45] vdd gnd cell_6t
Xbit_r46_c31 bl[31] br[31] wl[46] vdd gnd cell_6t
Xbit_r47_c31 bl[31] br[31] wl[47] vdd gnd cell_6t
Xbit_r48_c31 bl[31] br[31] wl[48] vdd gnd cell_6t
Xbit_r49_c31 bl[31] br[31] wl[49] vdd gnd cell_6t
Xbit_r50_c31 bl[31] br[31] wl[50] vdd gnd cell_6t
Xbit_r51_c31 bl[31] br[31] wl[51] vdd gnd cell_6t
Xbit_r52_c31 bl[31] br[31] wl[52] vdd gnd cell_6t
Xbit_r53_c31 bl[31] br[31] wl[53] vdd gnd cell_6t
Xbit_r54_c31 bl[31] br[31] wl[54] vdd gnd cell_6t
Xbit_r55_c31 bl[31] br[31] wl[55] vdd gnd cell_6t
Xbit_r56_c31 bl[31] br[31] wl[56] vdd gnd cell_6t
Xbit_r57_c31 bl[31] br[31] wl[57] vdd gnd cell_6t
Xbit_r58_c31 bl[31] br[31] wl[58] vdd gnd cell_6t
Xbit_r59_c31 bl[31] br[31] wl[59] vdd gnd cell_6t
Xbit_r60_c31 bl[31] br[31] wl[60] vdd gnd cell_6t
Xbit_r61_c31 bl[31] br[31] wl[61] vdd gnd cell_6t
Xbit_r62_c31 bl[31] br[31] wl[62] vdd gnd cell_6t
Xbit_r63_c31 bl[31] br[31] wl[63] vdd gnd cell_6t
Xbit_r64_c31 bl[31] br[31] wl[64] vdd gnd cell_6t
Xbit_r65_c31 bl[31] br[31] wl[65] vdd gnd cell_6t
Xbit_r66_c31 bl[31] br[31] wl[66] vdd gnd cell_6t
Xbit_r67_c31 bl[31] br[31] wl[67] vdd gnd cell_6t
Xbit_r68_c31 bl[31] br[31] wl[68] vdd gnd cell_6t
Xbit_r69_c31 bl[31] br[31] wl[69] vdd gnd cell_6t
Xbit_r70_c31 bl[31] br[31] wl[70] vdd gnd cell_6t
Xbit_r71_c31 bl[31] br[31] wl[71] vdd gnd cell_6t
Xbit_r72_c31 bl[31] br[31] wl[72] vdd gnd cell_6t
Xbit_r73_c31 bl[31] br[31] wl[73] vdd gnd cell_6t
Xbit_r74_c31 bl[31] br[31] wl[74] vdd gnd cell_6t
Xbit_r75_c31 bl[31] br[31] wl[75] vdd gnd cell_6t
Xbit_r76_c31 bl[31] br[31] wl[76] vdd gnd cell_6t
Xbit_r77_c31 bl[31] br[31] wl[77] vdd gnd cell_6t
Xbit_r78_c31 bl[31] br[31] wl[78] vdd gnd cell_6t
Xbit_r79_c31 bl[31] br[31] wl[79] vdd gnd cell_6t
Xbit_r80_c31 bl[31] br[31] wl[80] vdd gnd cell_6t
Xbit_r81_c31 bl[31] br[31] wl[81] vdd gnd cell_6t
Xbit_r82_c31 bl[31] br[31] wl[82] vdd gnd cell_6t
Xbit_r83_c31 bl[31] br[31] wl[83] vdd gnd cell_6t
Xbit_r84_c31 bl[31] br[31] wl[84] vdd gnd cell_6t
Xbit_r85_c31 bl[31] br[31] wl[85] vdd gnd cell_6t
Xbit_r86_c31 bl[31] br[31] wl[86] vdd gnd cell_6t
Xbit_r87_c31 bl[31] br[31] wl[87] vdd gnd cell_6t
Xbit_r88_c31 bl[31] br[31] wl[88] vdd gnd cell_6t
Xbit_r89_c31 bl[31] br[31] wl[89] vdd gnd cell_6t
Xbit_r90_c31 bl[31] br[31] wl[90] vdd gnd cell_6t
Xbit_r91_c31 bl[31] br[31] wl[91] vdd gnd cell_6t
Xbit_r92_c31 bl[31] br[31] wl[92] vdd gnd cell_6t
Xbit_r93_c31 bl[31] br[31] wl[93] vdd gnd cell_6t
Xbit_r94_c31 bl[31] br[31] wl[94] vdd gnd cell_6t
Xbit_r95_c31 bl[31] br[31] wl[95] vdd gnd cell_6t
Xbit_r96_c31 bl[31] br[31] wl[96] vdd gnd cell_6t
Xbit_r97_c31 bl[31] br[31] wl[97] vdd gnd cell_6t
Xbit_r98_c31 bl[31] br[31] wl[98] vdd gnd cell_6t
Xbit_r99_c31 bl[31] br[31] wl[99] vdd gnd cell_6t
Xbit_r100_c31 bl[31] br[31] wl[100] vdd gnd cell_6t
Xbit_r101_c31 bl[31] br[31] wl[101] vdd gnd cell_6t
Xbit_r102_c31 bl[31] br[31] wl[102] vdd gnd cell_6t
Xbit_r103_c31 bl[31] br[31] wl[103] vdd gnd cell_6t
Xbit_r104_c31 bl[31] br[31] wl[104] vdd gnd cell_6t
Xbit_r105_c31 bl[31] br[31] wl[105] vdd gnd cell_6t
Xbit_r106_c31 bl[31] br[31] wl[106] vdd gnd cell_6t
Xbit_r107_c31 bl[31] br[31] wl[107] vdd gnd cell_6t
Xbit_r108_c31 bl[31] br[31] wl[108] vdd gnd cell_6t
Xbit_r109_c31 bl[31] br[31] wl[109] vdd gnd cell_6t
Xbit_r110_c31 bl[31] br[31] wl[110] vdd gnd cell_6t
Xbit_r111_c31 bl[31] br[31] wl[111] vdd gnd cell_6t
Xbit_r112_c31 bl[31] br[31] wl[112] vdd gnd cell_6t
Xbit_r113_c31 bl[31] br[31] wl[113] vdd gnd cell_6t
Xbit_r114_c31 bl[31] br[31] wl[114] vdd gnd cell_6t
Xbit_r115_c31 bl[31] br[31] wl[115] vdd gnd cell_6t
Xbit_r116_c31 bl[31] br[31] wl[116] vdd gnd cell_6t
Xbit_r117_c31 bl[31] br[31] wl[117] vdd gnd cell_6t
Xbit_r118_c31 bl[31] br[31] wl[118] vdd gnd cell_6t
Xbit_r119_c31 bl[31] br[31] wl[119] vdd gnd cell_6t
Xbit_r120_c31 bl[31] br[31] wl[120] vdd gnd cell_6t
Xbit_r121_c31 bl[31] br[31] wl[121] vdd gnd cell_6t
Xbit_r122_c31 bl[31] br[31] wl[122] vdd gnd cell_6t
Xbit_r123_c31 bl[31] br[31] wl[123] vdd gnd cell_6t
Xbit_r124_c31 bl[31] br[31] wl[124] vdd gnd cell_6t
Xbit_r125_c31 bl[31] br[31] wl[125] vdd gnd cell_6t
Xbit_r126_c31 bl[31] br[31] wl[126] vdd gnd cell_6t
Xbit_r127_c31 bl[31] br[31] wl[127] vdd gnd cell_6t
Xbit_r128_c31 bl[31] br[31] wl[128] vdd gnd cell_6t
Xbit_r129_c31 bl[31] br[31] wl[129] vdd gnd cell_6t
Xbit_r130_c31 bl[31] br[31] wl[130] vdd gnd cell_6t
Xbit_r131_c31 bl[31] br[31] wl[131] vdd gnd cell_6t
Xbit_r132_c31 bl[31] br[31] wl[132] vdd gnd cell_6t
Xbit_r133_c31 bl[31] br[31] wl[133] vdd gnd cell_6t
Xbit_r134_c31 bl[31] br[31] wl[134] vdd gnd cell_6t
Xbit_r135_c31 bl[31] br[31] wl[135] vdd gnd cell_6t
Xbit_r136_c31 bl[31] br[31] wl[136] vdd gnd cell_6t
Xbit_r137_c31 bl[31] br[31] wl[137] vdd gnd cell_6t
Xbit_r138_c31 bl[31] br[31] wl[138] vdd gnd cell_6t
Xbit_r139_c31 bl[31] br[31] wl[139] vdd gnd cell_6t
Xbit_r140_c31 bl[31] br[31] wl[140] vdd gnd cell_6t
Xbit_r141_c31 bl[31] br[31] wl[141] vdd gnd cell_6t
Xbit_r142_c31 bl[31] br[31] wl[142] vdd gnd cell_6t
Xbit_r143_c31 bl[31] br[31] wl[143] vdd gnd cell_6t
Xbit_r144_c31 bl[31] br[31] wl[144] vdd gnd cell_6t
Xbit_r145_c31 bl[31] br[31] wl[145] vdd gnd cell_6t
Xbit_r146_c31 bl[31] br[31] wl[146] vdd gnd cell_6t
Xbit_r147_c31 bl[31] br[31] wl[147] vdd gnd cell_6t
Xbit_r148_c31 bl[31] br[31] wl[148] vdd gnd cell_6t
Xbit_r149_c31 bl[31] br[31] wl[149] vdd gnd cell_6t
Xbit_r150_c31 bl[31] br[31] wl[150] vdd gnd cell_6t
Xbit_r151_c31 bl[31] br[31] wl[151] vdd gnd cell_6t
Xbit_r152_c31 bl[31] br[31] wl[152] vdd gnd cell_6t
Xbit_r153_c31 bl[31] br[31] wl[153] vdd gnd cell_6t
Xbit_r154_c31 bl[31] br[31] wl[154] vdd gnd cell_6t
Xbit_r155_c31 bl[31] br[31] wl[155] vdd gnd cell_6t
Xbit_r156_c31 bl[31] br[31] wl[156] vdd gnd cell_6t
Xbit_r157_c31 bl[31] br[31] wl[157] vdd gnd cell_6t
Xbit_r158_c31 bl[31] br[31] wl[158] vdd gnd cell_6t
Xbit_r159_c31 bl[31] br[31] wl[159] vdd gnd cell_6t
Xbit_r160_c31 bl[31] br[31] wl[160] vdd gnd cell_6t
Xbit_r161_c31 bl[31] br[31] wl[161] vdd gnd cell_6t
Xbit_r162_c31 bl[31] br[31] wl[162] vdd gnd cell_6t
Xbit_r163_c31 bl[31] br[31] wl[163] vdd gnd cell_6t
Xbit_r164_c31 bl[31] br[31] wl[164] vdd gnd cell_6t
Xbit_r165_c31 bl[31] br[31] wl[165] vdd gnd cell_6t
Xbit_r166_c31 bl[31] br[31] wl[166] vdd gnd cell_6t
Xbit_r167_c31 bl[31] br[31] wl[167] vdd gnd cell_6t
Xbit_r168_c31 bl[31] br[31] wl[168] vdd gnd cell_6t
Xbit_r169_c31 bl[31] br[31] wl[169] vdd gnd cell_6t
Xbit_r170_c31 bl[31] br[31] wl[170] vdd gnd cell_6t
Xbit_r171_c31 bl[31] br[31] wl[171] vdd gnd cell_6t
Xbit_r172_c31 bl[31] br[31] wl[172] vdd gnd cell_6t
Xbit_r173_c31 bl[31] br[31] wl[173] vdd gnd cell_6t
Xbit_r174_c31 bl[31] br[31] wl[174] vdd gnd cell_6t
Xbit_r175_c31 bl[31] br[31] wl[175] vdd gnd cell_6t
Xbit_r176_c31 bl[31] br[31] wl[176] vdd gnd cell_6t
Xbit_r177_c31 bl[31] br[31] wl[177] vdd gnd cell_6t
Xbit_r178_c31 bl[31] br[31] wl[178] vdd gnd cell_6t
Xbit_r179_c31 bl[31] br[31] wl[179] vdd gnd cell_6t
Xbit_r180_c31 bl[31] br[31] wl[180] vdd gnd cell_6t
Xbit_r181_c31 bl[31] br[31] wl[181] vdd gnd cell_6t
Xbit_r182_c31 bl[31] br[31] wl[182] vdd gnd cell_6t
Xbit_r183_c31 bl[31] br[31] wl[183] vdd gnd cell_6t
Xbit_r184_c31 bl[31] br[31] wl[184] vdd gnd cell_6t
Xbit_r185_c31 bl[31] br[31] wl[185] vdd gnd cell_6t
Xbit_r186_c31 bl[31] br[31] wl[186] vdd gnd cell_6t
Xbit_r187_c31 bl[31] br[31] wl[187] vdd gnd cell_6t
Xbit_r188_c31 bl[31] br[31] wl[188] vdd gnd cell_6t
Xbit_r189_c31 bl[31] br[31] wl[189] vdd gnd cell_6t
Xbit_r190_c31 bl[31] br[31] wl[190] vdd gnd cell_6t
Xbit_r191_c31 bl[31] br[31] wl[191] vdd gnd cell_6t
Xbit_r192_c31 bl[31] br[31] wl[192] vdd gnd cell_6t
Xbit_r193_c31 bl[31] br[31] wl[193] vdd gnd cell_6t
Xbit_r194_c31 bl[31] br[31] wl[194] vdd gnd cell_6t
Xbit_r195_c31 bl[31] br[31] wl[195] vdd gnd cell_6t
Xbit_r196_c31 bl[31] br[31] wl[196] vdd gnd cell_6t
Xbit_r197_c31 bl[31] br[31] wl[197] vdd gnd cell_6t
Xbit_r198_c31 bl[31] br[31] wl[198] vdd gnd cell_6t
Xbit_r199_c31 bl[31] br[31] wl[199] vdd gnd cell_6t
Xbit_r200_c31 bl[31] br[31] wl[200] vdd gnd cell_6t
Xbit_r201_c31 bl[31] br[31] wl[201] vdd gnd cell_6t
Xbit_r202_c31 bl[31] br[31] wl[202] vdd gnd cell_6t
Xbit_r203_c31 bl[31] br[31] wl[203] vdd gnd cell_6t
Xbit_r204_c31 bl[31] br[31] wl[204] vdd gnd cell_6t
Xbit_r205_c31 bl[31] br[31] wl[205] vdd gnd cell_6t
Xbit_r206_c31 bl[31] br[31] wl[206] vdd gnd cell_6t
Xbit_r207_c31 bl[31] br[31] wl[207] vdd gnd cell_6t
Xbit_r208_c31 bl[31] br[31] wl[208] vdd gnd cell_6t
Xbit_r209_c31 bl[31] br[31] wl[209] vdd gnd cell_6t
Xbit_r210_c31 bl[31] br[31] wl[210] vdd gnd cell_6t
Xbit_r211_c31 bl[31] br[31] wl[211] vdd gnd cell_6t
Xbit_r212_c31 bl[31] br[31] wl[212] vdd gnd cell_6t
Xbit_r213_c31 bl[31] br[31] wl[213] vdd gnd cell_6t
Xbit_r214_c31 bl[31] br[31] wl[214] vdd gnd cell_6t
Xbit_r215_c31 bl[31] br[31] wl[215] vdd gnd cell_6t
Xbit_r216_c31 bl[31] br[31] wl[216] vdd gnd cell_6t
Xbit_r217_c31 bl[31] br[31] wl[217] vdd gnd cell_6t
Xbit_r218_c31 bl[31] br[31] wl[218] vdd gnd cell_6t
Xbit_r219_c31 bl[31] br[31] wl[219] vdd gnd cell_6t
Xbit_r220_c31 bl[31] br[31] wl[220] vdd gnd cell_6t
Xbit_r221_c31 bl[31] br[31] wl[221] vdd gnd cell_6t
Xbit_r222_c31 bl[31] br[31] wl[222] vdd gnd cell_6t
Xbit_r223_c31 bl[31] br[31] wl[223] vdd gnd cell_6t
Xbit_r224_c31 bl[31] br[31] wl[224] vdd gnd cell_6t
Xbit_r225_c31 bl[31] br[31] wl[225] vdd gnd cell_6t
Xbit_r226_c31 bl[31] br[31] wl[226] vdd gnd cell_6t
Xbit_r227_c31 bl[31] br[31] wl[227] vdd gnd cell_6t
Xbit_r228_c31 bl[31] br[31] wl[228] vdd gnd cell_6t
Xbit_r229_c31 bl[31] br[31] wl[229] vdd gnd cell_6t
Xbit_r230_c31 bl[31] br[31] wl[230] vdd gnd cell_6t
Xbit_r231_c31 bl[31] br[31] wl[231] vdd gnd cell_6t
Xbit_r232_c31 bl[31] br[31] wl[232] vdd gnd cell_6t
Xbit_r233_c31 bl[31] br[31] wl[233] vdd gnd cell_6t
Xbit_r234_c31 bl[31] br[31] wl[234] vdd gnd cell_6t
Xbit_r235_c31 bl[31] br[31] wl[235] vdd gnd cell_6t
Xbit_r236_c31 bl[31] br[31] wl[236] vdd gnd cell_6t
Xbit_r237_c31 bl[31] br[31] wl[237] vdd gnd cell_6t
Xbit_r238_c31 bl[31] br[31] wl[238] vdd gnd cell_6t
Xbit_r239_c31 bl[31] br[31] wl[239] vdd gnd cell_6t
Xbit_r240_c31 bl[31] br[31] wl[240] vdd gnd cell_6t
Xbit_r241_c31 bl[31] br[31] wl[241] vdd gnd cell_6t
Xbit_r242_c31 bl[31] br[31] wl[242] vdd gnd cell_6t
Xbit_r243_c31 bl[31] br[31] wl[243] vdd gnd cell_6t
Xbit_r244_c31 bl[31] br[31] wl[244] vdd gnd cell_6t
Xbit_r245_c31 bl[31] br[31] wl[245] vdd gnd cell_6t
Xbit_r246_c31 bl[31] br[31] wl[246] vdd gnd cell_6t
Xbit_r247_c31 bl[31] br[31] wl[247] vdd gnd cell_6t
Xbit_r248_c31 bl[31] br[31] wl[248] vdd gnd cell_6t
Xbit_r249_c31 bl[31] br[31] wl[249] vdd gnd cell_6t
Xbit_r250_c31 bl[31] br[31] wl[250] vdd gnd cell_6t
Xbit_r251_c31 bl[31] br[31] wl[251] vdd gnd cell_6t
Xbit_r252_c31 bl[31] br[31] wl[252] vdd gnd cell_6t
Xbit_r253_c31 bl[31] br[31] wl[253] vdd gnd cell_6t
Xbit_r254_c31 bl[31] br[31] wl[254] vdd gnd cell_6t
Xbit_r255_c31 bl[31] br[31] wl[255] vdd gnd cell_6t
Xbit_r0_c32 bl[32] br[32] wl[0] vdd gnd cell_6t
Xbit_r1_c32 bl[32] br[32] wl[1] vdd gnd cell_6t
Xbit_r2_c32 bl[32] br[32] wl[2] vdd gnd cell_6t
Xbit_r3_c32 bl[32] br[32] wl[3] vdd gnd cell_6t
Xbit_r4_c32 bl[32] br[32] wl[4] vdd gnd cell_6t
Xbit_r5_c32 bl[32] br[32] wl[5] vdd gnd cell_6t
Xbit_r6_c32 bl[32] br[32] wl[6] vdd gnd cell_6t
Xbit_r7_c32 bl[32] br[32] wl[7] vdd gnd cell_6t
Xbit_r8_c32 bl[32] br[32] wl[8] vdd gnd cell_6t
Xbit_r9_c32 bl[32] br[32] wl[9] vdd gnd cell_6t
Xbit_r10_c32 bl[32] br[32] wl[10] vdd gnd cell_6t
Xbit_r11_c32 bl[32] br[32] wl[11] vdd gnd cell_6t
Xbit_r12_c32 bl[32] br[32] wl[12] vdd gnd cell_6t
Xbit_r13_c32 bl[32] br[32] wl[13] vdd gnd cell_6t
Xbit_r14_c32 bl[32] br[32] wl[14] vdd gnd cell_6t
Xbit_r15_c32 bl[32] br[32] wl[15] vdd gnd cell_6t
Xbit_r16_c32 bl[32] br[32] wl[16] vdd gnd cell_6t
Xbit_r17_c32 bl[32] br[32] wl[17] vdd gnd cell_6t
Xbit_r18_c32 bl[32] br[32] wl[18] vdd gnd cell_6t
Xbit_r19_c32 bl[32] br[32] wl[19] vdd gnd cell_6t
Xbit_r20_c32 bl[32] br[32] wl[20] vdd gnd cell_6t
Xbit_r21_c32 bl[32] br[32] wl[21] vdd gnd cell_6t
Xbit_r22_c32 bl[32] br[32] wl[22] vdd gnd cell_6t
Xbit_r23_c32 bl[32] br[32] wl[23] vdd gnd cell_6t
Xbit_r24_c32 bl[32] br[32] wl[24] vdd gnd cell_6t
Xbit_r25_c32 bl[32] br[32] wl[25] vdd gnd cell_6t
Xbit_r26_c32 bl[32] br[32] wl[26] vdd gnd cell_6t
Xbit_r27_c32 bl[32] br[32] wl[27] vdd gnd cell_6t
Xbit_r28_c32 bl[32] br[32] wl[28] vdd gnd cell_6t
Xbit_r29_c32 bl[32] br[32] wl[29] vdd gnd cell_6t
Xbit_r30_c32 bl[32] br[32] wl[30] vdd gnd cell_6t
Xbit_r31_c32 bl[32] br[32] wl[31] vdd gnd cell_6t
Xbit_r32_c32 bl[32] br[32] wl[32] vdd gnd cell_6t
Xbit_r33_c32 bl[32] br[32] wl[33] vdd gnd cell_6t
Xbit_r34_c32 bl[32] br[32] wl[34] vdd gnd cell_6t
Xbit_r35_c32 bl[32] br[32] wl[35] vdd gnd cell_6t
Xbit_r36_c32 bl[32] br[32] wl[36] vdd gnd cell_6t
Xbit_r37_c32 bl[32] br[32] wl[37] vdd gnd cell_6t
Xbit_r38_c32 bl[32] br[32] wl[38] vdd gnd cell_6t
Xbit_r39_c32 bl[32] br[32] wl[39] vdd gnd cell_6t
Xbit_r40_c32 bl[32] br[32] wl[40] vdd gnd cell_6t
Xbit_r41_c32 bl[32] br[32] wl[41] vdd gnd cell_6t
Xbit_r42_c32 bl[32] br[32] wl[42] vdd gnd cell_6t
Xbit_r43_c32 bl[32] br[32] wl[43] vdd gnd cell_6t
Xbit_r44_c32 bl[32] br[32] wl[44] vdd gnd cell_6t
Xbit_r45_c32 bl[32] br[32] wl[45] vdd gnd cell_6t
Xbit_r46_c32 bl[32] br[32] wl[46] vdd gnd cell_6t
Xbit_r47_c32 bl[32] br[32] wl[47] vdd gnd cell_6t
Xbit_r48_c32 bl[32] br[32] wl[48] vdd gnd cell_6t
Xbit_r49_c32 bl[32] br[32] wl[49] vdd gnd cell_6t
Xbit_r50_c32 bl[32] br[32] wl[50] vdd gnd cell_6t
Xbit_r51_c32 bl[32] br[32] wl[51] vdd gnd cell_6t
Xbit_r52_c32 bl[32] br[32] wl[52] vdd gnd cell_6t
Xbit_r53_c32 bl[32] br[32] wl[53] vdd gnd cell_6t
Xbit_r54_c32 bl[32] br[32] wl[54] vdd gnd cell_6t
Xbit_r55_c32 bl[32] br[32] wl[55] vdd gnd cell_6t
Xbit_r56_c32 bl[32] br[32] wl[56] vdd gnd cell_6t
Xbit_r57_c32 bl[32] br[32] wl[57] vdd gnd cell_6t
Xbit_r58_c32 bl[32] br[32] wl[58] vdd gnd cell_6t
Xbit_r59_c32 bl[32] br[32] wl[59] vdd gnd cell_6t
Xbit_r60_c32 bl[32] br[32] wl[60] vdd gnd cell_6t
Xbit_r61_c32 bl[32] br[32] wl[61] vdd gnd cell_6t
Xbit_r62_c32 bl[32] br[32] wl[62] vdd gnd cell_6t
Xbit_r63_c32 bl[32] br[32] wl[63] vdd gnd cell_6t
Xbit_r64_c32 bl[32] br[32] wl[64] vdd gnd cell_6t
Xbit_r65_c32 bl[32] br[32] wl[65] vdd gnd cell_6t
Xbit_r66_c32 bl[32] br[32] wl[66] vdd gnd cell_6t
Xbit_r67_c32 bl[32] br[32] wl[67] vdd gnd cell_6t
Xbit_r68_c32 bl[32] br[32] wl[68] vdd gnd cell_6t
Xbit_r69_c32 bl[32] br[32] wl[69] vdd gnd cell_6t
Xbit_r70_c32 bl[32] br[32] wl[70] vdd gnd cell_6t
Xbit_r71_c32 bl[32] br[32] wl[71] vdd gnd cell_6t
Xbit_r72_c32 bl[32] br[32] wl[72] vdd gnd cell_6t
Xbit_r73_c32 bl[32] br[32] wl[73] vdd gnd cell_6t
Xbit_r74_c32 bl[32] br[32] wl[74] vdd gnd cell_6t
Xbit_r75_c32 bl[32] br[32] wl[75] vdd gnd cell_6t
Xbit_r76_c32 bl[32] br[32] wl[76] vdd gnd cell_6t
Xbit_r77_c32 bl[32] br[32] wl[77] vdd gnd cell_6t
Xbit_r78_c32 bl[32] br[32] wl[78] vdd gnd cell_6t
Xbit_r79_c32 bl[32] br[32] wl[79] vdd gnd cell_6t
Xbit_r80_c32 bl[32] br[32] wl[80] vdd gnd cell_6t
Xbit_r81_c32 bl[32] br[32] wl[81] vdd gnd cell_6t
Xbit_r82_c32 bl[32] br[32] wl[82] vdd gnd cell_6t
Xbit_r83_c32 bl[32] br[32] wl[83] vdd gnd cell_6t
Xbit_r84_c32 bl[32] br[32] wl[84] vdd gnd cell_6t
Xbit_r85_c32 bl[32] br[32] wl[85] vdd gnd cell_6t
Xbit_r86_c32 bl[32] br[32] wl[86] vdd gnd cell_6t
Xbit_r87_c32 bl[32] br[32] wl[87] vdd gnd cell_6t
Xbit_r88_c32 bl[32] br[32] wl[88] vdd gnd cell_6t
Xbit_r89_c32 bl[32] br[32] wl[89] vdd gnd cell_6t
Xbit_r90_c32 bl[32] br[32] wl[90] vdd gnd cell_6t
Xbit_r91_c32 bl[32] br[32] wl[91] vdd gnd cell_6t
Xbit_r92_c32 bl[32] br[32] wl[92] vdd gnd cell_6t
Xbit_r93_c32 bl[32] br[32] wl[93] vdd gnd cell_6t
Xbit_r94_c32 bl[32] br[32] wl[94] vdd gnd cell_6t
Xbit_r95_c32 bl[32] br[32] wl[95] vdd gnd cell_6t
Xbit_r96_c32 bl[32] br[32] wl[96] vdd gnd cell_6t
Xbit_r97_c32 bl[32] br[32] wl[97] vdd gnd cell_6t
Xbit_r98_c32 bl[32] br[32] wl[98] vdd gnd cell_6t
Xbit_r99_c32 bl[32] br[32] wl[99] vdd gnd cell_6t
Xbit_r100_c32 bl[32] br[32] wl[100] vdd gnd cell_6t
Xbit_r101_c32 bl[32] br[32] wl[101] vdd gnd cell_6t
Xbit_r102_c32 bl[32] br[32] wl[102] vdd gnd cell_6t
Xbit_r103_c32 bl[32] br[32] wl[103] vdd gnd cell_6t
Xbit_r104_c32 bl[32] br[32] wl[104] vdd gnd cell_6t
Xbit_r105_c32 bl[32] br[32] wl[105] vdd gnd cell_6t
Xbit_r106_c32 bl[32] br[32] wl[106] vdd gnd cell_6t
Xbit_r107_c32 bl[32] br[32] wl[107] vdd gnd cell_6t
Xbit_r108_c32 bl[32] br[32] wl[108] vdd gnd cell_6t
Xbit_r109_c32 bl[32] br[32] wl[109] vdd gnd cell_6t
Xbit_r110_c32 bl[32] br[32] wl[110] vdd gnd cell_6t
Xbit_r111_c32 bl[32] br[32] wl[111] vdd gnd cell_6t
Xbit_r112_c32 bl[32] br[32] wl[112] vdd gnd cell_6t
Xbit_r113_c32 bl[32] br[32] wl[113] vdd gnd cell_6t
Xbit_r114_c32 bl[32] br[32] wl[114] vdd gnd cell_6t
Xbit_r115_c32 bl[32] br[32] wl[115] vdd gnd cell_6t
Xbit_r116_c32 bl[32] br[32] wl[116] vdd gnd cell_6t
Xbit_r117_c32 bl[32] br[32] wl[117] vdd gnd cell_6t
Xbit_r118_c32 bl[32] br[32] wl[118] vdd gnd cell_6t
Xbit_r119_c32 bl[32] br[32] wl[119] vdd gnd cell_6t
Xbit_r120_c32 bl[32] br[32] wl[120] vdd gnd cell_6t
Xbit_r121_c32 bl[32] br[32] wl[121] vdd gnd cell_6t
Xbit_r122_c32 bl[32] br[32] wl[122] vdd gnd cell_6t
Xbit_r123_c32 bl[32] br[32] wl[123] vdd gnd cell_6t
Xbit_r124_c32 bl[32] br[32] wl[124] vdd gnd cell_6t
Xbit_r125_c32 bl[32] br[32] wl[125] vdd gnd cell_6t
Xbit_r126_c32 bl[32] br[32] wl[126] vdd gnd cell_6t
Xbit_r127_c32 bl[32] br[32] wl[127] vdd gnd cell_6t
Xbit_r128_c32 bl[32] br[32] wl[128] vdd gnd cell_6t
Xbit_r129_c32 bl[32] br[32] wl[129] vdd gnd cell_6t
Xbit_r130_c32 bl[32] br[32] wl[130] vdd gnd cell_6t
Xbit_r131_c32 bl[32] br[32] wl[131] vdd gnd cell_6t
Xbit_r132_c32 bl[32] br[32] wl[132] vdd gnd cell_6t
Xbit_r133_c32 bl[32] br[32] wl[133] vdd gnd cell_6t
Xbit_r134_c32 bl[32] br[32] wl[134] vdd gnd cell_6t
Xbit_r135_c32 bl[32] br[32] wl[135] vdd gnd cell_6t
Xbit_r136_c32 bl[32] br[32] wl[136] vdd gnd cell_6t
Xbit_r137_c32 bl[32] br[32] wl[137] vdd gnd cell_6t
Xbit_r138_c32 bl[32] br[32] wl[138] vdd gnd cell_6t
Xbit_r139_c32 bl[32] br[32] wl[139] vdd gnd cell_6t
Xbit_r140_c32 bl[32] br[32] wl[140] vdd gnd cell_6t
Xbit_r141_c32 bl[32] br[32] wl[141] vdd gnd cell_6t
Xbit_r142_c32 bl[32] br[32] wl[142] vdd gnd cell_6t
Xbit_r143_c32 bl[32] br[32] wl[143] vdd gnd cell_6t
Xbit_r144_c32 bl[32] br[32] wl[144] vdd gnd cell_6t
Xbit_r145_c32 bl[32] br[32] wl[145] vdd gnd cell_6t
Xbit_r146_c32 bl[32] br[32] wl[146] vdd gnd cell_6t
Xbit_r147_c32 bl[32] br[32] wl[147] vdd gnd cell_6t
Xbit_r148_c32 bl[32] br[32] wl[148] vdd gnd cell_6t
Xbit_r149_c32 bl[32] br[32] wl[149] vdd gnd cell_6t
Xbit_r150_c32 bl[32] br[32] wl[150] vdd gnd cell_6t
Xbit_r151_c32 bl[32] br[32] wl[151] vdd gnd cell_6t
Xbit_r152_c32 bl[32] br[32] wl[152] vdd gnd cell_6t
Xbit_r153_c32 bl[32] br[32] wl[153] vdd gnd cell_6t
Xbit_r154_c32 bl[32] br[32] wl[154] vdd gnd cell_6t
Xbit_r155_c32 bl[32] br[32] wl[155] vdd gnd cell_6t
Xbit_r156_c32 bl[32] br[32] wl[156] vdd gnd cell_6t
Xbit_r157_c32 bl[32] br[32] wl[157] vdd gnd cell_6t
Xbit_r158_c32 bl[32] br[32] wl[158] vdd gnd cell_6t
Xbit_r159_c32 bl[32] br[32] wl[159] vdd gnd cell_6t
Xbit_r160_c32 bl[32] br[32] wl[160] vdd gnd cell_6t
Xbit_r161_c32 bl[32] br[32] wl[161] vdd gnd cell_6t
Xbit_r162_c32 bl[32] br[32] wl[162] vdd gnd cell_6t
Xbit_r163_c32 bl[32] br[32] wl[163] vdd gnd cell_6t
Xbit_r164_c32 bl[32] br[32] wl[164] vdd gnd cell_6t
Xbit_r165_c32 bl[32] br[32] wl[165] vdd gnd cell_6t
Xbit_r166_c32 bl[32] br[32] wl[166] vdd gnd cell_6t
Xbit_r167_c32 bl[32] br[32] wl[167] vdd gnd cell_6t
Xbit_r168_c32 bl[32] br[32] wl[168] vdd gnd cell_6t
Xbit_r169_c32 bl[32] br[32] wl[169] vdd gnd cell_6t
Xbit_r170_c32 bl[32] br[32] wl[170] vdd gnd cell_6t
Xbit_r171_c32 bl[32] br[32] wl[171] vdd gnd cell_6t
Xbit_r172_c32 bl[32] br[32] wl[172] vdd gnd cell_6t
Xbit_r173_c32 bl[32] br[32] wl[173] vdd gnd cell_6t
Xbit_r174_c32 bl[32] br[32] wl[174] vdd gnd cell_6t
Xbit_r175_c32 bl[32] br[32] wl[175] vdd gnd cell_6t
Xbit_r176_c32 bl[32] br[32] wl[176] vdd gnd cell_6t
Xbit_r177_c32 bl[32] br[32] wl[177] vdd gnd cell_6t
Xbit_r178_c32 bl[32] br[32] wl[178] vdd gnd cell_6t
Xbit_r179_c32 bl[32] br[32] wl[179] vdd gnd cell_6t
Xbit_r180_c32 bl[32] br[32] wl[180] vdd gnd cell_6t
Xbit_r181_c32 bl[32] br[32] wl[181] vdd gnd cell_6t
Xbit_r182_c32 bl[32] br[32] wl[182] vdd gnd cell_6t
Xbit_r183_c32 bl[32] br[32] wl[183] vdd gnd cell_6t
Xbit_r184_c32 bl[32] br[32] wl[184] vdd gnd cell_6t
Xbit_r185_c32 bl[32] br[32] wl[185] vdd gnd cell_6t
Xbit_r186_c32 bl[32] br[32] wl[186] vdd gnd cell_6t
Xbit_r187_c32 bl[32] br[32] wl[187] vdd gnd cell_6t
Xbit_r188_c32 bl[32] br[32] wl[188] vdd gnd cell_6t
Xbit_r189_c32 bl[32] br[32] wl[189] vdd gnd cell_6t
Xbit_r190_c32 bl[32] br[32] wl[190] vdd gnd cell_6t
Xbit_r191_c32 bl[32] br[32] wl[191] vdd gnd cell_6t
Xbit_r192_c32 bl[32] br[32] wl[192] vdd gnd cell_6t
Xbit_r193_c32 bl[32] br[32] wl[193] vdd gnd cell_6t
Xbit_r194_c32 bl[32] br[32] wl[194] vdd gnd cell_6t
Xbit_r195_c32 bl[32] br[32] wl[195] vdd gnd cell_6t
Xbit_r196_c32 bl[32] br[32] wl[196] vdd gnd cell_6t
Xbit_r197_c32 bl[32] br[32] wl[197] vdd gnd cell_6t
Xbit_r198_c32 bl[32] br[32] wl[198] vdd gnd cell_6t
Xbit_r199_c32 bl[32] br[32] wl[199] vdd gnd cell_6t
Xbit_r200_c32 bl[32] br[32] wl[200] vdd gnd cell_6t
Xbit_r201_c32 bl[32] br[32] wl[201] vdd gnd cell_6t
Xbit_r202_c32 bl[32] br[32] wl[202] vdd gnd cell_6t
Xbit_r203_c32 bl[32] br[32] wl[203] vdd gnd cell_6t
Xbit_r204_c32 bl[32] br[32] wl[204] vdd gnd cell_6t
Xbit_r205_c32 bl[32] br[32] wl[205] vdd gnd cell_6t
Xbit_r206_c32 bl[32] br[32] wl[206] vdd gnd cell_6t
Xbit_r207_c32 bl[32] br[32] wl[207] vdd gnd cell_6t
Xbit_r208_c32 bl[32] br[32] wl[208] vdd gnd cell_6t
Xbit_r209_c32 bl[32] br[32] wl[209] vdd gnd cell_6t
Xbit_r210_c32 bl[32] br[32] wl[210] vdd gnd cell_6t
Xbit_r211_c32 bl[32] br[32] wl[211] vdd gnd cell_6t
Xbit_r212_c32 bl[32] br[32] wl[212] vdd gnd cell_6t
Xbit_r213_c32 bl[32] br[32] wl[213] vdd gnd cell_6t
Xbit_r214_c32 bl[32] br[32] wl[214] vdd gnd cell_6t
Xbit_r215_c32 bl[32] br[32] wl[215] vdd gnd cell_6t
Xbit_r216_c32 bl[32] br[32] wl[216] vdd gnd cell_6t
Xbit_r217_c32 bl[32] br[32] wl[217] vdd gnd cell_6t
Xbit_r218_c32 bl[32] br[32] wl[218] vdd gnd cell_6t
Xbit_r219_c32 bl[32] br[32] wl[219] vdd gnd cell_6t
Xbit_r220_c32 bl[32] br[32] wl[220] vdd gnd cell_6t
Xbit_r221_c32 bl[32] br[32] wl[221] vdd gnd cell_6t
Xbit_r222_c32 bl[32] br[32] wl[222] vdd gnd cell_6t
Xbit_r223_c32 bl[32] br[32] wl[223] vdd gnd cell_6t
Xbit_r224_c32 bl[32] br[32] wl[224] vdd gnd cell_6t
Xbit_r225_c32 bl[32] br[32] wl[225] vdd gnd cell_6t
Xbit_r226_c32 bl[32] br[32] wl[226] vdd gnd cell_6t
Xbit_r227_c32 bl[32] br[32] wl[227] vdd gnd cell_6t
Xbit_r228_c32 bl[32] br[32] wl[228] vdd gnd cell_6t
Xbit_r229_c32 bl[32] br[32] wl[229] vdd gnd cell_6t
Xbit_r230_c32 bl[32] br[32] wl[230] vdd gnd cell_6t
Xbit_r231_c32 bl[32] br[32] wl[231] vdd gnd cell_6t
Xbit_r232_c32 bl[32] br[32] wl[232] vdd gnd cell_6t
Xbit_r233_c32 bl[32] br[32] wl[233] vdd gnd cell_6t
Xbit_r234_c32 bl[32] br[32] wl[234] vdd gnd cell_6t
Xbit_r235_c32 bl[32] br[32] wl[235] vdd gnd cell_6t
Xbit_r236_c32 bl[32] br[32] wl[236] vdd gnd cell_6t
Xbit_r237_c32 bl[32] br[32] wl[237] vdd gnd cell_6t
Xbit_r238_c32 bl[32] br[32] wl[238] vdd gnd cell_6t
Xbit_r239_c32 bl[32] br[32] wl[239] vdd gnd cell_6t
Xbit_r240_c32 bl[32] br[32] wl[240] vdd gnd cell_6t
Xbit_r241_c32 bl[32] br[32] wl[241] vdd gnd cell_6t
Xbit_r242_c32 bl[32] br[32] wl[242] vdd gnd cell_6t
Xbit_r243_c32 bl[32] br[32] wl[243] vdd gnd cell_6t
Xbit_r244_c32 bl[32] br[32] wl[244] vdd gnd cell_6t
Xbit_r245_c32 bl[32] br[32] wl[245] vdd gnd cell_6t
Xbit_r246_c32 bl[32] br[32] wl[246] vdd gnd cell_6t
Xbit_r247_c32 bl[32] br[32] wl[247] vdd gnd cell_6t
Xbit_r248_c32 bl[32] br[32] wl[248] vdd gnd cell_6t
Xbit_r249_c32 bl[32] br[32] wl[249] vdd gnd cell_6t
Xbit_r250_c32 bl[32] br[32] wl[250] vdd gnd cell_6t
Xbit_r251_c32 bl[32] br[32] wl[251] vdd gnd cell_6t
Xbit_r252_c32 bl[32] br[32] wl[252] vdd gnd cell_6t
Xbit_r253_c32 bl[32] br[32] wl[253] vdd gnd cell_6t
Xbit_r254_c32 bl[32] br[32] wl[254] vdd gnd cell_6t
Xbit_r255_c32 bl[32] br[32] wl[255] vdd gnd cell_6t
Xbit_r0_c33 bl[33] br[33] wl[0] vdd gnd cell_6t
Xbit_r1_c33 bl[33] br[33] wl[1] vdd gnd cell_6t
Xbit_r2_c33 bl[33] br[33] wl[2] vdd gnd cell_6t
Xbit_r3_c33 bl[33] br[33] wl[3] vdd gnd cell_6t
Xbit_r4_c33 bl[33] br[33] wl[4] vdd gnd cell_6t
Xbit_r5_c33 bl[33] br[33] wl[5] vdd gnd cell_6t
Xbit_r6_c33 bl[33] br[33] wl[6] vdd gnd cell_6t
Xbit_r7_c33 bl[33] br[33] wl[7] vdd gnd cell_6t
Xbit_r8_c33 bl[33] br[33] wl[8] vdd gnd cell_6t
Xbit_r9_c33 bl[33] br[33] wl[9] vdd gnd cell_6t
Xbit_r10_c33 bl[33] br[33] wl[10] vdd gnd cell_6t
Xbit_r11_c33 bl[33] br[33] wl[11] vdd gnd cell_6t
Xbit_r12_c33 bl[33] br[33] wl[12] vdd gnd cell_6t
Xbit_r13_c33 bl[33] br[33] wl[13] vdd gnd cell_6t
Xbit_r14_c33 bl[33] br[33] wl[14] vdd gnd cell_6t
Xbit_r15_c33 bl[33] br[33] wl[15] vdd gnd cell_6t
Xbit_r16_c33 bl[33] br[33] wl[16] vdd gnd cell_6t
Xbit_r17_c33 bl[33] br[33] wl[17] vdd gnd cell_6t
Xbit_r18_c33 bl[33] br[33] wl[18] vdd gnd cell_6t
Xbit_r19_c33 bl[33] br[33] wl[19] vdd gnd cell_6t
Xbit_r20_c33 bl[33] br[33] wl[20] vdd gnd cell_6t
Xbit_r21_c33 bl[33] br[33] wl[21] vdd gnd cell_6t
Xbit_r22_c33 bl[33] br[33] wl[22] vdd gnd cell_6t
Xbit_r23_c33 bl[33] br[33] wl[23] vdd gnd cell_6t
Xbit_r24_c33 bl[33] br[33] wl[24] vdd gnd cell_6t
Xbit_r25_c33 bl[33] br[33] wl[25] vdd gnd cell_6t
Xbit_r26_c33 bl[33] br[33] wl[26] vdd gnd cell_6t
Xbit_r27_c33 bl[33] br[33] wl[27] vdd gnd cell_6t
Xbit_r28_c33 bl[33] br[33] wl[28] vdd gnd cell_6t
Xbit_r29_c33 bl[33] br[33] wl[29] vdd gnd cell_6t
Xbit_r30_c33 bl[33] br[33] wl[30] vdd gnd cell_6t
Xbit_r31_c33 bl[33] br[33] wl[31] vdd gnd cell_6t
Xbit_r32_c33 bl[33] br[33] wl[32] vdd gnd cell_6t
Xbit_r33_c33 bl[33] br[33] wl[33] vdd gnd cell_6t
Xbit_r34_c33 bl[33] br[33] wl[34] vdd gnd cell_6t
Xbit_r35_c33 bl[33] br[33] wl[35] vdd gnd cell_6t
Xbit_r36_c33 bl[33] br[33] wl[36] vdd gnd cell_6t
Xbit_r37_c33 bl[33] br[33] wl[37] vdd gnd cell_6t
Xbit_r38_c33 bl[33] br[33] wl[38] vdd gnd cell_6t
Xbit_r39_c33 bl[33] br[33] wl[39] vdd gnd cell_6t
Xbit_r40_c33 bl[33] br[33] wl[40] vdd gnd cell_6t
Xbit_r41_c33 bl[33] br[33] wl[41] vdd gnd cell_6t
Xbit_r42_c33 bl[33] br[33] wl[42] vdd gnd cell_6t
Xbit_r43_c33 bl[33] br[33] wl[43] vdd gnd cell_6t
Xbit_r44_c33 bl[33] br[33] wl[44] vdd gnd cell_6t
Xbit_r45_c33 bl[33] br[33] wl[45] vdd gnd cell_6t
Xbit_r46_c33 bl[33] br[33] wl[46] vdd gnd cell_6t
Xbit_r47_c33 bl[33] br[33] wl[47] vdd gnd cell_6t
Xbit_r48_c33 bl[33] br[33] wl[48] vdd gnd cell_6t
Xbit_r49_c33 bl[33] br[33] wl[49] vdd gnd cell_6t
Xbit_r50_c33 bl[33] br[33] wl[50] vdd gnd cell_6t
Xbit_r51_c33 bl[33] br[33] wl[51] vdd gnd cell_6t
Xbit_r52_c33 bl[33] br[33] wl[52] vdd gnd cell_6t
Xbit_r53_c33 bl[33] br[33] wl[53] vdd gnd cell_6t
Xbit_r54_c33 bl[33] br[33] wl[54] vdd gnd cell_6t
Xbit_r55_c33 bl[33] br[33] wl[55] vdd gnd cell_6t
Xbit_r56_c33 bl[33] br[33] wl[56] vdd gnd cell_6t
Xbit_r57_c33 bl[33] br[33] wl[57] vdd gnd cell_6t
Xbit_r58_c33 bl[33] br[33] wl[58] vdd gnd cell_6t
Xbit_r59_c33 bl[33] br[33] wl[59] vdd gnd cell_6t
Xbit_r60_c33 bl[33] br[33] wl[60] vdd gnd cell_6t
Xbit_r61_c33 bl[33] br[33] wl[61] vdd gnd cell_6t
Xbit_r62_c33 bl[33] br[33] wl[62] vdd gnd cell_6t
Xbit_r63_c33 bl[33] br[33] wl[63] vdd gnd cell_6t
Xbit_r64_c33 bl[33] br[33] wl[64] vdd gnd cell_6t
Xbit_r65_c33 bl[33] br[33] wl[65] vdd gnd cell_6t
Xbit_r66_c33 bl[33] br[33] wl[66] vdd gnd cell_6t
Xbit_r67_c33 bl[33] br[33] wl[67] vdd gnd cell_6t
Xbit_r68_c33 bl[33] br[33] wl[68] vdd gnd cell_6t
Xbit_r69_c33 bl[33] br[33] wl[69] vdd gnd cell_6t
Xbit_r70_c33 bl[33] br[33] wl[70] vdd gnd cell_6t
Xbit_r71_c33 bl[33] br[33] wl[71] vdd gnd cell_6t
Xbit_r72_c33 bl[33] br[33] wl[72] vdd gnd cell_6t
Xbit_r73_c33 bl[33] br[33] wl[73] vdd gnd cell_6t
Xbit_r74_c33 bl[33] br[33] wl[74] vdd gnd cell_6t
Xbit_r75_c33 bl[33] br[33] wl[75] vdd gnd cell_6t
Xbit_r76_c33 bl[33] br[33] wl[76] vdd gnd cell_6t
Xbit_r77_c33 bl[33] br[33] wl[77] vdd gnd cell_6t
Xbit_r78_c33 bl[33] br[33] wl[78] vdd gnd cell_6t
Xbit_r79_c33 bl[33] br[33] wl[79] vdd gnd cell_6t
Xbit_r80_c33 bl[33] br[33] wl[80] vdd gnd cell_6t
Xbit_r81_c33 bl[33] br[33] wl[81] vdd gnd cell_6t
Xbit_r82_c33 bl[33] br[33] wl[82] vdd gnd cell_6t
Xbit_r83_c33 bl[33] br[33] wl[83] vdd gnd cell_6t
Xbit_r84_c33 bl[33] br[33] wl[84] vdd gnd cell_6t
Xbit_r85_c33 bl[33] br[33] wl[85] vdd gnd cell_6t
Xbit_r86_c33 bl[33] br[33] wl[86] vdd gnd cell_6t
Xbit_r87_c33 bl[33] br[33] wl[87] vdd gnd cell_6t
Xbit_r88_c33 bl[33] br[33] wl[88] vdd gnd cell_6t
Xbit_r89_c33 bl[33] br[33] wl[89] vdd gnd cell_6t
Xbit_r90_c33 bl[33] br[33] wl[90] vdd gnd cell_6t
Xbit_r91_c33 bl[33] br[33] wl[91] vdd gnd cell_6t
Xbit_r92_c33 bl[33] br[33] wl[92] vdd gnd cell_6t
Xbit_r93_c33 bl[33] br[33] wl[93] vdd gnd cell_6t
Xbit_r94_c33 bl[33] br[33] wl[94] vdd gnd cell_6t
Xbit_r95_c33 bl[33] br[33] wl[95] vdd gnd cell_6t
Xbit_r96_c33 bl[33] br[33] wl[96] vdd gnd cell_6t
Xbit_r97_c33 bl[33] br[33] wl[97] vdd gnd cell_6t
Xbit_r98_c33 bl[33] br[33] wl[98] vdd gnd cell_6t
Xbit_r99_c33 bl[33] br[33] wl[99] vdd gnd cell_6t
Xbit_r100_c33 bl[33] br[33] wl[100] vdd gnd cell_6t
Xbit_r101_c33 bl[33] br[33] wl[101] vdd gnd cell_6t
Xbit_r102_c33 bl[33] br[33] wl[102] vdd gnd cell_6t
Xbit_r103_c33 bl[33] br[33] wl[103] vdd gnd cell_6t
Xbit_r104_c33 bl[33] br[33] wl[104] vdd gnd cell_6t
Xbit_r105_c33 bl[33] br[33] wl[105] vdd gnd cell_6t
Xbit_r106_c33 bl[33] br[33] wl[106] vdd gnd cell_6t
Xbit_r107_c33 bl[33] br[33] wl[107] vdd gnd cell_6t
Xbit_r108_c33 bl[33] br[33] wl[108] vdd gnd cell_6t
Xbit_r109_c33 bl[33] br[33] wl[109] vdd gnd cell_6t
Xbit_r110_c33 bl[33] br[33] wl[110] vdd gnd cell_6t
Xbit_r111_c33 bl[33] br[33] wl[111] vdd gnd cell_6t
Xbit_r112_c33 bl[33] br[33] wl[112] vdd gnd cell_6t
Xbit_r113_c33 bl[33] br[33] wl[113] vdd gnd cell_6t
Xbit_r114_c33 bl[33] br[33] wl[114] vdd gnd cell_6t
Xbit_r115_c33 bl[33] br[33] wl[115] vdd gnd cell_6t
Xbit_r116_c33 bl[33] br[33] wl[116] vdd gnd cell_6t
Xbit_r117_c33 bl[33] br[33] wl[117] vdd gnd cell_6t
Xbit_r118_c33 bl[33] br[33] wl[118] vdd gnd cell_6t
Xbit_r119_c33 bl[33] br[33] wl[119] vdd gnd cell_6t
Xbit_r120_c33 bl[33] br[33] wl[120] vdd gnd cell_6t
Xbit_r121_c33 bl[33] br[33] wl[121] vdd gnd cell_6t
Xbit_r122_c33 bl[33] br[33] wl[122] vdd gnd cell_6t
Xbit_r123_c33 bl[33] br[33] wl[123] vdd gnd cell_6t
Xbit_r124_c33 bl[33] br[33] wl[124] vdd gnd cell_6t
Xbit_r125_c33 bl[33] br[33] wl[125] vdd gnd cell_6t
Xbit_r126_c33 bl[33] br[33] wl[126] vdd gnd cell_6t
Xbit_r127_c33 bl[33] br[33] wl[127] vdd gnd cell_6t
Xbit_r128_c33 bl[33] br[33] wl[128] vdd gnd cell_6t
Xbit_r129_c33 bl[33] br[33] wl[129] vdd gnd cell_6t
Xbit_r130_c33 bl[33] br[33] wl[130] vdd gnd cell_6t
Xbit_r131_c33 bl[33] br[33] wl[131] vdd gnd cell_6t
Xbit_r132_c33 bl[33] br[33] wl[132] vdd gnd cell_6t
Xbit_r133_c33 bl[33] br[33] wl[133] vdd gnd cell_6t
Xbit_r134_c33 bl[33] br[33] wl[134] vdd gnd cell_6t
Xbit_r135_c33 bl[33] br[33] wl[135] vdd gnd cell_6t
Xbit_r136_c33 bl[33] br[33] wl[136] vdd gnd cell_6t
Xbit_r137_c33 bl[33] br[33] wl[137] vdd gnd cell_6t
Xbit_r138_c33 bl[33] br[33] wl[138] vdd gnd cell_6t
Xbit_r139_c33 bl[33] br[33] wl[139] vdd gnd cell_6t
Xbit_r140_c33 bl[33] br[33] wl[140] vdd gnd cell_6t
Xbit_r141_c33 bl[33] br[33] wl[141] vdd gnd cell_6t
Xbit_r142_c33 bl[33] br[33] wl[142] vdd gnd cell_6t
Xbit_r143_c33 bl[33] br[33] wl[143] vdd gnd cell_6t
Xbit_r144_c33 bl[33] br[33] wl[144] vdd gnd cell_6t
Xbit_r145_c33 bl[33] br[33] wl[145] vdd gnd cell_6t
Xbit_r146_c33 bl[33] br[33] wl[146] vdd gnd cell_6t
Xbit_r147_c33 bl[33] br[33] wl[147] vdd gnd cell_6t
Xbit_r148_c33 bl[33] br[33] wl[148] vdd gnd cell_6t
Xbit_r149_c33 bl[33] br[33] wl[149] vdd gnd cell_6t
Xbit_r150_c33 bl[33] br[33] wl[150] vdd gnd cell_6t
Xbit_r151_c33 bl[33] br[33] wl[151] vdd gnd cell_6t
Xbit_r152_c33 bl[33] br[33] wl[152] vdd gnd cell_6t
Xbit_r153_c33 bl[33] br[33] wl[153] vdd gnd cell_6t
Xbit_r154_c33 bl[33] br[33] wl[154] vdd gnd cell_6t
Xbit_r155_c33 bl[33] br[33] wl[155] vdd gnd cell_6t
Xbit_r156_c33 bl[33] br[33] wl[156] vdd gnd cell_6t
Xbit_r157_c33 bl[33] br[33] wl[157] vdd gnd cell_6t
Xbit_r158_c33 bl[33] br[33] wl[158] vdd gnd cell_6t
Xbit_r159_c33 bl[33] br[33] wl[159] vdd gnd cell_6t
Xbit_r160_c33 bl[33] br[33] wl[160] vdd gnd cell_6t
Xbit_r161_c33 bl[33] br[33] wl[161] vdd gnd cell_6t
Xbit_r162_c33 bl[33] br[33] wl[162] vdd gnd cell_6t
Xbit_r163_c33 bl[33] br[33] wl[163] vdd gnd cell_6t
Xbit_r164_c33 bl[33] br[33] wl[164] vdd gnd cell_6t
Xbit_r165_c33 bl[33] br[33] wl[165] vdd gnd cell_6t
Xbit_r166_c33 bl[33] br[33] wl[166] vdd gnd cell_6t
Xbit_r167_c33 bl[33] br[33] wl[167] vdd gnd cell_6t
Xbit_r168_c33 bl[33] br[33] wl[168] vdd gnd cell_6t
Xbit_r169_c33 bl[33] br[33] wl[169] vdd gnd cell_6t
Xbit_r170_c33 bl[33] br[33] wl[170] vdd gnd cell_6t
Xbit_r171_c33 bl[33] br[33] wl[171] vdd gnd cell_6t
Xbit_r172_c33 bl[33] br[33] wl[172] vdd gnd cell_6t
Xbit_r173_c33 bl[33] br[33] wl[173] vdd gnd cell_6t
Xbit_r174_c33 bl[33] br[33] wl[174] vdd gnd cell_6t
Xbit_r175_c33 bl[33] br[33] wl[175] vdd gnd cell_6t
Xbit_r176_c33 bl[33] br[33] wl[176] vdd gnd cell_6t
Xbit_r177_c33 bl[33] br[33] wl[177] vdd gnd cell_6t
Xbit_r178_c33 bl[33] br[33] wl[178] vdd gnd cell_6t
Xbit_r179_c33 bl[33] br[33] wl[179] vdd gnd cell_6t
Xbit_r180_c33 bl[33] br[33] wl[180] vdd gnd cell_6t
Xbit_r181_c33 bl[33] br[33] wl[181] vdd gnd cell_6t
Xbit_r182_c33 bl[33] br[33] wl[182] vdd gnd cell_6t
Xbit_r183_c33 bl[33] br[33] wl[183] vdd gnd cell_6t
Xbit_r184_c33 bl[33] br[33] wl[184] vdd gnd cell_6t
Xbit_r185_c33 bl[33] br[33] wl[185] vdd gnd cell_6t
Xbit_r186_c33 bl[33] br[33] wl[186] vdd gnd cell_6t
Xbit_r187_c33 bl[33] br[33] wl[187] vdd gnd cell_6t
Xbit_r188_c33 bl[33] br[33] wl[188] vdd gnd cell_6t
Xbit_r189_c33 bl[33] br[33] wl[189] vdd gnd cell_6t
Xbit_r190_c33 bl[33] br[33] wl[190] vdd gnd cell_6t
Xbit_r191_c33 bl[33] br[33] wl[191] vdd gnd cell_6t
Xbit_r192_c33 bl[33] br[33] wl[192] vdd gnd cell_6t
Xbit_r193_c33 bl[33] br[33] wl[193] vdd gnd cell_6t
Xbit_r194_c33 bl[33] br[33] wl[194] vdd gnd cell_6t
Xbit_r195_c33 bl[33] br[33] wl[195] vdd gnd cell_6t
Xbit_r196_c33 bl[33] br[33] wl[196] vdd gnd cell_6t
Xbit_r197_c33 bl[33] br[33] wl[197] vdd gnd cell_6t
Xbit_r198_c33 bl[33] br[33] wl[198] vdd gnd cell_6t
Xbit_r199_c33 bl[33] br[33] wl[199] vdd gnd cell_6t
Xbit_r200_c33 bl[33] br[33] wl[200] vdd gnd cell_6t
Xbit_r201_c33 bl[33] br[33] wl[201] vdd gnd cell_6t
Xbit_r202_c33 bl[33] br[33] wl[202] vdd gnd cell_6t
Xbit_r203_c33 bl[33] br[33] wl[203] vdd gnd cell_6t
Xbit_r204_c33 bl[33] br[33] wl[204] vdd gnd cell_6t
Xbit_r205_c33 bl[33] br[33] wl[205] vdd gnd cell_6t
Xbit_r206_c33 bl[33] br[33] wl[206] vdd gnd cell_6t
Xbit_r207_c33 bl[33] br[33] wl[207] vdd gnd cell_6t
Xbit_r208_c33 bl[33] br[33] wl[208] vdd gnd cell_6t
Xbit_r209_c33 bl[33] br[33] wl[209] vdd gnd cell_6t
Xbit_r210_c33 bl[33] br[33] wl[210] vdd gnd cell_6t
Xbit_r211_c33 bl[33] br[33] wl[211] vdd gnd cell_6t
Xbit_r212_c33 bl[33] br[33] wl[212] vdd gnd cell_6t
Xbit_r213_c33 bl[33] br[33] wl[213] vdd gnd cell_6t
Xbit_r214_c33 bl[33] br[33] wl[214] vdd gnd cell_6t
Xbit_r215_c33 bl[33] br[33] wl[215] vdd gnd cell_6t
Xbit_r216_c33 bl[33] br[33] wl[216] vdd gnd cell_6t
Xbit_r217_c33 bl[33] br[33] wl[217] vdd gnd cell_6t
Xbit_r218_c33 bl[33] br[33] wl[218] vdd gnd cell_6t
Xbit_r219_c33 bl[33] br[33] wl[219] vdd gnd cell_6t
Xbit_r220_c33 bl[33] br[33] wl[220] vdd gnd cell_6t
Xbit_r221_c33 bl[33] br[33] wl[221] vdd gnd cell_6t
Xbit_r222_c33 bl[33] br[33] wl[222] vdd gnd cell_6t
Xbit_r223_c33 bl[33] br[33] wl[223] vdd gnd cell_6t
Xbit_r224_c33 bl[33] br[33] wl[224] vdd gnd cell_6t
Xbit_r225_c33 bl[33] br[33] wl[225] vdd gnd cell_6t
Xbit_r226_c33 bl[33] br[33] wl[226] vdd gnd cell_6t
Xbit_r227_c33 bl[33] br[33] wl[227] vdd gnd cell_6t
Xbit_r228_c33 bl[33] br[33] wl[228] vdd gnd cell_6t
Xbit_r229_c33 bl[33] br[33] wl[229] vdd gnd cell_6t
Xbit_r230_c33 bl[33] br[33] wl[230] vdd gnd cell_6t
Xbit_r231_c33 bl[33] br[33] wl[231] vdd gnd cell_6t
Xbit_r232_c33 bl[33] br[33] wl[232] vdd gnd cell_6t
Xbit_r233_c33 bl[33] br[33] wl[233] vdd gnd cell_6t
Xbit_r234_c33 bl[33] br[33] wl[234] vdd gnd cell_6t
Xbit_r235_c33 bl[33] br[33] wl[235] vdd gnd cell_6t
Xbit_r236_c33 bl[33] br[33] wl[236] vdd gnd cell_6t
Xbit_r237_c33 bl[33] br[33] wl[237] vdd gnd cell_6t
Xbit_r238_c33 bl[33] br[33] wl[238] vdd gnd cell_6t
Xbit_r239_c33 bl[33] br[33] wl[239] vdd gnd cell_6t
Xbit_r240_c33 bl[33] br[33] wl[240] vdd gnd cell_6t
Xbit_r241_c33 bl[33] br[33] wl[241] vdd gnd cell_6t
Xbit_r242_c33 bl[33] br[33] wl[242] vdd gnd cell_6t
Xbit_r243_c33 bl[33] br[33] wl[243] vdd gnd cell_6t
Xbit_r244_c33 bl[33] br[33] wl[244] vdd gnd cell_6t
Xbit_r245_c33 bl[33] br[33] wl[245] vdd gnd cell_6t
Xbit_r246_c33 bl[33] br[33] wl[246] vdd gnd cell_6t
Xbit_r247_c33 bl[33] br[33] wl[247] vdd gnd cell_6t
Xbit_r248_c33 bl[33] br[33] wl[248] vdd gnd cell_6t
Xbit_r249_c33 bl[33] br[33] wl[249] vdd gnd cell_6t
Xbit_r250_c33 bl[33] br[33] wl[250] vdd gnd cell_6t
Xbit_r251_c33 bl[33] br[33] wl[251] vdd gnd cell_6t
Xbit_r252_c33 bl[33] br[33] wl[252] vdd gnd cell_6t
Xbit_r253_c33 bl[33] br[33] wl[253] vdd gnd cell_6t
Xbit_r254_c33 bl[33] br[33] wl[254] vdd gnd cell_6t
Xbit_r255_c33 bl[33] br[33] wl[255] vdd gnd cell_6t
Xbit_r0_c34 bl[34] br[34] wl[0] vdd gnd cell_6t
Xbit_r1_c34 bl[34] br[34] wl[1] vdd gnd cell_6t
Xbit_r2_c34 bl[34] br[34] wl[2] vdd gnd cell_6t
Xbit_r3_c34 bl[34] br[34] wl[3] vdd gnd cell_6t
Xbit_r4_c34 bl[34] br[34] wl[4] vdd gnd cell_6t
Xbit_r5_c34 bl[34] br[34] wl[5] vdd gnd cell_6t
Xbit_r6_c34 bl[34] br[34] wl[6] vdd gnd cell_6t
Xbit_r7_c34 bl[34] br[34] wl[7] vdd gnd cell_6t
Xbit_r8_c34 bl[34] br[34] wl[8] vdd gnd cell_6t
Xbit_r9_c34 bl[34] br[34] wl[9] vdd gnd cell_6t
Xbit_r10_c34 bl[34] br[34] wl[10] vdd gnd cell_6t
Xbit_r11_c34 bl[34] br[34] wl[11] vdd gnd cell_6t
Xbit_r12_c34 bl[34] br[34] wl[12] vdd gnd cell_6t
Xbit_r13_c34 bl[34] br[34] wl[13] vdd gnd cell_6t
Xbit_r14_c34 bl[34] br[34] wl[14] vdd gnd cell_6t
Xbit_r15_c34 bl[34] br[34] wl[15] vdd gnd cell_6t
Xbit_r16_c34 bl[34] br[34] wl[16] vdd gnd cell_6t
Xbit_r17_c34 bl[34] br[34] wl[17] vdd gnd cell_6t
Xbit_r18_c34 bl[34] br[34] wl[18] vdd gnd cell_6t
Xbit_r19_c34 bl[34] br[34] wl[19] vdd gnd cell_6t
Xbit_r20_c34 bl[34] br[34] wl[20] vdd gnd cell_6t
Xbit_r21_c34 bl[34] br[34] wl[21] vdd gnd cell_6t
Xbit_r22_c34 bl[34] br[34] wl[22] vdd gnd cell_6t
Xbit_r23_c34 bl[34] br[34] wl[23] vdd gnd cell_6t
Xbit_r24_c34 bl[34] br[34] wl[24] vdd gnd cell_6t
Xbit_r25_c34 bl[34] br[34] wl[25] vdd gnd cell_6t
Xbit_r26_c34 bl[34] br[34] wl[26] vdd gnd cell_6t
Xbit_r27_c34 bl[34] br[34] wl[27] vdd gnd cell_6t
Xbit_r28_c34 bl[34] br[34] wl[28] vdd gnd cell_6t
Xbit_r29_c34 bl[34] br[34] wl[29] vdd gnd cell_6t
Xbit_r30_c34 bl[34] br[34] wl[30] vdd gnd cell_6t
Xbit_r31_c34 bl[34] br[34] wl[31] vdd gnd cell_6t
Xbit_r32_c34 bl[34] br[34] wl[32] vdd gnd cell_6t
Xbit_r33_c34 bl[34] br[34] wl[33] vdd gnd cell_6t
Xbit_r34_c34 bl[34] br[34] wl[34] vdd gnd cell_6t
Xbit_r35_c34 bl[34] br[34] wl[35] vdd gnd cell_6t
Xbit_r36_c34 bl[34] br[34] wl[36] vdd gnd cell_6t
Xbit_r37_c34 bl[34] br[34] wl[37] vdd gnd cell_6t
Xbit_r38_c34 bl[34] br[34] wl[38] vdd gnd cell_6t
Xbit_r39_c34 bl[34] br[34] wl[39] vdd gnd cell_6t
Xbit_r40_c34 bl[34] br[34] wl[40] vdd gnd cell_6t
Xbit_r41_c34 bl[34] br[34] wl[41] vdd gnd cell_6t
Xbit_r42_c34 bl[34] br[34] wl[42] vdd gnd cell_6t
Xbit_r43_c34 bl[34] br[34] wl[43] vdd gnd cell_6t
Xbit_r44_c34 bl[34] br[34] wl[44] vdd gnd cell_6t
Xbit_r45_c34 bl[34] br[34] wl[45] vdd gnd cell_6t
Xbit_r46_c34 bl[34] br[34] wl[46] vdd gnd cell_6t
Xbit_r47_c34 bl[34] br[34] wl[47] vdd gnd cell_6t
Xbit_r48_c34 bl[34] br[34] wl[48] vdd gnd cell_6t
Xbit_r49_c34 bl[34] br[34] wl[49] vdd gnd cell_6t
Xbit_r50_c34 bl[34] br[34] wl[50] vdd gnd cell_6t
Xbit_r51_c34 bl[34] br[34] wl[51] vdd gnd cell_6t
Xbit_r52_c34 bl[34] br[34] wl[52] vdd gnd cell_6t
Xbit_r53_c34 bl[34] br[34] wl[53] vdd gnd cell_6t
Xbit_r54_c34 bl[34] br[34] wl[54] vdd gnd cell_6t
Xbit_r55_c34 bl[34] br[34] wl[55] vdd gnd cell_6t
Xbit_r56_c34 bl[34] br[34] wl[56] vdd gnd cell_6t
Xbit_r57_c34 bl[34] br[34] wl[57] vdd gnd cell_6t
Xbit_r58_c34 bl[34] br[34] wl[58] vdd gnd cell_6t
Xbit_r59_c34 bl[34] br[34] wl[59] vdd gnd cell_6t
Xbit_r60_c34 bl[34] br[34] wl[60] vdd gnd cell_6t
Xbit_r61_c34 bl[34] br[34] wl[61] vdd gnd cell_6t
Xbit_r62_c34 bl[34] br[34] wl[62] vdd gnd cell_6t
Xbit_r63_c34 bl[34] br[34] wl[63] vdd gnd cell_6t
Xbit_r64_c34 bl[34] br[34] wl[64] vdd gnd cell_6t
Xbit_r65_c34 bl[34] br[34] wl[65] vdd gnd cell_6t
Xbit_r66_c34 bl[34] br[34] wl[66] vdd gnd cell_6t
Xbit_r67_c34 bl[34] br[34] wl[67] vdd gnd cell_6t
Xbit_r68_c34 bl[34] br[34] wl[68] vdd gnd cell_6t
Xbit_r69_c34 bl[34] br[34] wl[69] vdd gnd cell_6t
Xbit_r70_c34 bl[34] br[34] wl[70] vdd gnd cell_6t
Xbit_r71_c34 bl[34] br[34] wl[71] vdd gnd cell_6t
Xbit_r72_c34 bl[34] br[34] wl[72] vdd gnd cell_6t
Xbit_r73_c34 bl[34] br[34] wl[73] vdd gnd cell_6t
Xbit_r74_c34 bl[34] br[34] wl[74] vdd gnd cell_6t
Xbit_r75_c34 bl[34] br[34] wl[75] vdd gnd cell_6t
Xbit_r76_c34 bl[34] br[34] wl[76] vdd gnd cell_6t
Xbit_r77_c34 bl[34] br[34] wl[77] vdd gnd cell_6t
Xbit_r78_c34 bl[34] br[34] wl[78] vdd gnd cell_6t
Xbit_r79_c34 bl[34] br[34] wl[79] vdd gnd cell_6t
Xbit_r80_c34 bl[34] br[34] wl[80] vdd gnd cell_6t
Xbit_r81_c34 bl[34] br[34] wl[81] vdd gnd cell_6t
Xbit_r82_c34 bl[34] br[34] wl[82] vdd gnd cell_6t
Xbit_r83_c34 bl[34] br[34] wl[83] vdd gnd cell_6t
Xbit_r84_c34 bl[34] br[34] wl[84] vdd gnd cell_6t
Xbit_r85_c34 bl[34] br[34] wl[85] vdd gnd cell_6t
Xbit_r86_c34 bl[34] br[34] wl[86] vdd gnd cell_6t
Xbit_r87_c34 bl[34] br[34] wl[87] vdd gnd cell_6t
Xbit_r88_c34 bl[34] br[34] wl[88] vdd gnd cell_6t
Xbit_r89_c34 bl[34] br[34] wl[89] vdd gnd cell_6t
Xbit_r90_c34 bl[34] br[34] wl[90] vdd gnd cell_6t
Xbit_r91_c34 bl[34] br[34] wl[91] vdd gnd cell_6t
Xbit_r92_c34 bl[34] br[34] wl[92] vdd gnd cell_6t
Xbit_r93_c34 bl[34] br[34] wl[93] vdd gnd cell_6t
Xbit_r94_c34 bl[34] br[34] wl[94] vdd gnd cell_6t
Xbit_r95_c34 bl[34] br[34] wl[95] vdd gnd cell_6t
Xbit_r96_c34 bl[34] br[34] wl[96] vdd gnd cell_6t
Xbit_r97_c34 bl[34] br[34] wl[97] vdd gnd cell_6t
Xbit_r98_c34 bl[34] br[34] wl[98] vdd gnd cell_6t
Xbit_r99_c34 bl[34] br[34] wl[99] vdd gnd cell_6t
Xbit_r100_c34 bl[34] br[34] wl[100] vdd gnd cell_6t
Xbit_r101_c34 bl[34] br[34] wl[101] vdd gnd cell_6t
Xbit_r102_c34 bl[34] br[34] wl[102] vdd gnd cell_6t
Xbit_r103_c34 bl[34] br[34] wl[103] vdd gnd cell_6t
Xbit_r104_c34 bl[34] br[34] wl[104] vdd gnd cell_6t
Xbit_r105_c34 bl[34] br[34] wl[105] vdd gnd cell_6t
Xbit_r106_c34 bl[34] br[34] wl[106] vdd gnd cell_6t
Xbit_r107_c34 bl[34] br[34] wl[107] vdd gnd cell_6t
Xbit_r108_c34 bl[34] br[34] wl[108] vdd gnd cell_6t
Xbit_r109_c34 bl[34] br[34] wl[109] vdd gnd cell_6t
Xbit_r110_c34 bl[34] br[34] wl[110] vdd gnd cell_6t
Xbit_r111_c34 bl[34] br[34] wl[111] vdd gnd cell_6t
Xbit_r112_c34 bl[34] br[34] wl[112] vdd gnd cell_6t
Xbit_r113_c34 bl[34] br[34] wl[113] vdd gnd cell_6t
Xbit_r114_c34 bl[34] br[34] wl[114] vdd gnd cell_6t
Xbit_r115_c34 bl[34] br[34] wl[115] vdd gnd cell_6t
Xbit_r116_c34 bl[34] br[34] wl[116] vdd gnd cell_6t
Xbit_r117_c34 bl[34] br[34] wl[117] vdd gnd cell_6t
Xbit_r118_c34 bl[34] br[34] wl[118] vdd gnd cell_6t
Xbit_r119_c34 bl[34] br[34] wl[119] vdd gnd cell_6t
Xbit_r120_c34 bl[34] br[34] wl[120] vdd gnd cell_6t
Xbit_r121_c34 bl[34] br[34] wl[121] vdd gnd cell_6t
Xbit_r122_c34 bl[34] br[34] wl[122] vdd gnd cell_6t
Xbit_r123_c34 bl[34] br[34] wl[123] vdd gnd cell_6t
Xbit_r124_c34 bl[34] br[34] wl[124] vdd gnd cell_6t
Xbit_r125_c34 bl[34] br[34] wl[125] vdd gnd cell_6t
Xbit_r126_c34 bl[34] br[34] wl[126] vdd gnd cell_6t
Xbit_r127_c34 bl[34] br[34] wl[127] vdd gnd cell_6t
Xbit_r128_c34 bl[34] br[34] wl[128] vdd gnd cell_6t
Xbit_r129_c34 bl[34] br[34] wl[129] vdd gnd cell_6t
Xbit_r130_c34 bl[34] br[34] wl[130] vdd gnd cell_6t
Xbit_r131_c34 bl[34] br[34] wl[131] vdd gnd cell_6t
Xbit_r132_c34 bl[34] br[34] wl[132] vdd gnd cell_6t
Xbit_r133_c34 bl[34] br[34] wl[133] vdd gnd cell_6t
Xbit_r134_c34 bl[34] br[34] wl[134] vdd gnd cell_6t
Xbit_r135_c34 bl[34] br[34] wl[135] vdd gnd cell_6t
Xbit_r136_c34 bl[34] br[34] wl[136] vdd gnd cell_6t
Xbit_r137_c34 bl[34] br[34] wl[137] vdd gnd cell_6t
Xbit_r138_c34 bl[34] br[34] wl[138] vdd gnd cell_6t
Xbit_r139_c34 bl[34] br[34] wl[139] vdd gnd cell_6t
Xbit_r140_c34 bl[34] br[34] wl[140] vdd gnd cell_6t
Xbit_r141_c34 bl[34] br[34] wl[141] vdd gnd cell_6t
Xbit_r142_c34 bl[34] br[34] wl[142] vdd gnd cell_6t
Xbit_r143_c34 bl[34] br[34] wl[143] vdd gnd cell_6t
Xbit_r144_c34 bl[34] br[34] wl[144] vdd gnd cell_6t
Xbit_r145_c34 bl[34] br[34] wl[145] vdd gnd cell_6t
Xbit_r146_c34 bl[34] br[34] wl[146] vdd gnd cell_6t
Xbit_r147_c34 bl[34] br[34] wl[147] vdd gnd cell_6t
Xbit_r148_c34 bl[34] br[34] wl[148] vdd gnd cell_6t
Xbit_r149_c34 bl[34] br[34] wl[149] vdd gnd cell_6t
Xbit_r150_c34 bl[34] br[34] wl[150] vdd gnd cell_6t
Xbit_r151_c34 bl[34] br[34] wl[151] vdd gnd cell_6t
Xbit_r152_c34 bl[34] br[34] wl[152] vdd gnd cell_6t
Xbit_r153_c34 bl[34] br[34] wl[153] vdd gnd cell_6t
Xbit_r154_c34 bl[34] br[34] wl[154] vdd gnd cell_6t
Xbit_r155_c34 bl[34] br[34] wl[155] vdd gnd cell_6t
Xbit_r156_c34 bl[34] br[34] wl[156] vdd gnd cell_6t
Xbit_r157_c34 bl[34] br[34] wl[157] vdd gnd cell_6t
Xbit_r158_c34 bl[34] br[34] wl[158] vdd gnd cell_6t
Xbit_r159_c34 bl[34] br[34] wl[159] vdd gnd cell_6t
Xbit_r160_c34 bl[34] br[34] wl[160] vdd gnd cell_6t
Xbit_r161_c34 bl[34] br[34] wl[161] vdd gnd cell_6t
Xbit_r162_c34 bl[34] br[34] wl[162] vdd gnd cell_6t
Xbit_r163_c34 bl[34] br[34] wl[163] vdd gnd cell_6t
Xbit_r164_c34 bl[34] br[34] wl[164] vdd gnd cell_6t
Xbit_r165_c34 bl[34] br[34] wl[165] vdd gnd cell_6t
Xbit_r166_c34 bl[34] br[34] wl[166] vdd gnd cell_6t
Xbit_r167_c34 bl[34] br[34] wl[167] vdd gnd cell_6t
Xbit_r168_c34 bl[34] br[34] wl[168] vdd gnd cell_6t
Xbit_r169_c34 bl[34] br[34] wl[169] vdd gnd cell_6t
Xbit_r170_c34 bl[34] br[34] wl[170] vdd gnd cell_6t
Xbit_r171_c34 bl[34] br[34] wl[171] vdd gnd cell_6t
Xbit_r172_c34 bl[34] br[34] wl[172] vdd gnd cell_6t
Xbit_r173_c34 bl[34] br[34] wl[173] vdd gnd cell_6t
Xbit_r174_c34 bl[34] br[34] wl[174] vdd gnd cell_6t
Xbit_r175_c34 bl[34] br[34] wl[175] vdd gnd cell_6t
Xbit_r176_c34 bl[34] br[34] wl[176] vdd gnd cell_6t
Xbit_r177_c34 bl[34] br[34] wl[177] vdd gnd cell_6t
Xbit_r178_c34 bl[34] br[34] wl[178] vdd gnd cell_6t
Xbit_r179_c34 bl[34] br[34] wl[179] vdd gnd cell_6t
Xbit_r180_c34 bl[34] br[34] wl[180] vdd gnd cell_6t
Xbit_r181_c34 bl[34] br[34] wl[181] vdd gnd cell_6t
Xbit_r182_c34 bl[34] br[34] wl[182] vdd gnd cell_6t
Xbit_r183_c34 bl[34] br[34] wl[183] vdd gnd cell_6t
Xbit_r184_c34 bl[34] br[34] wl[184] vdd gnd cell_6t
Xbit_r185_c34 bl[34] br[34] wl[185] vdd gnd cell_6t
Xbit_r186_c34 bl[34] br[34] wl[186] vdd gnd cell_6t
Xbit_r187_c34 bl[34] br[34] wl[187] vdd gnd cell_6t
Xbit_r188_c34 bl[34] br[34] wl[188] vdd gnd cell_6t
Xbit_r189_c34 bl[34] br[34] wl[189] vdd gnd cell_6t
Xbit_r190_c34 bl[34] br[34] wl[190] vdd gnd cell_6t
Xbit_r191_c34 bl[34] br[34] wl[191] vdd gnd cell_6t
Xbit_r192_c34 bl[34] br[34] wl[192] vdd gnd cell_6t
Xbit_r193_c34 bl[34] br[34] wl[193] vdd gnd cell_6t
Xbit_r194_c34 bl[34] br[34] wl[194] vdd gnd cell_6t
Xbit_r195_c34 bl[34] br[34] wl[195] vdd gnd cell_6t
Xbit_r196_c34 bl[34] br[34] wl[196] vdd gnd cell_6t
Xbit_r197_c34 bl[34] br[34] wl[197] vdd gnd cell_6t
Xbit_r198_c34 bl[34] br[34] wl[198] vdd gnd cell_6t
Xbit_r199_c34 bl[34] br[34] wl[199] vdd gnd cell_6t
Xbit_r200_c34 bl[34] br[34] wl[200] vdd gnd cell_6t
Xbit_r201_c34 bl[34] br[34] wl[201] vdd gnd cell_6t
Xbit_r202_c34 bl[34] br[34] wl[202] vdd gnd cell_6t
Xbit_r203_c34 bl[34] br[34] wl[203] vdd gnd cell_6t
Xbit_r204_c34 bl[34] br[34] wl[204] vdd gnd cell_6t
Xbit_r205_c34 bl[34] br[34] wl[205] vdd gnd cell_6t
Xbit_r206_c34 bl[34] br[34] wl[206] vdd gnd cell_6t
Xbit_r207_c34 bl[34] br[34] wl[207] vdd gnd cell_6t
Xbit_r208_c34 bl[34] br[34] wl[208] vdd gnd cell_6t
Xbit_r209_c34 bl[34] br[34] wl[209] vdd gnd cell_6t
Xbit_r210_c34 bl[34] br[34] wl[210] vdd gnd cell_6t
Xbit_r211_c34 bl[34] br[34] wl[211] vdd gnd cell_6t
Xbit_r212_c34 bl[34] br[34] wl[212] vdd gnd cell_6t
Xbit_r213_c34 bl[34] br[34] wl[213] vdd gnd cell_6t
Xbit_r214_c34 bl[34] br[34] wl[214] vdd gnd cell_6t
Xbit_r215_c34 bl[34] br[34] wl[215] vdd gnd cell_6t
Xbit_r216_c34 bl[34] br[34] wl[216] vdd gnd cell_6t
Xbit_r217_c34 bl[34] br[34] wl[217] vdd gnd cell_6t
Xbit_r218_c34 bl[34] br[34] wl[218] vdd gnd cell_6t
Xbit_r219_c34 bl[34] br[34] wl[219] vdd gnd cell_6t
Xbit_r220_c34 bl[34] br[34] wl[220] vdd gnd cell_6t
Xbit_r221_c34 bl[34] br[34] wl[221] vdd gnd cell_6t
Xbit_r222_c34 bl[34] br[34] wl[222] vdd gnd cell_6t
Xbit_r223_c34 bl[34] br[34] wl[223] vdd gnd cell_6t
Xbit_r224_c34 bl[34] br[34] wl[224] vdd gnd cell_6t
Xbit_r225_c34 bl[34] br[34] wl[225] vdd gnd cell_6t
Xbit_r226_c34 bl[34] br[34] wl[226] vdd gnd cell_6t
Xbit_r227_c34 bl[34] br[34] wl[227] vdd gnd cell_6t
Xbit_r228_c34 bl[34] br[34] wl[228] vdd gnd cell_6t
Xbit_r229_c34 bl[34] br[34] wl[229] vdd gnd cell_6t
Xbit_r230_c34 bl[34] br[34] wl[230] vdd gnd cell_6t
Xbit_r231_c34 bl[34] br[34] wl[231] vdd gnd cell_6t
Xbit_r232_c34 bl[34] br[34] wl[232] vdd gnd cell_6t
Xbit_r233_c34 bl[34] br[34] wl[233] vdd gnd cell_6t
Xbit_r234_c34 bl[34] br[34] wl[234] vdd gnd cell_6t
Xbit_r235_c34 bl[34] br[34] wl[235] vdd gnd cell_6t
Xbit_r236_c34 bl[34] br[34] wl[236] vdd gnd cell_6t
Xbit_r237_c34 bl[34] br[34] wl[237] vdd gnd cell_6t
Xbit_r238_c34 bl[34] br[34] wl[238] vdd gnd cell_6t
Xbit_r239_c34 bl[34] br[34] wl[239] vdd gnd cell_6t
Xbit_r240_c34 bl[34] br[34] wl[240] vdd gnd cell_6t
Xbit_r241_c34 bl[34] br[34] wl[241] vdd gnd cell_6t
Xbit_r242_c34 bl[34] br[34] wl[242] vdd gnd cell_6t
Xbit_r243_c34 bl[34] br[34] wl[243] vdd gnd cell_6t
Xbit_r244_c34 bl[34] br[34] wl[244] vdd gnd cell_6t
Xbit_r245_c34 bl[34] br[34] wl[245] vdd gnd cell_6t
Xbit_r246_c34 bl[34] br[34] wl[246] vdd gnd cell_6t
Xbit_r247_c34 bl[34] br[34] wl[247] vdd gnd cell_6t
Xbit_r248_c34 bl[34] br[34] wl[248] vdd gnd cell_6t
Xbit_r249_c34 bl[34] br[34] wl[249] vdd gnd cell_6t
Xbit_r250_c34 bl[34] br[34] wl[250] vdd gnd cell_6t
Xbit_r251_c34 bl[34] br[34] wl[251] vdd gnd cell_6t
Xbit_r252_c34 bl[34] br[34] wl[252] vdd gnd cell_6t
Xbit_r253_c34 bl[34] br[34] wl[253] vdd gnd cell_6t
Xbit_r254_c34 bl[34] br[34] wl[254] vdd gnd cell_6t
Xbit_r255_c34 bl[34] br[34] wl[255] vdd gnd cell_6t
Xbit_r0_c35 bl[35] br[35] wl[0] vdd gnd cell_6t
Xbit_r1_c35 bl[35] br[35] wl[1] vdd gnd cell_6t
Xbit_r2_c35 bl[35] br[35] wl[2] vdd gnd cell_6t
Xbit_r3_c35 bl[35] br[35] wl[3] vdd gnd cell_6t
Xbit_r4_c35 bl[35] br[35] wl[4] vdd gnd cell_6t
Xbit_r5_c35 bl[35] br[35] wl[5] vdd gnd cell_6t
Xbit_r6_c35 bl[35] br[35] wl[6] vdd gnd cell_6t
Xbit_r7_c35 bl[35] br[35] wl[7] vdd gnd cell_6t
Xbit_r8_c35 bl[35] br[35] wl[8] vdd gnd cell_6t
Xbit_r9_c35 bl[35] br[35] wl[9] vdd gnd cell_6t
Xbit_r10_c35 bl[35] br[35] wl[10] vdd gnd cell_6t
Xbit_r11_c35 bl[35] br[35] wl[11] vdd gnd cell_6t
Xbit_r12_c35 bl[35] br[35] wl[12] vdd gnd cell_6t
Xbit_r13_c35 bl[35] br[35] wl[13] vdd gnd cell_6t
Xbit_r14_c35 bl[35] br[35] wl[14] vdd gnd cell_6t
Xbit_r15_c35 bl[35] br[35] wl[15] vdd gnd cell_6t
Xbit_r16_c35 bl[35] br[35] wl[16] vdd gnd cell_6t
Xbit_r17_c35 bl[35] br[35] wl[17] vdd gnd cell_6t
Xbit_r18_c35 bl[35] br[35] wl[18] vdd gnd cell_6t
Xbit_r19_c35 bl[35] br[35] wl[19] vdd gnd cell_6t
Xbit_r20_c35 bl[35] br[35] wl[20] vdd gnd cell_6t
Xbit_r21_c35 bl[35] br[35] wl[21] vdd gnd cell_6t
Xbit_r22_c35 bl[35] br[35] wl[22] vdd gnd cell_6t
Xbit_r23_c35 bl[35] br[35] wl[23] vdd gnd cell_6t
Xbit_r24_c35 bl[35] br[35] wl[24] vdd gnd cell_6t
Xbit_r25_c35 bl[35] br[35] wl[25] vdd gnd cell_6t
Xbit_r26_c35 bl[35] br[35] wl[26] vdd gnd cell_6t
Xbit_r27_c35 bl[35] br[35] wl[27] vdd gnd cell_6t
Xbit_r28_c35 bl[35] br[35] wl[28] vdd gnd cell_6t
Xbit_r29_c35 bl[35] br[35] wl[29] vdd gnd cell_6t
Xbit_r30_c35 bl[35] br[35] wl[30] vdd gnd cell_6t
Xbit_r31_c35 bl[35] br[35] wl[31] vdd gnd cell_6t
Xbit_r32_c35 bl[35] br[35] wl[32] vdd gnd cell_6t
Xbit_r33_c35 bl[35] br[35] wl[33] vdd gnd cell_6t
Xbit_r34_c35 bl[35] br[35] wl[34] vdd gnd cell_6t
Xbit_r35_c35 bl[35] br[35] wl[35] vdd gnd cell_6t
Xbit_r36_c35 bl[35] br[35] wl[36] vdd gnd cell_6t
Xbit_r37_c35 bl[35] br[35] wl[37] vdd gnd cell_6t
Xbit_r38_c35 bl[35] br[35] wl[38] vdd gnd cell_6t
Xbit_r39_c35 bl[35] br[35] wl[39] vdd gnd cell_6t
Xbit_r40_c35 bl[35] br[35] wl[40] vdd gnd cell_6t
Xbit_r41_c35 bl[35] br[35] wl[41] vdd gnd cell_6t
Xbit_r42_c35 bl[35] br[35] wl[42] vdd gnd cell_6t
Xbit_r43_c35 bl[35] br[35] wl[43] vdd gnd cell_6t
Xbit_r44_c35 bl[35] br[35] wl[44] vdd gnd cell_6t
Xbit_r45_c35 bl[35] br[35] wl[45] vdd gnd cell_6t
Xbit_r46_c35 bl[35] br[35] wl[46] vdd gnd cell_6t
Xbit_r47_c35 bl[35] br[35] wl[47] vdd gnd cell_6t
Xbit_r48_c35 bl[35] br[35] wl[48] vdd gnd cell_6t
Xbit_r49_c35 bl[35] br[35] wl[49] vdd gnd cell_6t
Xbit_r50_c35 bl[35] br[35] wl[50] vdd gnd cell_6t
Xbit_r51_c35 bl[35] br[35] wl[51] vdd gnd cell_6t
Xbit_r52_c35 bl[35] br[35] wl[52] vdd gnd cell_6t
Xbit_r53_c35 bl[35] br[35] wl[53] vdd gnd cell_6t
Xbit_r54_c35 bl[35] br[35] wl[54] vdd gnd cell_6t
Xbit_r55_c35 bl[35] br[35] wl[55] vdd gnd cell_6t
Xbit_r56_c35 bl[35] br[35] wl[56] vdd gnd cell_6t
Xbit_r57_c35 bl[35] br[35] wl[57] vdd gnd cell_6t
Xbit_r58_c35 bl[35] br[35] wl[58] vdd gnd cell_6t
Xbit_r59_c35 bl[35] br[35] wl[59] vdd gnd cell_6t
Xbit_r60_c35 bl[35] br[35] wl[60] vdd gnd cell_6t
Xbit_r61_c35 bl[35] br[35] wl[61] vdd gnd cell_6t
Xbit_r62_c35 bl[35] br[35] wl[62] vdd gnd cell_6t
Xbit_r63_c35 bl[35] br[35] wl[63] vdd gnd cell_6t
Xbit_r64_c35 bl[35] br[35] wl[64] vdd gnd cell_6t
Xbit_r65_c35 bl[35] br[35] wl[65] vdd gnd cell_6t
Xbit_r66_c35 bl[35] br[35] wl[66] vdd gnd cell_6t
Xbit_r67_c35 bl[35] br[35] wl[67] vdd gnd cell_6t
Xbit_r68_c35 bl[35] br[35] wl[68] vdd gnd cell_6t
Xbit_r69_c35 bl[35] br[35] wl[69] vdd gnd cell_6t
Xbit_r70_c35 bl[35] br[35] wl[70] vdd gnd cell_6t
Xbit_r71_c35 bl[35] br[35] wl[71] vdd gnd cell_6t
Xbit_r72_c35 bl[35] br[35] wl[72] vdd gnd cell_6t
Xbit_r73_c35 bl[35] br[35] wl[73] vdd gnd cell_6t
Xbit_r74_c35 bl[35] br[35] wl[74] vdd gnd cell_6t
Xbit_r75_c35 bl[35] br[35] wl[75] vdd gnd cell_6t
Xbit_r76_c35 bl[35] br[35] wl[76] vdd gnd cell_6t
Xbit_r77_c35 bl[35] br[35] wl[77] vdd gnd cell_6t
Xbit_r78_c35 bl[35] br[35] wl[78] vdd gnd cell_6t
Xbit_r79_c35 bl[35] br[35] wl[79] vdd gnd cell_6t
Xbit_r80_c35 bl[35] br[35] wl[80] vdd gnd cell_6t
Xbit_r81_c35 bl[35] br[35] wl[81] vdd gnd cell_6t
Xbit_r82_c35 bl[35] br[35] wl[82] vdd gnd cell_6t
Xbit_r83_c35 bl[35] br[35] wl[83] vdd gnd cell_6t
Xbit_r84_c35 bl[35] br[35] wl[84] vdd gnd cell_6t
Xbit_r85_c35 bl[35] br[35] wl[85] vdd gnd cell_6t
Xbit_r86_c35 bl[35] br[35] wl[86] vdd gnd cell_6t
Xbit_r87_c35 bl[35] br[35] wl[87] vdd gnd cell_6t
Xbit_r88_c35 bl[35] br[35] wl[88] vdd gnd cell_6t
Xbit_r89_c35 bl[35] br[35] wl[89] vdd gnd cell_6t
Xbit_r90_c35 bl[35] br[35] wl[90] vdd gnd cell_6t
Xbit_r91_c35 bl[35] br[35] wl[91] vdd gnd cell_6t
Xbit_r92_c35 bl[35] br[35] wl[92] vdd gnd cell_6t
Xbit_r93_c35 bl[35] br[35] wl[93] vdd gnd cell_6t
Xbit_r94_c35 bl[35] br[35] wl[94] vdd gnd cell_6t
Xbit_r95_c35 bl[35] br[35] wl[95] vdd gnd cell_6t
Xbit_r96_c35 bl[35] br[35] wl[96] vdd gnd cell_6t
Xbit_r97_c35 bl[35] br[35] wl[97] vdd gnd cell_6t
Xbit_r98_c35 bl[35] br[35] wl[98] vdd gnd cell_6t
Xbit_r99_c35 bl[35] br[35] wl[99] vdd gnd cell_6t
Xbit_r100_c35 bl[35] br[35] wl[100] vdd gnd cell_6t
Xbit_r101_c35 bl[35] br[35] wl[101] vdd gnd cell_6t
Xbit_r102_c35 bl[35] br[35] wl[102] vdd gnd cell_6t
Xbit_r103_c35 bl[35] br[35] wl[103] vdd gnd cell_6t
Xbit_r104_c35 bl[35] br[35] wl[104] vdd gnd cell_6t
Xbit_r105_c35 bl[35] br[35] wl[105] vdd gnd cell_6t
Xbit_r106_c35 bl[35] br[35] wl[106] vdd gnd cell_6t
Xbit_r107_c35 bl[35] br[35] wl[107] vdd gnd cell_6t
Xbit_r108_c35 bl[35] br[35] wl[108] vdd gnd cell_6t
Xbit_r109_c35 bl[35] br[35] wl[109] vdd gnd cell_6t
Xbit_r110_c35 bl[35] br[35] wl[110] vdd gnd cell_6t
Xbit_r111_c35 bl[35] br[35] wl[111] vdd gnd cell_6t
Xbit_r112_c35 bl[35] br[35] wl[112] vdd gnd cell_6t
Xbit_r113_c35 bl[35] br[35] wl[113] vdd gnd cell_6t
Xbit_r114_c35 bl[35] br[35] wl[114] vdd gnd cell_6t
Xbit_r115_c35 bl[35] br[35] wl[115] vdd gnd cell_6t
Xbit_r116_c35 bl[35] br[35] wl[116] vdd gnd cell_6t
Xbit_r117_c35 bl[35] br[35] wl[117] vdd gnd cell_6t
Xbit_r118_c35 bl[35] br[35] wl[118] vdd gnd cell_6t
Xbit_r119_c35 bl[35] br[35] wl[119] vdd gnd cell_6t
Xbit_r120_c35 bl[35] br[35] wl[120] vdd gnd cell_6t
Xbit_r121_c35 bl[35] br[35] wl[121] vdd gnd cell_6t
Xbit_r122_c35 bl[35] br[35] wl[122] vdd gnd cell_6t
Xbit_r123_c35 bl[35] br[35] wl[123] vdd gnd cell_6t
Xbit_r124_c35 bl[35] br[35] wl[124] vdd gnd cell_6t
Xbit_r125_c35 bl[35] br[35] wl[125] vdd gnd cell_6t
Xbit_r126_c35 bl[35] br[35] wl[126] vdd gnd cell_6t
Xbit_r127_c35 bl[35] br[35] wl[127] vdd gnd cell_6t
Xbit_r128_c35 bl[35] br[35] wl[128] vdd gnd cell_6t
Xbit_r129_c35 bl[35] br[35] wl[129] vdd gnd cell_6t
Xbit_r130_c35 bl[35] br[35] wl[130] vdd gnd cell_6t
Xbit_r131_c35 bl[35] br[35] wl[131] vdd gnd cell_6t
Xbit_r132_c35 bl[35] br[35] wl[132] vdd gnd cell_6t
Xbit_r133_c35 bl[35] br[35] wl[133] vdd gnd cell_6t
Xbit_r134_c35 bl[35] br[35] wl[134] vdd gnd cell_6t
Xbit_r135_c35 bl[35] br[35] wl[135] vdd gnd cell_6t
Xbit_r136_c35 bl[35] br[35] wl[136] vdd gnd cell_6t
Xbit_r137_c35 bl[35] br[35] wl[137] vdd gnd cell_6t
Xbit_r138_c35 bl[35] br[35] wl[138] vdd gnd cell_6t
Xbit_r139_c35 bl[35] br[35] wl[139] vdd gnd cell_6t
Xbit_r140_c35 bl[35] br[35] wl[140] vdd gnd cell_6t
Xbit_r141_c35 bl[35] br[35] wl[141] vdd gnd cell_6t
Xbit_r142_c35 bl[35] br[35] wl[142] vdd gnd cell_6t
Xbit_r143_c35 bl[35] br[35] wl[143] vdd gnd cell_6t
Xbit_r144_c35 bl[35] br[35] wl[144] vdd gnd cell_6t
Xbit_r145_c35 bl[35] br[35] wl[145] vdd gnd cell_6t
Xbit_r146_c35 bl[35] br[35] wl[146] vdd gnd cell_6t
Xbit_r147_c35 bl[35] br[35] wl[147] vdd gnd cell_6t
Xbit_r148_c35 bl[35] br[35] wl[148] vdd gnd cell_6t
Xbit_r149_c35 bl[35] br[35] wl[149] vdd gnd cell_6t
Xbit_r150_c35 bl[35] br[35] wl[150] vdd gnd cell_6t
Xbit_r151_c35 bl[35] br[35] wl[151] vdd gnd cell_6t
Xbit_r152_c35 bl[35] br[35] wl[152] vdd gnd cell_6t
Xbit_r153_c35 bl[35] br[35] wl[153] vdd gnd cell_6t
Xbit_r154_c35 bl[35] br[35] wl[154] vdd gnd cell_6t
Xbit_r155_c35 bl[35] br[35] wl[155] vdd gnd cell_6t
Xbit_r156_c35 bl[35] br[35] wl[156] vdd gnd cell_6t
Xbit_r157_c35 bl[35] br[35] wl[157] vdd gnd cell_6t
Xbit_r158_c35 bl[35] br[35] wl[158] vdd gnd cell_6t
Xbit_r159_c35 bl[35] br[35] wl[159] vdd gnd cell_6t
Xbit_r160_c35 bl[35] br[35] wl[160] vdd gnd cell_6t
Xbit_r161_c35 bl[35] br[35] wl[161] vdd gnd cell_6t
Xbit_r162_c35 bl[35] br[35] wl[162] vdd gnd cell_6t
Xbit_r163_c35 bl[35] br[35] wl[163] vdd gnd cell_6t
Xbit_r164_c35 bl[35] br[35] wl[164] vdd gnd cell_6t
Xbit_r165_c35 bl[35] br[35] wl[165] vdd gnd cell_6t
Xbit_r166_c35 bl[35] br[35] wl[166] vdd gnd cell_6t
Xbit_r167_c35 bl[35] br[35] wl[167] vdd gnd cell_6t
Xbit_r168_c35 bl[35] br[35] wl[168] vdd gnd cell_6t
Xbit_r169_c35 bl[35] br[35] wl[169] vdd gnd cell_6t
Xbit_r170_c35 bl[35] br[35] wl[170] vdd gnd cell_6t
Xbit_r171_c35 bl[35] br[35] wl[171] vdd gnd cell_6t
Xbit_r172_c35 bl[35] br[35] wl[172] vdd gnd cell_6t
Xbit_r173_c35 bl[35] br[35] wl[173] vdd gnd cell_6t
Xbit_r174_c35 bl[35] br[35] wl[174] vdd gnd cell_6t
Xbit_r175_c35 bl[35] br[35] wl[175] vdd gnd cell_6t
Xbit_r176_c35 bl[35] br[35] wl[176] vdd gnd cell_6t
Xbit_r177_c35 bl[35] br[35] wl[177] vdd gnd cell_6t
Xbit_r178_c35 bl[35] br[35] wl[178] vdd gnd cell_6t
Xbit_r179_c35 bl[35] br[35] wl[179] vdd gnd cell_6t
Xbit_r180_c35 bl[35] br[35] wl[180] vdd gnd cell_6t
Xbit_r181_c35 bl[35] br[35] wl[181] vdd gnd cell_6t
Xbit_r182_c35 bl[35] br[35] wl[182] vdd gnd cell_6t
Xbit_r183_c35 bl[35] br[35] wl[183] vdd gnd cell_6t
Xbit_r184_c35 bl[35] br[35] wl[184] vdd gnd cell_6t
Xbit_r185_c35 bl[35] br[35] wl[185] vdd gnd cell_6t
Xbit_r186_c35 bl[35] br[35] wl[186] vdd gnd cell_6t
Xbit_r187_c35 bl[35] br[35] wl[187] vdd gnd cell_6t
Xbit_r188_c35 bl[35] br[35] wl[188] vdd gnd cell_6t
Xbit_r189_c35 bl[35] br[35] wl[189] vdd gnd cell_6t
Xbit_r190_c35 bl[35] br[35] wl[190] vdd gnd cell_6t
Xbit_r191_c35 bl[35] br[35] wl[191] vdd gnd cell_6t
Xbit_r192_c35 bl[35] br[35] wl[192] vdd gnd cell_6t
Xbit_r193_c35 bl[35] br[35] wl[193] vdd gnd cell_6t
Xbit_r194_c35 bl[35] br[35] wl[194] vdd gnd cell_6t
Xbit_r195_c35 bl[35] br[35] wl[195] vdd gnd cell_6t
Xbit_r196_c35 bl[35] br[35] wl[196] vdd gnd cell_6t
Xbit_r197_c35 bl[35] br[35] wl[197] vdd gnd cell_6t
Xbit_r198_c35 bl[35] br[35] wl[198] vdd gnd cell_6t
Xbit_r199_c35 bl[35] br[35] wl[199] vdd gnd cell_6t
Xbit_r200_c35 bl[35] br[35] wl[200] vdd gnd cell_6t
Xbit_r201_c35 bl[35] br[35] wl[201] vdd gnd cell_6t
Xbit_r202_c35 bl[35] br[35] wl[202] vdd gnd cell_6t
Xbit_r203_c35 bl[35] br[35] wl[203] vdd gnd cell_6t
Xbit_r204_c35 bl[35] br[35] wl[204] vdd gnd cell_6t
Xbit_r205_c35 bl[35] br[35] wl[205] vdd gnd cell_6t
Xbit_r206_c35 bl[35] br[35] wl[206] vdd gnd cell_6t
Xbit_r207_c35 bl[35] br[35] wl[207] vdd gnd cell_6t
Xbit_r208_c35 bl[35] br[35] wl[208] vdd gnd cell_6t
Xbit_r209_c35 bl[35] br[35] wl[209] vdd gnd cell_6t
Xbit_r210_c35 bl[35] br[35] wl[210] vdd gnd cell_6t
Xbit_r211_c35 bl[35] br[35] wl[211] vdd gnd cell_6t
Xbit_r212_c35 bl[35] br[35] wl[212] vdd gnd cell_6t
Xbit_r213_c35 bl[35] br[35] wl[213] vdd gnd cell_6t
Xbit_r214_c35 bl[35] br[35] wl[214] vdd gnd cell_6t
Xbit_r215_c35 bl[35] br[35] wl[215] vdd gnd cell_6t
Xbit_r216_c35 bl[35] br[35] wl[216] vdd gnd cell_6t
Xbit_r217_c35 bl[35] br[35] wl[217] vdd gnd cell_6t
Xbit_r218_c35 bl[35] br[35] wl[218] vdd gnd cell_6t
Xbit_r219_c35 bl[35] br[35] wl[219] vdd gnd cell_6t
Xbit_r220_c35 bl[35] br[35] wl[220] vdd gnd cell_6t
Xbit_r221_c35 bl[35] br[35] wl[221] vdd gnd cell_6t
Xbit_r222_c35 bl[35] br[35] wl[222] vdd gnd cell_6t
Xbit_r223_c35 bl[35] br[35] wl[223] vdd gnd cell_6t
Xbit_r224_c35 bl[35] br[35] wl[224] vdd gnd cell_6t
Xbit_r225_c35 bl[35] br[35] wl[225] vdd gnd cell_6t
Xbit_r226_c35 bl[35] br[35] wl[226] vdd gnd cell_6t
Xbit_r227_c35 bl[35] br[35] wl[227] vdd gnd cell_6t
Xbit_r228_c35 bl[35] br[35] wl[228] vdd gnd cell_6t
Xbit_r229_c35 bl[35] br[35] wl[229] vdd gnd cell_6t
Xbit_r230_c35 bl[35] br[35] wl[230] vdd gnd cell_6t
Xbit_r231_c35 bl[35] br[35] wl[231] vdd gnd cell_6t
Xbit_r232_c35 bl[35] br[35] wl[232] vdd gnd cell_6t
Xbit_r233_c35 bl[35] br[35] wl[233] vdd gnd cell_6t
Xbit_r234_c35 bl[35] br[35] wl[234] vdd gnd cell_6t
Xbit_r235_c35 bl[35] br[35] wl[235] vdd gnd cell_6t
Xbit_r236_c35 bl[35] br[35] wl[236] vdd gnd cell_6t
Xbit_r237_c35 bl[35] br[35] wl[237] vdd gnd cell_6t
Xbit_r238_c35 bl[35] br[35] wl[238] vdd gnd cell_6t
Xbit_r239_c35 bl[35] br[35] wl[239] vdd gnd cell_6t
Xbit_r240_c35 bl[35] br[35] wl[240] vdd gnd cell_6t
Xbit_r241_c35 bl[35] br[35] wl[241] vdd gnd cell_6t
Xbit_r242_c35 bl[35] br[35] wl[242] vdd gnd cell_6t
Xbit_r243_c35 bl[35] br[35] wl[243] vdd gnd cell_6t
Xbit_r244_c35 bl[35] br[35] wl[244] vdd gnd cell_6t
Xbit_r245_c35 bl[35] br[35] wl[245] vdd gnd cell_6t
Xbit_r246_c35 bl[35] br[35] wl[246] vdd gnd cell_6t
Xbit_r247_c35 bl[35] br[35] wl[247] vdd gnd cell_6t
Xbit_r248_c35 bl[35] br[35] wl[248] vdd gnd cell_6t
Xbit_r249_c35 bl[35] br[35] wl[249] vdd gnd cell_6t
Xbit_r250_c35 bl[35] br[35] wl[250] vdd gnd cell_6t
Xbit_r251_c35 bl[35] br[35] wl[251] vdd gnd cell_6t
Xbit_r252_c35 bl[35] br[35] wl[252] vdd gnd cell_6t
Xbit_r253_c35 bl[35] br[35] wl[253] vdd gnd cell_6t
Xbit_r254_c35 bl[35] br[35] wl[254] vdd gnd cell_6t
Xbit_r255_c35 bl[35] br[35] wl[255] vdd gnd cell_6t
Xbit_r0_c36 bl[36] br[36] wl[0] vdd gnd cell_6t
Xbit_r1_c36 bl[36] br[36] wl[1] vdd gnd cell_6t
Xbit_r2_c36 bl[36] br[36] wl[2] vdd gnd cell_6t
Xbit_r3_c36 bl[36] br[36] wl[3] vdd gnd cell_6t
Xbit_r4_c36 bl[36] br[36] wl[4] vdd gnd cell_6t
Xbit_r5_c36 bl[36] br[36] wl[5] vdd gnd cell_6t
Xbit_r6_c36 bl[36] br[36] wl[6] vdd gnd cell_6t
Xbit_r7_c36 bl[36] br[36] wl[7] vdd gnd cell_6t
Xbit_r8_c36 bl[36] br[36] wl[8] vdd gnd cell_6t
Xbit_r9_c36 bl[36] br[36] wl[9] vdd gnd cell_6t
Xbit_r10_c36 bl[36] br[36] wl[10] vdd gnd cell_6t
Xbit_r11_c36 bl[36] br[36] wl[11] vdd gnd cell_6t
Xbit_r12_c36 bl[36] br[36] wl[12] vdd gnd cell_6t
Xbit_r13_c36 bl[36] br[36] wl[13] vdd gnd cell_6t
Xbit_r14_c36 bl[36] br[36] wl[14] vdd gnd cell_6t
Xbit_r15_c36 bl[36] br[36] wl[15] vdd gnd cell_6t
Xbit_r16_c36 bl[36] br[36] wl[16] vdd gnd cell_6t
Xbit_r17_c36 bl[36] br[36] wl[17] vdd gnd cell_6t
Xbit_r18_c36 bl[36] br[36] wl[18] vdd gnd cell_6t
Xbit_r19_c36 bl[36] br[36] wl[19] vdd gnd cell_6t
Xbit_r20_c36 bl[36] br[36] wl[20] vdd gnd cell_6t
Xbit_r21_c36 bl[36] br[36] wl[21] vdd gnd cell_6t
Xbit_r22_c36 bl[36] br[36] wl[22] vdd gnd cell_6t
Xbit_r23_c36 bl[36] br[36] wl[23] vdd gnd cell_6t
Xbit_r24_c36 bl[36] br[36] wl[24] vdd gnd cell_6t
Xbit_r25_c36 bl[36] br[36] wl[25] vdd gnd cell_6t
Xbit_r26_c36 bl[36] br[36] wl[26] vdd gnd cell_6t
Xbit_r27_c36 bl[36] br[36] wl[27] vdd gnd cell_6t
Xbit_r28_c36 bl[36] br[36] wl[28] vdd gnd cell_6t
Xbit_r29_c36 bl[36] br[36] wl[29] vdd gnd cell_6t
Xbit_r30_c36 bl[36] br[36] wl[30] vdd gnd cell_6t
Xbit_r31_c36 bl[36] br[36] wl[31] vdd gnd cell_6t
Xbit_r32_c36 bl[36] br[36] wl[32] vdd gnd cell_6t
Xbit_r33_c36 bl[36] br[36] wl[33] vdd gnd cell_6t
Xbit_r34_c36 bl[36] br[36] wl[34] vdd gnd cell_6t
Xbit_r35_c36 bl[36] br[36] wl[35] vdd gnd cell_6t
Xbit_r36_c36 bl[36] br[36] wl[36] vdd gnd cell_6t
Xbit_r37_c36 bl[36] br[36] wl[37] vdd gnd cell_6t
Xbit_r38_c36 bl[36] br[36] wl[38] vdd gnd cell_6t
Xbit_r39_c36 bl[36] br[36] wl[39] vdd gnd cell_6t
Xbit_r40_c36 bl[36] br[36] wl[40] vdd gnd cell_6t
Xbit_r41_c36 bl[36] br[36] wl[41] vdd gnd cell_6t
Xbit_r42_c36 bl[36] br[36] wl[42] vdd gnd cell_6t
Xbit_r43_c36 bl[36] br[36] wl[43] vdd gnd cell_6t
Xbit_r44_c36 bl[36] br[36] wl[44] vdd gnd cell_6t
Xbit_r45_c36 bl[36] br[36] wl[45] vdd gnd cell_6t
Xbit_r46_c36 bl[36] br[36] wl[46] vdd gnd cell_6t
Xbit_r47_c36 bl[36] br[36] wl[47] vdd gnd cell_6t
Xbit_r48_c36 bl[36] br[36] wl[48] vdd gnd cell_6t
Xbit_r49_c36 bl[36] br[36] wl[49] vdd gnd cell_6t
Xbit_r50_c36 bl[36] br[36] wl[50] vdd gnd cell_6t
Xbit_r51_c36 bl[36] br[36] wl[51] vdd gnd cell_6t
Xbit_r52_c36 bl[36] br[36] wl[52] vdd gnd cell_6t
Xbit_r53_c36 bl[36] br[36] wl[53] vdd gnd cell_6t
Xbit_r54_c36 bl[36] br[36] wl[54] vdd gnd cell_6t
Xbit_r55_c36 bl[36] br[36] wl[55] vdd gnd cell_6t
Xbit_r56_c36 bl[36] br[36] wl[56] vdd gnd cell_6t
Xbit_r57_c36 bl[36] br[36] wl[57] vdd gnd cell_6t
Xbit_r58_c36 bl[36] br[36] wl[58] vdd gnd cell_6t
Xbit_r59_c36 bl[36] br[36] wl[59] vdd gnd cell_6t
Xbit_r60_c36 bl[36] br[36] wl[60] vdd gnd cell_6t
Xbit_r61_c36 bl[36] br[36] wl[61] vdd gnd cell_6t
Xbit_r62_c36 bl[36] br[36] wl[62] vdd gnd cell_6t
Xbit_r63_c36 bl[36] br[36] wl[63] vdd gnd cell_6t
Xbit_r64_c36 bl[36] br[36] wl[64] vdd gnd cell_6t
Xbit_r65_c36 bl[36] br[36] wl[65] vdd gnd cell_6t
Xbit_r66_c36 bl[36] br[36] wl[66] vdd gnd cell_6t
Xbit_r67_c36 bl[36] br[36] wl[67] vdd gnd cell_6t
Xbit_r68_c36 bl[36] br[36] wl[68] vdd gnd cell_6t
Xbit_r69_c36 bl[36] br[36] wl[69] vdd gnd cell_6t
Xbit_r70_c36 bl[36] br[36] wl[70] vdd gnd cell_6t
Xbit_r71_c36 bl[36] br[36] wl[71] vdd gnd cell_6t
Xbit_r72_c36 bl[36] br[36] wl[72] vdd gnd cell_6t
Xbit_r73_c36 bl[36] br[36] wl[73] vdd gnd cell_6t
Xbit_r74_c36 bl[36] br[36] wl[74] vdd gnd cell_6t
Xbit_r75_c36 bl[36] br[36] wl[75] vdd gnd cell_6t
Xbit_r76_c36 bl[36] br[36] wl[76] vdd gnd cell_6t
Xbit_r77_c36 bl[36] br[36] wl[77] vdd gnd cell_6t
Xbit_r78_c36 bl[36] br[36] wl[78] vdd gnd cell_6t
Xbit_r79_c36 bl[36] br[36] wl[79] vdd gnd cell_6t
Xbit_r80_c36 bl[36] br[36] wl[80] vdd gnd cell_6t
Xbit_r81_c36 bl[36] br[36] wl[81] vdd gnd cell_6t
Xbit_r82_c36 bl[36] br[36] wl[82] vdd gnd cell_6t
Xbit_r83_c36 bl[36] br[36] wl[83] vdd gnd cell_6t
Xbit_r84_c36 bl[36] br[36] wl[84] vdd gnd cell_6t
Xbit_r85_c36 bl[36] br[36] wl[85] vdd gnd cell_6t
Xbit_r86_c36 bl[36] br[36] wl[86] vdd gnd cell_6t
Xbit_r87_c36 bl[36] br[36] wl[87] vdd gnd cell_6t
Xbit_r88_c36 bl[36] br[36] wl[88] vdd gnd cell_6t
Xbit_r89_c36 bl[36] br[36] wl[89] vdd gnd cell_6t
Xbit_r90_c36 bl[36] br[36] wl[90] vdd gnd cell_6t
Xbit_r91_c36 bl[36] br[36] wl[91] vdd gnd cell_6t
Xbit_r92_c36 bl[36] br[36] wl[92] vdd gnd cell_6t
Xbit_r93_c36 bl[36] br[36] wl[93] vdd gnd cell_6t
Xbit_r94_c36 bl[36] br[36] wl[94] vdd gnd cell_6t
Xbit_r95_c36 bl[36] br[36] wl[95] vdd gnd cell_6t
Xbit_r96_c36 bl[36] br[36] wl[96] vdd gnd cell_6t
Xbit_r97_c36 bl[36] br[36] wl[97] vdd gnd cell_6t
Xbit_r98_c36 bl[36] br[36] wl[98] vdd gnd cell_6t
Xbit_r99_c36 bl[36] br[36] wl[99] vdd gnd cell_6t
Xbit_r100_c36 bl[36] br[36] wl[100] vdd gnd cell_6t
Xbit_r101_c36 bl[36] br[36] wl[101] vdd gnd cell_6t
Xbit_r102_c36 bl[36] br[36] wl[102] vdd gnd cell_6t
Xbit_r103_c36 bl[36] br[36] wl[103] vdd gnd cell_6t
Xbit_r104_c36 bl[36] br[36] wl[104] vdd gnd cell_6t
Xbit_r105_c36 bl[36] br[36] wl[105] vdd gnd cell_6t
Xbit_r106_c36 bl[36] br[36] wl[106] vdd gnd cell_6t
Xbit_r107_c36 bl[36] br[36] wl[107] vdd gnd cell_6t
Xbit_r108_c36 bl[36] br[36] wl[108] vdd gnd cell_6t
Xbit_r109_c36 bl[36] br[36] wl[109] vdd gnd cell_6t
Xbit_r110_c36 bl[36] br[36] wl[110] vdd gnd cell_6t
Xbit_r111_c36 bl[36] br[36] wl[111] vdd gnd cell_6t
Xbit_r112_c36 bl[36] br[36] wl[112] vdd gnd cell_6t
Xbit_r113_c36 bl[36] br[36] wl[113] vdd gnd cell_6t
Xbit_r114_c36 bl[36] br[36] wl[114] vdd gnd cell_6t
Xbit_r115_c36 bl[36] br[36] wl[115] vdd gnd cell_6t
Xbit_r116_c36 bl[36] br[36] wl[116] vdd gnd cell_6t
Xbit_r117_c36 bl[36] br[36] wl[117] vdd gnd cell_6t
Xbit_r118_c36 bl[36] br[36] wl[118] vdd gnd cell_6t
Xbit_r119_c36 bl[36] br[36] wl[119] vdd gnd cell_6t
Xbit_r120_c36 bl[36] br[36] wl[120] vdd gnd cell_6t
Xbit_r121_c36 bl[36] br[36] wl[121] vdd gnd cell_6t
Xbit_r122_c36 bl[36] br[36] wl[122] vdd gnd cell_6t
Xbit_r123_c36 bl[36] br[36] wl[123] vdd gnd cell_6t
Xbit_r124_c36 bl[36] br[36] wl[124] vdd gnd cell_6t
Xbit_r125_c36 bl[36] br[36] wl[125] vdd gnd cell_6t
Xbit_r126_c36 bl[36] br[36] wl[126] vdd gnd cell_6t
Xbit_r127_c36 bl[36] br[36] wl[127] vdd gnd cell_6t
Xbit_r128_c36 bl[36] br[36] wl[128] vdd gnd cell_6t
Xbit_r129_c36 bl[36] br[36] wl[129] vdd gnd cell_6t
Xbit_r130_c36 bl[36] br[36] wl[130] vdd gnd cell_6t
Xbit_r131_c36 bl[36] br[36] wl[131] vdd gnd cell_6t
Xbit_r132_c36 bl[36] br[36] wl[132] vdd gnd cell_6t
Xbit_r133_c36 bl[36] br[36] wl[133] vdd gnd cell_6t
Xbit_r134_c36 bl[36] br[36] wl[134] vdd gnd cell_6t
Xbit_r135_c36 bl[36] br[36] wl[135] vdd gnd cell_6t
Xbit_r136_c36 bl[36] br[36] wl[136] vdd gnd cell_6t
Xbit_r137_c36 bl[36] br[36] wl[137] vdd gnd cell_6t
Xbit_r138_c36 bl[36] br[36] wl[138] vdd gnd cell_6t
Xbit_r139_c36 bl[36] br[36] wl[139] vdd gnd cell_6t
Xbit_r140_c36 bl[36] br[36] wl[140] vdd gnd cell_6t
Xbit_r141_c36 bl[36] br[36] wl[141] vdd gnd cell_6t
Xbit_r142_c36 bl[36] br[36] wl[142] vdd gnd cell_6t
Xbit_r143_c36 bl[36] br[36] wl[143] vdd gnd cell_6t
Xbit_r144_c36 bl[36] br[36] wl[144] vdd gnd cell_6t
Xbit_r145_c36 bl[36] br[36] wl[145] vdd gnd cell_6t
Xbit_r146_c36 bl[36] br[36] wl[146] vdd gnd cell_6t
Xbit_r147_c36 bl[36] br[36] wl[147] vdd gnd cell_6t
Xbit_r148_c36 bl[36] br[36] wl[148] vdd gnd cell_6t
Xbit_r149_c36 bl[36] br[36] wl[149] vdd gnd cell_6t
Xbit_r150_c36 bl[36] br[36] wl[150] vdd gnd cell_6t
Xbit_r151_c36 bl[36] br[36] wl[151] vdd gnd cell_6t
Xbit_r152_c36 bl[36] br[36] wl[152] vdd gnd cell_6t
Xbit_r153_c36 bl[36] br[36] wl[153] vdd gnd cell_6t
Xbit_r154_c36 bl[36] br[36] wl[154] vdd gnd cell_6t
Xbit_r155_c36 bl[36] br[36] wl[155] vdd gnd cell_6t
Xbit_r156_c36 bl[36] br[36] wl[156] vdd gnd cell_6t
Xbit_r157_c36 bl[36] br[36] wl[157] vdd gnd cell_6t
Xbit_r158_c36 bl[36] br[36] wl[158] vdd gnd cell_6t
Xbit_r159_c36 bl[36] br[36] wl[159] vdd gnd cell_6t
Xbit_r160_c36 bl[36] br[36] wl[160] vdd gnd cell_6t
Xbit_r161_c36 bl[36] br[36] wl[161] vdd gnd cell_6t
Xbit_r162_c36 bl[36] br[36] wl[162] vdd gnd cell_6t
Xbit_r163_c36 bl[36] br[36] wl[163] vdd gnd cell_6t
Xbit_r164_c36 bl[36] br[36] wl[164] vdd gnd cell_6t
Xbit_r165_c36 bl[36] br[36] wl[165] vdd gnd cell_6t
Xbit_r166_c36 bl[36] br[36] wl[166] vdd gnd cell_6t
Xbit_r167_c36 bl[36] br[36] wl[167] vdd gnd cell_6t
Xbit_r168_c36 bl[36] br[36] wl[168] vdd gnd cell_6t
Xbit_r169_c36 bl[36] br[36] wl[169] vdd gnd cell_6t
Xbit_r170_c36 bl[36] br[36] wl[170] vdd gnd cell_6t
Xbit_r171_c36 bl[36] br[36] wl[171] vdd gnd cell_6t
Xbit_r172_c36 bl[36] br[36] wl[172] vdd gnd cell_6t
Xbit_r173_c36 bl[36] br[36] wl[173] vdd gnd cell_6t
Xbit_r174_c36 bl[36] br[36] wl[174] vdd gnd cell_6t
Xbit_r175_c36 bl[36] br[36] wl[175] vdd gnd cell_6t
Xbit_r176_c36 bl[36] br[36] wl[176] vdd gnd cell_6t
Xbit_r177_c36 bl[36] br[36] wl[177] vdd gnd cell_6t
Xbit_r178_c36 bl[36] br[36] wl[178] vdd gnd cell_6t
Xbit_r179_c36 bl[36] br[36] wl[179] vdd gnd cell_6t
Xbit_r180_c36 bl[36] br[36] wl[180] vdd gnd cell_6t
Xbit_r181_c36 bl[36] br[36] wl[181] vdd gnd cell_6t
Xbit_r182_c36 bl[36] br[36] wl[182] vdd gnd cell_6t
Xbit_r183_c36 bl[36] br[36] wl[183] vdd gnd cell_6t
Xbit_r184_c36 bl[36] br[36] wl[184] vdd gnd cell_6t
Xbit_r185_c36 bl[36] br[36] wl[185] vdd gnd cell_6t
Xbit_r186_c36 bl[36] br[36] wl[186] vdd gnd cell_6t
Xbit_r187_c36 bl[36] br[36] wl[187] vdd gnd cell_6t
Xbit_r188_c36 bl[36] br[36] wl[188] vdd gnd cell_6t
Xbit_r189_c36 bl[36] br[36] wl[189] vdd gnd cell_6t
Xbit_r190_c36 bl[36] br[36] wl[190] vdd gnd cell_6t
Xbit_r191_c36 bl[36] br[36] wl[191] vdd gnd cell_6t
Xbit_r192_c36 bl[36] br[36] wl[192] vdd gnd cell_6t
Xbit_r193_c36 bl[36] br[36] wl[193] vdd gnd cell_6t
Xbit_r194_c36 bl[36] br[36] wl[194] vdd gnd cell_6t
Xbit_r195_c36 bl[36] br[36] wl[195] vdd gnd cell_6t
Xbit_r196_c36 bl[36] br[36] wl[196] vdd gnd cell_6t
Xbit_r197_c36 bl[36] br[36] wl[197] vdd gnd cell_6t
Xbit_r198_c36 bl[36] br[36] wl[198] vdd gnd cell_6t
Xbit_r199_c36 bl[36] br[36] wl[199] vdd gnd cell_6t
Xbit_r200_c36 bl[36] br[36] wl[200] vdd gnd cell_6t
Xbit_r201_c36 bl[36] br[36] wl[201] vdd gnd cell_6t
Xbit_r202_c36 bl[36] br[36] wl[202] vdd gnd cell_6t
Xbit_r203_c36 bl[36] br[36] wl[203] vdd gnd cell_6t
Xbit_r204_c36 bl[36] br[36] wl[204] vdd gnd cell_6t
Xbit_r205_c36 bl[36] br[36] wl[205] vdd gnd cell_6t
Xbit_r206_c36 bl[36] br[36] wl[206] vdd gnd cell_6t
Xbit_r207_c36 bl[36] br[36] wl[207] vdd gnd cell_6t
Xbit_r208_c36 bl[36] br[36] wl[208] vdd gnd cell_6t
Xbit_r209_c36 bl[36] br[36] wl[209] vdd gnd cell_6t
Xbit_r210_c36 bl[36] br[36] wl[210] vdd gnd cell_6t
Xbit_r211_c36 bl[36] br[36] wl[211] vdd gnd cell_6t
Xbit_r212_c36 bl[36] br[36] wl[212] vdd gnd cell_6t
Xbit_r213_c36 bl[36] br[36] wl[213] vdd gnd cell_6t
Xbit_r214_c36 bl[36] br[36] wl[214] vdd gnd cell_6t
Xbit_r215_c36 bl[36] br[36] wl[215] vdd gnd cell_6t
Xbit_r216_c36 bl[36] br[36] wl[216] vdd gnd cell_6t
Xbit_r217_c36 bl[36] br[36] wl[217] vdd gnd cell_6t
Xbit_r218_c36 bl[36] br[36] wl[218] vdd gnd cell_6t
Xbit_r219_c36 bl[36] br[36] wl[219] vdd gnd cell_6t
Xbit_r220_c36 bl[36] br[36] wl[220] vdd gnd cell_6t
Xbit_r221_c36 bl[36] br[36] wl[221] vdd gnd cell_6t
Xbit_r222_c36 bl[36] br[36] wl[222] vdd gnd cell_6t
Xbit_r223_c36 bl[36] br[36] wl[223] vdd gnd cell_6t
Xbit_r224_c36 bl[36] br[36] wl[224] vdd gnd cell_6t
Xbit_r225_c36 bl[36] br[36] wl[225] vdd gnd cell_6t
Xbit_r226_c36 bl[36] br[36] wl[226] vdd gnd cell_6t
Xbit_r227_c36 bl[36] br[36] wl[227] vdd gnd cell_6t
Xbit_r228_c36 bl[36] br[36] wl[228] vdd gnd cell_6t
Xbit_r229_c36 bl[36] br[36] wl[229] vdd gnd cell_6t
Xbit_r230_c36 bl[36] br[36] wl[230] vdd gnd cell_6t
Xbit_r231_c36 bl[36] br[36] wl[231] vdd gnd cell_6t
Xbit_r232_c36 bl[36] br[36] wl[232] vdd gnd cell_6t
Xbit_r233_c36 bl[36] br[36] wl[233] vdd gnd cell_6t
Xbit_r234_c36 bl[36] br[36] wl[234] vdd gnd cell_6t
Xbit_r235_c36 bl[36] br[36] wl[235] vdd gnd cell_6t
Xbit_r236_c36 bl[36] br[36] wl[236] vdd gnd cell_6t
Xbit_r237_c36 bl[36] br[36] wl[237] vdd gnd cell_6t
Xbit_r238_c36 bl[36] br[36] wl[238] vdd gnd cell_6t
Xbit_r239_c36 bl[36] br[36] wl[239] vdd gnd cell_6t
Xbit_r240_c36 bl[36] br[36] wl[240] vdd gnd cell_6t
Xbit_r241_c36 bl[36] br[36] wl[241] vdd gnd cell_6t
Xbit_r242_c36 bl[36] br[36] wl[242] vdd gnd cell_6t
Xbit_r243_c36 bl[36] br[36] wl[243] vdd gnd cell_6t
Xbit_r244_c36 bl[36] br[36] wl[244] vdd gnd cell_6t
Xbit_r245_c36 bl[36] br[36] wl[245] vdd gnd cell_6t
Xbit_r246_c36 bl[36] br[36] wl[246] vdd gnd cell_6t
Xbit_r247_c36 bl[36] br[36] wl[247] vdd gnd cell_6t
Xbit_r248_c36 bl[36] br[36] wl[248] vdd gnd cell_6t
Xbit_r249_c36 bl[36] br[36] wl[249] vdd gnd cell_6t
Xbit_r250_c36 bl[36] br[36] wl[250] vdd gnd cell_6t
Xbit_r251_c36 bl[36] br[36] wl[251] vdd gnd cell_6t
Xbit_r252_c36 bl[36] br[36] wl[252] vdd gnd cell_6t
Xbit_r253_c36 bl[36] br[36] wl[253] vdd gnd cell_6t
Xbit_r254_c36 bl[36] br[36] wl[254] vdd gnd cell_6t
Xbit_r255_c36 bl[36] br[36] wl[255] vdd gnd cell_6t
Xbit_r0_c37 bl[37] br[37] wl[0] vdd gnd cell_6t
Xbit_r1_c37 bl[37] br[37] wl[1] vdd gnd cell_6t
Xbit_r2_c37 bl[37] br[37] wl[2] vdd gnd cell_6t
Xbit_r3_c37 bl[37] br[37] wl[3] vdd gnd cell_6t
Xbit_r4_c37 bl[37] br[37] wl[4] vdd gnd cell_6t
Xbit_r5_c37 bl[37] br[37] wl[5] vdd gnd cell_6t
Xbit_r6_c37 bl[37] br[37] wl[6] vdd gnd cell_6t
Xbit_r7_c37 bl[37] br[37] wl[7] vdd gnd cell_6t
Xbit_r8_c37 bl[37] br[37] wl[8] vdd gnd cell_6t
Xbit_r9_c37 bl[37] br[37] wl[9] vdd gnd cell_6t
Xbit_r10_c37 bl[37] br[37] wl[10] vdd gnd cell_6t
Xbit_r11_c37 bl[37] br[37] wl[11] vdd gnd cell_6t
Xbit_r12_c37 bl[37] br[37] wl[12] vdd gnd cell_6t
Xbit_r13_c37 bl[37] br[37] wl[13] vdd gnd cell_6t
Xbit_r14_c37 bl[37] br[37] wl[14] vdd gnd cell_6t
Xbit_r15_c37 bl[37] br[37] wl[15] vdd gnd cell_6t
Xbit_r16_c37 bl[37] br[37] wl[16] vdd gnd cell_6t
Xbit_r17_c37 bl[37] br[37] wl[17] vdd gnd cell_6t
Xbit_r18_c37 bl[37] br[37] wl[18] vdd gnd cell_6t
Xbit_r19_c37 bl[37] br[37] wl[19] vdd gnd cell_6t
Xbit_r20_c37 bl[37] br[37] wl[20] vdd gnd cell_6t
Xbit_r21_c37 bl[37] br[37] wl[21] vdd gnd cell_6t
Xbit_r22_c37 bl[37] br[37] wl[22] vdd gnd cell_6t
Xbit_r23_c37 bl[37] br[37] wl[23] vdd gnd cell_6t
Xbit_r24_c37 bl[37] br[37] wl[24] vdd gnd cell_6t
Xbit_r25_c37 bl[37] br[37] wl[25] vdd gnd cell_6t
Xbit_r26_c37 bl[37] br[37] wl[26] vdd gnd cell_6t
Xbit_r27_c37 bl[37] br[37] wl[27] vdd gnd cell_6t
Xbit_r28_c37 bl[37] br[37] wl[28] vdd gnd cell_6t
Xbit_r29_c37 bl[37] br[37] wl[29] vdd gnd cell_6t
Xbit_r30_c37 bl[37] br[37] wl[30] vdd gnd cell_6t
Xbit_r31_c37 bl[37] br[37] wl[31] vdd gnd cell_6t
Xbit_r32_c37 bl[37] br[37] wl[32] vdd gnd cell_6t
Xbit_r33_c37 bl[37] br[37] wl[33] vdd gnd cell_6t
Xbit_r34_c37 bl[37] br[37] wl[34] vdd gnd cell_6t
Xbit_r35_c37 bl[37] br[37] wl[35] vdd gnd cell_6t
Xbit_r36_c37 bl[37] br[37] wl[36] vdd gnd cell_6t
Xbit_r37_c37 bl[37] br[37] wl[37] vdd gnd cell_6t
Xbit_r38_c37 bl[37] br[37] wl[38] vdd gnd cell_6t
Xbit_r39_c37 bl[37] br[37] wl[39] vdd gnd cell_6t
Xbit_r40_c37 bl[37] br[37] wl[40] vdd gnd cell_6t
Xbit_r41_c37 bl[37] br[37] wl[41] vdd gnd cell_6t
Xbit_r42_c37 bl[37] br[37] wl[42] vdd gnd cell_6t
Xbit_r43_c37 bl[37] br[37] wl[43] vdd gnd cell_6t
Xbit_r44_c37 bl[37] br[37] wl[44] vdd gnd cell_6t
Xbit_r45_c37 bl[37] br[37] wl[45] vdd gnd cell_6t
Xbit_r46_c37 bl[37] br[37] wl[46] vdd gnd cell_6t
Xbit_r47_c37 bl[37] br[37] wl[47] vdd gnd cell_6t
Xbit_r48_c37 bl[37] br[37] wl[48] vdd gnd cell_6t
Xbit_r49_c37 bl[37] br[37] wl[49] vdd gnd cell_6t
Xbit_r50_c37 bl[37] br[37] wl[50] vdd gnd cell_6t
Xbit_r51_c37 bl[37] br[37] wl[51] vdd gnd cell_6t
Xbit_r52_c37 bl[37] br[37] wl[52] vdd gnd cell_6t
Xbit_r53_c37 bl[37] br[37] wl[53] vdd gnd cell_6t
Xbit_r54_c37 bl[37] br[37] wl[54] vdd gnd cell_6t
Xbit_r55_c37 bl[37] br[37] wl[55] vdd gnd cell_6t
Xbit_r56_c37 bl[37] br[37] wl[56] vdd gnd cell_6t
Xbit_r57_c37 bl[37] br[37] wl[57] vdd gnd cell_6t
Xbit_r58_c37 bl[37] br[37] wl[58] vdd gnd cell_6t
Xbit_r59_c37 bl[37] br[37] wl[59] vdd gnd cell_6t
Xbit_r60_c37 bl[37] br[37] wl[60] vdd gnd cell_6t
Xbit_r61_c37 bl[37] br[37] wl[61] vdd gnd cell_6t
Xbit_r62_c37 bl[37] br[37] wl[62] vdd gnd cell_6t
Xbit_r63_c37 bl[37] br[37] wl[63] vdd gnd cell_6t
Xbit_r64_c37 bl[37] br[37] wl[64] vdd gnd cell_6t
Xbit_r65_c37 bl[37] br[37] wl[65] vdd gnd cell_6t
Xbit_r66_c37 bl[37] br[37] wl[66] vdd gnd cell_6t
Xbit_r67_c37 bl[37] br[37] wl[67] vdd gnd cell_6t
Xbit_r68_c37 bl[37] br[37] wl[68] vdd gnd cell_6t
Xbit_r69_c37 bl[37] br[37] wl[69] vdd gnd cell_6t
Xbit_r70_c37 bl[37] br[37] wl[70] vdd gnd cell_6t
Xbit_r71_c37 bl[37] br[37] wl[71] vdd gnd cell_6t
Xbit_r72_c37 bl[37] br[37] wl[72] vdd gnd cell_6t
Xbit_r73_c37 bl[37] br[37] wl[73] vdd gnd cell_6t
Xbit_r74_c37 bl[37] br[37] wl[74] vdd gnd cell_6t
Xbit_r75_c37 bl[37] br[37] wl[75] vdd gnd cell_6t
Xbit_r76_c37 bl[37] br[37] wl[76] vdd gnd cell_6t
Xbit_r77_c37 bl[37] br[37] wl[77] vdd gnd cell_6t
Xbit_r78_c37 bl[37] br[37] wl[78] vdd gnd cell_6t
Xbit_r79_c37 bl[37] br[37] wl[79] vdd gnd cell_6t
Xbit_r80_c37 bl[37] br[37] wl[80] vdd gnd cell_6t
Xbit_r81_c37 bl[37] br[37] wl[81] vdd gnd cell_6t
Xbit_r82_c37 bl[37] br[37] wl[82] vdd gnd cell_6t
Xbit_r83_c37 bl[37] br[37] wl[83] vdd gnd cell_6t
Xbit_r84_c37 bl[37] br[37] wl[84] vdd gnd cell_6t
Xbit_r85_c37 bl[37] br[37] wl[85] vdd gnd cell_6t
Xbit_r86_c37 bl[37] br[37] wl[86] vdd gnd cell_6t
Xbit_r87_c37 bl[37] br[37] wl[87] vdd gnd cell_6t
Xbit_r88_c37 bl[37] br[37] wl[88] vdd gnd cell_6t
Xbit_r89_c37 bl[37] br[37] wl[89] vdd gnd cell_6t
Xbit_r90_c37 bl[37] br[37] wl[90] vdd gnd cell_6t
Xbit_r91_c37 bl[37] br[37] wl[91] vdd gnd cell_6t
Xbit_r92_c37 bl[37] br[37] wl[92] vdd gnd cell_6t
Xbit_r93_c37 bl[37] br[37] wl[93] vdd gnd cell_6t
Xbit_r94_c37 bl[37] br[37] wl[94] vdd gnd cell_6t
Xbit_r95_c37 bl[37] br[37] wl[95] vdd gnd cell_6t
Xbit_r96_c37 bl[37] br[37] wl[96] vdd gnd cell_6t
Xbit_r97_c37 bl[37] br[37] wl[97] vdd gnd cell_6t
Xbit_r98_c37 bl[37] br[37] wl[98] vdd gnd cell_6t
Xbit_r99_c37 bl[37] br[37] wl[99] vdd gnd cell_6t
Xbit_r100_c37 bl[37] br[37] wl[100] vdd gnd cell_6t
Xbit_r101_c37 bl[37] br[37] wl[101] vdd gnd cell_6t
Xbit_r102_c37 bl[37] br[37] wl[102] vdd gnd cell_6t
Xbit_r103_c37 bl[37] br[37] wl[103] vdd gnd cell_6t
Xbit_r104_c37 bl[37] br[37] wl[104] vdd gnd cell_6t
Xbit_r105_c37 bl[37] br[37] wl[105] vdd gnd cell_6t
Xbit_r106_c37 bl[37] br[37] wl[106] vdd gnd cell_6t
Xbit_r107_c37 bl[37] br[37] wl[107] vdd gnd cell_6t
Xbit_r108_c37 bl[37] br[37] wl[108] vdd gnd cell_6t
Xbit_r109_c37 bl[37] br[37] wl[109] vdd gnd cell_6t
Xbit_r110_c37 bl[37] br[37] wl[110] vdd gnd cell_6t
Xbit_r111_c37 bl[37] br[37] wl[111] vdd gnd cell_6t
Xbit_r112_c37 bl[37] br[37] wl[112] vdd gnd cell_6t
Xbit_r113_c37 bl[37] br[37] wl[113] vdd gnd cell_6t
Xbit_r114_c37 bl[37] br[37] wl[114] vdd gnd cell_6t
Xbit_r115_c37 bl[37] br[37] wl[115] vdd gnd cell_6t
Xbit_r116_c37 bl[37] br[37] wl[116] vdd gnd cell_6t
Xbit_r117_c37 bl[37] br[37] wl[117] vdd gnd cell_6t
Xbit_r118_c37 bl[37] br[37] wl[118] vdd gnd cell_6t
Xbit_r119_c37 bl[37] br[37] wl[119] vdd gnd cell_6t
Xbit_r120_c37 bl[37] br[37] wl[120] vdd gnd cell_6t
Xbit_r121_c37 bl[37] br[37] wl[121] vdd gnd cell_6t
Xbit_r122_c37 bl[37] br[37] wl[122] vdd gnd cell_6t
Xbit_r123_c37 bl[37] br[37] wl[123] vdd gnd cell_6t
Xbit_r124_c37 bl[37] br[37] wl[124] vdd gnd cell_6t
Xbit_r125_c37 bl[37] br[37] wl[125] vdd gnd cell_6t
Xbit_r126_c37 bl[37] br[37] wl[126] vdd gnd cell_6t
Xbit_r127_c37 bl[37] br[37] wl[127] vdd gnd cell_6t
Xbit_r128_c37 bl[37] br[37] wl[128] vdd gnd cell_6t
Xbit_r129_c37 bl[37] br[37] wl[129] vdd gnd cell_6t
Xbit_r130_c37 bl[37] br[37] wl[130] vdd gnd cell_6t
Xbit_r131_c37 bl[37] br[37] wl[131] vdd gnd cell_6t
Xbit_r132_c37 bl[37] br[37] wl[132] vdd gnd cell_6t
Xbit_r133_c37 bl[37] br[37] wl[133] vdd gnd cell_6t
Xbit_r134_c37 bl[37] br[37] wl[134] vdd gnd cell_6t
Xbit_r135_c37 bl[37] br[37] wl[135] vdd gnd cell_6t
Xbit_r136_c37 bl[37] br[37] wl[136] vdd gnd cell_6t
Xbit_r137_c37 bl[37] br[37] wl[137] vdd gnd cell_6t
Xbit_r138_c37 bl[37] br[37] wl[138] vdd gnd cell_6t
Xbit_r139_c37 bl[37] br[37] wl[139] vdd gnd cell_6t
Xbit_r140_c37 bl[37] br[37] wl[140] vdd gnd cell_6t
Xbit_r141_c37 bl[37] br[37] wl[141] vdd gnd cell_6t
Xbit_r142_c37 bl[37] br[37] wl[142] vdd gnd cell_6t
Xbit_r143_c37 bl[37] br[37] wl[143] vdd gnd cell_6t
Xbit_r144_c37 bl[37] br[37] wl[144] vdd gnd cell_6t
Xbit_r145_c37 bl[37] br[37] wl[145] vdd gnd cell_6t
Xbit_r146_c37 bl[37] br[37] wl[146] vdd gnd cell_6t
Xbit_r147_c37 bl[37] br[37] wl[147] vdd gnd cell_6t
Xbit_r148_c37 bl[37] br[37] wl[148] vdd gnd cell_6t
Xbit_r149_c37 bl[37] br[37] wl[149] vdd gnd cell_6t
Xbit_r150_c37 bl[37] br[37] wl[150] vdd gnd cell_6t
Xbit_r151_c37 bl[37] br[37] wl[151] vdd gnd cell_6t
Xbit_r152_c37 bl[37] br[37] wl[152] vdd gnd cell_6t
Xbit_r153_c37 bl[37] br[37] wl[153] vdd gnd cell_6t
Xbit_r154_c37 bl[37] br[37] wl[154] vdd gnd cell_6t
Xbit_r155_c37 bl[37] br[37] wl[155] vdd gnd cell_6t
Xbit_r156_c37 bl[37] br[37] wl[156] vdd gnd cell_6t
Xbit_r157_c37 bl[37] br[37] wl[157] vdd gnd cell_6t
Xbit_r158_c37 bl[37] br[37] wl[158] vdd gnd cell_6t
Xbit_r159_c37 bl[37] br[37] wl[159] vdd gnd cell_6t
Xbit_r160_c37 bl[37] br[37] wl[160] vdd gnd cell_6t
Xbit_r161_c37 bl[37] br[37] wl[161] vdd gnd cell_6t
Xbit_r162_c37 bl[37] br[37] wl[162] vdd gnd cell_6t
Xbit_r163_c37 bl[37] br[37] wl[163] vdd gnd cell_6t
Xbit_r164_c37 bl[37] br[37] wl[164] vdd gnd cell_6t
Xbit_r165_c37 bl[37] br[37] wl[165] vdd gnd cell_6t
Xbit_r166_c37 bl[37] br[37] wl[166] vdd gnd cell_6t
Xbit_r167_c37 bl[37] br[37] wl[167] vdd gnd cell_6t
Xbit_r168_c37 bl[37] br[37] wl[168] vdd gnd cell_6t
Xbit_r169_c37 bl[37] br[37] wl[169] vdd gnd cell_6t
Xbit_r170_c37 bl[37] br[37] wl[170] vdd gnd cell_6t
Xbit_r171_c37 bl[37] br[37] wl[171] vdd gnd cell_6t
Xbit_r172_c37 bl[37] br[37] wl[172] vdd gnd cell_6t
Xbit_r173_c37 bl[37] br[37] wl[173] vdd gnd cell_6t
Xbit_r174_c37 bl[37] br[37] wl[174] vdd gnd cell_6t
Xbit_r175_c37 bl[37] br[37] wl[175] vdd gnd cell_6t
Xbit_r176_c37 bl[37] br[37] wl[176] vdd gnd cell_6t
Xbit_r177_c37 bl[37] br[37] wl[177] vdd gnd cell_6t
Xbit_r178_c37 bl[37] br[37] wl[178] vdd gnd cell_6t
Xbit_r179_c37 bl[37] br[37] wl[179] vdd gnd cell_6t
Xbit_r180_c37 bl[37] br[37] wl[180] vdd gnd cell_6t
Xbit_r181_c37 bl[37] br[37] wl[181] vdd gnd cell_6t
Xbit_r182_c37 bl[37] br[37] wl[182] vdd gnd cell_6t
Xbit_r183_c37 bl[37] br[37] wl[183] vdd gnd cell_6t
Xbit_r184_c37 bl[37] br[37] wl[184] vdd gnd cell_6t
Xbit_r185_c37 bl[37] br[37] wl[185] vdd gnd cell_6t
Xbit_r186_c37 bl[37] br[37] wl[186] vdd gnd cell_6t
Xbit_r187_c37 bl[37] br[37] wl[187] vdd gnd cell_6t
Xbit_r188_c37 bl[37] br[37] wl[188] vdd gnd cell_6t
Xbit_r189_c37 bl[37] br[37] wl[189] vdd gnd cell_6t
Xbit_r190_c37 bl[37] br[37] wl[190] vdd gnd cell_6t
Xbit_r191_c37 bl[37] br[37] wl[191] vdd gnd cell_6t
Xbit_r192_c37 bl[37] br[37] wl[192] vdd gnd cell_6t
Xbit_r193_c37 bl[37] br[37] wl[193] vdd gnd cell_6t
Xbit_r194_c37 bl[37] br[37] wl[194] vdd gnd cell_6t
Xbit_r195_c37 bl[37] br[37] wl[195] vdd gnd cell_6t
Xbit_r196_c37 bl[37] br[37] wl[196] vdd gnd cell_6t
Xbit_r197_c37 bl[37] br[37] wl[197] vdd gnd cell_6t
Xbit_r198_c37 bl[37] br[37] wl[198] vdd gnd cell_6t
Xbit_r199_c37 bl[37] br[37] wl[199] vdd gnd cell_6t
Xbit_r200_c37 bl[37] br[37] wl[200] vdd gnd cell_6t
Xbit_r201_c37 bl[37] br[37] wl[201] vdd gnd cell_6t
Xbit_r202_c37 bl[37] br[37] wl[202] vdd gnd cell_6t
Xbit_r203_c37 bl[37] br[37] wl[203] vdd gnd cell_6t
Xbit_r204_c37 bl[37] br[37] wl[204] vdd gnd cell_6t
Xbit_r205_c37 bl[37] br[37] wl[205] vdd gnd cell_6t
Xbit_r206_c37 bl[37] br[37] wl[206] vdd gnd cell_6t
Xbit_r207_c37 bl[37] br[37] wl[207] vdd gnd cell_6t
Xbit_r208_c37 bl[37] br[37] wl[208] vdd gnd cell_6t
Xbit_r209_c37 bl[37] br[37] wl[209] vdd gnd cell_6t
Xbit_r210_c37 bl[37] br[37] wl[210] vdd gnd cell_6t
Xbit_r211_c37 bl[37] br[37] wl[211] vdd gnd cell_6t
Xbit_r212_c37 bl[37] br[37] wl[212] vdd gnd cell_6t
Xbit_r213_c37 bl[37] br[37] wl[213] vdd gnd cell_6t
Xbit_r214_c37 bl[37] br[37] wl[214] vdd gnd cell_6t
Xbit_r215_c37 bl[37] br[37] wl[215] vdd gnd cell_6t
Xbit_r216_c37 bl[37] br[37] wl[216] vdd gnd cell_6t
Xbit_r217_c37 bl[37] br[37] wl[217] vdd gnd cell_6t
Xbit_r218_c37 bl[37] br[37] wl[218] vdd gnd cell_6t
Xbit_r219_c37 bl[37] br[37] wl[219] vdd gnd cell_6t
Xbit_r220_c37 bl[37] br[37] wl[220] vdd gnd cell_6t
Xbit_r221_c37 bl[37] br[37] wl[221] vdd gnd cell_6t
Xbit_r222_c37 bl[37] br[37] wl[222] vdd gnd cell_6t
Xbit_r223_c37 bl[37] br[37] wl[223] vdd gnd cell_6t
Xbit_r224_c37 bl[37] br[37] wl[224] vdd gnd cell_6t
Xbit_r225_c37 bl[37] br[37] wl[225] vdd gnd cell_6t
Xbit_r226_c37 bl[37] br[37] wl[226] vdd gnd cell_6t
Xbit_r227_c37 bl[37] br[37] wl[227] vdd gnd cell_6t
Xbit_r228_c37 bl[37] br[37] wl[228] vdd gnd cell_6t
Xbit_r229_c37 bl[37] br[37] wl[229] vdd gnd cell_6t
Xbit_r230_c37 bl[37] br[37] wl[230] vdd gnd cell_6t
Xbit_r231_c37 bl[37] br[37] wl[231] vdd gnd cell_6t
Xbit_r232_c37 bl[37] br[37] wl[232] vdd gnd cell_6t
Xbit_r233_c37 bl[37] br[37] wl[233] vdd gnd cell_6t
Xbit_r234_c37 bl[37] br[37] wl[234] vdd gnd cell_6t
Xbit_r235_c37 bl[37] br[37] wl[235] vdd gnd cell_6t
Xbit_r236_c37 bl[37] br[37] wl[236] vdd gnd cell_6t
Xbit_r237_c37 bl[37] br[37] wl[237] vdd gnd cell_6t
Xbit_r238_c37 bl[37] br[37] wl[238] vdd gnd cell_6t
Xbit_r239_c37 bl[37] br[37] wl[239] vdd gnd cell_6t
Xbit_r240_c37 bl[37] br[37] wl[240] vdd gnd cell_6t
Xbit_r241_c37 bl[37] br[37] wl[241] vdd gnd cell_6t
Xbit_r242_c37 bl[37] br[37] wl[242] vdd gnd cell_6t
Xbit_r243_c37 bl[37] br[37] wl[243] vdd gnd cell_6t
Xbit_r244_c37 bl[37] br[37] wl[244] vdd gnd cell_6t
Xbit_r245_c37 bl[37] br[37] wl[245] vdd gnd cell_6t
Xbit_r246_c37 bl[37] br[37] wl[246] vdd gnd cell_6t
Xbit_r247_c37 bl[37] br[37] wl[247] vdd gnd cell_6t
Xbit_r248_c37 bl[37] br[37] wl[248] vdd gnd cell_6t
Xbit_r249_c37 bl[37] br[37] wl[249] vdd gnd cell_6t
Xbit_r250_c37 bl[37] br[37] wl[250] vdd gnd cell_6t
Xbit_r251_c37 bl[37] br[37] wl[251] vdd gnd cell_6t
Xbit_r252_c37 bl[37] br[37] wl[252] vdd gnd cell_6t
Xbit_r253_c37 bl[37] br[37] wl[253] vdd gnd cell_6t
Xbit_r254_c37 bl[37] br[37] wl[254] vdd gnd cell_6t
Xbit_r255_c37 bl[37] br[37] wl[255] vdd gnd cell_6t
Xbit_r0_c38 bl[38] br[38] wl[0] vdd gnd cell_6t
Xbit_r1_c38 bl[38] br[38] wl[1] vdd gnd cell_6t
Xbit_r2_c38 bl[38] br[38] wl[2] vdd gnd cell_6t
Xbit_r3_c38 bl[38] br[38] wl[3] vdd gnd cell_6t
Xbit_r4_c38 bl[38] br[38] wl[4] vdd gnd cell_6t
Xbit_r5_c38 bl[38] br[38] wl[5] vdd gnd cell_6t
Xbit_r6_c38 bl[38] br[38] wl[6] vdd gnd cell_6t
Xbit_r7_c38 bl[38] br[38] wl[7] vdd gnd cell_6t
Xbit_r8_c38 bl[38] br[38] wl[8] vdd gnd cell_6t
Xbit_r9_c38 bl[38] br[38] wl[9] vdd gnd cell_6t
Xbit_r10_c38 bl[38] br[38] wl[10] vdd gnd cell_6t
Xbit_r11_c38 bl[38] br[38] wl[11] vdd gnd cell_6t
Xbit_r12_c38 bl[38] br[38] wl[12] vdd gnd cell_6t
Xbit_r13_c38 bl[38] br[38] wl[13] vdd gnd cell_6t
Xbit_r14_c38 bl[38] br[38] wl[14] vdd gnd cell_6t
Xbit_r15_c38 bl[38] br[38] wl[15] vdd gnd cell_6t
Xbit_r16_c38 bl[38] br[38] wl[16] vdd gnd cell_6t
Xbit_r17_c38 bl[38] br[38] wl[17] vdd gnd cell_6t
Xbit_r18_c38 bl[38] br[38] wl[18] vdd gnd cell_6t
Xbit_r19_c38 bl[38] br[38] wl[19] vdd gnd cell_6t
Xbit_r20_c38 bl[38] br[38] wl[20] vdd gnd cell_6t
Xbit_r21_c38 bl[38] br[38] wl[21] vdd gnd cell_6t
Xbit_r22_c38 bl[38] br[38] wl[22] vdd gnd cell_6t
Xbit_r23_c38 bl[38] br[38] wl[23] vdd gnd cell_6t
Xbit_r24_c38 bl[38] br[38] wl[24] vdd gnd cell_6t
Xbit_r25_c38 bl[38] br[38] wl[25] vdd gnd cell_6t
Xbit_r26_c38 bl[38] br[38] wl[26] vdd gnd cell_6t
Xbit_r27_c38 bl[38] br[38] wl[27] vdd gnd cell_6t
Xbit_r28_c38 bl[38] br[38] wl[28] vdd gnd cell_6t
Xbit_r29_c38 bl[38] br[38] wl[29] vdd gnd cell_6t
Xbit_r30_c38 bl[38] br[38] wl[30] vdd gnd cell_6t
Xbit_r31_c38 bl[38] br[38] wl[31] vdd gnd cell_6t
Xbit_r32_c38 bl[38] br[38] wl[32] vdd gnd cell_6t
Xbit_r33_c38 bl[38] br[38] wl[33] vdd gnd cell_6t
Xbit_r34_c38 bl[38] br[38] wl[34] vdd gnd cell_6t
Xbit_r35_c38 bl[38] br[38] wl[35] vdd gnd cell_6t
Xbit_r36_c38 bl[38] br[38] wl[36] vdd gnd cell_6t
Xbit_r37_c38 bl[38] br[38] wl[37] vdd gnd cell_6t
Xbit_r38_c38 bl[38] br[38] wl[38] vdd gnd cell_6t
Xbit_r39_c38 bl[38] br[38] wl[39] vdd gnd cell_6t
Xbit_r40_c38 bl[38] br[38] wl[40] vdd gnd cell_6t
Xbit_r41_c38 bl[38] br[38] wl[41] vdd gnd cell_6t
Xbit_r42_c38 bl[38] br[38] wl[42] vdd gnd cell_6t
Xbit_r43_c38 bl[38] br[38] wl[43] vdd gnd cell_6t
Xbit_r44_c38 bl[38] br[38] wl[44] vdd gnd cell_6t
Xbit_r45_c38 bl[38] br[38] wl[45] vdd gnd cell_6t
Xbit_r46_c38 bl[38] br[38] wl[46] vdd gnd cell_6t
Xbit_r47_c38 bl[38] br[38] wl[47] vdd gnd cell_6t
Xbit_r48_c38 bl[38] br[38] wl[48] vdd gnd cell_6t
Xbit_r49_c38 bl[38] br[38] wl[49] vdd gnd cell_6t
Xbit_r50_c38 bl[38] br[38] wl[50] vdd gnd cell_6t
Xbit_r51_c38 bl[38] br[38] wl[51] vdd gnd cell_6t
Xbit_r52_c38 bl[38] br[38] wl[52] vdd gnd cell_6t
Xbit_r53_c38 bl[38] br[38] wl[53] vdd gnd cell_6t
Xbit_r54_c38 bl[38] br[38] wl[54] vdd gnd cell_6t
Xbit_r55_c38 bl[38] br[38] wl[55] vdd gnd cell_6t
Xbit_r56_c38 bl[38] br[38] wl[56] vdd gnd cell_6t
Xbit_r57_c38 bl[38] br[38] wl[57] vdd gnd cell_6t
Xbit_r58_c38 bl[38] br[38] wl[58] vdd gnd cell_6t
Xbit_r59_c38 bl[38] br[38] wl[59] vdd gnd cell_6t
Xbit_r60_c38 bl[38] br[38] wl[60] vdd gnd cell_6t
Xbit_r61_c38 bl[38] br[38] wl[61] vdd gnd cell_6t
Xbit_r62_c38 bl[38] br[38] wl[62] vdd gnd cell_6t
Xbit_r63_c38 bl[38] br[38] wl[63] vdd gnd cell_6t
Xbit_r64_c38 bl[38] br[38] wl[64] vdd gnd cell_6t
Xbit_r65_c38 bl[38] br[38] wl[65] vdd gnd cell_6t
Xbit_r66_c38 bl[38] br[38] wl[66] vdd gnd cell_6t
Xbit_r67_c38 bl[38] br[38] wl[67] vdd gnd cell_6t
Xbit_r68_c38 bl[38] br[38] wl[68] vdd gnd cell_6t
Xbit_r69_c38 bl[38] br[38] wl[69] vdd gnd cell_6t
Xbit_r70_c38 bl[38] br[38] wl[70] vdd gnd cell_6t
Xbit_r71_c38 bl[38] br[38] wl[71] vdd gnd cell_6t
Xbit_r72_c38 bl[38] br[38] wl[72] vdd gnd cell_6t
Xbit_r73_c38 bl[38] br[38] wl[73] vdd gnd cell_6t
Xbit_r74_c38 bl[38] br[38] wl[74] vdd gnd cell_6t
Xbit_r75_c38 bl[38] br[38] wl[75] vdd gnd cell_6t
Xbit_r76_c38 bl[38] br[38] wl[76] vdd gnd cell_6t
Xbit_r77_c38 bl[38] br[38] wl[77] vdd gnd cell_6t
Xbit_r78_c38 bl[38] br[38] wl[78] vdd gnd cell_6t
Xbit_r79_c38 bl[38] br[38] wl[79] vdd gnd cell_6t
Xbit_r80_c38 bl[38] br[38] wl[80] vdd gnd cell_6t
Xbit_r81_c38 bl[38] br[38] wl[81] vdd gnd cell_6t
Xbit_r82_c38 bl[38] br[38] wl[82] vdd gnd cell_6t
Xbit_r83_c38 bl[38] br[38] wl[83] vdd gnd cell_6t
Xbit_r84_c38 bl[38] br[38] wl[84] vdd gnd cell_6t
Xbit_r85_c38 bl[38] br[38] wl[85] vdd gnd cell_6t
Xbit_r86_c38 bl[38] br[38] wl[86] vdd gnd cell_6t
Xbit_r87_c38 bl[38] br[38] wl[87] vdd gnd cell_6t
Xbit_r88_c38 bl[38] br[38] wl[88] vdd gnd cell_6t
Xbit_r89_c38 bl[38] br[38] wl[89] vdd gnd cell_6t
Xbit_r90_c38 bl[38] br[38] wl[90] vdd gnd cell_6t
Xbit_r91_c38 bl[38] br[38] wl[91] vdd gnd cell_6t
Xbit_r92_c38 bl[38] br[38] wl[92] vdd gnd cell_6t
Xbit_r93_c38 bl[38] br[38] wl[93] vdd gnd cell_6t
Xbit_r94_c38 bl[38] br[38] wl[94] vdd gnd cell_6t
Xbit_r95_c38 bl[38] br[38] wl[95] vdd gnd cell_6t
Xbit_r96_c38 bl[38] br[38] wl[96] vdd gnd cell_6t
Xbit_r97_c38 bl[38] br[38] wl[97] vdd gnd cell_6t
Xbit_r98_c38 bl[38] br[38] wl[98] vdd gnd cell_6t
Xbit_r99_c38 bl[38] br[38] wl[99] vdd gnd cell_6t
Xbit_r100_c38 bl[38] br[38] wl[100] vdd gnd cell_6t
Xbit_r101_c38 bl[38] br[38] wl[101] vdd gnd cell_6t
Xbit_r102_c38 bl[38] br[38] wl[102] vdd gnd cell_6t
Xbit_r103_c38 bl[38] br[38] wl[103] vdd gnd cell_6t
Xbit_r104_c38 bl[38] br[38] wl[104] vdd gnd cell_6t
Xbit_r105_c38 bl[38] br[38] wl[105] vdd gnd cell_6t
Xbit_r106_c38 bl[38] br[38] wl[106] vdd gnd cell_6t
Xbit_r107_c38 bl[38] br[38] wl[107] vdd gnd cell_6t
Xbit_r108_c38 bl[38] br[38] wl[108] vdd gnd cell_6t
Xbit_r109_c38 bl[38] br[38] wl[109] vdd gnd cell_6t
Xbit_r110_c38 bl[38] br[38] wl[110] vdd gnd cell_6t
Xbit_r111_c38 bl[38] br[38] wl[111] vdd gnd cell_6t
Xbit_r112_c38 bl[38] br[38] wl[112] vdd gnd cell_6t
Xbit_r113_c38 bl[38] br[38] wl[113] vdd gnd cell_6t
Xbit_r114_c38 bl[38] br[38] wl[114] vdd gnd cell_6t
Xbit_r115_c38 bl[38] br[38] wl[115] vdd gnd cell_6t
Xbit_r116_c38 bl[38] br[38] wl[116] vdd gnd cell_6t
Xbit_r117_c38 bl[38] br[38] wl[117] vdd gnd cell_6t
Xbit_r118_c38 bl[38] br[38] wl[118] vdd gnd cell_6t
Xbit_r119_c38 bl[38] br[38] wl[119] vdd gnd cell_6t
Xbit_r120_c38 bl[38] br[38] wl[120] vdd gnd cell_6t
Xbit_r121_c38 bl[38] br[38] wl[121] vdd gnd cell_6t
Xbit_r122_c38 bl[38] br[38] wl[122] vdd gnd cell_6t
Xbit_r123_c38 bl[38] br[38] wl[123] vdd gnd cell_6t
Xbit_r124_c38 bl[38] br[38] wl[124] vdd gnd cell_6t
Xbit_r125_c38 bl[38] br[38] wl[125] vdd gnd cell_6t
Xbit_r126_c38 bl[38] br[38] wl[126] vdd gnd cell_6t
Xbit_r127_c38 bl[38] br[38] wl[127] vdd gnd cell_6t
Xbit_r128_c38 bl[38] br[38] wl[128] vdd gnd cell_6t
Xbit_r129_c38 bl[38] br[38] wl[129] vdd gnd cell_6t
Xbit_r130_c38 bl[38] br[38] wl[130] vdd gnd cell_6t
Xbit_r131_c38 bl[38] br[38] wl[131] vdd gnd cell_6t
Xbit_r132_c38 bl[38] br[38] wl[132] vdd gnd cell_6t
Xbit_r133_c38 bl[38] br[38] wl[133] vdd gnd cell_6t
Xbit_r134_c38 bl[38] br[38] wl[134] vdd gnd cell_6t
Xbit_r135_c38 bl[38] br[38] wl[135] vdd gnd cell_6t
Xbit_r136_c38 bl[38] br[38] wl[136] vdd gnd cell_6t
Xbit_r137_c38 bl[38] br[38] wl[137] vdd gnd cell_6t
Xbit_r138_c38 bl[38] br[38] wl[138] vdd gnd cell_6t
Xbit_r139_c38 bl[38] br[38] wl[139] vdd gnd cell_6t
Xbit_r140_c38 bl[38] br[38] wl[140] vdd gnd cell_6t
Xbit_r141_c38 bl[38] br[38] wl[141] vdd gnd cell_6t
Xbit_r142_c38 bl[38] br[38] wl[142] vdd gnd cell_6t
Xbit_r143_c38 bl[38] br[38] wl[143] vdd gnd cell_6t
Xbit_r144_c38 bl[38] br[38] wl[144] vdd gnd cell_6t
Xbit_r145_c38 bl[38] br[38] wl[145] vdd gnd cell_6t
Xbit_r146_c38 bl[38] br[38] wl[146] vdd gnd cell_6t
Xbit_r147_c38 bl[38] br[38] wl[147] vdd gnd cell_6t
Xbit_r148_c38 bl[38] br[38] wl[148] vdd gnd cell_6t
Xbit_r149_c38 bl[38] br[38] wl[149] vdd gnd cell_6t
Xbit_r150_c38 bl[38] br[38] wl[150] vdd gnd cell_6t
Xbit_r151_c38 bl[38] br[38] wl[151] vdd gnd cell_6t
Xbit_r152_c38 bl[38] br[38] wl[152] vdd gnd cell_6t
Xbit_r153_c38 bl[38] br[38] wl[153] vdd gnd cell_6t
Xbit_r154_c38 bl[38] br[38] wl[154] vdd gnd cell_6t
Xbit_r155_c38 bl[38] br[38] wl[155] vdd gnd cell_6t
Xbit_r156_c38 bl[38] br[38] wl[156] vdd gnd cell_6t
Xbit_r157_c38 bl[38] br[38] wl[157] vdd gnd cell_6t
Xbit_r158_c38 bl[38] br[38] wl[158] vdd gnd cell_6t
Xbit_r159_c38 bl[38] br[38] wl[159] vdd gnd cell_6t
Xbit_r160_c38 bl[38] br[38] wl[160] vdd gnd cell_6t
Xbit_r161_c38 bl[38] br[38] wl[161] vdd gnd cell_6t
Xbit_r162_c38 bl[38] br[38] wl[162] vdd gnd cell_6t
Xbit_r163_c38 bl[38] br[38] wl[163] vdd gnd cell_6t
Xbit_r164_c38 bl[38] br[38] wl[164] vdd gnd cell_6t
Xbit_r165_c38 bl[38] br[38] wl[165] vdd gnd cell_6t
Xbit_r166_c38 bl[38] br[38] wl[166] vdd gnd cell_6t
Xbit_r167_c38 bl[38] br[38] wl[167] vdd gnd cell_6t
Xbit_r168_c38 bl[38] br[38] wl[168] vdd gnd cell_6t
Xbit_r169_c38 bl[38] br[38] wl[169] vdd gnd cell_6t
Xbit_r170_c38 bl[38] br[38] wl[170] vdd gnd cell_6t
Xbit_r171_c38 bl[38] br[38] wl[171] vdd gnd cell_6t
Xbit_r172_c38 bl[38] br[38] wl[172] vdd gnd cell_6t
Xbit_r173_c38 bl[38] br[38] wl[173] vdd gnd cell_6t
Xbit_r174_c38 bl[38] br[38] wl[174] vdd gnd cell_6t
Xbit_r175_c38 bl[38] br[38] wl[175] vdd gnd cell_6t
Xbit_r176_c38 bl[38] br[38] wl[176] vdd gnd cell_6t
Xbit_r177_c38 bl[38] br[38] wl[177] vdd gnd cell_6t
Xbit_r178_c38 bl[38] br[38] wl[178] vdd gnd cell_6t
Xbit_r179_c38 bl[38] br[38] wl[179] vdd gnd cell_6t
Xbit_r180_c38 bl[38] br[38] wl[180] vdd gnd cell_6t
Xbit_r181_c38 bl[38] br[38] wl[181] vdd gnd cell_6t
Xbit_r182_c38 bl[38] br[38] wl[182] vdd gnd cell_6t
Xbit_r183_c38 bl[38] br[38] wl[183] vdd gnd cell_6t
Xbit_r184_c38 bl[38] br[38] wl[184] vdd gnd cell_6t
Xbit_r185_c38 bl[38] br[38] wl[185] vdd gnd cell_6t
Xbit_r186_c38 bl[38] br[38] wl[186] vdd gnd cell_6t
Xbit_r187_c38 bl[38] br[38] wl[187] vdd gnd cell_6t
Xbit_r188_c38 bl[38] br[38] wl[188] vdd gnd cell_6t
Xbit_r189_c38 bl[38] br[38] wl[189] vdd gnd cell_6t
Xbit_r190_c38 bl[38] br[38] wl[190] vdd gnd cell_6t
Xbit_r191_c38 bl[38] br[38] wl[191] vdd gnd cell_6t
Xbit_r192_c38 bl[38] br[38] wl[192] vdd gnd cell_6t
Xbit_r193_c38 bl[38] br[38] wl[193] vdd gnd cell_6t
Xbit_r194_c38 bl[38] br[38] wl[194] vdd gnd cell_6t
Xbit_r195_c38 bl[38] br[38] wl[195] vdd gnd cell_6t
Xbit_r196_c38 bl[38] br[38] wl[196] vdd gnd cell_6t
Xbit_r197_c38 bl[38] br[38] wl[197] vdd gnd cell_6t
Xbit_r198_c38 bl[38] br[38] wl[198] vdd gnd cell_6t
Xbit_r199_c38 bl[38] br[38] wl[199] vdd gnd cell_6t
Xbit_r200_c38 bl[38] br[38] wl[200] vdd gnd cell_6t
Xbit_r201_c38 bl[38] br[38] wl[201] vdd gnd cell_6t
Xbit_r202_c38 bl[38] br[38] wl[202] vdd gnd cell_6t
Xbit_r203_c38 bl[38] br[38] wl[203] vdd gnd cell_6t
Xbit_r204_c38 bl[38] br[38] wl[204] vdd gnd cell_6t
Xbit_r205_c38 bl[38] br[38] wl[205] vdd gnd cell_6t
Xbit_r206_c38 bl[38] br[38] wl[206] vdd gnd cell_6t
Xbit_r207_c38 bl[38] br[38] wl[207] vdd gnd cell_6t
Xbit_r208_c38 bl[38] br[38] wl[208] vdd gnd cell_6t
Xbit_r209_c38 bl[38] br[38] wl[209] vdd gnd cell_6t
Xbit_r210_c38 bl[38] br[38] wl[210] vdd gnd cell_6t
Xbit_r211_c38 bl[38] br[38] wl[211] vdd gnd cell_6t
Xbit_r212_c38 bl[38] br[38] wl[212] vdd gnd cell_6t
Xbit_r213_c38 bl[38] br[38] wl[213] vdd gnd cell_6t
Xbit_r214_c38 bl[38] br[38] wl[214] vdd gnd cell_6t
Xbit_r215_c38 bl[38] br[38] wl[215] vdd gnd cell_6t
Xbit_r216_c38 bl[38] br[38] wl[216] vdd gnd cell_6t
Xbit_r217_c38 bl[38] br[38] wl[217] vdd gnd cell_6t
Xbit_r218_c38 bl[38] br[38] wl[218] vdd gnd cell_6t
Xbit_r219_c38 bl[38] br[38] wl[219] vdd gnd cell_6t
Xbit_r220_c38 bl[38] br[38] wl[220] vdd gnd cell_6t
Xbit_r221_c38 bl[38] br[38] wl[221] vdd gnd cell_6t
Xbit_r222_c38 bl[38] br[38] wl[222] vdd gnd cell_6t
Xbit_r223_c38 bl[38] br[38] wl[223] vdd gnd cell_6t
Xbit_r224_c38 bl[38] br[38] wl[224] vdd gnd cell_6t
Xbit_r225_c38 bl[38] br[38] wl[225] vdd gnd cell_6t
Xbit_r226_c38 bl[38] br[38] wl[226] vdd gnd cell_6t
Xbit_r227_c38 bl[38] br[38] wl[227] vdd gnd cell_6t
Xbit_r228_c38 bl[38] br[38] wl[228] vdd gnd cell_6t
Xbit_r229_c38 bl[38] br[38] wl[229] vdd gnd cell_6t
Xbit_r230_c38 bl[38] br[38] wl[230] vdd gnd cell_6t
Xbit_r231_c38 bl[38] br[38] wl[231] vdd gnd cell_6t
Xbit_r232_c38 bl[38] br[38] wl[232] vdd gnd cell_6t
Xbit_r233_c38 bl[38] br[38] wl[233] vdd gnd cell_6t
Xbit_r234_c38 bl[38] br[38] wl[234] vdd gnd cell_6t
Xbit_r235_c38 bl[38] br[38] wl[235] vdd gnd cell_6t
Xbit_r236_c38 bl[38] br[38] wl[236] vdd gnd cell_6t
Xbit_r237_c38 bl[38] br[38] wl[237] vdd gnd cell_6t
Xbit_r238_c38 bl[38] br[38] wl[238] vdd gnd cell_6t
Xbit_r239_c38 bl[38] br[38] wl[239] vdd gnd cell_6t
Xbit_r240_c38 bl[38] br[38] wl[240] vdd gnd cell_6t
Xbit_r241_c38 bl[38] br[38] wl[241] vdd gnd cell_6t
Xbit_r242_c38 bl[38] br[38] wl[242] vdd gnd cell_6t
Xbit_r243_c38 bl[38] br[38] wl[243] vdd gnd cell_6t
Xbit_r244_c38 bl[38] br[38] wl[244] vdd gnd cell_6t
Xbit_r245_c38 bl[38] br[38] wl[245] vdd gnd cell_6t
Xbit_r246_c38 bl[38] br[38] wl[246] vdd gnd cell_6t
Xbit_r247_c38 bl[38] br[38] wl[247] vdd gnd cell_6t
Xbit_r248_c38 bl[38] br[38] wl[248] vdd gnd cell_6t
Xbit_r249_c38 bl[38] br[38] wl[249] vdd gnd cell_6t
Xbit_r250_c38 bl[38] br[38] wl[250] vdd gnd cell_6t
Xbit_r251_c38 bl[38] br[38] wl[251] vdd gnd cell_6t
Xbit_r252_c38 bl[38] br[38] wl[252] vdd gnd cell_6t
Xbit_r253_c38 bl[38] br[38] wl[253] vdd gnd cell_6t
Xbit_r254_c38 bl[38] br[38] wl[254] vdd gnd cell_6t
Xbit_r255_c38 bl[38] br[38] wl[255] vdd gnd cell_6t
Xbit_r0_c39 bl[39] br[39] wl[0] vdd gnd cell_6t
Xbit_r1_c39 bl[39] br[39] wl[1] vdd gnd cell_6t
Xbit_r2_c39 bl[39] br[39] wl[2] vdd gnd cell_6t
Xbit_r3_c39 bl[39] br[39] wl[3] vdd gnd cell_6t
Xbit_r4_c39 bl[39] br[39] wl[4] vdd gnd cell_6t
Xbit_r5_c39 bl[39] br[39] wl[5] vdd gnd cell_6t
Xbit_r6_c39 bl[39] br[39] wl[6] vdd gnd cell_6t
Xbit_r7_c39 bl[39] br[39] wl[7] vdd gnd cell_6t
Xbit_r8_c39 bl[39] br[39] wl[8] vdd gnd cell_6t
Xbit_r9_c39 bl[39] br[39] wl[9] vdd gnd cell_6t
Xbit_r10_c39 bl[39] br[39] wl[10] vdd gnd cell_6t
Xbit_r11_c39 bl[39] br[39] wl[11] vdd gnd cell_6t
Xbit_r12_c39 bl[39] br[39] wl[12] vdd gnd cell_6t
Xbit_r13_c39 bl[39] br[39] wl[13] vdd gnd cell_6t
Xbit_r14_c39 bl[39] br[39] wl[14] vdd gnd cell_6t
Xbit_r15_c39 bl[39] br[39] wl[15] vdd gnd cell_6t
Xbit_r16_c39 bl[39] br[39] wl[16] vdd gnd cell_6t
Xbit_r17_c39 bl[39] br[39] wl[17] vdd gnd cell_6t
Xbit_r18_c39 bl[39] br[39] wl[18] vdd gnd cell_6t
Xbit_r19_c39 bl[39] br[39] wl[19] vdd gnd cell_6t
Xbit_r20_c39 bl[39] br[39] wl[20] vdd gnd cell_6t
Xbit_r21_c39 bl[39] br[39] wl[21] vdd gnd cell_6t
Xbit_r22_c39 bl[39] br[39] wl[22] vdd gnd cell_6t
Xbit_r23_c39 bl[39] br[39] wl[23] vdd gnd cell_6t
Xbit_r24_c39 bl[39] br[39] wl[24] vdd gnd cell_6t
Xbit_r25_c39 bl[39] br[39] wl[25] vdd gnd cell_6t
Xbit_r26_c39 bl[39] br[39] wl[26] vdd gnd cell_6t
Xbit_r27_c39 bl[39] br[39] wl[27] vdd gnd cell_6t
Xbit_r28_c39 bl[39] br[39] wl[28] vdd gnd cell_6t
Xbit_r29_c39 bl[39] br[39] wl[29] vdd gnd cell_6t
Xbit_r30_c39 bl[39] br[39] wl[30] vdd gnd cell_6t
Xbit_r31_c39 bl[39] br[39] wl[31] vdd gnd cell_6t
Xbit_r32_c39 bl[39] br[39] wl[32] vdd gnd cell_6t
Xbit_r33_c39 bl[39] br[39] wl[33] vdd gnd cell_6t
Xbit_r34_c39 bl[39] br[39] wl[34] vdd gnd cell_6t
Xbit_r35_c39 bl[39] br[39] wl[35] vdd gnd cell_6t
Xbit_r36_c39 bl[39] br[39] wl[36] vdd gnd cell_6t
Xbit_r37_c39 bl[39] br[39] wl[37] vdd gnd cell_6t
Xbit_r38_c39 bl[39] br[39] wl[38] vdd gnd cell_6t
Xbit_r39_c39 bl[39] br[39] wl[39] vdd gnd cell_6t
Xbit_r40_c39 bl[39] br[39] wl[40] vdd gnd cell_6t
Xbit_r41_c39 bl[39] br[39] wl[41] vdd gnd cell_6t
Xbit_r42_c39 bl[39] br[39] wl[42] vdd gnd cell_6t
Xbit_r43_c39 bl[39] br[39] wl[43] vdd gnd cell_6t
Xbit_r44_c39 bl[39] br[39] wl[44] vdd gnd cell_6t
Xbit_r45_c39 bl[39] br[39] wl[45] vdd gnd cell_6t
Xbit_r46_c39 bl[39] br[39] wl[46] vdd gnd cell_6t
Xbit_r47_c39 bl[39] br[39] wl[47] vdd gnd cell_6t
Xbit_r48_c39 bl[39] br[39] wl[48] vdd gnd cell_6t
Xbit_r49_c39 bl[39] br[39] wl[49] vdd gnd cell_6t
Xbit_r50_c39 bl[39] br[39] wl[50] vdd gnd cell_6t
Xbit_r51_c39 bl[39] br[39] wl[51] vdd gnd cell_6t
Xbit_r52_c39 bl[39] br[39] wl[52] vdd gnd cell_6t
Xbit_r53_c39 bl[39] br[39] wl[53] vdd gnd cell_6t
Xbit_r54_c39 bl[39] br[39] wl[54] vdd gnd cell_6t
Xbit_r55_c39 bl[39] br[39] wl[55] vdd gnd cell_6t
Xbit_r56_c39 bl[39] br[39] wl[56] vdd gnd cell_6t
Xbit_r57_c39 bl[39] br[39] wl[57] vdd gnd cell_6t
Xbit_r58_c39 bl[39] br[39] wl[58] vdd gnd cell_6t
Xbit_r59_c39 bl[39] br[39] wl[59] vdd gnd cell_6t
Xbit_r60_c39 bl[39] br[39] wl[60] vdd gnd cell_6t
Xbit_r61_c39 bl[39] br[39] wl[61] vdd gnd cell_6t
Xbit_r62_c39 bl[39] br[39] wl[62] vdd gnd cell_6t
Xbit_r63_c39 bl[39] br[39] wl[63] vdd gnd cell_6t
Xbit_r64_c39 bl[39] br[39] wl[64] vdd gnd cell_6t
Xbit_r65_c39 bl[39] br[39] wl[65] vdd gnd cell_6t
Xbit_r66_c39 bl[39] br[39] wl[66] vdd gnd cell_6t
Xbit_r67_c39 bl[39] br[39] wl[67] vdd gnd cell_6t
Xbit_r68_c39 bl[39] br[39] wl[68] vdd gnd cell_6t
Xbit_r69_c39 bl[39] br[39] wl[69] vdd gnd cell_6t
Xbit_r70_c39 bl[39] br[39] wl[70] vdd gnd cell_6t
Xbit_r71_c39 bl[39] br[39] wl[71] vdd gnd cell_6t
Xbit_r72_c39 bl[39] br[39] wl[72] vdd gnd cell_6t
Xbit_r73_c39 bl[39] br[39] wl[73] vdd gnd cell_6t
Xbit_r74_c39 bl[39] br[39] wl[74] vdd gnd cell_6t
Xbit_r75_c39 bl[39] br[39] wl[75] vdd gnd cell_6t
Xbit_r76_c39 bl[39] br[39] wl[76] vdd gnd cell_6t
Xbit_r77_c39 bl[39] br[39] wl[77] vdd gnd cell_6t
Xbit_r78_c39 bl[39] br[39] wl[78] vdd gnd cell_6t
Xbit_r79_c39 bl[39] br[39] wl[79] vdd gnd cell_6t
Xbit_r80_c39 bl[39] br[39] wl[80] vdd gnd cell_6t
Xbit_r81_c39 bl[39] br[39] wl[81] vdd gnd cell_6t
Xbit_r82_c39 bl[39] br[39] wl[82] vdd gnd cell_6t
Xbit_r83_c39 bl[39] br[39] wl[83] vdd gnd cell_6t
Xbit_r84_c39 bl[39] br[39] wl[84] vdd gnd cell_6t
Xbit_r85_c39 bl[39] br[39] wl[85] vdd gnd cell_6t
Xbit_r86_c39 bl[39] br[39] wl[86] vdd gnd cell_6t
Xbit_r87_c39 bl[39] br[39] wl[87] vdd gnd cell_6t
Xbit_r88_c39 bl[39] br[39] wl[88] vdd gnd cell_6t
Xbit_r89_c39 bl[39] br[39] wl[89] vdd gnd cell_6t
Xbit_r90_c39 bl[39] br[39] wl[90] vdd gnd cell_6t
Xbit_r91_c39 bl[39] br[39] wl[91] vdd gnd cell_6t
Xbit_r92_c39 bl[39] br[39] wl[92] vdd gnd cell_6t
Xbit_r93_c39 bl[39] br[39] wl[93] vdd gnd cell_6t
Xbit_r94_c39 bl[39] br[39] wl[94] vdd gnd cell_6t
Xbit_r95_c39 bl[39] br[39] wl[95] vdd gnd cell_6t
Xbit_r96_c39 bl[39] br[39] wl[96] vdd gnd cell_6t
Xbit_r97_c39 bl[39] br[39] wl[97] vdd gnd cell_6t
Xbit_r98_c39 bl[39] br[39] wl[98] vdd gnd cell_6t
Xbit_r99_c39 bl[39] br[39] wl[99] vdd gnd cell_6t
Xbit_r100_c39 bl[39] br[39] wl[100] vdd gnd cell_6t
Xbit_r101_c39 bl[39] br[39] wl[101] vdd gnd cell_6t
Xbit_r102_c39 bl[39] br[39] wl[102] vdd gnd cell_6t
Xbit_r103_c39 bl[39] br[39] wl[103] vdd gnd cell_6t
Xbit_r104_c39 bl[39] br[39] wl[104] vdd gnd cell_6t
Xbit_r105_c39 bl[39] br[39] wl[105] vdd gnd cell_6t
Xbit_r106_c39 bl[39] br[39] wl[106] vdd gnd cell_6t
Xbit_r107_c39 bl[39] br[39] wl[107] vdd gnd cell_6t
Xbit_r108_c39 bl[39] br[39] wl[108] vdd gnd cell_6t
Xbit_r109_c39 bl[39] br[39] wl[109] vdd gnd cell_6t
Xbit_r110_c39 bl[39] br[39] wl[110] vdd gnd cell_6t
Xbit_r111_c39 bl[39] br[39] wl[111] vdd gnd cell_6t
Xbit_r112_c39 bl[39] br[39] wl[112] vdd gnd cell_6t
Xbit_r113_c39 bl[39] br[39] wl[113] vdd gnd cell_6t
Xbit_r114_c39 bl[39] br[39] wl[114] vdd gnd cell_6t
Xbit_r115_c39 bl[39] br[39] wl[115] vdd gnd cell_6t
Xbit_r116_c39 bl[39] br[39] wl[116] vdd gnd cell_6t
Xbit_r117_c39 bl[39] br[39] wl[117] vdd gnd cell_6t
Xbit_r118_c39 bl[39] br[39] wl[118] vdd gnd cell_6t
Xbit_r119_c39 bl[39] br[39] wl[119] vdd gnd cell_6t
Xbit_r120_c39 bl[39] br[39] wl[120] vdd gnd cell_6t
Xbit_r121_c39 bl[39] br[39] wl[121] vdd gnd cell_6t
Xbit_r122_c39 bl[39] br[39] wl[122] vdd gnd cell_6t
Xbit_r123_c39 bl[39] br[39] wl[123] vdd gnd cell_6t
Xbit_r124_c39 bl[39] br[39] wl[124] vdd gnd cell_6t
Xbit_r125_c39 bl[39] br[39] wl[125] vdd gnd cell_6t
Xbit_r126_c39 bl[39] br[39] wl[126] vdd gnd cell_6t
Xbit_r127_c39 bl[39] br[39] wl[127] vdd gnd cell_6t
Xbit_r128_c39 bl[39] br[39] wl[128] vdd gnd cell_6t
Xbit_r129_c39 bl[39] br[39] wl[129] vdd gnd cell_6t
Xbit_r130_c39 bl[39] br[39] wl[130] vdd gnd cell_6t
Xbit_r131_c39 bl[39] br[39] wl[131] vdd gnd cell_6t
Xbit_r132_c39 bl[39] br[39] wl[132] vdd gnd cell_6t
Xbit_r133_c39 bl[39] br[39] wl[133] vdd gnd cell_6t
Xbit_r134_c39 bl[39] br[39] wl[134] vdd gnd cell_6t
Xbit_r135_c39 bl[39] br[39] wl[135] vdd gnd cell_6t
Xbit_r136_c39 bl[39] br[39] wl[136] vdd gnd cell_6t
Xbit_r137_c39 bl[39] br[39] wl[137] vdd gnd cell_6t
Xbit_r138_c39 bl[39] br[39] wl[138] vdd gnd cell_6t
Xbit_r139_c39 bl[39] br[39] wl[139] vdd gnd cell_6t
Xbit_r140_c39 bl[39] br[39] wl[140] vdd gnd cell_6t
Xbit_r141_c39 bl[39] br[39] wl[141] vdd gnd cell_6t
Xbit_r142_c39 bl[39] br[39] wl[142] vdd gnd cell_6t
Xbit_r143_c39 bl[39] br[39] wl[143] vdd gnd cell_6t
Xbit_r144_c39 bl[39] br[39] wl[144] vdd gnd cell_6t
Xbit_r145_c39 bl[39] br[39] wl[145] vdd gnd cell_6t
Xbit_r146_c39 bl[39] br[39] wl[146] vdd gnd cell_6t
Xbit_r147_c39 bl[39] br[39] wl[147] vdd gnd cell_6t
Xbit_r148_c39 bl[39] br[39] wl[148] vdd gnd cell_6t
Xbit_r149_c39 bl[39] br[39] wl[149] vdd gnd cell_6t
Xbit_r150_c39 bl[39] br[39] wl[150] vdd gnd cell_6t
Xbit_r151_c39 bl[39] br[39] wl[151] vdd gnd cell_6t
Xbit_r152_c39 bl[39] br[39] wl[152] vdd gnd cell_6t
Xbit_r153_c39 bl[39] br[39] wl[153] vdd gnd cell_6t
Xbit_r154_c39 bl[39] br[39] wl[154] vdd gnd cell_6t
Xbit_r155_c39 bl[39] br[39] wl[155] vdd gnd cell_6t
Xbit_r156_c39 bl[39] br[39] wl[156] vdd gnd cell_6t
Xbit_r157_c39 bl[39] br[39] wl[157] vdd gnd cell_6t
Xbit_r158_c39 bl[39] br[39] wl[158] vdd gnd cell_6t
Xbit_r159_c39 bl[39] br[39] wl[159] vdd gnd cell_6t
Xbit_r160_c39 bl[39] br[39] wl[160] vdd gnd cell_6t
Xbit_r161_c39 bl[39] br[39] wl[161] vdd gnd cell_6t
Xbit_r162_c39 bl[39] br[39] wl[162] vdd gnd cell_6t
Xbit_r163_c39 bl[39] br[39] wl[163] vdd gnd cell_6t
Xbit_r164_c39 bl[39] br[39] wl[164] vdd gnd cell_6t
Xbit_r165_c39 bl[39] br[39] wl[165] vdd gnd cell_6t
Xbit_r166_c39 bl[39] br[39] wl[166] vdd gnd cell_6t
Xbit_r167_c39 bl[39] br[39] wl[167] vdd gnd cell_6t
Xbit_r168_c39 bl[39] br[39] wl[168] vdd gnd cell_6t
Xbit_r169_c39 bl[39] br[39] wl[169] vdd gnd cell_6t
Xbit_r170_c39 bl[39] br[39] wl[170] vdd gnd cell_6t
Xbit_r171_c39 bl[39] br[39] wl[171] vdd gnd cell_6t
Xbit_r172_c39 bl[39] br[39] wl[172] vdd gnd cell_6t
Xbit_r173_c39 bl[39] br[39] wl[173] vdd gnd cell_6t
Xbit_r174_c39 bl[39] br[39] wl[174] vdd gnd cell_6t
Xbit_r175_c39 bl[39] br[39] wl[175] vdd gnd cell_6t
Xbit_r176_c39 bl[39] br[39] wl[176] vdd gnd cell_6t
Xbit_r177_c39 bl[39] br[39] wl[177] vdd gnd cell_6t
Xbit_r178_c39 bl[39] br[39] wl[178] vdd gnd cell_6t
Xbit_r179_c39 bl[39] br[39] wl[179] vdd gnd cell_6t
Xbit_r180_c39 bl[39] br[39] wl[180] vdd gnd cell_6t
Xbit_r181_c39 bl[39] br[39] wl[181] vdd gnd cell_6t
Xbit_r182_c39 bl[39] br[39] wl[182] vdd gnd cell_6t
Xbit_r183_c39 bl[39] br[39] wl[183] vdd gnd cell_6t
Xbit_r184_c39 bl[39] br[39] wl[184] vdd gnd cell_6t
Xbit_r185_c39 bl[39] br[39] wl[185] vdd gnd cell_6t
Xbit_r186_c39 bl[39] br[39] wl[186] vdd gnd cell_6t
Xbit_r187_c39 bl[39] br[39] wl[187] vdd gnd cell_6t
Xbit_r188_c39 bl[39] br[39] wl[188] vdd gnd cell_6t
Xbit_r189_c39 bl[39] br[39] wl[189] vdd gnd cell_6t
Xbit_r190_c39 bl[39] br[39] wl[190] vdd gnd cell_6t
Xbit_r191_c39 bl[39] br[39] wl[191] vdd gnd cell_6t
Xbit_r192_c39 bl[39] br[39] wl[192] vdd gnd cell_6t
Xbit_r193_c39 bl[39] br[39] wl[193] vdd gnd cell_6t
Xbit_r194_c39 bl[39] br[39] wl[194] vdd gnd cell_6t
Xbit_r195_c39 bl[39] br[39] wl[195] vdd gnd cell_6t
Xbit_r196_c39 bl[39] br[39] wl[196] vdd gnd cell_6t
Xbit_r197_c39 bl[39] br[39] wl[197] vdd gnd cell_6t
Xbit_r198_c39 bl[39] br[39] wl[198] vdd gnd cell_6t
Xbit_r199_c39 bl[39] br[39] wl[199] vdd gnd cell_6t
Xbit_r200_c39 bl[39] br[39] wl[200] vdd gnd cell_6t
Xbit_r201_c39 bl[39] br[39] wl[201] vdd gnd cell_6t
Xbit_r202_c39 bl[39] br[39] wl[202] vdd gnd cell_6t
Xbit_r203_c39 bl[39] br[39] wl[203] vdd gnd cell_6t
Xbit_r204_c39 bl[39] br[39] wl[204] vdd gnd cell_6t
Xbit_r205_c39 bl[39] br[39] wl[205] vdd gnd cell_6t
Xbit_r206_c39 bl[39] br[39] wl[206] vdd gnd cell_6t
Xbit_r207_c39 bl[39] br[39] wl[207] vdd gnd cell_6t
Xbit_r208_c39 bl[39] br[39] wl[208] vdd gnd cell_6t
Xbit_r209_c39 bl[39] br[39] wl[209] vdd gnd cell_6t
Xbit_r210_c39 bl[39] br[39] wl[210] vdd gnd cell_6t
Xbit_r211_c39 bl[39] br[39] wl[211] vdd gnd cell_6t
Xbit_r212_c39 bl[39] br[39] wl[212] vdd gnd cell_6t
Xbit_r213_c39 bl[39] br[39] wl[213] vdd gnd cell_6t
Xbit_r214_c39 bl[39] br[39] wl[214] vdd gnd cell_6t
Xbit_r215_c39 bl[39] br[39] wl[215] vdd gnd cell_6t
Xbit_r216_c39 bl[39] br[39] wl[216] vdd gnd cell_6t
Xbit_r217_c39 bl[39] br[39] wl[217] vdd gnd cell_6t
Xbit_r218_c39 bl[39] br[39] wl[218] vdd gnd cell_6t
Xbit_r219_c39 bl[39] br[39] wl[219] vdd gnd cell_6t
Xbit_r220_c39 bl[39] br[39] wl[220] vdd gnd cell_6t
Xbit_r221_c39 bl[39] br[39] wl[221] vdd gnd cell_6t
Xbit_r222_c39 bl[39] br[39] wl[222] vdd gnd cell_6t
Xbit_r223_c39 bl[39] br[39] wl[223] vdd gnd cell_6t
Xbit_r224_c39 bl[39] br[39] wl[224] vdd gnd cell_6t
Xbit_r225_c39 bl[39] br[39] wl[225] vdd gnd cell_6t
Xbit_r226_c39 bl[39] br[39] wl[226] vdd gnd cell_6t
Xbit_r227_c39 bl[39] br[39] wl[227] vdd gnd cell_6t
Xbit_r228_c39 bl[39] br[39] wl[228] vdd gnd cell_6t
Xbit_r229_c39 bl[39] br[39] wl[229] vdd gnd cell_6t
Xbit_r230_c39 bl[39] br[39] wl[230] vdd gnd cell_6t
Xbit_r231_c39 bl[39] br[39] wl[231] vdd gnd cell_6t
Xbit_r232_c39 bl[39] br[39] wl[232] vdd gnd cell_6t
Xbit_r233_c39 bl[39] br[39] wl[233] vdd gnd cell_6t
Xbit_r234_c39 bl[39] br[39] wl[234] vdd gnd cell_6t
Xbit_r235_c39 bl[39] br[39] wl[235] vdd gnd cell_6t
Xbit_r236_c39 bl[39] br[39] wl[236] vdd gnd cell_6t
Xbit_r237_c39 bl[39] br[39] wl[237] vdd gnd cell_6t
Xbit_r238_c39 bl[39] br[39] wl[238] vdd gnd cell_6t
Xbit_r239_c39 bl[39] br[39] wl[239] vdd gnd cell_6t
Xbit_r240_c39 bl[39] br[39] wl[240] vdd gnd cell_6t
Xbit_r241_c39 bl[39] br[39] wl[241] vdd gnd cell_6t
Xbit_r242_c39 bl[39] br[39] wl[242] vdd gnd cell_6t
Xbit_r243_c39 bl[39] br[39] wl[243] vdd gnd cell_6t
Xbit_r244_c39 bl[39] br[39] wl[244] vdd gnd cell_6t
Xbit_r245_c39 bl[39] br[39] wl[245] vdd gnd cell_6t
Xbit_r246_c39 bl[39] br[39] wl[246] vdd gnd cell_6t
Xbit_r247_c39 bl[39] br[39] wl[247] vdd gnd cell_6t
Xbit_r248_c39 bl[39] br[39] wl[248] vdd gnd cell_6t
Xbit_r249_c39 bl[39] br[39] wl[249] vdd gnd cell_6t
Xbit_r250_c39 bl[39] br[39] wl[250] vdd gnd cell_6t
Xbit_r251_c39 bl[39] br[39] wl[251] vdd gnd cell_6t
Xbit_r252_c39 bl[39] br[39] wl[252] vdd gnd cell_6t
Xbit_r253_c39 bl[39] br[39] wl[253] vdd gnd cell_6t
Xbit_r254_c39 bl[39] br[39] wl[254] vdd gnd cell_6t
Xbit_r255_c39 bl[39] br[39] wl[255] vdd gnd cell_6t
Xbit_r0_c40 bl[40] br[40] wl[0] vdd gnd cell_6t
Xbit_r1_c40 bl[40] br[40] wl[1] vdd gnd cell_6t
Xbit_r2_c40 bl[40] br[40] wl[2] vdd gnd cell_6t
Xbit_r3_c40 bl[40] br[40] wl[3] vdd gnd cell_6t
Xbit_r4_c40 bl[40] br[40] wl[4] vdd gnd cell_6t
Xbit_r5_c40 bl[40] br[40] wl[5] vdd gnd cell_6t
Xbit_r6_c40 bl[40] br[40] wl[6] vdd gnd cell_6t
Xbit_r7_c40 bl[40] br[40] wl[7] vdd gnd cell_6t
Xbit_r8_c40 bl[40] br[40] wl[8] vdd gnd cell_6t
Xbit_r9_c40 bl[40] br[40] wl[9] vdd gnd cell_6t
Xbit_r10_c40 bl[40] br[40] wl[10] vdd gnd cell_6t
Xbit_r11_c40 bl[40] br[40] wl[11] vdd gnd cell_6t
Xbit_r12_c40 bl[40] br[40] wl[12] vdd gnd cell_6t
Xbit_r13_c40 bl[40] br[40] wl[13] vdd gnd cell_6t
Xbit_r14_c40 bl[40] br[40] wl[14] vdd gnd cell_6t
Xbit_r15_c40 bl[40] br[40] wl[15] vdd gnd cell_6t
Xbit_r16_c40 bl[40] br[40] wl[16] vdd gnd cell_6t
Xbit_r17_c40 bl[40] br[40] wl[17] vdd gnd cell_6t
Xbit_r18_c40 bl[40] br[40] wl[18] vdd gnd cell_6t
Xbit_r19_c40 bl[40] br[40] wl[19] vdd gnd cell_6t
Xbit_r20_c40 bl[40] br[40] wl[20] vdd gnd cell_6t
Xbit_r21_c40 bl[40] br[40] wl[21] vdd gnd cell_6t
Xbit_r22_c40 bl[40] br[40] wl[22] vdd gnd cell_6t
Xbit_r23_c40 bl[40] br[40] wl[23] vdd gnd cell_6t
Xbit_r24_c40 bl[40] br[40] wl[24] vdd gnd cell_6t
Xbit_r25_c40 bl[40] br[40] wl[25] vdd gnd cell_6t
Xbit_r26_c40 bl[40] br[40] wl[26] vdd gnd cell_6t
Xbit_r27_c40 bl[40] br[40] wl[27] vdd gnd cell_6t
Xbit_r28_c40 bl[40] br[40] wl[28] vdd gnd cell_6t
Xbit_r29_c40 bl[40] br[40] wl[29] vdd gnd cell_6t
Xbit_r30_c40 bl[40] br[40] wl[30] vdd gnd cell_6t
Xbit_r31_c40 bl[40] br[40] wl[31] vdd gnd cell_6t
Xbit_r32_c40 bl[40] br[40] wl[32] vdd gnd cell_6t
Xbit_r33_c40 bl[40] br[40] wl[33] vdd gnd cell_6t
Xbit_r34_c40 bl[40] br[40] wl[34] vdd gnd cell_6t
Xbit_r35_c40 bl[40] br[40] wl[35] vdd gnd cell_6t
Xbit_r36_c40 bl[40] br[40] wl[36] vdd gnd cell_6t
Xbit_r37_c40 bl[40] br[40] wl[37] vdd gnd cell_6t
Xbit_r38_c40 bl[40] br[40] wl[38] vdd gnd cell_6t
Xbit_r39_c40 bl[40] br[40] wl[39] vdd gnd cell_6t
Xbit_r40_c40 bl[40] br[40] wl[40] vdd gnd cell_6t
Xbit_r41_c40 bl[40] br[40] wl[41] vdd gnd cell_6t
Xbit_r42_c40 bl[40] br[40] wl[42] vdd gnd cell_6t
Xbit_r43_c40 bl[40] br[40] wl[43] vdd gnd cell_6t
Xbit_r44_c40 bl[40] br[40] wl[44] vdd gnd cell_6t
Xbit_r45_c40 bl[40] br[40] wl[45] vdd gnd cell_6t
Xbit_r46_c40 bl[40] br[40] wl[46] vdd gnd cell_6t
Xbit_r47_c40 bl[40] br[40] wl[47] vdd gnd cell_6t
Xbit_r48_c40 bl[40] br[40] wl[48] vdd gnd cell_6t
Xbit_r49_c40 bl[40] br[40] wl[49] vdd gnd cell_6t
Xbit_r50_c40 bl[40] br[40] wl[50] vdd gnd cell_6t
Xbit_r51_c40 bl[40] br[40] wl[51] vdd gnd cell_6t
Xbit_r52_c40 bl[40] br[40] wl[52] vdd gnd cell_6t
Xbit_r53_c40 bl[40] br[40] wl[53] vdd gnd cell_6t
Xbit_r54_c40 bl[40] br[40] wl[54] vdd gnd cell_6t
Xbit_r55_c40 bl[40] br[40] wl[55] vdd gnd cell_6t
Xbit_r56_c40 bl[40] br[40] wl[56] vdd gnd cell_6t
Xbit_r57_c40 bl[40] br[40] wl[57] vdd gnd cell_6t
Xbit_r58_c40 bl[40] br[40] wl[58] vdd gnd cell_6t
Xbit_r59_c40 bl[40] br[40] wl[59] vdd gnd cell_6t
Xbit_r60_c40 bl[40] br[40] wl[60] vdd gnd cell_6t
Xbit_r61_c40 bl[40] br[40] wl[61] vdd gnd cell_6t
Xbit_r62_c40 bl[40] br[40] wl[62] vdd gnd cell_6t
Xbit_r63_c40 bl[40] br[40] wl[63] vdd gnd cell_6t
Xbit_r64_c40 bl[40] br[40] wl[64] vdd gnd cell_6t
Xbit_r65_c40 bl[40] br[40] wl[65] vdd gnd cell_6t
Xbit_r66_c40 bl[40] br[40] wl[66] vdd gnd cell_6t
Xbit_r67_c40 bl[40] br[40] wl[67] vdd gnd cell_6t
Xbit_r68_c40 bl[40] br[40] wl[68] vdd gnd cell_6t
Xbit_r69_c40 bl[40] br[40] wl[69] vdd gnd cell_6t
Xbit_r70_c40 bl[40] br[40] wl[70] vdd gnd cell_6t
Xbit_r71_c40 bl[40] br[40] wl[71] vdd gnd cell_6t
Xbit_r72_c40 bl[40] br[40] wl[72] vdd gnd cell_6t
Xbit_r73_c40 bl[40] br[40] wl[73] vdd gnd cell_6t
Xbit_r74_c40 bl[40] br[40] wl[74] vdd gnd cell_6t
Xbit_r75_c40 bl[40] br[40] wl[75] vdd gnd cell_6t
Xbit_r76_c40 bl[40] br[40] wl[76] vdd gnd cell_6t
Xbit_r77_c40 bl[40] br[40] wl[77] vdd gnd cell_6t
Xbit_r78_c40 bl[40] br[40] wl[78] vdd gnd cell_6t
Xbit_r79_c40 bl[40] br[40] wl[79] vdd gnd cell_6t
Xbit_r80_c40 bl[40] br[40] wl[80] vdd gnd cell_6t
Xbit_r81_c40 bl[40] br[40] wl[81] vdd gnd cell_6t
Xbit_r82_c40 bl[40] br[40] wl[82] vdd gnd cell_6t
Xbit_r83_c40 bl[40] br[40] wl[83] vdd gnd cell_6t
Xbit_r84_c40 bl[40] br[40] wl[84] vdd gnd cell_6t
Xbit_r85_c40 bl[40] br[40] wl[85] vdd gnd cell_6t
Xbit_r86_c40 bl[40] br[40] wl[86] vdd gnd cell_6t
Xbit_r87_c40 bl[40] br[40] wl[87] vdd gnd cell_6t
Xbit_r88_c40 bl[40] br[40] wl[88] vdd gnd cell_6t
Xbit_r89_c40 bl[40] br[40] wl[89] vdd gnd cell_6t
Xbit_r90_c40 bl[40] br[40] wl[90] vdd gnd cell_6t
Xbit_r91_c40 bl[40] br[40] wl[91] vdd gnd cell_6t
Xbit_r92_c40 bl[40] br[40] wl[92] vdd gnd cell_6t
Xbit_r93_c40 bl[40] br[40] wl[93] vdd gnd cell_6t
Xbit_r94_c40 bl[40] br[40] wl[94] vdd gnd cell_6t
Xbit_r95_c40 bl[40] br[40] wl[95] vdd gnd cell_6t
Xbit_r96_c40 bl[40] br[40] wl[96] vdd gnd cell_6t
Xbit_r97_c40 bl[40] br[40] wl[97] vdd gnd cell_6t
Xbit_r98_c40 bl[40] br[40] wl[98] vdd gnd cell_6t
Xbit_r99_c40 bl[40] br[40] wl[99] vdd gnd cell_6t
Xbit_r100_c40 bl[40] br[40] wl[100] vdd gnd cell_6t
Xbit_r101_c40 bl[40] br[40] wl[101] vdd gnd cell_6t
Xbit_r102_c40 bl[40] br[40] wl[102] vdd gnd cell_6t
Xbit_r103_c40 bl[40] br[40] wl[103] vdd gnd cell_6t
Xbit_r104_c40 bl[40] br[40] wl[104] vdd gnd cell_6t
Xbit_r105_c40 bl[40] br[40] wl[105] vdd gnd cell_6t
Xbit_r106_c40 bl[40] br[40] wl[106] vdd gnd cell_6t
Xbit_r107_c40 bl[40] br[40] wl[107] vdd gnd cell_6t
Xbit_r108_c40 bl[40] br[40] wl[108] vdd gnd cell_6t
Xbit_r109_c40 bl[40] br[40] wl[109] vdd gnd cell_6t
Xbit_r110_c40 bl[40] br[40] wl[110] vdd gnd cell_6t
Xbit_r111_c40 bl[40] br[40] wl[111] vdd gnd cell_6t
Xbit_r112_c40 bl[40] br[40] wl[112] vdd gnd cell_6t
Xbit_r113_c40 bl[40] br[40] wl[113] vdd gnd cell_6t
Xbit_r114_c40 bl[40] br[40] wl[114] vdd gnd cell_6t
Xbit_r115_c40 bl[40] br[40] wl[115] vdd gnd cell_6t
Xbit_r116_c40 bl[40] br[40] wl[116] vdd gnd cell_6t
Xbit_r117_c40 bl[40] br[40] wl[117] vdd gnd cell_6t
Xbit_r118_c40 bl[40] br[40] wl[118] vdd gnd cell_6t
Xbit_r119_c40 bl[40] br[40] wl[119] vdd gnd cell_6t
Xbit_r120_c40 bl[40] br[40] wl[120] vdd gnd cell_6t
Xbit_r121_c40 bl[40] br[40] wl[121] vdd gnd cell_6t
Xbit_r122_c40 bl[40] br[40] wl[122] vdd gnd cell_6t
Xbit_r123_c40 bl[40] br[40] wl[123] vdd gnd cell_6t
Xbit_r124_c40 bl[40] br[40] wl[124] vdd gnd cell_6t
Xbit_r125_c40 bl[40] br[40] wl[125] vdd gnd cell_6t
Xbit_r126_c40 bl[40] br[40] wl[126] vdd gnd cell_6t
Xbit_r127_c40 bl[40] br[40] wl[127] vdd gnd cell_6t
Xbit_r128_c40 bl[40] br[40] wl[128] vdd gnd cell_6t
Xbit_r129_c40 bl[40] br[40] wl[129] vdd gnd cell_6t
Xbit_r130_c40 bl[40] br[40] wl[130] vdd gnd cell_6t
Xbit_r131_c40 bl[40] br[40] wl[131] vdd gnd cell_6t
Xbit_r132_c40 bl[40] br[40] wl[132] vdd gnd cell_6t
Xbit_r133_c40 bl[40] br[40] wl[133] vdd gnd cell_6t
Xbit_r134_c40 bl[40] br[40] wl[134] vdd gnd cell_6t
Xbit_r135_c40 bl[40] br[40] wl[135] vdd gnd cell_6t
Xbit_r136_c40 bl[40] br[40] wl[136] vdd gnd cell_6t
Xbit_r137_c40 bl[40] br[40] wl[137] vdd gnd cell_6t
Xbit_r138_c40 bl[40] br[40] wl[138] vdd gnd cell_6t
Xbit_r139_c40 bl[40] br[40] wl[139] vdd gnd cell_6t
Xbit_r140_c40 bl[40] br[40] wl[140] vdd gnd cell_6t
Xbit_r141_c40 bl[40] br[40] wl[141] vdd gnd cell_6t
Xbit_r142_c40 bl[40] br[40] wl[142] vdd gnd cell_6t
Xbit_r143_c40 bl[40] br[40] wl[143] vdd gnd cell_6t
Xbit_r144_c40 bl[40] br[40] wl[144] vdd gnd cell_6t
Xbit_r145_c40 bl[40] br[40] wl[145] vdd gnd cell_6t
Xbit_r146_c40 bl[40] br[40] wl[146] vdd gnd cell_6t
Xbit_r147_c40 bl[40] br[40] wl[147] vdd gnd cell_6t
Xbit_r148_c40 bl[40] br[40] wl[148] vdd gnd cell_6t
Xbit_r149_c40 bl[40] br[40] wl[149] vdd gnd cell_6t
Xbit_r150_c40 bl[40] br[40] wl[150] vdd gnd cell_6t
Xbit_r151_c40 bl[40] br[40] wl[151] vdd gnd cell_6t
Xbit_r152_c40 bl[40] br[40] wl[152] vdd gnd cell_6t
Xbit_r153_c40 bl[40] br[40] wl[153] vdd gnd cell_6t
Xbit_r154_c40 bl[40] br[40] wl[154] vdd gnd cell_6t
Xbit_r155_c40 bl[40] br[40] wl[155] vdd gnd cell_6t
Xbit_r156_c40 bl[40] br[40] wl[156] vdd gnd cell_6t
Xbit_r157_c40 bl[40] br[40] wl[157] vdd gnd cell_6t
Xbit_r158_c40 bl[40] br[40] wl[158] vdd gnd cell_6t
Xbit_r159_c40 bl[40] br[40] wl[159] vdd gnd cell_6t
Xbit_r160_c40 bl[40] br[40] wl[160] vdd gnd cell_6t
Xbit_r161_c40 bl[40] br[40] wl[161] vdd gnd cell_6t
Xbit_r162_c40 bl[40] br[40] wl[162] vdd gnd cell_6t
Xbit_r163_c40 bl[40] br[40] wl[163] vdd gnd cell_6t
Xbit_r164_c40 bl[40] br[40] wl[164] vdd gnd cell_6t
Xbit_r165_c40 bl[40] br[40] wl[165] vdd gnd cell_6t
Xbit_r166_c40 bl[40] br[40] wl[166] vdd gnd cell_6t
Xbit_r167_c40 bl[40] br[40] wl[167] vdd gnd cell_6t
Xbit_r168_c40 bl[40] br[40] wl[168] vdd gnd cell_6t
Xbit_r169_c40 bl[40] br[40] wl[169] vdd gnd cell_6t
Xbit_r170_c40 bl[40] br[40] wl[170] vdd gnd cell_6t
Xbit_r171_c40 bl[40] br[40] wl[171] vdd gnd cell_6t
Xbit_r172_c40 bl[40] br[40] wl[172] vdd gnd cell_6t
Xbit_r173_c40 bl[40] br[40] wl[173] vdd gnd cell_6t
Xbit_r174_c40 bl[40] br[40] wl[174] vdd gnd cell_6t
Xbit_r175_c40 bl[40] br[40] wl[175] vdd gnd cell_6t
Xbit_r176_c40 bl[40] br[40] wl[176] vdd gnd cell_6t
Xbit_r177_c40 bl[40] br[40] wl[177] vdd gnd cell_6t
Xbit_r178_c40 bl[40] br[40] wl[178] vdd gnd cell_6t
Xbit_r179_c40 bl[40] br[40] wl[179] vdd gnd cell_6t
Xbit_r180_c40 bl[40] br[40] wl[180] vdd gnd cell_6t
Xbit_r181_c40 bl[40] br[40] wl[181] vdd gnd cell_6t
Xbit_r182_c40 bl[40] br[40] wl[182] vdd gnd cell_6t
Xbit_r183_c40 bl[40] br[40] wl[183] vdd gnd cell_6t
Xbit_r184_c40 bl[40] br[40] wl[184] vdd gnd cell_6t
Xbit_r185_c40 bl[40] br[40] wl[185] vdd gnd cell_6t
Xbit_r186_c40 bl[40] br[40] wl[186] vdd gnd cell_6t
Xbit_r187_c40 bl[40] br[40] wl[187] vdd gnd cell_6t
Xbit_r188_c40 bl[40] br[40] wl[188] vdd gnd cell_6t
Xbit_r189_c40 bl[40] br[40] wl[189] vdd gnd cell_6t
Xbit_r190_c40 bl[40] br[40] wl[190] vdd gnd cell_6t
Xbit_r191_c40 bl[40] br[40] wl[191] vdd gnd cell_6t
Xbit_r192_c40 bl[40] br[40] wl[192] vdd gnd cell_6t
Xbit_r193_c40 bl[40] br[40] wl[193] vdd gnd cell_6t
Xbit_r194_c40 bl[40] br[40] wl[194] vdd gnd cell_6t
Xbit_r195_c40 bl[40] br[40] wl[195] vdd gnd cell_6t
Xbit_r196_c40 bl[40] br[40] wl[196] vdd gnd cell_6t
Xbit_r197_c40 bl[40] br[40] wl[197] vdd gnd cell_6t
Xbit_r198_c40 bl[40] br[40] wl[198] vdd gnd cell_6t
Xbit_r199_c40 bl[40] br[40] wl[199] vdd gnd cell_6t
Xbit_r200_c40 bl[40] br[40] wl[200] vdd gnd cell_6t
Xbit_r201_c40 bl[40] br[40] wl[201] vdd gnd cell_6t
Xbit_r202_c40 bl[40] br[40] wl[202] vdd gnd cell_6t
Xbit_r203_c40 bl[40] br[40] wl[203] vdd gnd cell_6t
Xbit_r204_c40 bl[40] br[40] wl[204] vdd gnd cell_6t
Xbit_r205_c40 bl[40] br[40] wl[205] vdd gnd cell_6t
Xbit_r206_c40 bl[40] br[40] wl[206] vdd gnd cell_6t
Xbit_r207_c40 bl[40] br[40] wl[207] vdd gnd cell_6t
Xbit_r208_c40 bl[40] br[40] wl[208] vdd gnd cell_6t
Xbit_r209_c40 bl[40] br[40] wl[209] vdd gnd cell_6t
Xbit_r210_c40 bl[40] br[40] wl[210] vdd gnd cell_6t
Xbit_r211_c40 bl[40] br[40] wl[211] vdd gnd cell_6t
Xbit_r212_c40 bl[40] br[40] wl[212] vdd gnd cell_6t
Xbit_r213_c40 bl[40] br[40] wl[213] vdd gnd cell_6t
Xbit_r214_c40 bl[40] br[40] wl[214] vdd gnd cell_6t
Xbit_r215_c40 bl[40] br[40] wl[215] vdd gnd cell_6t
Xbit_r216_c40 bl[40] br[40] wl[216] vdd gnd cell_6t
Xbit_r217_c40 bl[40] br[40] wl[217] vdd gnd cell_6t
Xbit_r218_c40 bl[40] br[40] wl[218] vdd gnd cell_6t
Xbit_r219_c40 bl[40] br[40] wl[219] vdd gnd cell_6t
Xbit_r220_c40 bl[40] br[40] wl[220] vdd gnd cell_6t
Xbit_r221_c40 bl[40] br[40] wl[221] vdd gnd cell_6t
Xbit_r222_c40 bl[40] br[40] wl[222] vdd gnd cell_6t
Xbit_r223_c40 bl[40] br[40] wl[223] vdd gnd cell_6t
Xbit_r224_c40 bl[40] br[40] wl[224] vdd gnd cell_6t
Xbit_r225_c40 bl[40] br[40] wl[225] vdd gnd cell_6t
Xbit_r226_c40 bl[40] br[40] wl[226] vdd gnd cell_6t
Xbit_r227_c40 bl[40] br[40] wl[227] vdd gnd cell_6t
Xbit_r228_c40 bl[40] br[40] wl[228] vdd gnd cell_6t
Xbit_r229_c40 bl[40] br[40] wl[229] vdd gnd cell_6t
Xbit_r230_c40 bl[40] br[40] wl[230] vdd gnd cell_6t
Xbit_r231_c40 bl[40] br[40] wl[231] vdd gnd cell_6t
Xbit_r232_c40 bl[40] br[40] wl[232] vdd gnd cell_6t
Xbit_r233_c40 bl[40] br[40] wl[233] vdd gnd cell_6t
Xbit_r234_c40 bl[40] br[40] wl[234] vdd gnd cell_6t
Xbit_r235_c40 bl[40] br[40] wl[235] vdd gnd cell_6t
Xbit_r236_c40 bl[40] br[40] wl[236] vdd gnd cell_6t
Xbit_r237_c40 bl[40] br[40] wl[237] vdd gnd cell_6t
Xbit_r238_c40 bl[40] br[40] wl[238] vdd gnd cell_6t
Xbit_r239_c40 bl[40] br[40] wl[239] vdd gnd cell_6t
Xbit_r240_c40 bl[40] br[40] wl[240] vdd gnd cell_6t
Xbit_r241_c40 bl[40] br[40] wl[241] vdd gnd cell_6t
Xbit_r242_c40 bl[40] br[40] wl[242] vdd gnd cell_6t
Xbit_r243_c40 bl[40] br[40] wl[243] vdd gnd cell_6t
Xbit_r244_c40 bl[40] br[40] wl[244] vdd gnd cell_6t
Xbit_r245_c40 bl[40] br[40] wl[245] vdd gnd cell_6t
Xbit_r246_c40 bl[40] br[40] wl[246] vdd gnd cell_6t
Xbit_r247_c40 bl[40] br[40] wl[247] vdd gnd cell_6t
Xbit_r248_c40 bl[40] br[40] wl[248] vdd gnd cell_6t
Xbit_r249_c40 bl[40] br[40] wl[249] vdd gnd cell_6t
Xbit_r250_c40 bl[40] br[40] wl[250] vdd gnd cell_6t
Xbit_r251_c40 bl[40] br[40] wl[251] vdd gnd cell_6t
Xbit_r252_c40 bl[40] br[40] wl[252] vdd gnd cell_6t
Xbit_r253_c40 bl[40] br[40] wl[253] vdd gnd cell_6t
Xbit_r254_c40 bl[40] br[40] wl[254] vdd gnd cell_6t
Xbit_r255_c40 bl[40] br[40] wl[255] vdd gnd cell_6t
Xbit_r0_c41 bl[41] br[41] wl[0] vdd gnd cell_6t
Xbit_r1_c41 bl[41] br[41] wl[1] vdd gnd cell_6t
Xbit_r2_c41 bl[41] br[41] wl[2] vdd gnd cell_6t
Xbit_r3_c41 bl[41] br[41] wl[3] vdd gnd cell_6t
Xbit_r4_c41 bl[41] br[41] wl[4] vdd gnd cell_6t
Xbit_r5_c41 bl[41] br[41] wl[5] vdd gnd cell_6t
Xbit_r6_c41 bl[41] br[41] wl[6] vdd gnd cell_6t
Xbit_r7_c41 bl[41] br[41] wl[7] vdd gnd cell_6t
Xbit_r8_c41 bl[41] br[41] wl[8] vdd gnd cell_6t
Xbit_r9_c41 bl[41] br[41] wl[9] vdd gnd cell_6t
Xbit_r10_c41 bl[41] br[41] wl[10] vdd gnd cell_6t
Xbit_r11_c41 bl[41] br[41] wl[11] vdd gnd cell_6t
Xbit_r12_c41 bl[41] br[41] wl[12] vdd gnd cell_6t
Xbit_r13_c41 bl[41] br[41] wl[13] vdd gnd cell_6t
Xbit_r14_c41 bl[41] br[41] wl[14] vdd gnd cell_6t
Xbit_r15_c41 bl[41] br[41] wl[15] vdd gnd cell_6t
Xbit_r16_c41 bl[41] br[41] wl[16] vdd gnd cell_6t
Xbit_r17_c41 bl[41] br[41] wl[17] vdd gnd cell_6t
Xbit_r18_c41 bl[41] br[41] wl[18] vdd gnd cell_6t
Xbit_r19_c41 bl[41] br[41] wl[19] vdd gnd cell_6t
Xbit_r20_c41 bl[41] br[41] wl[20] vdd gnd cell_6t
Xbit_r21_c41 bl[41] br[41] wl[21] vdd gnd cell_6t
Xbit_r22_c41 bl[41] br[41] wl[22] vdd gnd cell_6t
Xbit_r23_c41 bl[41] br[41] wl[23] vdd gnd cell_6t
Xbit_r24_c41 bl[41] br[41] wl[24] vdd gnd cell_6t
Xbit_r25_c41 bl[41] br[41] wl[25] vdd gnd cell_6t
Xbit_r26_c41 bl[41] br[41] wl[26] vdd gnd cell_6t
Xbit_r27_c41 bl[41] br[41] wl[27] vdd gnd cell_6t
Xbit_r28_c41 bl[41] br[41] wl[28] vdd gnd cell_6t
Xbit_r29_c41 bl[41] br[41] wl[29] vdd gnd cell_6t
Xbit_r30_c41 bl[41] br[41] wl[30] vdd gnd cell_6t
Xbit_r31_c41 bl[41] br[41] wl[31] vdd gnd cell_6t
Xbit_r32_c41 bl[41] br[41] wl[32] vdd gnd cell_6t
Xbit_r33_c41 bl[41] br[41] wl[33] vdd gnd cell_6t
Xbit_r34_c41 bl[41] br[41] wl[34] vdd gnd cell_6t
Xbit_r35_c41 bl[41] br[41] wl[35] vdd gnd cell_6t
Xbit_r36_c41 bl[41] br[41] wl[36] vdd gnd cell_6t
Xbit_r37_c41 bl[41] br[41] wl[37] vdd gnd cell_6t
Xbit_r38_c41 bl[41] br[41] wl[38] vdd gnd cell_6t
Xbit_r39_c41 bl[41] br[41] wl[39] vdd gnd cell_6t
Xbit_r40_c41 bl[41] br[41] wl[40] vdd gnd cell_6t
Xbit_r41_c41 bl[41] br[41] wl[41] vdd gnd cell_6t
Xbit_r42_c41 bl[41] br[41] wl[42] vdd gnd cell_6t
Xbit_r43_c41 bl[41] br[41] wl[43] vdd gnd cell_6t
Xbit_r44_c41 bl[41] br[41] wl[44] vdd gnd cell_6t
Xbit_r45_c41 bl[41] br[41] wl[45] vdd gnd cell_6t
Xbit_r46_c41 bl[41] br[41] wl[46] vdd gnd cell_6t
Xbit_r47_c41 bl[41] br[41] wl[47] vdd gnd cell_6t
Xbit_r48_c41 bl[41] br[41] wl[48] vdd gnd cell_6t
Xbit_r49_c41 bl[41] br[41] wl[49] vdd gnd cell_6t
Xbit_r50_c41 bl[41] br[41] wl[50] vdd gnd cell_6t
Xbit_r51_c41 bl[41] br[41] wl[51] vdd gnd cell_6t
Xbit_r52_c41 bl[41] br[41] wl[52] vdd gnd cell_6t
Xbit_r53_c41 bl[41] br[41] wl[53] vdd gnd cell_6t
Xbit_r54_c41 bl[41] br[41] wl[54] vdd gnd cell_6t
Xbit_r55_c41 bl[41] br[41] wl[55] vdd gnd cell_6t
Xbit_r56_c41 bl[41] br[41] wl[56] vdd gnd cell_6t
Xbit_r57_c41 bl[41] br[41] wl[57] vdd gnd cell_6t
Xbit_r58_c41 bl[41] br[41] wl[58] vdd gnd cell_6t
Xbit_r59_c41 bl[41] br[41] wl[59] vdd gnd cell_6t
Xbit_r60_c41 bl[41] br[41] wl[60] vdd gnd cell_6t
Xbit_r61_c41 bl[41] br[41] wl[61] vdd gnd cell_6t
Xbit_r62_c41 bl[41] br[41] wl[62] vdd gnd cell_6t
Xbit_r63_c41 bl[41] br[41] wl[63] vdd gnd cell_6t
Xbit_r64_c41 bl[41] br[41] wl[64] vdd gnd cell_6t
Xbit_r65_c41 bl[41] br[41] wl[65] vdd gnd cell_6t
Xbit_r66_c41 bl[41] br[41] wl[66] vdd gnd cell_6t
Xbit_r67_c41 bl[41] br[41] wl[67] vdd gnd cell_6t
Xbit_r68_c41 bl[41] br[41] wl[68] vdd gnd cell_6t
Xbit_r69_c41 bl[41] br[41] wl[69] vdd gnd cell_6t
Xbit_r70_c41 bl[41] br[41] wl[70] vdd gnd cell_6t
Xbit_r71_c41 bl[41] br[41] wl[71] vdd gnd cell_6t
Xbit_r72_c41 bl[41] br[41] wl[72] vdd gnd cell_6t
Xbit_r73_c41 bl[41] br[41] wl[73] vdd gnd cell_6t
Xbit_r74_c41 bl[41] br[41] wl[74] vdd gnd cell_6t
Xbit_r75_c41 bl[41] br[41] wl[75] vdd gnd cell_6t
Xbit_r76_c41 bl[41] br[41] wl[76] vdd gnd cell_6t
Xbit_r77_c41 bl[41] br[41] wl[77] vdd gnd cell_6t
Xbit_r78_c41 bl[41] br[41] wl[78] vdd gnd cell_6t
Xbit_r79_c41 bl[41] br[41] wl[79] vdd gnd cell_6t
Xbit_r80_c41 bl[41] br[41] wl[80] vdd gnd cell_6t
Xbit_r81_c41 bl[41] br[41] wl[81] vdd gnd cell_6t
Xbit_r82_c41 bl[41] br[41] wl[82] vdd gnd cell_6t
Xbit_r83_c41 bl[41] br[41] wl[83] vdd gnd cell_6t
Xbit_r84_c41 bl[41] br[41] wl[84] vdd gnd cell_6t
Xbit_r85_c41 bl[41] br[41] wl[85] vdd gnd cell_6t
Xbit_r86_c41 bl[41] br[41] wl[86] vdd gnd cell_6t
Xbit_r87_c41 bl[41] br[41] wl[87] vdd gnd cell_6t
Xbit_r88_c41 bl[41] br[41] wl[88] vdd gnd cell_6t
Xbit_r89_c41 bl[41] br[41] wl[89] vdd gnd cell_6t
Xbit_r90_c41 bl[41] br[41] wl[90] vdd gnd cell_6t
Xbit_r91_c41 bl[41] br[41] wl[91] vdd gnd cell_6t
Xbit_r92_c41 bl[41] br[41] wl[92] vdd gnd cell_6t
Xbit_r93_c41 bl[41] br[41] wl[93] vdd gnd cell_6t
Xbit_r94_c41 bl[41] br[41] wl[94] vdd gnd cell_6t
Xbit_r95_c41 bl[41] br[41] wl[95] vdd gnd cell_6t
Xbit_r96_c41 bl[41] br[41] wl[96] vdd gnd cell_6t
Xbit_r97_c41 bl[41] br[41] wl[97] vdd gnd cell_6t
Xbit_r98_c41 bl[41] br[41] wl[98] vdd gnd cell_6t
Xbit_r99_c41 bl[41] br[41] wl[99] vdd gnd cell_6t
Xbit_r100_c41 bl[41] br[41] wl[100] vdd gnd cell_6t
Xbit_r101_c41 bl[41] br[41] wl[101] vdd gnd cell_6t
Xbit_r102_c41 bl[41] br[41] wl[102] vdd gnd cell_6t
Xbit_r103_c41 bl[41] br[41] wl[103] vdd gnd cell_6t
Xbit_r104_c41 bl[41] br[41] wl[104] vdd gnd cell_6t
Xbit_r105_c41 bl[41] br[41] wl[105] vdd gnd cell_6t
Xbit_r106_c41 bl[41] br[41] wl[106] vdd gnd cell_6t
Xbit_r107_c41 bl[41] br[41] wl[107] vdd gnd cell_6t
Xbit_r108_c41 bl[41] br[41] wl[108] vdd gnd cell_6t
Xbit_r109_c41 bl[41] br[41] wl[109] vdd gnd cell_6t
Xbit_r110_c41 bl[41] br[41] wl[110] vdd gnd cell_6t
Xbit_r111_c41 bl[41] br[41] wl[111] vdd gnd cell_6t
Xbit_r112_c41 bl[41] br[41] wl[112] vdd gnd cell_6t
Xbit_r113_c41 bl[41] br[41] wl[113] vdd gnd cell_6t
Xbit_r114_c41 bl[41] br[41] wl[114] vdd gnd cell_6t
Xbit_r115_c41 bl[41] br[41] wl[115] vdd gnd cell_6t
Xbit_r116_c41 bl[41] br[41] wl[116] vdd gnd cell_6t
Xbit_r117_c41 bl[41] br[41] wl[117] vdd gnd cell_6t
Xbit_r118_c41 bl[41] br[41] wl[118] vdd gnd cell_6t
Xbit_r119_c41 bl[41] br[41] wl[119] vdd gnd cell_6t
Xbit_r120_c41 bl[41] br[41] wl[120] vdd gnd cell_6t
Xbit_r121_c41 bl[41] br[41] wl[121] vdd gnd cell_6t
Xbit_r122_c41 bl[41] br[41] wl[122] vdd gnd cell_6t
Xbit_r123_c41 bl[41] br[41] wl[123] vdd gnd cell_6t
Xbit_r124_c41 bl[41] br[41] wl[124] vdd gnd cell_6t
Xbit_r125_c41 bl[41] br[41] wl[125] vdd gnd cell_6t
Xbit_r126_c41 bl[41] br[41] wl[126] vdd gnd cell_6t
Xbit_r127_c41 bl[41] br[41] wl[127] vdd gnd cell_6t
Xbit_r128_c41 bl[41] br[41] wl[128] vdd gnd cell_6t
Xbit_r129_c41 bl[41] br[41] wl[129] vdd gnd cell_6t
Xbit_r130_c41 bl[41] br[41] wl[130] vdd gnd cell_6t
Xbit_r131_c41 bl[41] br[41] wl[131] vdd gnd cell_6t
Xbit_r132_c41 bl[41] br[41] wl[132] vdd gnd cell_6t
Xbit_r133_c41 bl[41] br[41] wl[133] vdd gnd cell_6t
Xbit_r134_c41 bl[41] br[41] wl[134] vdd gnd cell_6t
Xbit_r135_c41 bl[41] br[41] wl[135] vdd gnd cell_6t
Xbit_r136_c41 bl[41] br[41] wl[136] vdd gnd cell_6t
Xbit_r137_c41 bl[41] br[41] wl[137] vdd gnd cell_6t
Xbit_r138_c41 bl[41] br[41] wl[138] vdd gnd cell_6t
Xbit_r139_c41 bl[41] br[41] wl[139] vdd gnd cell_6t
Xbit_r140_c41 bl[41] br[41] wl[140] vdd gnd cell_6t
Xbit_r141_c41 bl[41] br[41] wl[141] vdd gnd cell_6t
Xbit_r142_c41 bl[41] br[41] wl[142] vdd gnd cell_6t
Xbit_r143_c41 bl[41] br[41] wl[143] vdd gnd cell_6t
Xbit_r144_c41 bl[41] br[41] wl[144] vdd gnd cell_6t
Xbit_r145_c41 bl[41] br[41] wl[145] vdd gnd cell_6t
Xbit_r146_c41 bl[41] br[41] wl[146] vdd gnd cell_6t
Xbit_r147_c41 bl[41] br[41] wl[147] vdd gnd cell_6t
Xbit_r148_c41 bl[41] br[41] wl[148] vdd gnd cell_6t
Xbit_r149_c41 bl[41] br[41] wl[149] vdd gnd cell_6t
Xbit_r150_c41 bl[41] br[41] wl[150] vdd gnd cell_6t
Xbit_r151_c41 bl[41] br[41] wl[151] vdd gnd cell_6t
Xbit_r152_c41 bl[41] br[41] wl[152] vdd gnd cell_6t
Xbit_r153_c41 bl[41] br[41] wl[153] vdd gnd cell_6t
Xbit_r154_c41 bl[41] br[41] wl[154] vdd gnd cell_6t
Xbit_r155_c41 bl[41] br[41] wl[155] vdd gnd cell_6t
Xbit_r156_c41 bl[41] br[41] wl[156] vdd gnd cell_6t
Xbit_r157_c41 bl[41] br[41] wl[157] vdd gnd cell_6t
Xbit_r158_c41 bl[41] br[41] wl[158] vdd gnd cell_6t
Xbit_r159_c41 bl[41] br[41] wl[159] vdd gnd cell_6t
Xbit_r160_c41 bl[41] br[41] wl[160] vdd gnd cell_6t
Xbit_r161_c41 bl[41] br[41] wl[161] vdd gnd cell_6t
Xbit_r162_c41 bl[41] br[41] wl[162] vdd gnd cell_6t
Xbit_r163_c41 bl[41] br[41] wl[163] vdd gnd cell_6t
Xbit_r164_c41 bl[41] br[41] wl[164] vdd gnd cell_6t
Xbit_r165_c41 bl[41] br[41] wl[165] vdd gnd cell_6t
Xbit_r166_c41 bl[41] br[41] wl[166] vdd gnd cell_6t
Xbit_r167_c41 bl[41] br[41] wl[167] vdd gnd cell_6t
Xbit_r168_c41 bl[41] br[41] wl[168] vdd gnd cell_6t
Xbit_r169_c41 bl[41] br[41] wl[169] vdd gnd cell_6t
Xbit_r170_c41 bl[41] br[41] wl[170] vdd gnd cell_6t
Xbit_r171_c41 bl[41] br[41] wl[171] vdd gnd cell_6t
Xbit_r172_c41 bl[41] br[41] wl[172] vdd gnd cell_6t
Xbit_r173_c41 bl[41] br[41] wl[173] vdd gnd cell_6t
Xbit_r174_c41 bl[41] br[41] wl[174] vdd gnd cell_6t
Xbit_r175_c41 bl[41] br[41] wl[175] vdd gnd cell_6t
Xbit_r176_c41 bl[41] br[41] wl[176] vdd gnd cell_6t
Xbit_r177_c41 bl[41] br[41] wl[177] vdd gnd cell_6t
Xbit_r178_c41 bl[41] br[41] wl[178] vdd gnd cell_6t
Xbit_r179_c41 bl[41] br[41] wl[179] vdd gnd cell_6t
Xbit_r180_c41 bl[41] br[41] wl[180] vdd gnd cell_6t
Xbit_r181_c41 bl[41] br[41] wl[181] vdd gnd cell_6t
Xbit_r182_c41 bl[41] br[41] wl[182] vdd gnd cell_6t
Xbit_r183_c41 bl[41] br[41] wl[183] vdd gnd cell_6t
Xbit_r184_c41 bl[41] br[41] wl[184] vdd gnd cell_6t
Xbit_r185_c41 bl[41] br[41] wl[185] vdd gnd cell_6t
Xbit_r186_c41 bl[41] br[41] wl[186] vdd gnd cell_6t
Xbit_r187_c41 bl[41] br[41] wl[187] vdd gnd cell_6t
Xbit_r188_c41 bl[41] br[41] wl[188] vdd gnd cell_6t
Xbit_r189_c41 bl[41] br[41] wl[189] vdd gnd cell_6t
Xbit_r190_c41 bl[41] br[41] wl[190] vdd gnd cell_6t
Xbit_r191_c41 bl[41] br[41] wl[191] vdd gnd cell_6t
Xbit_r192_c41 bl[41] br[41] wl[192] vdd gnd cell_6t
Xbit_r193_c41 bl[41] br[41] wl[193] vdd gnd cell_6t
Xbit_r194_c41 bl[41] br[41] wl[194] vdd gnd cell_6t
Xbit_r195_c41 bl[41] br[41] wl[195] vdd gnd cell_6t
Xbit_r196_c41 bl[41] br[41] wl[196] vdd gnd cell_6t
Xbit_r197_c41 bl[41] br[41] wl[197] vdd gnd cell_6t
Xbit_r198_c41 bl[41] br[41] wl[198] vdd gnd cell_6t
Xbit_r199_c41 bl[41] br[41] wl[199] vdd gnd cell_6t
Xbit_r200_c41 bl[41] br[41] wl[200] vdd gnd cell_6t
Xbit_r201_c41 bl[41] br[41] wl[201] vdd gnd cell_6t
Xbit_r202_c41 bl[41] br[41] wl[202] vdd gnd cell_6t
Xbit_r203_c41 bl[41] br[41] wl[203] vdd gnd cell_6t
Xbit_r204_c41 bl[41] br[41] wl[204] vdd gnd cell_6t
Xbit_r205_c41 bl[41] br[41] wl[205] vdd gnd cell_6t
Xbit_r206_c41 bl[41] br[41] wl[206] vdd gnd cell_6t
Xbit_r207_c41 bl[41] br[41] wl[207] vdd gnd cell_6t
Xbit_r208_c41 bl[41] br[41] wl[208] vdd gnd cell_6t
Xbit_r209_c41 bl[41] br[41] wl[209] vdd gnd cell_6t
Xbit_r210_c41 bl[41] br[41] wl[210] vdd gnd cell_6t
Xbit_r211_c41 bl[41] br[41] wl[211] vdd gnd cell_6t
Xbit_r212_c41 bl[41] br[41] wl[212] vdd gnd cell_6t
Xbit_r213_c41 bl[41] br[41] wl[213] vdd gnd cell_6t
Xbit_r214_c41 bl[41] br[41] wl[214] vdd gnd cell_6t
Xbit_r215_c41 bl[41] br[41] wl[215] vdd gnd cell_6t
Xbit_r216_c41 bl[41] br[41] wl[216] vdd gnd cell_6t
Xbit_r217_c41 bl[41] br[41] wl[217] vdd gnd cell_6t
Xbit_r218_c41 bl[41] br[41] wl[218] vdd gnd cell_6t
Xbit_r219_c41 bl[41] br[41] wl[219] vdd gnd cell_6t
Xbit_r220_c41 bl[41] br[41] wl[220] vdd gnd cell_6t
Xbit_r221_c41 bl[41] br[41] wl[221] vdd gnd cell_6t
Xbit_r222_c41 bl[41] br[41] wl[222] vdd gnd cell_6t
Xbit_r223_c41 bl[41] br[41] wl[223] vdd gnd cell_6t
Xbit_r224_c41 bl[41] br[41] wl[224] vdd gnd cell_6t
Xbit_r225_c41 bl[41] br[41] wl[225] vdd gnd cell_6t
Xbit_r226_c41 bl[41] br[41] wl[226] vdd gnd cell_6t
Xbit_r227_c41 bl[41] br[41] wl[227] vdd gnd cell_6t
Xbit_r228_c41 bl[41] br[41] wl[228] vdd gnd cell_6t
Xbit_r229_c41 bl[41] br[41] wl[229] vdd gnd cell_6t
Xbit_r230_c41 bl[41] br[41] wl[230] vdd gnd cell_6t
Xbit_r231_c41 bl[41] br[41] wl[231] vdd gnd cell_6t
Xbit_r232_c41 bl[41] br[41] wl[232] vdd gnd cell_6t
Xbit_r233_c41 bl[41] br[41] wl[233] vdd gnd cell_6t
Xbit_r234_c41 bl[41] br[41] wl[234] vdd gnd cell_6t
Xbit_r235_c41 bl[41] br[41] wl[235] vdd gnd cell_6t
Xbit_r236_c41 bl[41] br[41] wl[236] vdd gnd cell_6t
Xbit_r237_c41 bl[41] br[41] wl[237] vdd gnd cell_6t
Xbit_r238_c41 bl[41] br[41] wl[238] vdd gnd cell_6t
Xbit_r239_c41 bl[41] br[41] wl[239] vdd gnd cell_6t
Xbit_r240_c41 bl[41] br[41] wl[240] vdd gnd cell_6t
Xbit_r241_c41 bl[41] br[41] wl[241] vdd gnd cell_6t
Xbit_r242_c41 bl[41] br[41] wl[242] vdd gnd cell_6t
Xbit_r243_c41 bl[41] br[41] wl[243] vdd gnd cell_6t
Xbit_r244_c41 bl[41] br[41] wl[244] vdd gnd cell_6t
Xbit_r245_c41 bl[41] br[41] wl[245] vdd gnd cell_6t
Xbit_r246_c41 bl[41] br[41] wl[246] vdd gnd cell_6t
Xbit_r247_c41 bl[41] br[41] wl[247] vdd gnd cell_6t
Xbit_r248_c41 bl[41] br[41] wl[248] vdd gnd cell_6t
Xbit_r249_c41 bl[41] br[41] wl[249] vdd gnd cell_6t
Xbit_r250_c41 bl[41] br[41] wl[250] vdd gnd cell_6t
Xbit_r251_c41 bl[41] br[41] wl[251] vdd gnd cell_6t
Xbit_r252_c41 bl[41] br[41] wl[252] vdd gnd cell_6t
Xbit_r253_c41 bl[41] br[41] wl[253] vdd gnd cell_6t
Xbit_r254_c41 bl[41] br[41] wl[254] vdd gnd cell_6t
Xbit_r255_c41 bl[41] br[41] wl[255] vdd gnd cell_6t
Xbit_r0_c42 bl[42] br[42] wl[0] vdd gnd cell_6t
Xbit_r1_c42 bl[42] br[42] wl[1] vdd gnd cell_6t
Xbit_r2_c42 bl[42] br[42] wl[2] vdd gnd cell_6t
Xbit_r3_c42 bl[42] br[42] wl[3] vdd gnd cell_6t
Xbit_r4_c42 bl[42] br[42] wl[4] vdd gnd cell_6t
Xbit_r5_c42 bl[42] br[42] wl[5] vdd gnd cell_6t
Xbit_r6_c42 bl[42] br[42] wl[6] vdd gnd cell_6t
Xbit_r7_c42 bl[42] br[42] wl[7] vdd gnd cell_6t
Xbit_r8_c42 bl[42] br[42] wl[8] vdd gnd cell_6t
Xbit_r9_c42 bl[42] br[42] wl[9] vdd gnd cell_6t
Xbit_r10_c42 bl[42] br[42] wl[10] vdd gnd cell_6t
Xbit_r11_c42 bl[42] br[42] wl[11] vdd gnd cell_6t
Xbit_r12_c42 bl[42] br[42] wl[12] vdd gnd cell_6t
Xbit_r13_c42 bl[42] br[42] wl[13] vdd gnd cell_6t
Xbit_r14_c42 bl[42] br[42] wl[14] vdd gnd cell_6t
Xbit_r15_c42 bl[42] br[42] wl[15] vdd gnd cell_6t
Xbit_r16_c42 bl[42] br[42] wl[16] vdd gnd cell_6t
Xbit_r17_c42 bl[42] br[42] wl[17] vdd gnd cell_6t
Xbit_r18_c42 bl[42] br[42] wl[18] vdd gnd cell_6t
Xbit_r19_c42 bl[42] br[42] wl[19] vdd gnd cell_6t
Xbit_r20_c42 bl[42] br[42] wl[20] vdd gnd cell_6t
Xbit_r21_c42 bl[42] br[42] wl[21] vdd gnd cell_6t
Xbit_r22_c42 bl[42] br[42] wl[22] vdd gnd cell_6t
Xbit_r23_c42 bl[42] br[42] wl[23] vdd gnd cell_6t
Xbit_r24_c42 bl[42] br[42] wl[24] vdd gnd cell_6t
Xbit_r25_c42 bl[42] br[42] wl[25] vdd gnd cell_6t
Xbit_r26_c42 bl[42] br[42] wl[26] vdd gnd cell_6t
Xbit_r27_c42 bl[42] br[42] wl[27] vdd gnd cell_6t
Xbit_r28_c42 bl[42] br[42] wl[28] vdd gnd cell_6t
Xbit_r29_c42 bl[42] br[42] wl[29] vdd gnd cell_6t
Xbit_r30_c42 bl[42] br[42] wl[30] vdd gnd cell_6t
Xbit_r31_c42 bl[42] br[42] wl[31] vdd gnd cell_6t
Xbit_r32_c42 bl[42] br[42] wl[32] vdd gnd cell_6t
Xbit_r33_c42 bl[42] br[42] wl[33] vdd gnd cell_6t
Xbit_r34_c42 bl[42] br[42] wl[34] vdd gnd cell_6t
Xbit_r35_c42 bl[42] br[42] wl[35] vdd gnd cell_6t
Xbit_r36_c42 bl[42] br[42] wl[36] vdd gnd cell_6t
Xbit_r37_c42 bl[42] br[42] wl[37] vdd gnd cell_6t
Xbit_r38_c42 bl[42] br[42] wl[38] vdd gnd cell_6t
Xbit_r39_c42 bl[42] br[42] wl[39] vdd gnd cell_6t
Xbit_r40_c42 bl[42] br[42] wl[40] vdd gnd cell_6t
Xbit_r41_c42 bl[42] br[42] wl[41] vdd gnd cell_6t
Xbit_r42_c42 bl[42] br[42] wl[42] vdd gnd cell_6t
Xbit_r43_c42 bl[42] br[42] wl[43] vdd gnd cell_6t
Xbit_r44_c42 bl[42] br[42] wl[44] vdd gnd cell_6t
Xbit_r45_c42 bl[42] br[42] wl[45] vdd gnd cell_6t
Xbit_r46_c42 bl[42] br[42] wl[46] vdd gnd cell_6t
Xbit_r47_c42 bl[42] br[42] wl[47] vdd gnd cell_6t
Xbit_r48_c42 bl[42] br[42] wl[48] vdd gnd cell_6t
Xbit_r49_c42 bl[42] br[42] wl[49] vdd gnd cell_6t
Xbit_r50_c42 bl[42] br[42] wl[50] vdd gnd cell_6t
Xbit_r51_c42 bl[42] br[42] wl[51] vdd gnd cell_6t
Xbit_r52_c42 bl[42] br[42] wl[52] vdd gnd cell_6t
Xbit_r53_c42 bl[42] br[42] wl[53] vdd gnd cell_6t
Xbit_r54_c42 bl[42] br[42] wl[54] vdd gnd cell_6t
Xbit_r55_c42 bl[42] br[42] wl[55] vdd gnd cell_6t
Xbit_r56_c42 bl[42] br[42] wl[56] vdd gnd cell_6t
Xbit_r57_c42 bl[42] br[42] wl[57] vdd gnd cell_6t
Xbit_r58_c42 bl[42] br[42] wl[58] vdd gnd cell_6t
Xbit_r59_c42 bl[42] br[42] wl[59] vdd gnd cell_6t
Xbit_r60_c42 bl[42] br[42] wl[60] vdd gnd cell_6t
Xbit_r61_c42 bl[42] br[42] wl[61] vdd gnd cell_6t
Xbit_r62_c42 bl[42] br[42] wl[62] vdd gnd cell_6t
Xbit_r63_c42 bl[42] br[42] wl[63] vdd gnd cell_6t
Xbit_r64_c42 bl[42] br[42] wl[64] vdd gnd cell_6t
Xbit_r65_c42 bl[42] br[42] wl[65] vdd gnd cell_6t
Xbit_r66_c42 bl[42] br[42] wl[66] vdd gnd cell_6t
Xbit_r67_c42 bl[42] br[42] wl[67] vdd gnd cell_6t
Xbit_r68_c42 bl[42] br[42] wl[68] vdd gnd cell_6t
Xbit_r69_c42 bl[42] br[42] wl[69] vdd gnd cell_6t
Xbit_r70_c42 bl[42] br[42] wl[70] vdd gnd cell_6t
Xbit_r71_c42 bl[42] br[42] wl[71] vdd gnd cell_6t
Xbit_r72_c42 bl[42] br[42] wl[72] vdd gnd cell_6t
Xbit_r73_c42 bl[42] br[42] wl[73] vdd gnd cell_6t
Xbit_r74_c42 bl[42] br[42] wl[74] vdd gnd cell_6t
Xbit_r75_c42 bl[42] br[42] wl[75] vdd gnd cell_6t
Xbit_r76_c42 bl[42] br[42] wl[76] vdd gnd cell_6t
Xbit_r77_c42 bl[42] br[42] wl[77] vdd gnd cell_6t
Xbit_r78_c42 bl[42] br[42] wl[78] vdd gnd cell_6t
Xbit_r79_c42 bl[42] br[42] wl[79] vdd gnd cell_6t
Xbit_r80_c42 bl[42] br[42] wl[80] vdd gnd cell_6t
Xbit_r81_c42 bl[42] br[42] wl[81] vdd gnd cell_6t
Xbit_r82_c42 bl[42] br[42] wl[82] vdd gnd cell_6t
Xbit_r83_c42 bl[42] br[42] wl[83] vdd gnd cell_6t
Xbit_r84_c42 bl[42] br[42] wl[84] vdd gnd cell_6t
Xbit_r85_c42 bl[42] br[42] wl[85] vdd gnd cell_6t
Xbit_r86_c42 bl[42] br[42] wl[86] vdd gnd cell_6t
Xbit_r87_c42 bl[42] br[42] wl[87] vdd gnd cell_6t
Xbit_r88_c42 bl[42] br[42] wl[88] vdd gnd cell_6t
Xbit_r89_c42 bl[42] br[42] wl[89] vdd gnd cell_6t
Xbit_r90_c42 bl[42] br[42] wl[90] vdd gnd cell_6t
Xbit_r91_c42 bl[42] br[42] wl[91] vdd gnd cell_6t
Xbit_r92_c42 bl[42] br[42] wl[92] vdd gnd cell_6t
Xbit_r93_c42 bl[42] br[42] wl[93] vdd gnd cell_6t
Xbit_r94_c42 bl[42] br[42] wl[94] vdd gnd cell_6t
Xbit_r95_c42 bl[42] br[42] wl[95] vdd gnd cell_6t
Xbit_r96_c42 bl[42] br[42] wl[96] vdd gnd cell_6t
Xbit_r97_c42 bl[42] br[42] wl[97] vdd gnd cell_6t
Xbit_r98_c42 bl[42] br[42] wl[98] vdd gnd cell_6t
Xbit_r99_c42 bl[42] br[42] wl[99] vdd gnd cell_6t
Xbit_r100_c42 bl[42] br[42] wl[100] vdd gnd cell_6t
Xbit_r101_c42 bl[42] br[42] wl[101] vdd gnd cell_6t
Xbit_r102_c42 bl[42] br[42] wl[102] vdd gnd cell_6t
Xbit_r103_c42 bl[42] br[42] wl[103] vdd gnd cell_6t
Xbit_r104_c42 bl[42] br[42] wl[104] vdd gnd cell_6t
Xbit_r105_c42 bl[42] br[42] wl[105] vdd gnd cell_6t
Xbit_r106_c42 bl[42] br[42] wl[106] vdd gnd cell_6t
Xbit_r107_c42 bl[42] br[42] wl[107] vdd gnd cell_6t
Xbit_r108_c42 bl[42] br[42] wl[108] vdd gnd cell_6t
Xbit_r109_c42 bl[42] br[42] wl[109] vdd gnd cell_6t
Xbit_r110_c42 bl[42] br[42] wl[110] vdd gnd cell_6t
Xbit_r111_c42 bl[42] br[42] wl[111] vdd gnd cell_6t
Xbit_r112_c42 bl[42] br[42] wl[112] vdd gnd cell_6t
Xbit_r113_c42 bl[42] br[42] wl[113] vdd gnd cell_6t
Xbit_r114_c42 bl[42] br[42] wl[114] vdd gnd cell_6t
Xbit_r115_c42 bl[42] br[42] wl[115] vdd gnd cell_6t
Xbit_r116_c42 bl[42] br[42] wl[116] vdd gnd cell_6t
Xbit_r117_c42 bl[42] br[42] wl[117] vdd gnd cell_6t
Xbit_r118_c42 bl[42] br[42] wl[118] vdd gnd cell_6t
Xbit_r119_c42 bl[42] br[42] wl[119] vdd gnd cell_6t
Xbit_r120_c42 bl[42] br[42] wl[120] vdd gnd cell_6t
Xbit_r121_c42 bl[42] br[42] wl[121] vdd gnd cell_6t
Xbit_r122_c42 bl[42] br[42] wl[122] vdd gnd cell_6t
Xbit_r123_c42 bl[42] br[42] wl[123] vdd gnd cell_6t
Xbit_r124_c42 bl[42] br[42] wl[124] vdd gnd cell_6t
Xbit_r125_c42 bl[42] br[42] wl[125] vdd gnd cell_6t
Xbit_r126_c42 bl[42] br[42] wl[126] vdd gnd cell_6t
Xbit_r127_c42 bl[42] br[42] wl[127] vdd gnd cell_6t
Xbit_r128_c42 bl[42] br[42] wl[128] vdd gnd cell_6t
Xbit_r129_c42 bl[42] br[42] wl[129] vdd gnd cell_6t
Xbit_r130_c42 bl[42] br[42] wl[130] vdd gnd cell_6t
Xbit_r131_c42 bl[42] br[42] wl[131] vdd gnd cell_6t
Xbit_r132_c42 bl[42] br[42] wl[132] vdd gnd cell_6t
Xbit_r133_c42 bl[42] br[42] wl[133] vdd gnd cell_6t
Xbit_r134_c42 bl[42] br[42] wl[134] vdd gnd cell_6t
Xbit_r135_c42 bl[42] br[42] wl[135] vdd gnd cell_6t
Xbit_r136_c42 bl[42] br[42] wl[136] vdd gnd cell_6t
Xbit_r137_c42 bl[42] br[42] wl[137] vdd gnd cell_6t
Xbit_r138_c42 bl[42] br[42] wl[138] vdd gnd cell_6t
Xbit_r139_c42 bl[42] br[42] wl[139] vdd gnd cell_6t
Xbit_r140_c42 bl[42] br[42] wl[140] vdd gnd cell_6t
Xbit_r141_c42 bl[42] br[42] wl[141] vdd gnd cell_6t
Xbit_r142_c42 bl[42] br[42] wl[142] vdd gnd cell_6t
Xbit_r143_c42 bl[42] br[42] wl[143] vdd gnd cell_6t
Xbit_r144_c42 bl[42] br[42] wl[144] vdd gnd cell_6t
Xbit_r145_c42 bl[42] br[42] wl[145] vdd gnd cell_6t
Xbit_r146_c42 bl[42] br[42] wl[146] vdd gnd cell_6t
Xbit_r147_c42 bl[42] br[42] wl[147] vdd gnd cell_6t
Xbit_r148_c42 bl[42] br[42] wl[148] vdd gnd cell_6t
Xbit_r149_c42 bl[42] br[42] wl[149] vdd gnd cell_6t
Xbit_r150_c42 bl[42] br[42] wl[150] vdd gnd cell_6t
Xbit_r151_c42 bl[42] br[42] wl[151] vdd gnd cell_6t
Xbit_r152_c42 bl[42] br[42] wl[152] vdd gnd cell_6t
Xbit_r153_c42 bl[42] br[42] wl[153] vdd gnd cell_6t
Xbit_r154_c42 bl[42] br[42] wl[154] vdd gnd cell_6t
Xbit_r155_c42 bl[42] br[42] wl[155] vdd gnd cell_6t
Xbit_r156_c42 bl[42] br[42] wl[156] vdd gnd cell_6t
Xbit_r157_c42 bl[42] br[42] wl[157] vdd gnd cell_6t
Xbit_r158_c42 bl[42] br[42] wl[158] vdd gnd cell_6t
Xbit_r159_c42 bl[42] br[42] wl[159] vdd gnd cell_6t
Xbit_r160_c42 bl[42] br[42] wl[160] vdd gnd cell_6t
Xbit_r161_c42 bl[42] br[42] wl[161] vdd gnd cell_6t
Xbit_r162_c42 bl[42] br[42] wl[162] vdd gnd cell_6t
Xbit_r163_c42 bl[42] br[42] wl[163] vdd gnd cell_6t
Xbit_r164_c42 bl[42] br[42] wl[164] vdd gnd cell_6t
Xbit_r165_c42 bl[42] br[42] wl[165] vdd gnd cell_6t
Xbit_r166_c42 bl[42] br[42] wl[166] vdd gnd cell_6t
Xbit_r167_c42 bl[42] br[42] wl[167] vdd gnd cell_6t
Xbit_r168_c42 bl[42] br[42] wl[168] vdd gnd cell_6t
Xbit_r169_c42 bl[42] br[42] wl[169] vdd gnd cell_6t
Xbit_r170_c42 bl[42] br[42] wl[170] vdd gnd cell_6t
Xbit_r171_c42 bl[42] br[42] wl[171] vdd gnd cell_6t
Xbit_r172_c42 bl[42] br[42] wl[172] vdd gnd cell_6t
Xbit_r173_c42 bl[42] br[42] wl[173] vdd gnd cell_6t
Xbit_r174_c42 bl[42] br[42] wl[174] vdd gnd cell_6t
Xbit_r175_c42 bl[42] br[42] wl[175] vdd gnd cell_6t
Xbit_r176_c42 bl[42] br[42] wl[176] vdd gnd cell_6t
Xbit_r177_c42 bl[42] br[42] wl[177] vdd gnd cell_6t
Xbit_r178_c42 bl[42] br[42] wl[178] vdd gnd cell_6t
Xbit_r179_c42 bl[42] br[42] wl[179] vdd gnd cell_6t
Xbit_r180_c42 bl[42] br[42] wl[180] vdd gnd cell_6t
Xbit_r181_c42 bl[42] br[42] wl[181] vdd gnd cell_6t
Xbit_r182_c42 bl[42] br[42] wl[182] vdd gnd cell_6t
Xbit_r183_c42 bl[42] br[42] wl[183] vdd gnd cell_6t
Xbit_r184_c42 bl[42] br[42] wl[184] vdd gnd cell_6t
Xbit_r185_c42 bl[42] br[42] wl[185] vdd gnd cell_6t
Xbit_r186_c42 bl[42] br[42] wl[186] vdd gnd cell_6t
Xbit_r187_c42 bl[42] br[42] wl[187] vdd gnd cell_6t
Xbit_r188_c42 bl[42] br[42] wl[188] vdd gnd cell_6t
Xbit_r189_c42 bl[42] br[42] wl[189] vdd gnd cell_6t
Xbit_r190_c42 bl[42] br[42] wl[190] vdd gnd cell_6t
Xbit_r191_c42 bl[42] br[42] wl[191] vdd gnd cell_6t
Xbit_r192_c42 bl[42] br[42] wl[192] vdd gnd cell_6t
Xbit_r193_c42 bl[42] br[42] wl[193] vdd gnd cell_6t
Xbit_r194_c42 bl[42] br[42] wl[194] vdd gnd cell_6t
Xbit_r195_c42 bl[42] br[42] wl[195] vdd gnd cell_6t
Xbit_r196_c42 bl[42] br[42] wl[196] vdd gnd cell_6t
Xbit_r197_c42 bl[42] br[42] wl[197] vdd gnd cell_6t
Xbit_r198_c42 bl[42] br[42] wl[198] vdd gnd cell_6t
Xbit_r199_c42 bl[42] br[42] wl[199] vdd gnd cell_6t
Xbit_r200_c42 bl[42] br[42] wl[200] vdd gnd cell_6t
Xbit_r201_c42 bl[42] br[42] wl[201] vdd gnd cell_6t
Xbit_r202_c42 bl[42] br[42] wl[202] vdd gnd cell_6t
Xbit_r203_c42 bl[42] br[42] wl[203] vdd gnd cell_6t
Xbit_r204_c42 bl[42] br[42] wl[204] vdd gnd cell_6t
Xbit_r205_c42 bl[42] br[42] wl[205] vdd gnd cell_6t
Xbit_r206_c42 bl[42] br[42] wl[206] vdd gnd cell_6t
Xbit_r207_c42 bl[42] br[42] wl[207] vdd gnd cell_6t
Xbit_r208_c42 bl[42] br[42] wl[208] vdd gnd cell_6t
Xbit_r209_c42 bl[42] br[42] wl[209] vdd gnd cell_6t
Xbit_r210_c42 bl[42] br[42] wl[210] vdd gnd cell_6t
Xbit_r211_c42 bl[42] br[42] wl[211] vdd gnd cell_6t
Xbit_r212_c42 bl[42] br[42] wl[212] vdd gnd cell_6t
Xbit_r213_c42 bl[42] br[42] wl[213] vdd gnd cell_6t
Xbit_r214_c42 bl[42] br[42] wl[214] vdd gnd cell_6t
Xbit_r215_c42 bl[42] br[42] wl[215] vdd gnd cell_6t
Xbit_r216_c42 bl[42] br[42] wl[216] vdd gnd cell_6t
Xbit_r217_c42 bl[42] br[42] wl[217] vdd gnd cell_6t
Xbit_r218_c42 bl[42] br[42] wl[218] vdd gnd cell_6t
Xbit_r219_c42 bl[42] br[42] wl[219] vdd gnd cell_6t
Xbit_r220_c42 bl[42] br[42] wl[220] vdd gnd cell_6t
Xbit_r221_c42 bl[42] br[42] wl[221] vdd gnd cell_6t
Xbit_r222_c42 bl[42] br[42] wl[222] vdd gnd cell_6t
Xbit_r223_c42 bl[42] br[42] wl[223] vdd gnd cell_6t
Xbit_r224_c42 bl[42] br[42] wl[224] vdd gnd cell_6t
Xbit_r225_c42 bl[42] br[42] wl[225] vdd gnd cell_6t
Xbit_r226_c42 bl[42] br[42] wl[226] vdd gnd cell_6t
Xbit_r227_c42 bl[42] br[42] wl[227] vdd gnd cell_6t
Xbit_r228_c42 bl[42] br[42] wl[228] vdd gnd cell_6t
Xbit_r229_c42 bl[42] br[42] wl[229] vdd gnd cell_6t
Xbit_r230_c42 bl[42] br[42] wl[230] vdd gnd cell_6t
Xbit_r231_c42 bl[42] br[42] wl[231] vdd gnd cell_6t
Xbit_r232_c42 bl[42] br[42] wl[232] vdd gnd cell_6t
Xbit_r233_c42 bl[42] br[42] wl[233] vdd gnd cell_6t
Xbit_r234_c42 bl[42] br[42] wl[234] vdd gnd cell_6t
Xbit_r235_c42 bl[42] br[42] wl[235] vdd gnd cell_6t
Xbit_r236_c42 bl[42] br[42] wl[236] vdd gnd cell_6t
Xbit_r237_c42 bl[42] br[42] wl[237] vdd gnd cell_6t
Xbit_r238_c42 bl[42] br[42] wl[238] vdd gnd cell_6t
Xbit_r239_c42 bl[42] br[42] wl[239] vdd gnd cell_6t
Xbit_r240_c42 bl[42] br[42] wl[240] vdd gnd cell_6t
Xbit_r241_c42 bl[42] br[42] wl[241] vdd gnd cell_6t
Xbit_r242_c42 bl[42] br[42] wl[242] vdd gnd cell_6t
Xbit_r243_c42 bl[42] br[42] wl[243] vdd gnd cell_6t
Xbit_r244_c42 bl[42] br[42] wl[244] vdd gnd cell_6t
Xbit_r245_c42 bl[42] br[42] wl[245] vdd gnd cell_6t
Xbit_r246_c42 bl[42] br[42] wl[246] vdd gnd cell_6t
Xbit_r247_c42 bl[42] br[42] wl[247] vdd gnd cell_6t
Xbit_r248_c42 bl[42] br[42] wl[248] vdd gnd cell_6t
Xbit_r249_c42 bl[42] br[42] wl[249] vdd gnd cell_6t
Xbit_r250_c42 bl[42] br[42] wl[250] vdd gnd cell_6t
Xbit_r251_c42 bl[42] br[42] wl[251] vdd gnd cell_6t
Xbit_r252_c42 bl[42] br[42] wl[252] vdd gnd cell_6t
Xbit_r253_c42 bl[42] br[42] wl[253] vdd gnd cell_6t
Xbit_r254_c42 bl[42] br[42] wl[254] vdd gnd cell_6t
Xbit_r255_c42 bl[42] br[42] wl[255] vdd gnd cell_6t
Xbit_r0_c43 bl[43] br[43] wl[0] vdd gnd cell_6t
Xbit_r1_c43 bl[43] br[43] wl[1] vdd gnd cell_6t
Xbit_r2_c43 bl[43] br[43] wl[2] vdd gnd cell_6t
Xbit_r3_c43 bl[43] br[43] wl[3] vdd gnd cell_6t
Xbit_r4_c43 bl[43] br[43] wl[4] vdd gnd cell_6t
Xbit_r5_c43 bl[43] br[43] wl[5] vdd gnd cell_6t
Xbit_r6_c43 bl[43] br[43] wl[6] vdd gnd cell_6t
Xbit_r7_c43 bl[43] br[43] wl[7] vdd gnd cell_6t
Xbit_r8_c43 bl[43] br[43] wl[8] vdd gnd cell_6t
Xbit_r9_c43 bl[43] br[43] wl[9] vdd gnd cell_6t
Xbit_r10_c43 bl[43] br[43] wl[10] vdd gnd cell_6t
Xbit_r11_c43 bl[43] br[43] wl[11] vdd gnd cell_6t
Xbit_r12_c43 bl[43] br[43] wl[12] vdd gnd cell_6t
Xbit_r13_c43 bl[43] br[43] wl[13] vdd gnd cell_6t
Xbit_r14_c43 bl[43] br[43] wl[14] vdd gnd cell_6t
Xbit_r15_c43 bl[43] br[43] wl[15] vdd gnd cell_6t
Xbit_r16_c43 bl[43] br[43] wl[16] vdd gnd cell_6t
Xbit_r17_c43 bl[43] br[43] wl[17] vdd gnd cell_6t
Xbit_r18_c43 bl[43] br[43] wl[18] vdd gnd cell_6t
Xbit_r19_c43 bl[43] br[43] wl[19] vdd gnd cell_6t
Xbit_r20_c43 bl[43] br[43] wl[20] vdd gnd cell_6t
Xbit_r21_c43 bl[43] br[43] wl[21] vdd gnd cell_6t
Xbit_r22_c43 bl[43] br[43] wl[22] vdd gnd cell_6t
Xbit_r23_c43 bl[43] br[43] wl[23] vdd gnd cell_6t
Xbit_r24_c43 bl[43] br[43] wl[24] vdd gnd cell_6t
Xbit_r25_c43 bl[43] br[43] wl[25] vdd gnd cell_6t
Xbit_r26_c43 bl[43] br[43] wl[26] vdd gnd cell_6t
Xbit_r27_c43 bl[43] br[43] wl[27] vdd gnd cell_6t
Xbit_r28_c43 bl[43] br[43] wl[28] vdd gnd cell_6t
Xbit_r29_c43 bl[43] br[43] wl[29] vdd gnd cell_6t
Xbit_r30_c43 bl[43] br[43] wl[30] vdd gnd cell_6t
Xbit_r31_c43 bl[43] br[43] wl[31] vdd gnd cell_6t
Xbit_r32_c43 bl[43] br[43] wl[32] vdd gnd cell_6t
Xbit_r33_c43 bl[43] br[43] wl[33] vdd gnd cell_6t
Xbit_r34_c43 bl[43] br[43] wl[34] vdd gnd cell_6t
Xbit_r35_c43 bl[43] br[43] wl[35] vdd gnd cell_6t
Xbit_r36_c43 bl[43] br[43] wl[36] vdd gnd cell_6t
Xbit_r37_c43 bl[43] br[43] wl[37] vdd gnd cell_6t
Xbit_r38_c43 bl[43] br[43] wl[38] vdd gnd cell_6t
Xbit_r39_c43 bl[43] br[43] wl[39] vdd gnd cell_6t
Xbit_r40_c43 bl[43] br[43] wl[40] vdd gnd cell_6t
Xbit_r41_c43 bl[43] br[43] wl[41] vdd gnd cell_6t
Xbit_r42_c43 bl[43] br[43] wl[42] vdd gnd cell_6t
Xbit_r43_c43 bl[43] br[43] wl[43] vdd gnd cell_6t
Xbit_r44_c43 bl[43] br[43] wl[44] vdd gnd cell_6t
Xbit_r45_c43 bl[43] br[43] wl[45] vdd gnd cell_6t
Xbit_r46_c43 bl[43] br[43] wl[46] vdd gnd cell_6t
Xbit_r47_c43 bl[43] br[43] wl[47] vdd gnd cell_6t
Xbit_r48_c43 bl[43] br[43] wl[48] vdd gnd cell_6t
Xbit_r49_c43 bl[43] br[43] wl[49] vdd gnd cell_6t
Xbit_r50_c43 bl[43] br[43] wl[50] vdd gnd cell_6t
Xbit_r51_c43 bl[43] br[43] wl[51] vdd gnd cell_6t
Xbit_r52_c43 bl[43] br[43] wl[52] vdd gnd cell_6t
Xbit_r53_c43 bl[43] br[43] wl[53] vdd gnd cell_6t
Xbit_r54_c43 bl[43] br[43] wl[54] vdd gnd cell_6t
Xbit_r55_c43 bl[43] br[43] wl[55] vdd gnd cell_6t
Xbit_r56_c43 bl[43] br[43] wl[56] vdd gnd cell_6t
Xbit_r57_c43 bl[43] br[43] wl[57] vdd gnd cell_6t
Xbit_r58_c43 bl[43] br[43] wl[58] vdd gnd cell_6t
Xbit_r59_c43 bl[43] br[43] wl[59] vdd gnd cell_6t
Xbit_r60_c43 bl[43] br[43] wl[60] vdd gnd cell_6t
Xbit_r61_c43 bl[43] br[43] wl[61] vdd gnd cell_6t
Xbit_r62_c43 bl[43] br[43] wl[62] vdd gnd cell_6t
Xbit_r63_c43 bl[43] br[43] wl[63] vdd gnd cell_6t
Xbit_r64_c43 bl[43] br[43] wl[64] vdd gnd cell_6t
Xbit_r65_c43 bl[43] br[43] wl[65] vdd gnd cell_6t
Xbit_r66_c43 bl[43] br[43] wl[66] vdd gnd cell_6t
Xbit_r67_c43 bl[43] br[43] wl[67] vdd gnd cell_6t
Xbit_r68_c43 bl[43] br[43] wl[68] vdd gnd cell_6t
Xbit_r69_c43 bl[43] br[43] wl[69] vdd gnd cell_6t
Xbit_r70_c43 bl[43] br[43] wl[70] vdd gnd cell_6t
Xbit_r71_c43 bl[43] br[43] wl[71] vdd gnd cell_6t
Xbit_r72_c43 bl[43] br[43] wl[72] vdd gnd cell_6t
Xbit_r73_c43 bl[43] br[43] wl[73] vdd gnd cell_6t
Xbit_r74_c43 bl[43] br[43] wl[74] vdd gnd cell_6t
Xbit_r75_c43 bl[43] br[43] wl[75] vdd gnd cell_6t
Xbit_r76_c43 bl[43] br[43] wl[76] vdd gnd cell_6t
Xbit_r77_c43 bl[43] br[43] wl[77] vdd gnd cell_6t
Xbit_r78_c43 bl[43] br[43] wl[78] vdd gnd cell_6t
Xbit_r79_c43 bl[43] br[43] wl[79] vdd gnd cell_6t
Xbit_r80_c43 bl[43] br[43] wl[80] vdd gnd cell_6t
Xbit_r81_c43 bl[43] br[43] wl[81] vdd gnd cell_6t
Xbit_r82_c43 bl[43] br[43] wl[82] vdd gnd cell_6t
Xbit_r83_c43 bl[43] br[43] wl[83] vdd gnd cell_6t
Xbit_r84_c43 bl[43] br[43] wl[84] vdd gnd cell_6t
Xbit_r85_c43 bl[43] br[43] wl[85] vdd gnd cell_6t
Xbit_r86_c43 bl[43] br[43] wl[86] vdd gnd cell_6t
Xbit_r87_c43 bl[43] br[43] wl[87] vdd gnd cell_6t
Xbit_r88_c43 bl[43] br[43] wl[88] vdd gnd cell_6t
Xbit_r89_c43 bl[43] br[43] wl[89] vdd gnd cell_6t
Xbit_r90_c43 bl[43] br[43] wl[90] vdd gnd cell_6t
Xbit_r91_c43 bl[43] br[43] wl[91] vdd gnd cell_6t
Xbit_r92_c43 bl[43] br[43] wl[92] vdd gnd cell_6t
Xbit_r93_c43 bl[43] br[43] wl[93] vdd gnd cell_6t
Xbit_r94_c43 bl[43] br[43] wl[94] vdd gnd cell_6t
Xbit_r95_c43 bl[43] br[43] wl[95] vdd gnd cell_6t
Xbit_r96_c43 bl[43] br[43] wl[96] vdd gnd cell_6t
Xbit_r97_c43 bl[43] br[43] wl[97] vdd gnd cell_6t
Xbit_r98_c43 bl[43] br[43] wl[98] vdd gnd cell_6t
Xbit_r99_c43 bl[43] br[43] wl[99] vdd gnd cell_6t
Xbit_r100_c43 bl[43] br[43] wl[100] vdd gnd cell_6t
Xbit_r101_c43 bl[43] br[43] wl[101] vdd gnd cell_6t
Xbit_r102_c43 bl[43] br[43] wl[102] vdd gnd cell_6t
Xbit_r103_c43 bl[43] br[43] wl[103] vdd gnd cell_6t
Xbit_r104_c43 bl[43] br[43] wl[104] vdd gnd cell_6t
Xbit_r105_c43 bl[43] br[43] wl[105] vdd gnd cell_6t
Xbit_r106_c43 bl[43] br[43] wl[106] vdd gnd cell_6t
Xbit_r107_c43 bl[43] br[43] wl[107] vdd gnd cell_6t
Xbit_r108_c43 bl[43] br[43] wl[108] vdd gnd cell_6t
Xbit_r109_c43 bl[43] br[43] wl[109] vdd gnd cell_6t
Xbit_r110_c43 bl[43] br[43] wl[110] vdd gnd cell_6t
Xbit_r111_c43 bl[43] br[43] wl[111] vdd gnd cell_6t
Xbit_r112_c43 bl[43] br[43] wl[112] vdd gnd cell_6t
Xbit_r113_c43 bl[43] br[43] wl[113] vdd gnd cell_6t
Xbit_r114_c43 bl[43] br[43] wl[114] vdd gnd cell_6t
Xbit_r115_c43 bl[43] br[43] wl[115] vdd gnd cell_6t
Xbit_r116_c43 bl[43] br[43] wl[116] vdd gnd cell_6t
Xbit_r117_c43 bl[43] br[43] wl[117] vdd gnd cell_6t
Xbit_r118_c43 bl[43] br[43] wl[118] vdd gnd cell_6t
Xbit_r119_c43 bl[43] br[43] wl[119] vdd gnd cell_6t
Xbit_r120_c43 bl[43] br[43] wl[120] vdd gnd cell_6t
Xbit_r121_c43 bl[43] br[43] wl[121] vdd gnd cell_6t
Xbit_r122_c43 bl[43] br[43] wl[122] vdd gnd cell_6t
Xbit_r123_c43 bl[43] br[43] wl[123] vdd gnd cell_6t
Xbit_r124_c43 bl[43] br[43] wl[124] vdd gnd cell_6t
Xbit_r125_c43 bl[43] br[43] wl[125] vdd gnd cell_6t
Xbit_r126_c43 bl[43] br[43] wl[126] vdd gnd cell_6t
Xbit_r127_c43 bl[43] br[43] wl[127] vdd gnd cell_6t
Xbit_r128_c43 bl[43] br[43] wl[128] vdd gnd cell_6t
Xbit_r129_c43 bl[43] br[43] wl[129] vdd gnd cell_6t
Xbit_r130_c43 bl[43] br[43] wl[130] vdd gnd cell_6t
Xbit_r131_c43 bl[43] br[43] wl[131] vdd gnd cell_6t
Xbit_r132_c43 bl[43] br[43] wl[132] vdd gnd cell_6t
Xbit_r133_c43 bl[43] br[43] wl[133] vdd gnd cell_6t
Xbit_r134_c43 bl[43] br[43] wl[134] vdd gnd cell_6t
Xbit_r135_c43 bl[43] br[43] wl[135] vdd gnd cell_6t
Xbit_r136_c43 bl[43] br[43] wl[136] vdd gnd cell_6t
Xbit_r137_c43 bl[43] br[43] wl[137] vdd gnd cell_6t
Xbit_r138_c43 bl[43] br[43] wl[138] vdd gnd cell_6t
Xbit_r139_c43 bl[43] br[43] wl[139] vdd gnd cell_6t
Xbit_r140_c43 bl[43] br[43] wl[140] vdd gnd cell_6t
Xbit_r141_c43 bl[43] br[43] wl[141] vdd gnd cell_6t
Xbit_r142_c43 bl[43] br[43] wl[142] vdd gnd cell_6t
Xbit_r143_c43 bl[43] br[43] wl[143] vdd gnd cell_6t
Xbit_r144_c43 bl[43] br[43] wl[144] vdd gnd cell_6t
Xbit_r145_c43 bl[43] br[43] wl[145] vdd gnd cell_6t
Xbit_r146_c43 bl[43] br[43] wl[146] vdd gnd cell_6t
Xbit_r147_c43 bl[43] br[43] wl[147] vdd gnd cell_6t
Xbit_r148_c43 bl[43] br[43] wl[148] vdd gnd cell_6t
Xbit_r149_c43 bl[43] br[43] wl[149] vdd gnd cell_6t
Xbit_r150_c43 bl[43] br[43] wl[150] vdd gnd cell_6t
Xbit_r151_c43 bl[43] br[43] wl[151] vdd gnd cell_6t
Xbit_r152_c43 bl[43] br[43] wl[152] vdd gnd cell_6t
Xbit_r153_c43 bl[43] br[43] wl[153] vdd gnd cell_6t
Xbit_r154_c43 bl[43] br[43] wl[154] vdd gnd cell_6t
Xbit_r155_c43 bl[43] br[43] wl[155] vdd gnd cell_6t
Xbit_r156_c43 bl[43] br[43] wl[156] vdd gnd cell_6t
Xbit_r157_c43 bl[43] br[43] wl[157] vdd gnd cell_6t
Xbit_r158_c43 bl[43] br[43] wl[158] vdd gnd cell_6t
Xbit_r159_c43 bl[43] br[43] wl[159] vdd gnd cell_6t
Xbit_r160_c43 bl[43] br[43] wl[160] vdd gnd cell_6t
Xbit_r161_c43 bl[43] br[43] wl[161] vdd gnd cell_6t
Xbit_r162_c43 bl[43] br[43] wl[162] vdd gnd cell_6t
Xbit_r163_c43 bl[43] br[43] wl[163] vdd gnd cell_6t
Xbit_r164_c43 bl[43] br[43] wl[164] vdd gnd cell_6t
Xbit_r165_c43 bl[43] br[43] wl[165] vdd gnd cell_6t
Xbit_r166_c43 bl[43] br[43] wl[166] vdd gnd cell_6t
Xbit_r167_c43 bl[43] br[43] wl[167] vdd gnd cell_6t
Xbit_r168_c43 bl[43] br[43] wl[168] vdd gnd cell_6t
Xbit_r169_c43 bl[43] br[43] wl[169] vdd gnd cell_6t
Xbit_r170_c43 bl[43] br[43] wl[170] vdd gnd cell_6t
Xbit_r171_c43 bl[43] br[43] wl[171] vdd gnd cell_6t
Xbit_r172_c43 bl[43] br[43] wl[172] vdd gnd cell_6t
Xbit_r173_c43 bl[43] br[43] wl[173] vdd gnd cell_6t
Xbit_r174_c43 bl[43] br[43] wl[174] vdd gnd cell_6t
Xbit_r175_c43 bl[43] br[43] wl[175] vdd gnd cell_6t
Xbit_r176_c43 bl[43] br[43] wl[176] vdd gnd cell_6t
Xbit_r177_c43 bl[43] br[43] wl[177] vdd gnd cell_6t
Xbit_r178_c43 bl[43] br[43] wl[178] vdd gnd cell_6t
Xbit_r179_c43 bl[43] br[43] wl[179] vdd gnd cell_6t
Xbit_r180_c43 bl[43] br[43] wl[180] vdd gnd cell_6t
Xbit_r181_c43 bl[43] br[43] wl[181] vdd gnd cell_6t
Xbit_r182_c43 bl[43] br[43] wl[182] vdd gnd cell_6t
Xbit_r183_c43 bl[43] br[43] wl[183] vdd gnd cell_6t
Xbit_r184_c43 bl[43] br[43] wl[184] vdd gnd cell_6t
Xbit_r185_c43 bl[43] br[43] wl[185] vdd gnd cell_6t
Xbit_r186_c43 bl[43] br[43] wl[186] vdd gnd cell_6t
Xbit_r187_c43 bl[43] br[43] wl[187] vdd gnd cell_6t
Xbit_r188_c43 bl[43] br[43] wl[188] vdd gnd cell_6t
Xbit_r189_c43 bl[43] br[43] wl[189] vdd gnd cell_6t
Xbit_r190_c43 bl[43] br[43] wl[190] vdd gnd cell_6t
Xbit_r191_c43 bl[43] br[43] wl[191] vdd gnd cell_6t
Xbit_r192_c43 bl[43] br[43] wl[192] vdd gnd cell_6t
Xbit_r193_c43 bl[43] br[43] wl[193] vdd gnd cell_6t
Xbit_r194_c43 bl[43] br[43] wl[194] vdd gnd cell_6t
Xbit_r195_c43 bl[43] br[43] wl[195] vdd gnd cell_6t
Xbit_r196_c43 bl[43] br[43] wl[196] vdd gnd cell_6t
Xbit_r197_c43 bl[43] br[43] wl[197] vdd gnd cell_6t
Xbit_r198_c43 bl[43] br[43] wl[198] vdd gnd cell_6t
Xbit_r199_c43 bl[43] br[43] wl[199] vdd gnd cell_6t
Xbit_r200_c43 bl[43] br[43] wl[200] vdd gnd cell_6t
Xbit_r201_c43 bl[43] br[43] wl[201] vdd gnd cell_6t
Xbit_r202_c43 bl[43] br[43] wl[202] vdd gnd cell_6t
Xbit_r203_c43 bl[43] br[43] wl[203] vdd gnd cell_6t
Xbit_r204_c43 bl[43] br[43] wl[204] vdd gnd cell_6t
Xbit_r205_c43 bl[43] br[43] wl[205] vdd gnd cell_6t
Xbit_r206_c43 bl[43] br[43] wl[206] vdd gnd cell_6t
Xbit_r207_c43 bl[43] br[43] wl[207] vdd gnd cell_6t
Xbit_r208_c43 bl[43] br[43] wl[208] vdd gnd cell_6t
Xbit_r209_c43 bl[43] br[43] wl[209] vdd gnd cell_6t
Xbit_r210_c43 bl[43] br[43] wl[210] vdd gnd cell_6t
Xbit_r211_c43 bl[43] br[43] wl[211] vdd gnd cell_6t
Xbit_r212_c43 bl[43] br[43] wl[212] vdd gnd cell_6t
Xbit_r213_c43 bl[43] br[43] wl[213] vdd gnd cell_6t
Xbit_r214_c43 bl[43] br[43] wl[214] vdd gnd cell_6t
Xbit_r215_c43 bl[43] br[43] wl[215] vdd gnd cell_6t
Xbit_r216_c43 bl[43] br[43] wl[216] vdd gnd cell_6t
Xbit_r217_c43 bl[43] br[43] wl[217] vdd gnd cell_6t
Xbit_r218_c43 bl[43] br[43] wl[218] vdd gnd cell_6t
Xbit_r219_c43 bl[43] br[43] wl[219] vdd gnd cell_6t
Xbit_r220_c43 bl[43] br[43] wl[220] vdd gnd cell_6t
Xbit_r221_c43 bl[43] br[43] wl[221] vdd gnd cell_6t
Xbit_r222_c43 bl[43] br[43] wl[222] vdd gnd cell_6t
Xbit_r223_c43 bl[43] br[43] wl[223] vdd gnd cell_6t
Xbit_r224_c43 bl[43] br[43] wl[224] vdd gnd cell_6t
Xbit_r225_c43 bl[43] br[43] wl[225] vdd gnd cell_6t
Xbit_r226_c43 bl[43] br[43] wl[226] vdd gnd cell_6t
Xbit_r227_c43 bl[43] br[43] wl[227] vdd gnd cell_6t
Xbit_r228_c43 bl[43] br[43] wl[228] vdd gnd cell_6t
Xbit_r229_c43 bl[43] br[43] wl[229] vdd gnd cell_6t
Xbit_r230_c43 bl[43] br[43] wl[230] vdd gnd cell_6t
Xbit_r231_c43 bl[43] br[43] wl[231] vdd gnd cell_6t
Xbit_r232_c43 bl[43] br[43] wl[232] vdd gnd cell_6t
Xbit_r233_c43 bl[43] br[43] wl[233] vdd gnd cell_6t
Xbit_r234_c43 bl[43] br[43] wl[234] vdd gnd cell_6t
Xbit_r235_c43 bl[43] br[43] wl[235] vdd gnd cell_6t
Xbit_r236_c43 bl[43] br[43] wl[236] vdd gnd cell_6t
Xbit_r237_c43 bl[43] br[43] wl[237] vdd gnd cell_6t
Xbit_r238_c43 bl[43] br[43] wl[238] vdd gnd cell_6t
Xbit_r239_c43 bl[43] br[43] wl[239] vdd gnd cell_6t
Xbit_r240_c43 bl[43] br[43] wl[240] vdd gnd cell_6t
Xbit_r241_c43 bl[43] br[43] wl[241] vdd gnd cell_6t
Xbit_r242_c43 bl[43] br[43] wl[242] vdd gnd cell_6t
Xbit_r243_c43 bl[43] br[43] wl[243] vdd gnd cell_6t
Xbit_r244_c43 bl[43] br[43] wl[244] vdd gnd cell_6t
Xbit_r245_c43 bl[43] br[43] wl[245] vdd gnd cell_6t
Xbit_r246_c43 bl[43] br[43] wl[246] vdd gnd cell_6t
Xbit_r247_c43 bl[43] br[43] wl[247] vdd gnd cell_6t
Xbit_r248_c43 bl[43] br[43] wl[248] vdd gnd cell_6t
Xbit_r249_c43 bl[43] br[43] wl[249] vdd gnd cell_6t
Xbit_r250_c43 bl[43] br[43] wl[250] vdd gnd cell_6t
Xbit_r251_c43 bl[43] br[43] wl[251] vdd gnd cell_6t
Xbit_r252_c43 bl[43] br[43] wl[252] vdd gnd cell_6t
Xbit_r253_c43 bl[43] br[43] wl[253] vdd gnd cell_6t
Xbit_r254_c43 bl[43] br[43] wl[254] vdd gnd cell_6t
Xbit_r255_c43 bl[43] br[43] wl[255] vdd gnd cell_6t
Xbit_r0_c44 bl[44] br[44] wl[0] vdd gnd cell_6t
Xbit_r1_c44 bl[44] br[44] wl[1] vdd gnd cell_6t
Xbit_r2_c44 bl[44] br[44] wl[2] vdd gnd cell_6t
Xbit_r3_c44 bl[44] br[44] wl[3] vdd gnd cell_6t
Xbit_r4_c44 bl[44] br[44] wl[4] vdd gnd cell_6t
Xbit_r5_c44 bl[44] br[44] wl[5] vdd gnd cell_6t
Xbit_r6_c44 bl[44] br[44] wl[6] vdd gnd cell_6t
Xbit_r7_c44 bl[44] br[44] wl[7] vdd gnd cell_6t
Xbit_r8_c44 bl[44] br[44] wl[8] vdd gnd cell_6t
Xbit_r9_c44 bl[44] br[44] wl[9] vdd gnd cell_6t
Xbit_r10_c44 bl[44] br[44] wl[10] vdd gnd cell_6t
Xbit_r11_c44 bl[44] br[44] wl[11] vdd gnd cell_6t
Xbit_r12_c44 bl[44] br[44] wl[12] vdd gnd cell_6t
Xbit_r13_c44 bl[44] br[44] wl[13] vdd gnd cell_6t
Xbit_r14_c44 bl[44] br[44] wl[14] vdd gnd cell_6t
Xbit_r15_c44 bl[44] br[44] wl[15] vdd gnd cell_6t
Xbit_r16_c44 bl[44] br[44] wl[16] vdd gnd cell_6t
Xbit_r17_c44 bl[44] br[44] wl[17] vdd gnd cell_6t
Xbit_r18_c44 bl[44] br[44] wl[18] vdd gnd cell_6t
Xbit_r19_c44 bl[44] br[44] wl[19] vdd gnd cell_6t
Xbit_r20_c44 bl[44] br[44] wl[20] vdd gnd cell_6t
Xbit_r21_c44 bl[44] br[44] wl[21] vdd gnd cell_6t
Xbit_r22_c44 bl[44] br[44] wl[22] vdd gnd cell_6t
Xbit_r23_c44 bl[44] br[44] wl[23] vdd gnd cell_6t
Xbit_r24_c44 bl[44] br[44] wl[24] vdd gnd cell_6t
Xbit_r25_c44 bl[44] br[44] wl[25] vdd gnd cell_6t
Xbit_r26_c44 bl[44] br[44] wl[26] vdd gnd cell_6t
Xbit_r27_c44 bl[44] br[44] wl[27] vdd gnd cell_6t
Xbit_r28_c44 bl[44] br[44] wl[28] vdd gnd cell_6t
Xbit_r29_c44 bl[44] br[44] wl[29] vdd gnd cell_6t
Xbit_r30_c44 bl[44] br[44] wl[30] vdd gnd cell_6t
Xbit_r31_c44 bl[44] br[44] wl[31] vdd gnd cell_6t
Xbit_r32_c44 bl[44] br[44] wl[32] vdd gnd cell_6t
Xbit_r33_c44 bl[44] br[44] wl[33] vdd gnd cell_6t
Xbit_r34_c44 bl[44] br[44] wl[34] vdd gnd cell_6t
Xbit_r35_c44 bl[44] br[44] wl[35] vdd gnd cell_6t
Xbit_r36_c44 bl[44] br[44] wl[36] vdd gnd cell_6t
Xbit_r37_c44 bl[44] br[44] wl[37] vdd gnd cell_6t
Xbit_r38_c44 bl[44] br[44] wl[38] vdd gnd cell_6t
Xbit_r39_c44 bl[44] br[44] wl[39] vdd gnd cell_6t
Xbit_r40_c44 bl[44] br[44] wl[40] vdd gnd cell_6t
Xbit_r41_c44 bl[44] br[44] wl[41] vdd gnd cell_6t
Xbit_r42_c44 bl[44] br[44] wl[42] vdd gnd cell_6t
Xbit_r43_c44 bl[44] br[44] wl[43] vdd gnd cell_6t
Xbit_r44_c44 bl[44] br[44] wl[44] vdd gnd cell_6t
Xbit_r45_c44 bl[44] br[44] wl[45] vdd gnd cell_6t
Xbit_r46_c44 bl[44] br[44] wl[46] vdd gnd cell_6t
Xbit_r47_c44 bl[44] br[44] wl[47] vdd gnd cell_6t
Xbit_r48_c44 bl[44] br[44] wl[48] vdd gnd cell_6t
Xbit_r49_c44 bl[44] br[44] wl[49] vdd gnd cell_6t
Xbit_r50_c44 bl[44] br[44] wl[50] vdd gnd cell_6t
Xbit_r51_c44 bl[44] br[44] wl[51] vdd gnd cell_6t
Xbit_r52_c44 bl[44] br[44] wl[52] vdd gnd cell_6t
Xbit_r53_c44 bl[44] br[44] wl[53] vdd gnd cell_6t
Xbit_r54_c44 bl[44] br[44] wl[54] vdd gnd cell_6t
Xbit_r55_c44 bl[44] br[44] wl[55] vdd gnd cell_6t
Xbit_r56_c44 bl[44] br[44] wl[56] vdd gnd cell_6t
Xbit_r57_c44 bl[44] br[44] wl[57] vdd gnd cell_6t
Xbit_r58_c44 bl[44] br[44] wl[58] vdd gnd cell_6t
Xbit_r59_c44 bl[44] br[44] wl[59] vdd gnd cell_6t
Xbit_r60_c44 bl[44] br[44] wl[60] vdd gnd cell_6t
Xbit_r61_c44 bl[44] br[44] wl[61] vdd gnd cell_6t
Xbit_r62_c44 bl[44] br[44] wl[62] vdd gnd cell_6t
Xbit_r63_c44 bl[44] br[44] wl[63] vdd gnd cell_6t
Xbit_r64_c44 bl[44] br[44] wl[64] vdd gnd cell_6t
Xbit_r65_c44 bl[44] br[44] wl[65] vdd gnd cell_6t
Xbit_r66_c44 bl[44] br[44] wl[66] vdd gnd cell_6t
Xbit_r67_c44 bl[44] br[44] wl[67] vdd gnd cell_6t
Xbit_r68_c44 bl[44] br[44] wl[68] vdd gnd cell_6t
Xbit_r69_c44 bl[44] br[44] wl[69] vdd gnd cell_6t
Xbit_r70_c44 bl[44] br[44] wl[70] vdd gnd cell_6t
Xbit_r71_c44 bl[44] br[44] wl[71] vdd gnd cell_6t
Xbit_r72_c44 bl[44] br[44] wl[72] vdd gnd cell_6t
Xbit_r73_c44 bl[44] br[44] wl[73] vdd gnd cell_6t
Xbit_r74_c44 bl[44] br[44] wl[74] vdd gnd cell_6t
Xbit_r75_c44 bl[44] br[44] wl[75] vdd gnd cell_6t
Xbit_r76_c44 bl[44] br[44] wl[76] vdd gnd cell_6t
Xbit_r77_c44 bl[44] br[44] wl[77] vdd gnd cell_6t
Xbit_r78_c44 bl[44] br[44] wl[78] vdd gnd cell_6t
Xbit_r79_c44 bl[44] br[44] wl[79] vdd gnd cell_6t
Xbit_r80_c44 bl[44] br[44] wl[80] vdd gnd cell_6t
Xbit_r81_c44 bl[44] br[44] wl[81] vdd gnd cell_6t
Xbit_r82_c44 bl[44] br[44] wl[82] vdd gnd cell_6t
Xbit_r83_c44 bl[44] br[44] wl[83] vdd gnd cell_6t
Xbit_r84_c44 bl[44] br[44] wl[84] vdd gnd cell_6t
Xbit_r85_c44 bl[44] br[44] wl[85] vdd gnd cell_6t
Xbit_r86_c44 bl[44] br[44] wl[86] vdd gnd cell_6t
Xbit_r87_c44 bl[44] br[44] wl[87] vdd gnd cell_6t
Xbit_r88_c44 bl[44] br[44] wl[88] vdd gnd cell_6t
Xbit_r89_c44 bl[44] br[44] wl[89] vdd gnd cell_6t
Xbit_r90_c44 bl[44] br[44] wl[90] vdd gnd cell_6t
Xbit_r91_c44 bl[44] br[44] wl[91] vdd gnd cell_6t
Xbit_r92_c44 bl[44] br[44] wl[92] vdd gnd cell_6t
Xbit_r93_c44 bl[44] br[44] wl[93] vdd gnd cell_6t
Xbit_r94_c44 bl[44] br[44] wl[94] vdd gnd cell_6t
Xbit_r95_c44 bl[44] br[44] wl[95] vdd gnd cell_6t
Xbit_r96_c44 bl[44] br[44] wl[96] vdd gnd cell_6t
Xbit_r97_c44 bl[44] br[44] wl[97] vdd gnd cell_6t
Xbit_r98_c44 bl[44] br[44] wl[98] vdd gnd cell_6t
Xbit_r99_c44 bl[44] br[44] wl[99] vdd gnd cell_6t
Xbit_r100_c44 bl[44] br[44] wl[100] vdd gnd cell_6t
Xbit_r101_c44 bl[44] br[44] wl[101] vdd gnd cell_6t
Xbit_r102_c44 bl[44] br[44] wl[102] vdd gnd cell_6t
Xbit_r103_c44 bl[44] br[44] wl[103] vdd gnd cell_6t
Xbit_r104_c44 bl[44] br[44] wl[104] vdd gnd cell_6t
Xbit_r105_c44 bl[44] br[44] wl[105] vdd gnd cell_6t
Xbit_r106_c44 bl[44] br[44] wl[106] vdd gnd cell_6t
Xbit_r107_c44 bl[44] br[44] wl[107] vdd gnd cell_6t
Xbit_r108_c44 bl[44] br[44] wl[108] vdd gnd cell_6t
Xbit_r109_c44 bl[44] br[44] wl[109] vdd gnd cell_6t
Xbit_r110_c44 bl[44] br[44] wl[110] vdd gnd cell_6t
Xbit_r111_c44 bl[44] br[44] wl[111] vdd gnd cell_6t
Xbit_r112_c44 bl[44] br[44] wl[112] vdd gnd cell_6t
Xbit_r113_c44 bl[44] br[44] wl[113] vdd gnd cell_6t
Xbit_r114_c44 bl[44] br[44] wl[114] vdd gnd cell_6t
Xbit_r115_c44 bl[44] br[44] wl[115] vdd gnd cell_6t
Xbit_r116_c44 bl[44] br[44] wl[116] vdd gnd cell_6t
Xbit_r117_c44 bl[44] br[44] wl[117] vdd gnd cell_6t
Xbit_r118_c44 bl[44] br[44] wl[118] vdd gnd cell_6t
Xbit_r119_c44 bl[44] br[44] wl[119] vdd gnd cell_6t
Xbit_r120_c44 bl[44] br[44] wl[120] vdd gnd cell_6t
Xbit_r121_c44 bl[44] br[44] wl[121] vdd gnd cell_6t
Xbit_r122_c44 bl[44] br[44] wl[122] vdd gnd cell_6t
Xbit_r123_c44 bl[44] br[44] wl[123] vdd gnd cell_6t
Xbit_r124_c44 bl[44] br[44] wl[124] vdd gnd cell_6t
Xbit_r125_c44 bl[44] br[44] wl[125] vdd gnd cell_6t
Xbit_r126_c44 bl[44] br[44] wl[126] vdd gnd cell_6t
Xbit_r127_c44 bl[44] br[44] wl[127] vdd gnd cell_6t
Xbit_r128_c44 bl[44] br[44] wl[128] vdd gnd cell_6t
Xbit_r129_c44 bl[44] br[44] wl[129] vdd gnd cell_6t
Xbit_r130_c44 bl[44] br[44] wl[130] vdd gnd cell_6t
Xbit_r131_c44 bl[44] br[44] wl[131] vdd gnd cell_6t
Xbit_r132_c44 bl[44] br[44] wl[132] vdd gnd cell_6t
Xbit_r133_c44 bl[44] br[44] wl[133] vdd gnd cell_6t
Xbit_r134_c44 bl[44] br[44] wl[134] vdd gnd cell_6t
Xbit_r135_c44 bl[44] br[44] wl[135] vdd gnd cell_6t
Xbit_r136_c44 bl[44] br[44] wl[136] vdd gnd cell_6t
Xbit_r137_c44 bl[44] br[44] wl[137] vdd gnd cell_6t
Xbit_r138_c44 bl[44] br[44] wl[138] vdd gnd cell_6t
Xbit_r139_c44 bl[44] br[44] wl[139] vdd gnd cell_6t
Xbit_r140_c44 bl[44] br[44] wl[140] vdd gnd cell_6t
Xbit_r141_c44 bl[44] br[44] wl[141] vdd gnd cell_6t
Xbit_r142_c44 bl[44] br[44] wl[142] vdd gnd cell_6t
Xbit_r143_c44 bl[44] br[44] wl[143] vdd gnd cell_6t
Xbit_r144_c44 bl[44] br[44] wl[144] vdd gnd cell_6t
Xbit_r145_c44 bl[44] br[44] wl[145] vdd gnd cell_6t
Xbit_r146_c44 bl[44] br[44] wl[146] vdd gnd cell_6t
Xbit_r147_c44 bl[44] br[44] wl[147] vdd gnd cell_6t
Xbit_r148_c44 bl[44] br[44] wl[148] vdd gnd cell_6t
Xbit_r149_c44 bl[44] br[44] wl[149] vdd gnd cell_6t
Xbit_r150_c44 bl[44] br[44] wl[150] vdd gnd cell_6t
Xbit_r151_c44 bl[44] br[44] wl[151] vdd gnd cell_6t
Xbit_r152_c44 bl[44] br[44] wl[152] vdd gnd cell_6t
Xbit_r153_c44 bl[44] br[44] wl[153] vdd gnd cell_6t
Xbit_r154_c44 bl[44] br[44] wl[154] vdd gnd cell_6t
Xbit_r155_c44 bl[44] br[44] wl[155] vdd gnd cell_6t
Xbit_r156_c44 bl[44] br[44] wl[156] vdd gnd cell_6t
Xbit_r157_c44 bl[44] br[44] wl[157] vdd gnd cell_6t
Xbit_r158_c44 bl[44] br[44] wl[158] vdd gnd cell_6t
Xbit_r159_c44 bl[44] br[44] wl[159] vdd gnd cell_6t
Xbit_r160_c44 bl[44] br[44] wl[160] vdd gnd cell_6t
Xbit_r161_c44 bl[44] br[44] wl[161] vdd gnd cell_6t
Xbit_r162_c44 bl[44] br[44] wl[162] vdd gnd cell_6t
Xbit_r163_c44 bl[44] br[44] wl[163] vdd gnd cell_6t
Xbit_r164_c44 bl[44] br[44] wl[164] vdd gnd cell_6t
Xbit_r165_c44 bl[44] br[44] wl[165] vdd gnd cell_6t
Xbit_r166_c44 bl[44] br[44] wl[166] vdd gnd cell_6t
Xbit_r167_c44 bl[44] br[44] wl[167] vdd gnd cell_6t
Xbit_r168_c44 bl[44] br[44] wl[168] vdd gnd cell_6t
Xbit_r169_c44 bl[44] br[44] wl[169] vdd gnd cell_6t
Xbit_r170_c44 bl[44] br[44] wl[170] vdd gnd cell_6t
Xbit_r171_c44 bl[44] br[44] wl[171] vdd gnd cell_6t
Xbit_r172_c44 bl[44] br[44] wl[172] vdd gnd cell_6t
Xbit_r173_c44 bl[44] br[44] wl[173] vdd gnd cell_6t
Xbit_r174_c44 bl[44] br[44] wl[174] vdd gnd cell_6t
Xbit_r175_c44 bl[44] br[44] wl[175] vdd gnd cell_6t
Xbit_r176_c44 bl[44] br[44] wl[176] vdd gnd cell_6t
Xbit_r177_c44 bl[44] br[44] wl[177] vdd gnd cell_6t
Xbit_r178_c44 bl[44] br[44] wl[178] vdd gnd cell_6t
Xbit_r179_c44 bl[44] br[44] wl[179] vdd gnd cell_6t
Xbit_r180_c44 bl[44] br[44] wl[180] vdd gnd cell_6t
Xbit_r181_c44 bl[44] br[44] wl[181] vdd gnd cell_6t
Xbit_r182_c44 bl[44] br[44] wl[182] vdd gnd cell_6t
Xbit_r183_c44 bl[44] br[44] wl[183] vdd gnd cell_6t
Xbit_r184_c44 bl[44] br[44] wl[184] vdd gnd cell_6t
Xbit_r185_c44 bl[44] br[44] wl[185] vdd gnd cell_6t
Xbit_r186_c44 bl[44] br[44] wl[186] vdd gnd cell_6t
Xbit_r187_c44 bl[44] br[44] wl[187] vdd gnd cell_6t
Xbit_r188_c44 bl[44] br[44] wl[188] vdd gnd cell_6t
Xbit_r189_c44 bl[44] br[44] wl[189] vdd gnd cell_6t
Xbit_r190_c44 bl[44] br[44] wl[190] vdd gnd cell_6t
Xbit_r191_c44 bl[44] br[44] wl[191] vdd gnd cell_6t
Xbit_r192_c44 bl[44] br[44] wl[192] vdd gnd cell_6t
Xbit_r193_c44 bl[44] br[44] wl[193] vdd gnd cell_6t
Xbit_r194_c44 bl[44] br[44] wl[194] vdd gnd cell_6t
Xbit_r195_c44 bl[44] br[44] wl[195] vdd gnd cell_6t
Xbit_r196_c44 bl[44] br[44] wl[196] vdd gnd cell_6t
Xbit_r197_c44 bl[44] br[44] wl[197] vdd gnd cell_6t
Xbit_r198_c44 bl[44] br[44] wl[198] vdd gnd cell_6t
Xbit_r199_c44 bl[44] br[44] wl[199] vdd gnd cell_6t
Xbit_r200_c44 bl[44] br[44] wl[200] vdd gnd cell_6t
Xbit_r201_c44 bl[44] br[44] wl[201] vdd gnd cell_6t
Xbit_r202_c44 bl[44] br[44] wl[202] vdd gnd cell_6t
Xbit_r203_c44 bl[44] br[44] wl[203] vdd gnd cell_6t
Xbit_r204_c44 bl[44] br[44] wl[204] vdd gnd cell_6t
Xbit_r205_c44 bl[44] br[44] wl[205] vdd gnd cell_6t
Xbit_r206_c44 bl[44] br[44] wl[206] vdd gnd cell_6t
Xbit_r207_c44 bl[44] br[44] wl[207] vdd gnd cell_6t
Xbit_r208_c44 bl[44] br[44] wl[208] vdd gnd cell_6t
Xbit_r209_c44 bl[44] br[44] wl[209] vdd gnd cell_6t
Xbit_r210_c44 bl[44] br[44] wl[210] vdd gnd cell_6t
Xbit_r211_c44 bl[44] br[44] wl[211] vdd gnd cell_6t
Xbit_r212_c44 bl[44] br[44] wl[212] vdd gnd cell_6t
Xbit_r213_c44 bl[44] br[44] wl[213] vdd gnd cell_6t
Xbit_r214_c44 bl[44] br[44] wl[214] vdd gnd cell_6t
Xbit_r215_c44 bl[44] br[44] wl[215] vdd gnd cell_6t
Xbit_r216_c44 bl[44] br[44] wl[216] vdd gnd cell_6t
Xbit_r217_c44 bl[44] br[44] wl[217] vdd gnd cell_6t
Xbit_r218_c44 bl[44] br[44] wl[218] vdd gnd cell_6t
Xbit_r219_c44 bl[44] br[44] wl[219] vdd gnd cell_6t
Xbit_r220_c44 bl[44] br[44] wl[220] vdd gnd cell_6t
Xbit_r221_c44 bl[44] br[44] wl[221] vdd gnd cell_6t
Xbit_r222_c44 bl[44] br[44] wl[222] vdd gnd cell_6t
Xbit_r223_c44 bl[44] br[44] wl[223] vdd gnd cell_6t
Xbit_r224_c44 bl[44] br[44] wl[224] vdd gnd cell_6t
Xbit_r225_c44 bl[44] br[44] wl[225] vdd gnd cell_6t
Xbit_r226_c44 bl[44] br[44] wl[226] vdd gnd cell_6t
Xbit_r227_c44 bl[44] br[44] wl[227] vdd gnd cell_6t
Xbit_r228_c44 bl[44] br[44] wl[228] vdd gnd cell_6t
Xbit_r229_c44 bl[44] br[44] wl[229] vdd gnd cell_6t
Xbit_r230_c44 bl[44] br[44] wl[230] vdd gnd cell_6t
Xbit_r231_c44 bl[44] br[44] wl[231] vdd gnd cell_6t
Xbit_r232_c44 bl[44] br[44] wl[232] vdd gnd cell_6t
Xbit_r233_c44 bl[44] br[44] wl[233] vdd gnd cell_6t
Xbit_r234_c44 bl[44] br[44] wl[234] vdd gnd cell_6t
Xbit_r235_c44 bl[44] br[44] wl[235] vdd gnd cell_6t
Xbit_r236_c44 bl[44] br[44] wl[236] vdd gnd cell_6t
Xbit_r237_c44 bl[44] br[44] wl[237] vdd gnd cell_6t
Xbit_r238_c44 bl[44] br[44] wl[238] vdd gnd cell_6t
Xbit_r239_c44 bl[44] br[44] wl[239] vdd gnd cell_6t
Xbit_r240_c44 bl[44] br[44] wl[240] vdd gnd cell_6t
Xbit_r241_c44 bl[44] br[44] wl[241] vdd gnd cell_6t
Xbit_r242_c44 bl[44] br[44] wl[242] vdd gnd cell_6t
Xbit_r243_c44 bl[44] br[44] wl[243] vdd gnd cell_6t
Xbit_r244_c44 bl[44] br[44] wl[244] vdd gnd cell_6t
Xbit_r245_c44 bl[44] br[44] wl[245] vdd gnd cell_6t
Xbit_r246_c44 bl[44] br[44] wl[246] vdd gnd cell_6t
Xbit_r247_c44 bl[44] br[44] wl[247] vdd gnd cell_6t
Xbit_r248_c44 bl[44] br[44] wl[248] vdd gnd cell_6t
Xbit_r249_c44 bl[44] br[44] wl[249] vdd gnd cell_6t
Xbit_r250_c44 bl[44] br[44] wl[250] vdd gnd cell_6t
Xbit_r251_c44 bl[44] br[44] wl[251] vdd gnd cell_6t
Xbit_r252_c44 bl[44] br[44] wl[252] vdd gnd cell_6t
Xbit_r253_c44 bl[44] br[44] wl[253] vdd gnd cell_6t
Xbit_r254_c44 bl[44] br[44] wl[254] vdd gnd cell_6t
Xbit_r255_c44 bl[44] br[44] wl[255] vdd gnd cell_6t
Xbit_r0_c45 bl[45] br[45] wl[0] vdd gnd cell_6t
Xbit_r1_c45 bl[45] br[45] wl[1] vdd gnd cell_6t
Xbit_r2_c45 bl[45] br[45] wl[2] vdd gnd cell_6t
Xbit_r3_c45 bl[45] br[45] wl[3] vdd gnd cell_6t
Xbit_r4_c45 bl[45] br[45] wl[4] vdd gnd cell_6t
Xbit_r5_c45 bl[45] br[45] wl[5] vdd gnd cell_6t
Xbit_r6_c45 bl[45] br[45] wl[6] vdd gnd cell_6t
Xbit_r7_c45 bl[45] br[45] wl[7] vdd gnd cell_6t
Xbit_r8_c45 bl[45] br[45] wl[8] vdd gnd cell_6t
Xbit_r9_c45 bl[45] br[45] wl[9] vdd gnd cell_6t
Xbit_r10_c45 bl[45] br[45] wl[10] vdd gnd cell_6t
Xbit_r11_c45 bl[45] br[45] wl[11] vdd gnd cell_6t
Xbit_r12_c45 bl[45] br[45] wl[12] vdd gnd cell_6t
Xbit_r13_c45 bl[45] br[45] wl[13] vdd gnd cell_6t
Xbit_r14_c45 bl[45] br[45] wl[14] vdd gnd cell_6t
Xbit_r15_c45 bl[45] br[45] wl[15] vdd gnd cell_6t
Xbit_r16_c45 bl[45] br[45] wl[16] vdd gnd cell_6t
Xbit_r17_c45 bl[45] br[45] wl[17] vdd gnd cell_6t
Xbit_r18_c45 bl[45] br[45] wl[18] vdd gnd cell_6t
Xbit_r19_c45 bl[45] br[45] wl[19] vdd gnd cell_6t
Xbit_r20_c45 bl[45] br[45] wl[20] vdd gnd cell_6t
Xbit_r21_c45 bl[45] br[45] wl[21] vdd gnd cell_6t
Xbit_r22_c45 bl[45] br[45] wl[22] vdd gnd cell_6t
Xbit_r23_c45 bl[45] br[45] wl[23] vdd gnd cell_6t
Xbit_r24_c45 bl[45] br[45] wl[24] vdd gnd cell_6t
Xbit_r25_c45 bl[45] br[45] wl[25] vdd gnd cell_6t
Xbit_r26_c45 bl[45] br[45] wl[26] vdd gnd cell_6t
Xbit_r27_c45 bl[45] br[45] wl[27] vdd gnd cell_6t
Xbit_r28_c45 bl[45] br[45] wl[28] vdd gnd cell_6t
Xbit_r29_c45 bl[45] br[45] wl[29] vdd gnd cell_6t
Xbit_r30_c45 bl[45] br[45] wl[30] vdd gnd cell_6t
Xbit_r31_c45 bl[45] br[45] wl[31] vdd gnd cell_6t
Xbit_r32_c45 bl[45] br[45] wl[32] vdd gnd cell_6t
Xbit_r33_c45 bl[45] br[45] wl[33] vdd gnd cell_6t
Xbit_r34_c45 bl[45] br[45] wl[34] vdd gnd cell_6t
Xbit_r35_c45 bl[45] br[45] wl[35] vdd gnd cell_6t
Xbit_r36_c45 bl[45] br[45] wl[36] vdd gnd cell_6t
Xbit_r37_c45 bl[45] br[45] wl[37] vdd gnd cell_6t
Xbit_r38_c45 bl[45] br[45] wl[38] vdd gnd cell_6t
Xbit_r39_c45 bl[45] br[45] wl[39] vdd gnd cell_6t
Xbit_r40_c45 bl[45] br[45] wl[40] vdd gnd cell_6t
Xbit_r41_c45 bl[45] br[45] wl[41] vdd gnd cell_6t
Xbit_r42_c45 bl[45] br[45] wl[42] vdd gnd cell_6t
Xbit_r43_c45 bl[45] br[45] wl[43] vdd gnd cell_6t
Xbit_r44_c45 bl[45] br[45] wl[44] vdd gnd cell_6t
Xbit_r45_c45 bl[45] br[45] wl[45] vdd gnd cell_6t
Xbit_r46_c45 bl[45] br[45] wl[46] vdd gnd cell_6t
Xbit_r47_c45 bl[45] br[45] wl[47] vdd gnd cell_6t
Xbit_r48_c45 bl[45] br[45] wl[48] vdd gnd cell_6t
Xbit_r49_c45 bl[45] br[45] wl[49] vdd gnd cell_6t
Xbit_r50_c45 bl[45] br[45] wl[50] vdd gnd cell_6t
Xbit_r51_c45 bl[45] br[45] wl[51] vdd gnd cell_6t
Xbit_r52_c45 bl[45] br[45] wl[52] vdd gnd cell_6t
Xbit_r53_c45 bl[45] br[45] wl[53] vdd gnd cell_6t
Xbit_r54_c45 bl[45] br[45] wl[54] vdd gnd cell_6t
Xbit_r55_c45 bl[45] br[45] wl[55] vdd gnd cell_6t
Xbit_r56_c45 bl[45] br[45] wl[56] vdd gnd cell_6t
Xbit_r57_c45 bl[45] br[45] wl[57] vdd gnd cell_6t
Xbit_r58_c45 bl[45] br[45] wl[58] vdd gnd cell_6t
Xbit_r59_c45 bl[45] br[45] wl[59] vdd gnd cell_6t
Xbit_r60_c45 bl[45] br[45] wl[60] vdd gnd cell_6t
Xbit_r61_c45 bl[45] br[45] wl[61] vdd gnd cell_6t
Xbit_r62_c45 bl[45] br[45] wl[62] vdd gnd cell_6t
Xbit_r63_c45 bl[45] br[45] wl[63] vdd gnd cell_6t
Xbit_r64_c45 bl[45] br[45] wl[64] vdd gnd cell_6t
Xbit_r65_c45 bl[45] br[45] wl[65] vdd gnd cell_6t
Xbit_r66_c45 bl[45] br[45] wl[66] vdd gnd cell_6t
Xbit_r67_c45 bl[45] br[45] wl[67] vdd gnd cell_6t
Xbit_r68_c45 bl[45] br[45] wl[68] vdd gnd cell_6t
Xbit_r69_c45 bl[45] br[45] wl[69] vdd gnd cell_6t
Xbit_r70_c45 bl[45] br[45] wl[70] vdd gnd cell_6t
Xbit_r71_c45 bl[45] br[45] wl[71] vdd gnd cell_6t
Xbit_r72_c45 bl[45] br[45] wl[72] vdd gnd cell_6t
Xbit_r73_c45 bl[45] br[45] wl[73] vdd gnd cell_6t
Xbit_r74_c45 bl[45] br[45] wl[74] vdd gnd cell_6t
Xbit_r75_c45 bl[45] br[45] wl[75] vdd gnd cell_6t
Xbit_r76_c45 bl[45] br[45] wl[76] vdd gnd cell_6t
Xbit_r77_c45 bl[45] br[45] wl[77] vdd gnd cell_6t
Xbit_r78_c45 bl[45] br[45] wl[78] vdd gnd cell_6t
Xbit_r79_c45 bl[45] br[45] wl[79] vdd gnd cell_6t
Xbit_r80_c45 bl[45] br[45] wl[80] vdd gnd cell_6t
Xbit_r81_c45 bl[45] br[45] wl[81] vdd gnd cell_6t
Xbit_r82_c45 bl[45] br[45] wl[82] vdd gnd cell_6t
Xbit_r83_c45 bl[45] br[45] wl[83] vdd gnd cell_6t
Xbit_r84_c45 bl[45] br[45] wl[84] vdd gnd cell_6t
Xbit_r85_c45 bl[45] br[45] wl[85] vdd gnd cell_6t
Xbit_r86_c45 bl[45] br[45] wl[86] vdd gnd cell_6t
Xbit_r87_c45 bl[45] br[45] wl[87] vdd gnd cell_6t
Xbit_r88_c45 bl[45] br[45] wl[88] vdd gnd cell_6t
Xbit_r89_c45 bl[45] br[45] wl[89] vdd gnd cell_6t
Xbit_r90_c45 bl[45] br[45] wl[90] vdd gnd cell_6t
Xbit_r91_c45 bl[45] br[45] wl[91] vdd gnd cell_6t
Xbit_r92_c45 bl[45] br[45] wl[92] vdd gnd cell_6t
Xbit_r93_c45 bl[45] br[45] wl[93] vdd gnd cell_6t
Xbit_r94_c45 bl[45] br[45] wl[94] vdd gnd cell_6t
Xbit_r95_c45 bl[45] br[45] wl[95] vdd gnd cell_6t
Xbit_r96_c45 bl[45] br[45] wl[96] vdd gnd cell_6t
Xbit_r97_c45 bl[45] br[45] wl[97] vdd gnd cell_6t
Xbit_r98_c45 bl[45] br[45] wl[98] vdd gnd cell_6t
Xbit_r99_c45 bl[45] br[45] wl[99] vdd gnd cell_6t
Xbit_r100_c45 bl[45] br[45] wl[100] vdd gnd cell_6t
Xbit_r101_c45 bl[45] br[45] wl[101] vdd gnd cell_6t
Xbit_r102_c45 bl[45] br[45] wl[102] vdd gnd cell_6t
Xbit_r103_c45 bl[45] br[45] wl[103] vdd gnd cell_6t
Xbit_r104_c45 bl[45] br[45] wl[104] vdd gnd cell_6t
Xbit_r105_c45 bl[45] br[45] wl[105] vdd gnd cell_6t
Xbit_r106_c45 bl[45] br[45] wl[106] vdd gnd cell_6t
Xbit_r107_c45 bl[45] br[45] wl[107] vdd gnd cell_6t
Xbit_r108_c45 bl[45] br[45] wl[108] vdd gnd cell_6t
Xbit_r109_c45 bl[45] br[45] wl[109] vdd gnd cell_6t
Xbit_r110_c45 bl[45] br[45] wl[110] vdd gnd cell_6t
Xbit_r111_c45 bl[45] br[45] wl[111] vdd gnd cell_6t
Xbit_r112_c45 bl[45] br[45] wl[112] vdd gnd cell_6t
Xbit_r113_c45 bl[45] br[45] wl[113] vdd gnd cell_6t
Xbit_r114_c45 bl[45] br[45] wl[114] vdd gnd cell_6t
Xbit_r115_c45 bl[45] br[45] wl[115] vdd gnd cell_6t
Xbit_r116_c45 bl[45] br[45] wl[116] vdd gnd cell_6t
Xbit_r117_c45 bl[45] br[45] wl[117] vdd gnd cell_6t
Xbit_r118_c45 bl[45] br[45] wl[118] vdd gnd cell_6t
Xbit_r119_c45 bl[45] br[45] wl[119] vdd gnd cell_6t
Xbit_r120_c45 bl[45] br[45] wl[120] vdd gnd cell_6t
Xbit_r121_c45 bl[45] br[45] wl[121] vdd gnd cell_6t
Xbit_r122_c45 bl[45] br[45] wl[122] vdd gnd cell_6t
Xbit_r123_c45 bl[45] br[45] wl[123] vdd gnd cell_6t
Xbit_r124_c45 bl[45] br[45] wl[124] vdd gnd cell_6t
Xbit_r125_c45 bl[45] br[45] wl[125] vdd gnd cell_6t
Xbit_r126_c45 bl[45] br[45] wl[126] vdd gnd cell_6t
Xbit_r127_c45 bl[45] br[45] wl[127] vdd gnd cell_6t
Xbit_r128_c45 bl[45] br[45] wl[128] vdd gnd cell_6t
Xbit_r129_c45 bl[45] br[45] wl[129] vdd gnd cell_6t
Xbit_r130_c45 bl[45] br[45] wl[130] vdd gnd cell_6t
Xbit_r131_c45 bl[45] br[45] wl[131] vdd gnd cell_6t
Xbit_r132_c45 bl[45] br[45] wl[132] vdd gnd cell_6t
Xbit_r133_c45 bl[45] br[45] wl[133] vdd gnd cell_6t
Xbit_r134_c45 bl[45] br[45] wl[134] vdd gnd cell_6t
Xbit_r135_c45 bl[45] br[45] wl[135] vdd gnd cell_6t
Xbit_r136_c45 bl[45] br[45] wl[136] vdd gnd cell_6t
Xbit_r137_c45 bl[45] br[45] wl[137] vdd gnd cell_6t
Xbit_r138_c45 bl[45] br[45] wl[138] vdd gnd cell_6t
Xbit_r139_c45 bl[45] br[45] wl[139] vdd gnd cell_6t
Xbit_r140_c45 bl[45] br[45] wl[140] vdd gnd cell_6t
Xbit_r141_c45 bl[45] br[45] wl[141] vdd gnd cell_6t
Xbit_r142_c45 bl[45] br[45] wl[142] vdd gnd cell_6t
Xbit_r143_c45 bl[45] br[45] wl[143] vdd gnd cell_6t
Xbit_r144_c45 bl[45] br[45] wl[144] vdd gnd cell_6t
Xbit_r145_c45 bl[45] br[45] wl[145] vdd gnd cell_6t
Xbit_r146_c45 bl[45] br[45] wl[146] vdd gnd cell_6t
Xbit_r147_c45 bl[45] br[45] wl[147] vdd gnd cell_6t
Xbit_r148_c45 bl[45] br[45] wl[148] vdd gnd cell_6t
Xbit_r149_c45 bl[45] br[45] wl[149] vdd gnd cell_6t
Xbit_r150_c45 bl[45] br[45] wl[150] vdd gnd cell_6t
Xbit_r151_c45 bl[45] br[45] wl[151] vdd gnd cell_6t
Xbit_r152_c45 bl[45] br[45] wl[152] vdd gnd cell_6t
Xbit_r153_c45 bl[45] br[45] wl[153] vdd gnd cell_6t
Xbit_r154_c45 bl[45] br[45] wl[154] vdd gnd cell_6t
Xbit_r155_c45 bl[45] br[45] wl[155] vdd gnd cell_6t
Xbit_r156_c45 bl[45] br[45] wl[156] vdd gnd cell_6t
Xbit_r157_c45 bl[45] br[45] wl[157] vdd gnd cell_6t
Xbit_r158_c45 bl[45] br[45] wl[158] vdd gnd cell_6t
Xbit_r159_c45 bl[45] br[45] wl[159] vdd gnd cell_6t
Xbit_r160_c45 bl[45] br[45] wl[160] vdd gnd cell_6t
Xbit_r161_c45 bl[45] br[45] wl[161] vdd gnd cell_6t
Xbit_r162_c45 bl[45] br[45] wl[162] vdd gnd cell_6t
Xbit_r163_c45 bl[45] br[45] wl[163] vdd gnd cell_6t
Xbit_r164_c45 bl[45] br[45] wl[164] vdd gnd cell_6t
Xbit_r165_c45 bl[45] br[45] wl[165] vdd gnd cell_6t
Xbit_r166_c45 bl[45] br[45] wl[166] vdd gnd cell_6t
Xbit_r167_c45 bl[45] br[45] wl[167] vdd gnd cell_6t
Xbit_r168_c45 bl[45] br[45] wl[168] vdd gnd cell_6t
Xbit_r169_c45 bl[45] br[45] wl[169] vdd gnd cell_6t
Xbit_r170_c45 bl[45] br[45] wl[170] vdd gnd cell_6t
Xbit_r171_c45 bl[45] br[45] wl[171] vdd gnd cell_6t
Xbit_r172_c45 bl[45] br[45] wl[172] vdd gnd cell_6t
Xbit_r173_c45 bl[45] br[45] wl[173] vdd gnd cell_6t
Xbit_r174_c45 bl[45] br[45] wl[174] vdd gnd cell_6t
Xbit_r175_c45 bl[45] br[45] wl[175] vdd gnd cell_6t
Xbit_r176_c45 bl[45] br[45] wl[176] vdd gnd cell_6t
Xbit_r177_c45 bl[45] br[45] wl[177] vdd gnd cell_6t
Xbit_r178_c45 bl[45] br[45] wl[178] vdd gnd cell_6t
Xbit_r179_c45 bl[45] br[45] wl[179] vdd gnd cell_6t
Xbit_r180_c45 bl[45] br[45] wl[180] vdd gnd cell_6t
Xbit_r181_c45 bl[45] br[45] wl[181] vdd gnd cell_6t
Xbit_r182_c45 bl[45] br[45] wl[182] vdd gnd cell_6t
Xbit_r183_c45 bl[45] br[45] wl[183] vdd gnd cell_6t
Xbit_r184_c45 bl[45] br[45] wl[184] vdd gnd cell_6t
Xbit_r185_c45 bl[45] br[45] wl[185] vdd gnd cell_6t
Xbit_r186_c45 bl[45] br[45] wl[186] vdd gnd cell_6t
Xbit_r187_c45 bl[45] br[45] wl[187] vdd gnd cell_6t
Xbit_r188_c45 bl[45] br[45] wl[188] vdd gnd cell_6t
Xbit_r189_c45 bl[45] br[45] wl[189] vdd gnd cell_6t
Xbit_r190_c45 bl[45] br[45] wl[190] vdd gnd cell_6t
Xbit_r191_c45 bl[45] br[45] wl[191] vdd gnd cell_6t
Xbit_r192_c45 bl[45] br[45] wl[192] vdd gnd cell_6t
Xbit_r193_c45 bl[45] br[45] wl[193] vdd gnd cell_6t
Xbit_r194_c45 bl[45] br[45] wl[194] vdd gnd cell_6t
Xbit_r195_c45 bl[45] br[45] wl[195] vdd gnd cell_6t
Xbit_r196_c45 bl[45] br[45] wl[196] vdd gnd cell_6t
Xbit_r197_c45 bl[45] br[45] wl[197] vdd gnd cell_6t
Xbit_r198_c45 bl[45] br[45] wl[198] vdd gnd cell_6t
Xbit_r199_c45 bl[45] br[45] wl[199] vdd gnd cell_6t
Xbit_r200_c45 bl[45] br[45] wl[200] vdd gnd cell_6t
Xbit_r201_c45 bl[45] br[45] wl[201] vdd gnd cell_6t
Xbit_r202_c45 bl[45] br[45] wl[202] vdd gnd cell_6t
Xbit_r203_c45 bl[45] br[45] wl[203] vdd gnd cell_6t
Xbit_r204_c45 bl[45] br[45] wl[204] vdd gnd cell_6t
Xbit_r205_c45 bl[45] br[45] wl[205] vdd gnd cell_6t
Xbit_r206_c45 bl[45] br[45] wl[206] vdd gnd cell_6t
Xbit_r207_c45 bl[45] br[45] wl[207] vdd gnd cell_6t
Xbit_r208_c45 bl[45] br[45] wl[208] vdd gnd cell_6t
Xbit_r209_c45 bl[45] br[45] wl[209] vdd gnd cell_6t
Xbit_r210_c45 bl[45] br[45] wl[210] vdd gnd cell_6t
Xbit_r211_c45 bl[45] br[45] wl[211] vdd gnd cell_6t
Xbit_r212_c45 bl[45] br[45] wl[212] vdd gnd cell_6t
Xbit_r213_c45 bl[45] br[45] wl[213] vdd gnd cell_6t
Xbit_r214_c45 bl[45] br[45] wl[214] vdd gnd cell_6t
Xbit_r215_c45 bl[45] br[45] wl[215] vdd gnd cell_6t
Xbit_r216_c45 bl[45] br[45] wl[216] vdd gnd cell_6t
Xbit_r217_c45 bl[45] br[45] wl[217] vdd gnd cell_6t
Xbit_r218_c45 bl[45] br[45] wl[218] vdd gnd cell_6t
Xbit_r219_c45 bl[45] br[45] wl[219] vdd gnd cell_6t
Xbit_r220_c45 bl[45] br[45] wl[220] vdd gnd cell_6t
Xbit_r221_c45 bl[45] br[45] wl[221] vdd gnd cell_6t
Xbit_r222_c45 bl[45] br[45] wl[222] vdd gnd cell_6t
Xbit_r223_c45 bl[45] br[45] wl[223] vdd gnd cell_6t
Xbit_r224_c45 bl[45] br[45] wl[224] vdd gnd cell_6t
Xbit_r225_c45 bl[45] br[45] wl[225] vdd gnd cell_6t
Xbit_r226_c45 bl[45] br[45] wl[226] vdd gnd cell_6t
Xbit_r227_c45 bl[45] br[45] wl[227] vdd gnd cell_6t
Xbit_r228_c45 bl[45] br[45] wl[228] vdd gnd cell_6t
Xbit_r229_c45 bl[45] br[45] wl[229] vdd gnd cell_6t
Xbit_r230_c45 bl[45] br[45] wl[230] vdd gnd cell_6t
Xbit_r231_c45 bl[45] br[45] wl[231] vdd gnd cell_6t
Xbit_r232_c45 bl[45] br[45] wl[232] vdd gnd cell_6t
Xbit_r233_c45 bl[45] br[45] wl[233] vdd gnd cell_6t
Xbit_r234_c45 bl[45] br[45] wl[234] vdd gnd cell_6t
Xbit_r235_c45 bl[45] br[45] wl[235] vdd gnd cell_6t
Xbit_r236_c45 bl[45] br[45] wl[236] vdd gnd cell_6t
Xbit_r237_c45 bl[45] br[45] wl[237] vdd gnd cell_6t
Xbit_r238_c45 bl[45] br[45] wl[238] vdd gnd cell_6t
Xbit_r239_c45 bl[45] br[45] wl[239] vdd gnd cell_6t
Xbit_r240_c45 bl[45] br[45] wl[240] vdd gnd cell_6t
Xbit_r241_c45 bl[45] br[45] wl[241] vdd gnd cell_6t
Xbit_r242_c45 bl[45] br[45] wl[242] vdd gnd cell_6t
Xbit_r243_c45 bl[45] br[45] wl[243] vdd gnd cell_6t
Xbit_r244_c45 bl[45] br[45] wl[244] vdd gnd cell_6t
Xbit_r245_c45 bl[45] br[45] wl[245] vdd gnd cell_6t
Xbit_r246_c45 bl[45] br[45] wl[246] vdd gnd cell_6t
Xbit_r247_c45 bl[45] br[45] wl[247] vdd gnd cell_6t
Xbit_r248_c45 bl[45] br[45] wl[248] vdd gnd cell_6t
Xbit_r249_c45 bl[45] br[45] wl[249] vdd gnd cell_6t
Xbit_r250_c45 bl[45] br[45] wl[250] vdd gnd cell_6t
Xbit_r251_c45 bl[45] br[45] wl[251] vdd gnd cell_6t
Xbit_r252_c45 bl[45] br[45] wl[252] vdd gnd cell_6t
Xbit_r253_c45 bl[45] br[45] wl[253] vdd gnd cell_6t
Xbit_r254_c45 bl[45] br[45] wl[254] vdd gnd cell_6t
Xbit_r255_c45 bl[45] br[45] wl[255] vdd gnd cell_6t
Xbit_r0_c46 bl[46] br[46] wl[0] vdd gnd cell_6t
Xbit_r1_c46 bl[46] br[46] wl[1] vdd gnd cell_6t
Xbit_r2_c46 bl[46] br[46] wl[2] vdd gnd cell_6t
Xbit_r3_c46 bl[46] br[46] wl[3] vdd gnd cell_6t
Xbit_r4_c46 bl[46] br[46] wl[4] vdd gnd cell_6t
Xbit_r5_c46 bl[46] br[46] wl[5] vdd gnd cell_6t
Xbit_r6_c46 bl[46] br[46] wl[6] vdd gnd cell_6t
Xbit_r7_c46 bl[46] br[46] wl[7] vdd gnd cell_6t
Xbit_r8_c46 bl[46] br[46] wl[8] vdd gnd cell_6t
Xbit_r9_c46 bl[46] br[46] wl[9] vdd gnd cell_6t
Xbit_r10_c46 bl[46] br[46] wl[10] vdd gnd cell_6t
Xbit_r11_c46 bl[46] br[46] wl[11] vdd gnd cell_6t
Xbit_r12_c46 bl[46] br[46] wl[12] vdd gnd cell_6t
Xbit_r13_c46 bl[46] br[46] wl[13] vdd gnd cell_6t
Xbit_r14_c46 bl[46] br[46] wl[14] vdd gnd cell_6t
Xbit_r15_c46 bl[46] br[46] wl[15] vdd gnd cell_6t
Xbit_r16_c46 bl[46] br[46] wl[16] vdd gnd cell_6t
Xbit_r17_c46 bl[46] br[46] wl[17] vdd gnd cell_6t
Xbit_r18_c46 bl[46] br[46] wl[18] vdd gnd cell_6t
Xbit_r19_c46 bl[46] br[46] wl[19] vdd gnd cell_6t
Xbit_r20_c46 bl[46] br[46] wl[20] vdd gnd cell_6t
Xbit_r21_c46 bl[46] br[46] wl[21] vdd gnd cell_6t
Xbit_r22_c46 bl[46] br[46] wl[22] vdd gnd cell_6t
Xbit_r23_c46 bl[46] br[46] wl[23] vdd gnd cell_6t
Xbit_r24_c46 bl[46] br[46] wl[24] vdd gnd cell_6t
Xbit_r25_c46 bl[46] br[46] wl[25] vdd gnd cell_6t
Xbit_r26_c46 bl[46] br[46] wl[26] vdd gnd cell_6t
Xbit_r27_c46 bl[46] br[46] wl[27] vdd gnd cell_6t
Xbit_r28_c46 bl[46] br[46] wl[28] vdd gnd cell_6t
Xbit_r29_c46 bl[46] br[46] wl[29] vdd gnd cell_6t
Xbit_r30_c46 bl[46] br[46] wl[30] vdd gnd cell_6t
Xbit_r31_c46 bl[46] br[46] wl[31] vdd gnd cell_6t
Xbit_r32_c46 bl[46] br[46] wl[32] vdd gnd cell_6t
Xbit_r33_c46 bl[46] br[46] wl[33] vdd gnd cell_6t
Xbit_r34_c46 bl[46] br[46] wl[34] vdd gnd cell_6t
Xbit_r35_c46 bl[46] br[46] wl[35] vdd gnd cell_6t
Xbit_r36_c46 bl[46] br[46] wl[36] vdd gnd cell_6t
Xbit_r37_c46 bl[46] br[46] wl[37] vdd gnd cell_6t
Xbit_r38_c46 bl[46] br[46] wl[38] vdd gnd cell_6t
Xbit_r39_c46 bl[46] br[46] wl[39] vdd gnd cell_6t
Xbit_r40_c46 bl[46] br[46] wl[40] vdd gnd cell_6t
Xbit_r41_c46 bl[46] br[46] wl[41] vdd gnd cell_6t
Xbit_r42_c46 bl[46] br[46] wl[42] vdd gnd cell_6t
Xbit_r43_c46 bl[46] br[46] wl[43] vdd gnd cell_6t
Xbit_r44_c46 bl[46] br[46] wl[44] vdd gnd cell_6t
Xbit_r45_c46 bl[46] br[46] wl[45] vdd gnd cell_6t
Xbit_r46_c46 bl[46] br[46] wl[46] vdd gnd cell_6t
Xbit_r47_c46 bl[46] br[46] wl[47] vdd gnd cell_6t
Xbit_r48_c46 bl[46] br[46] wl[48] vdd gnd cell_6t
Xbit_r49_c46 bl[46] br[46] wl[49] vdd gnd cell_6t
Xbit_r50_c46 bl[46] br[46] wl[50] vdd gnd cell_6t
Xbit_r51_c46 bl[46] br[46] wl[51] vdd gnd cell_6t
Xbit_r52_c46 bl[46] br[46] wl[52] vdd gnd cell_6t
Xbit_r53_c46 bl[46] br[46] wl[53] vdd gnd cell_6t
Xbit_r54_c46 bl[46] br[46] wl[54] vdd gnd cell_6t
Xbit_r55_c46 bl[46] br[46] wl[55] vdd gnd cell_6t
Xbit_r56_c46 bl[46] br[46] wl[56] vdd gnd cell_6t
Xbit_r57_c46 bl[46] br[46] wl[57] vdd gnd cell_6t
Xbit_r58_c46 bl[46] br[46] wl[58] vdd gnd cell_6t
Xbit_r59_c46 bl[46] br[46] wl[59] vdd gnd cell_6t
Xbit_r60_c46 bl[46] br[46] wl[60] vdd gnd cell_6t
Xbit_r61_c46 bl[46] br[46] wl[61] vdd gnd cell_6t
Xbit_r62_c46 bl[46] br[46] wl[62] vdd gnd cell_6t
Xbit_r63_c46 bl[46] br[46] wl[63] vdd gnd cell_6t
Xbit_r64_c46 bl[46] br[46] wl[64] vdd gnd cell_6t
Xbit_r65_c46 bl[46] br[46] wl[65] vdd gnd cell_6t
Xbit_r66_c46 bl[46] br[46] wl[66] vdd gnd cell_6t
Xbit_r67_c46 bl[46] br[46] wl[67] vdd gnd cell_6t
Xbit_r68_c46 bl[46] br[46] wl[68] vdd gnd cell_6t
Xbit_r69_c46 bl[46] br[46] wl[69] vdd gnd cell_6t
Xbit_r70_c46 bl[46] br[46] wl[70] vdd gnd cell_6t
Xbit_r71_c46 bl[46] br[46] wl[71] vdd gnd cell_6t
Xbit_r72_c46 bl[46] br[46] wl[72] vdd gnd cell_6t
Xbit_r73_c46 bl[46] br[46] wl[73] vdd gnd cell_6t
Xbit_r74_c46 bl[46] br[46] wl[74] vdd gnd cell_6t
Xbit_r75_c46 bl[46] br[46] wl[75] vdd gnd cell_6t
Xbit_r76_c46 bl[46] br[46] wl[76] vdd gnd cell_6t
Xbit_r77_c46 bl[46] br[46] wl[77] vdd gnd cell_6t
Xbit_r78_c46 bl[46] br[46] wl[78] vdd gnd cell_6t
Xbit_r79_c46 bl[46] br[46] wl[79] vdd gnd cell_6t
Xbit_r80_c46 bl[46] br[46] wl[80] vdd gnd cell_6t
Xbit_r81_c46 bl[46] br[46] wl[81] vdd gnd cell_6t
Xbit_r82_c46 bl[46] br[46] wl[82] vdd gnd cell_6t
Xbit_r83_c46 bl[46] br[46] wl[83] vdd gnd cell_6t
Xbit_r84_c46 bl[46] br[46] wl[84] vdd gnd cell_6t
Xbit_r85_c46 bl[46] br[46] wl[85] vdd gnd cell_6t
Xbit_r86_c46 bl[46] br[46] wl[86] vdd gnd cell_6t
Xbit_r87_c46 bl[46] br[46] wl[87] vdd gnd cell_6t
Xbit_r88_c46 bl[46] br[46] wl[88] vdd gnd cell_6t
Xbit_r89_c46 bl[46] br[46] wl[89] vdd gnd cell_6t
Xbit_r90_c46 bl[46] br[46] wl[90] vdd gnd cell_6t
Xbit_r91_c46 bl[46] br[46] wl[91] vdd gnd cell_6t
Xbit_r92_c46 bl[46] br[46] wl[92] vdd gnd cell_6t
Xbit_r93_c46 bl[46] br[46] wl[93] vdd gnd cell_6t
Xbit_r94_c46 bl[46] br[46] wl[94] vdd gnd cell_6t
Xbit_r95_c46 bl[46] br[46] wl[95] vdd gnd cell_6t
Xbit_r96_c46 bl[46] br[46] wl[96] vdd gnd cell_6t
Xbit_r97_c46 bl[46] br[46] wl[97] vdd gnd cell_6t
Xbit_r98_c46 bl[46] br[46] wl[98] vdd gnd cell_6t
Xbit_r99_c46 bl[46] br[46] wl[99] vdd gnd cell_6t
Xbit_r100_c46 bl[46] br[46] wl[100] vdd gnd cell_6t
Xbit_r101_c46 bl[46] br[46] wl[101] vdd gnd cell_6t
Xbit_r102_c46 bl[46] br[46] wl[102] vdd gnd cell_6t
Xbit_r103_c46 bl[46] br[46] wl[103] vdd gnd cell_6t
Xbit_r104_c46 bl[46] br[46] wl[104] vdd gnd cell_6t
Xbit_r105_c46 bl[46] br[46] wl[105] vdd gnd cell_6t
Xbit_r106_c46 bl[46] br[46] wl[106] vdd gnd cell_6t
Xbit_r107_c46 bl[46] br[46] wl[107] vdd gnd cell_6t
Xbit_r108_c46 bl[46] br[46] wl[108] vdd gnd cell_6t
Xbit_r109_c46 bl[46] br[46] wl[109] vdd gnd cell_6t
Xbit_r110_c46 bl[46] br[46] wl[110] vdd gnd cell_6t
Xbit_r111_c46 bl[46] br[46] wl[111] vdd gnd cell_6t
Xbit_r112_c46 bl[46] br[46] wl[112] vdd gnd cell_6t
Xbit_r113_c46 bl[46] br[46] wl[113] vdd gnd cell_6t
Xbit_r114_c46 bl[46] br[46] wl[114] vdd gnd cell_6t
Xbit_r115_c46 bl[46] br[46] wl[115] vdd gnd cell_6t
Xbit_r116_c46 bl[46] br[46] wl[116] vdd gnd cell_6t
Xbit_r117_c46 bl[46] br[46] wl[117] vdd gnd cell_6t
Xbit_r118_c46 bl[46] br[46] wl[118] vdd gnd cell_6t
Xbit_r119_c46 bl[46] br[46] wl[119] vdd gnd cell_6t
Xbit_r120_c46 bl[46] br[46] wl[120] vdd gnd cell_6t
Xbit_r121_c46 bl[46] br[46] wl[121] vdd gnd cell_6t
Xbit_r122_c46 bl[46] br[46] wl[122] vdd gnd cell_6t
Xbit_r123_c46 bl[46] br[46] wl[123] vdd gnd cell_6t
Xbit_r124_c46 bl[46] br[46] wl[124] vdd gnd cell_6t
Xbit_r125_c46 bl[46] br[46] wl[125] vdd gnd cell_6t
Xbit_r126_c46 bl[46] br[46] wl[126] vdd gnd cell_6t
Xbit_r127_c46 bl[46] br[46] wl[127] vdd gnd cell_6t
Xbit_r128_c46 bl[46] br[46] wl[128] vdd gnd cell_6t
Xbit_r129_c46 bl[46] br[46] wl[129] vdd gnd cell_6t
Xbit_r130_c46 bl[46] br[46] wl[130] vdd gnd cell_6t
Xbit_r131_c46 bl[46] br[46] wl[131] vdd gnd cell_6t
Xbit_r132_c46 bl[46] br[46] wl[132] vdd gnd cell_6t
Xbit_r133_c46 bl[46] br[46] wl[133] vdd gnd cell_6t
Xbit_r134_c46 bl[46] br[46] wl[134] vdd gnd cell_6t
Xbit_r135_c46 bl[46] br[46] wl[135] vdd gnd cell_6t
Xbit_r136_c46 bl[46] br[46] wl[136] vdd gnd cell_6t
Xbit_r137_c46 bl[46] br[46] wl[137] vdd gnd cell_6t
Xbit_r138_c46 bl[46] br[46] wl[138] vdd gnd cell_6t
Xbit_r139_c46 bl[46] br[46] wl[139] vdd gnd cell_6t
Xbit_r140_c46 bl[46] br[46] wl[140] vdd gnd cell_6t
Xbit_r141_c46 bl[46] br[46] wl[141] vdd gnd cell_6t
Xbit_r142_c46 bl[46] br[46] wl[142] vdd gnd cell_6t
Xbit_r143_c46 bl[46] br[46] wl[143] vdd gnd cell_6t
Xbit_r144_c46 bl[46] br[46] wl[144] vdd gnd cell_6t
Xbit_r145_c46 bl[46] br[46] wl[145] vdd gnd cell_6t
Xbit_r146_c46 bl[46] br[46] wl[146] vdd gnd cell_6t
Xbit_r147_c46 bl[46] br[46] wl[147] vdd gnd cell_6t
Xbit_r148_c46 bl[46] br[46] wl[148] vdd gnd cell_6t
Xbit_r149_c46 bl[46] br[46] wl[149] vdd gnd cell_6t
Xbit_r150_c46 bl[46] br[46] wl[150] vdd gnd cell_6t
Xbit_r151_c46 bl[46] br[46] wl[151] vdd gnd cell_6t
Xbit_r152_c46 bl[46] br[46] wl[152] vdd gnd cell_6t
Xbit_r153_c46 bl[46] br[46] wl[153] vdd gnd cell_6t
Xbit_r154_c46 bl[46] br[46] wl[154] vdd gnd cell_6t
Xbit_r155_c46 bl[46] br[46] wl[155] vdd gnd cell_6t
Xbit_r156_c46 bl[46] br[46] wl[156] vdd gnd cell_6t
Xbit_r157_c46 bl[46] br[46] wl[157] vdd gnd cell_6t
Xbit_r158_c46 bl[46] br[46] wl[158] vdd gnd cell_6t
Xbit_r159_c46 bl[46] br[46] wl[159] vdd gnd cell_6t
Xbit_r160_c46 bl[46] br[46] wl[160] vdd gnd cell_6t
Xbit_r161_c46 bl[46] br[46] wl[161] vdd gnd cell_6t
Xbit_r162_c46 bl[46] br[46] wl[162] vdd gnd cell_6t
Xbit_r163_c46 bl[46] br[46] wl[163] vdd gnd cell_6t
Xbit_r164_c46 bl[46] br[46] wl[164] vdd gnd cell_6t
Xbit_r165_c46 bl[46] br[46] wl[165] vdd gnd cell_6t
Xbit_r166_c46 bl[46] br[46] wl[166] vdd gnd cell_6t
Xbit_r167_c46 bl[46] br[46] wl[167] vdd gnd cell_6t
Xbit_r168_c46 bl[46] br[46] wl[168] vdd gnd cell_6t
Xbit_r169_c46 bl[46] br[46] wl[169] vdd gnd cell_6t
Xbit_r170_c46 bl[46] br[46] wl[170] vdd gnd cell_6t
Xbit_r171_c46 bl[46] br[46] wl[171] vdd gnd cell_6t
Xbit_r172_c46 bl[46] br[46] wl[172] vdd gnd cell_6t
Xbit_r173_c46 bl[46] br[46] wl[173] vdd gnd cell_6t
Xbit_r174_c46 bl[46] br[46] wl[174] vdd gnd cell_6t
Xbit_r175_c46 bl[46] br[46] wl[175] vdd gnd cell_6t
Xbit_r176_c46 bl[46] br[46] wl[176] vdd gnd cell_6t
Xbit_r177_c46 bl[46] br[46] wl[177] vdd gnd cell_6t
Xbit_r178_c46 bl[46] br[46] wl[178] vdd gnd cell_6t
Xbit_r179_c46 bl[46] br[46] wl[179] vdd gnd cell_6t
Xbit_r180_c46 bl[46] br[46] wl[180] vdd gnd cell_6t
Xbit_r181_c46 bl[46] br[46] wl[181] vdd gnd cell_6t
Xbit_r182_c46 bl[46] br[46] wl[182] vdd gnd cell_6t
Xbit_r183_c46 bl[46] br[46] wl[183] vdd gnd cell_6t
Xbit_r184_c46 bl[46] br[46] wl[184] vdd gnd cell_6t
Xbit_r185_c46 bl[46] br[46] wl[185] vdd gnd cell_6t
Xbit_r186_c46 bl[46] br[46] wl[186] vdd gnd cell_6t
Xbit_r187_c46 bl[46] br[46] wl[187] vdd gnd cell_6t
Xbit_r188_c46 bl[46] br[46] wl[188] vdd gnd cell_6t
Xbit_r189_c46 bl[46] br[46] wl[189] vdd gnd cell_6t
Xbit_r190_c46 bl[46] br[46] wl[190] vdd gnd cell_6t
Xbit_r191_c46 bl[46] br[46] wl[191] vdd gnd cell_6t
Xbit_r192_c46 bl[46] br[46] wl[192] vdd gnd cell_6t
Xbit_r193_c46 bl[46] br[46] wl[193] vdd gnd cell_6t
Xbit_r194_c46 bl[46] br[46] wl[194] vdd gnd cell_6t
Xbit_r195_c46 bl[46] br[46] wl[195] vdd gnd cell_6t
Xbit_r196_c46 bl[46] br[46] wl[196] vdd gnd cell_6t
Xbit_r197_c46 bl[46] br[46] wl[197] vdd gnd cell_6t
Xbit_r198_c46 bl[46] br[46] wl[198] vdd gnd cell_6t
Xbit_r199_c46 bl[46] br[46] wl[199] vdd gnd cell_6t
Xbit_r200_c46 bl[46] br[46] wl[200] vdd gnd cell_6t
Xbit_r201_c46 bl[46] br[46] wl[201] vdd gnd cell_6t
Xbit_r202_c46 bl[46] br[46] wl[202] vdd gnd cell_6t
Xbit_r203_c46 bl[46] br[46] wl[203] vdd gnd cell_6t
Xbit_r204_c46 bl[46] br[46] wl[204] vdd gnd cell_6t
Xbit_r205_c46 bl[46] br[46] wl[205] vdd gnd cell_6t
Xbit_r206_c46 bl[46] br[46] wl[206] vdd gnd cell_6t
Xbit_r207_c46 bl[46] br[46] wl[207] vdd gnd cell_6t
Xbit_r208_c46 bl[46] br[46] wl[208] vdd gnd cell_6t
Xbit_r209_c46 bl[46] br[46] wl[209] vdd gnd cell_6t
Xbit_r210_c46 bl[46] br[46] wl[210] vdd gnd cell_6t
Xbit_r211_c46 bl[46] br[46] wl[211] vdd gnd cell_6t
Xbit_r212_c46 bl[46] br[46] wl[212] vdd gnd cell_6t
Xbit_r213_c46 bl[46] br[46] wl[213] vdd gnd cell_6t
Xbit_r214_c46 bl[46] br[46] wl[214] vdd gnd cell_6t
Xbit_r215_c46 bl[46] br[46] wl[215] vdd gnd cell_6t
Xbit_r216_c46 bl[46] br[46] wl[216] vdd gnd cell_6t
Xbit_r217_c46 bl[46] br[46] wl[217] vdd gnd cell_6t
Xbit_r218_c46 bl[46] br[46] wl[218] vdd gnd cell_6t
Xbit_r219_c46 bl[46] br[46] wl[219] vdd gnd cell_6t
Xbit_r220_c46 bl[46] br[46] wl[220] vdd gnd cell_6t
Xbit_r221_c46 bl[46] br[46] wl[221] vdd gnd cell_6t
Xbit_r222_c46 bl[46] br[46] wl[222] vdd gnd cell_6t
Xbit_r223_c46 bl[46] br[46] wl[223] vdd gnd cell_6t
Xbit_r224_c46 bl[46] br[46] wl[224] vdd gnd cell_6t
Xbit_r225_c46 bl[46] br[46] wl[225] vdd gnd cell_6t
Xbit_r226_c46 bl[46] br[46] wl[226] vdd gnd cell_6t
Xbit_r227_c46 bl[46] br[46] wl[227] vdd gnd cell_6t
Xbit_r228_c46 bl[46] br[46] wl[228] vdd gnd cell_6t
Xbit_r229_c46 bl[46] br[46] wl[229] vdd gnd cell_6t
Xbit_r230_c46 bl[46] br[46] wl[230] vdd gnd cell_6t
Xbit_r231_c46 bl[46] br[46] wl[231] vdd gnd cell_6t
Xbit_r232_c46 bl[46] br[46] wl[232] vdd gnd cell_6t
Xbit_r233_c46 bl[46] br[46] wl[233] vdd gnd cell_6t
Xbit_r234_c46 bl[46] br[46] wl[234] vdd gnd cell_6t
Xbit_r235_c46 bl[46] br[46] wl[235] vdd gnd cell_6t
Xbit_r236_c46 bl[46] br[46] wl[236] vdd gnd cell_6t
Xbit_r237_c46 bl[46] br[46] wl[237] vdd gnd cell_6t
Xbit_r238_c46 bl[46] br[46] wl[238] vdd gnd cell_6t
Xbit_r239_c46 bl[46] br[46] wl[239] vdd gnd cell_6t
Xbit_r240_c46 bl[46] br[46] wl[240] vdd gnd cell_6t
Xbit_r241_c46 bl[46] br[46] wl[241] vdd gnd cell_6t
Xbit_r242_c46 bl[46] br[46] wl[242] vdd gnd cell_6t
Xbit_r243_c46 bl[46] br[46] wl[243] vdd gnd cell_6t
Xbit_r244_c46 bl[46] br[46] wl[244] vdd gnd cell_6t
Xbit_r245_c46 bl[46] br[46] wl[245] vdd gnd cell_6t
Xbit_r246_c46 bl[46] br[46] wl[246] vdd gnd cell_6t
Xbit_r247_c46 bl[46] br[46] wl[247] vdd gnd cell_6t
Xbit_r248_c46 bl[46] br[46] wl[248] vdd gnd cell_6t
Xbit_r249_c46 bl[46] br[46] wl[249] vdd gnd cell_6t
Xbit_r250_c46 bl[46] br[46] wl[250] vdd gnd cell_6t
Xbit_r251_c46 bl[46] br[46] wl[251] vdd gnd cell_6t
Xbit_r252_c46 bl[46] br[46] wl[252] vdd gnd cell_6t
Xbit_r253_c46 bl[46] br[46] wl[253] vdd gnd cell_6t
Xbit_r254_c46 bl[46] br[46] wl[254] vdd gnd cell_6t
Xbit_r255_c46 bl[46] br[46] wl[255] vdd gnd cell_6t
Xbit_r0_c47 bl[47] br[47] wl[0] vdd gnd cell_6t
Xbit_r1_c47 bl[47] br[47] wl[1] vdd gnd cell_6t
Xbit_r2_c47 bl[47] br[47] wl[2] vdd gnd cell_6t
Xbit_r3_c47 bl[47] br[47] wl[3] vdd gnd cell_6t
Xbit_r4_c47 bl[47] br[47] wl[4] vdd gnd cell_6t
Xbit_r5_c47 bl[47] br[47] wl[5] vdd gnd cell_6t
Xbit_r6_c47 bl[47] br[47] wl[6] vdd gnd cell_6t
Xbit_r7_c47 bl[47] br[47] wl[7] vdd gnd cell_6t
Xbit_r8_c47 bl[47] br[47] wl[8] vdd gnd cell_6t
Xbit_r9_c47 bl[47] br[47] wl[9] vdd gnd cell_6t
Xbit_r10_c47 bl[47] br[47] wl[10] vdd gnd cell_6t
Xbit_r11_c47 bl[47] br[47] wl[11] vdd gnd cell_6t
Xbit_r12_c47 bl[47] br[47] wl[12] vdd gnd cell_6t
Xbit_r13_c47 bl[47] br[47] wl[13] vdd gnd cell_6t
Xbit_r14_c47 bl[47] br[47] wl[14] vdd gnd cell_6t
Xbit_r15_c47 bl[47] br[47] wl[15] vdd gnd cell_6t
Xbit_r16_c47 bl[47] br[47] wl[16] vdd gnd cell_6t
Xbit_r17_c47 bl[47] br[47] wl[17] vdd gnd cell_6t
Xbit_r18_c47 bl[47] br[47] wl[18] vdd gnd cell_6t
Xbit_r19_c47 bl[47] br[47] wl[19] vdd gnd cell_6t
Xbit_r20_c47 bl[47] br[47] wl[20] vdd gnd cell_6t
Xbit_r21_c47 bl[47] br[47] wl[21] vdd gnd cell_6t
Xbit_r22_c47 bl[47] br[47] wl[22] vdd gnd cell_6t
Xbit_r23_c47 bl[47] br[47] wl[23] vdd gnd cell_6t
Xbit_r24_c47 bl[47] br[47] wl[24] vdd gnd cell_6t
Xbit_r25_c47 bl[47] br[47] wl[25] vdd gnd cell_6t
Xbit_r26_c47 bl[47] br[47] wl[26] vdd gnd cell_6t
Xbit_r27_c47 bl[47] br[47] wl[27] vdd gnd cell_6t
Xbit_r28_c47 bl[47] br[47] wl[28] vdd gnd cell_6t
Xbit_r29_c47 bl[47] br[47] wl[29] vdd gnd cell_6t
Xbit_r30_c47 bl[47] br[47] wl[30] vdd gnd cell_6t
Xbit_r31_c47 bl[47] br[47] wl[31] vdd gnd cell_6t
Xbit_r32_c47 bl[47] br[47] wl[32] vdd gnd cell_6t
Xbit_r33_c47 bl[47] br[47] wl[33] vdd gnd cell_6t
Xbit_r34_c47 bl[47] br[47] wl[34] vdd gnd cell_6t
Xbit_r35_c47 bl[47] br[47] wl[35] vdd gnd cell_6t
Xbit_r36_c47 bl[47] br[47] wl[36] vdd gnd cell_6t
Xbit_r37_c47 bl[47] br[47] wl[37] vdd gnd cell_6t
Xbit_r38_c47 bl[47] br[47] wl[38] vdd gnd cell_6t
Xbit_r39_c47 bl[47] br[47] wl[39] vdd gnd cell_6t
Xbit_r40_c47 bl[47] br[47] wl[40] vdd gnd cell_6t
Xbit_r41_c47 bl[47] br[47] wl[41] vdd gnd cell_6t
Xbit_r42_c47 bl[47] br[47] wl[42] vdd gnd cell_6t
Xbit_r43_c47 bl[47] br[47] wl[43] vdd gnd cell_6t
Xbit_r44_c47 bl[47] br[47] wl[44] vdd gnd cell_6t
Xbit_r45_c47 bl[47] br[47] wl[45] vdd gnd cell_6t
Xbit_r46_c47 bl[47] br[47] wl[46] vdd gnd cell_6t
Xbit_r47_c47 bl[47] br[47] wl[47] vdd gnd cell_6t
Xbit_r48_c47 bl[47] br[47] wl[48] vdd gnd cell_6t
Xbit_r49_c47 bl[47] br[47] wl[49] vdd gnd cell_6t
Xbit_r50_c47 bl[47] br[47] wl[50] vdd gnd cell_6t
Xbit_r51_c47 bl[47] br[47] wl[51] vdd gnd cell_6t
Xbit_r52_c47 bl[47] br[47] wl[52] vdd gnd cell_6t
Xbit_r53_c47 bl[47] br[47] wl[53] vdd gnd cell_6t
Xbit_r54_c47 bl[47] br[47] wl[54] vdd gnd cell_6t
Xbit_r55_c47 bl[47] br[47] wl[55] vdd gnd cell_6t
Xbit_r56_c47 bl[47] br[47] wl[56] vdd gnd cell_6t
Xbit_r57_c47 bl[47] br[47] wl[57] vdd gnd cell_6t
Xbit_r58_c47 bl[47] br[47] wl[58] vdd gnd cell_6t
Xbit_r59_c47 bl[47] br[47] wl[59] vdd gnd cell_6t
Xbit_r60_c47 bl[47] br[47] wl[60] vdd gnd cell_6t
Xbit_r61_c47 bl[47] br[47] wl[61] vdd gnd cell_6t
Xbit_r62_c47 bl[47] br[47] wl[62] vdd gnd cell_6t
Xbit_r63_c47 bl[47] br[47] wl[63] vdd gnd cell_6t
Xbit_r64_c47 bl[47] br[47] wl[64] vdd gnd cell_6t
Xbit_r65_c47 bl[47] br[47] wl[65] vdd gnd cell_6t
Xbit_r66_c47 bl[47] br[47] wl[66] vdd gnd cell_6t
Xbit_r67_c47 bl[47] br[47] wl[67] vdd gnd cell_6t
Xbit_r68_c47 bl[47] br[47] wl[68] vdd gnd cell_6t
Xbit_r69_c47 bl[47] br[47] wl[69] vdd gnd cell_6t
Xbit_r70_c47 bl[47] br[47] wl[70] vdd gnd cell_6t
Xbit_r71_c47 bl[47] br[47] wl[71] vdd gnd cell_6t
Xbit_r72_c47 bl[47] br[47] wl[72] vdd gnd cell_6t
Xbit_r73_c47 bl[47] br[47] wl[73] vdd gnd cell_6t
Xbit_r74_c47 bl[47] br[47] wl[74] vdd gnd cell_6t
Xbit_r75_c47 bl[47] br[47] wl[75] vdd gnd cell_6t
Xbit_r76_c47 bl[47] br[47] wl[76] vdd gnd cell_6t
Xbit_r77_c47 bl[47] br[47] wl[77] vdd gnd cell_6t
Xbit_r78_c47 bl[47] br[47] wl[78] vdd gnd cell_6t
Xbit_r79_c47 bl[47] br[47] wl[79] vdd gnd cell_6t
Xbit_r80_c47 bl[47] br[47] wl[80] vdd gnd cell_6t
Xbit_r81_c47 bl[47] br[47] wl[81] vdd gnd cell_6t
Xbit_r82_c47 bl[47] br[47] wl[82] vdd gnd cell_6t
Xbit_r83_c47 bl[47] br[47] wl[83] vdd gnd cell_6t
Xbit_r84_c47 bl[47] br[47] wl[84] vdd gnd cell_6t
Xbit_r85_c47 bl[47] br[47] wl[85] vdd gnd cell_6t
Xbit_r86_c47 bl[47] br[47] wl[86] vdd gnd cell_6t
Xbit_r87_c47 bl[47] br[47] wl[87] vdd gnd cell_6t
Xbit_r88_c47 bl[47] br[47] wl[88] vdd gnd cell_6t
Xbit_r89_c47 bl[47] br[47] wl[89] vdd gnd cell_6t
Xbit_r90_c47 bl[47] br[47] wl[90] vdd gnd cell_6t
Xbit_r91_c47 bl[47] br[47] wl[91] vdd gnd cell_6t
Xbit_r92_c47 bl[47] br[47] wl[92] vdd gnd cell_6t
Xbit_r93_c47 bl[47] br[47] wl[93] vdd gnd cell_6t
Xbit_r94_c47 bl[47] br[47] wl[94] vdd gnd cell_6t
Xbit_r95_c47 bl[47] br[47] wl[95] vdd gnd cell_6t
Xbit_r96_c47 bl[47] br[47] wl[96] vdd gnd cell_6t
Xbit_r97_c47 bl[47] br[47] wl[97] vdd gnd cell_6t
Xbit_r98_c47 bl[47] br[47] wl[98] vdd gnd cell_6t
Xbit_r99_c47 bl[47] br[47] wl[99] vdd gnd cell_6t
Xbit_r100_c47 bl[47] br[47] wl[100] vdd gnd cell_6t
Xbit_r101_c47 bl[47] br[47] wl[101] vdd gnd cell_6t
Xbit_r102_c47 bl[47] br[47] wl[102] vdd gnd cell_6t
Xbit_r103_c47 bl[47] br[47] wl[103] vdd gnd cell_6t
Xbit_r104_c47 bl[47] br[47] wl[104] vdd gnd cell_6t
Xbit_r105_c47 bl[47] br[47] wl[105] vdd gnd cell_6t
Xbit_r106_c47 bl[47] br[47] wl[106] vdd gnd cell_6t
Xbit_r107_c47 bl[47] br[47] wl[107] vdd gnd cell_6t
Xbit_r108_c47 bl[47] br[47] wl[108] vdd gnd cell_6t
Xbit_r109_c47 bl[47] br[47] wl[109] vdd gnd cell_6t
Xbit_r110_c47 bl[47] br[47] wl[110] vdd gnd cell_6t
Xbit_r111_c47 bl[47] br[47] wl[111] vdd gnd cell_6t
Xbit_r112_c47 bl[47] br[47] wl[112] vdd gnd cell_6t
Xbit_r113_c47 bl[47] br[47] wl[113] vdd gnd cell_6t
Xbit_r114_c47 bl[47] br[47] wl[114] vdd gnd cell_6t
Xbit_r115_c47 bl[47] br[47] wl[115] vdd gnd cell_6t
Xbit_r116_c47 bl[47] br[47] wl[116] vdd gnd cell_6t
Xbit_r117_c47 bl[47] br[47] wl[117] vdd gnd cell_6t
Xbit_r118_c47 bl[47] br[47] wl[118] vdd gnd cell_6t
Xbit_r119_c47 bl[47] br[47] wl[119] vdd gnd cell_6t
Xbit_r120_c47 bl[47] br[47] wl[120] vdd gnd cell_6t
Xbit_r121_c47 bl[47] br[47] wl[121] vdd gnd cell_6t
Xbit_r122_c47 bl[47] br[47] wl[122] vdd gnd cell_6t
Xbit_r123_c47 bl[47] br[47] wl[123] vdd gnd cell_6t
Xbit_r124_c47 bl[47] br[47] wl[124] vdd gnd cell_6t
Xbit_r125_c47 bl[47] br[47] wl[125] vdd gnd cell_6t
Xbit_r126_c47 bl[47] br[47] wl[126] vdd gnd cell_6t
Xbit_r127_c47 bl[47] br[47] wl[127] vdd gnd cell_6t
Xbit_r128_c47 bl[47] br[47] wl[128] vdd gnd cell_6t
Xbit_r129_c47 bl[47] br[47] wl[129] vdd gnd cell_6t
Xbit_r130_c47 bl[47] br[47] wl[130] vdd gnd cell_6t
Xbit_r131_c47 bl[47] br[47] wl[131] vdd gnd cell_6t
Xbit_r132_c47 bl[47] br[47] wl[132] vdd gnd cell_6t
Xbit_r133_c47 bl[47] br[47] wl[133] vdd gnd cell_6t
Xbit_r134_c47 bl[47] br[47] wl[134] vdd gnd cell_6t
Xbit_r135_c47 bl[47] br[47] wl[135] vdd gnd cell_6t
Xbit_r136_c47 bl[47] br[47] wl[136] vdd gnd cell_6t
Xbit_r137_c47 bl[47] br[47] wl[137] vdd gnd cell_6t
Xbit_r138_c47 bl[47] br[47] wl[138] vdd gnd cell_6t
Xbit_r139_c47 bl[47] br[47] wl[139] vdd gnd cell_6t
Xbit_r140_c47 bl[47] br[47] wl[140] vdd gnd cell_6t
Xbit_r141_c47 bl[47] br[47] wl[141] vdd gnd cell_6t
Xbit_r142_c47 bl[47] br[47] wl[142] vdd gnd cell_6t
Xbit_r143_c47 bl[47] br[47] wl[143] vdd gnd cell_6t
Xbit_r144_c47 bl[47] br[47] wl[144] vdd gnd cell_6t
Xbit_r145_c47 bl[47] br[47] wl[145] vdd gnd cell_6t
Xbit_r146_c47 bl[47] br[47] wl[146] vdd gnd cell_6t
Xbit_r147_c47 bl[47] br[47] wl[147] vdd gnd cell_6t
Xbit_r148_c47 bl[47] br[47] wl[148] vdd gnd cell_6t
Xbit_r149_c47 bl[47] br[47] wl[149] vdd gnd cell_6t
Xbit_r150_c47 bl[47] br[47] wl[150] vdd gnd cell_6t
Xbit_r151_c47 bl[47] br[47] wl[151] vdd gnd cell_6t
Xbit_r152_c47 bl[47] br[47] wl[152] vdd gnd cell_6t
Xbit_r153_c47 bl[47] br[47] wl[153] vdd gnd cell_6t
Xbit_r154_c47 bl[47] br[47] wl[154] vdd gnd cell_6t
Xbit_r155_c47 bl[47] br[47] wl[155] vdd gnd cell_6t
Xbit_r156_c47 bl[47] br[47] wl[156] vdd gnd cell_6t
Xbit_r157_c47 bl[47] br[47] wl[157] vdd gnd cell_6t
Xbit_r158_c47 bl[47] br[47] wl[158] vdd gnd cell_6t
Xbit_r159_c47 bl[47] br[47] wl[159] vdd gnd cell_6t
Xbit_r160_c47 bl[47] br[47] wl[160] vdd gnd cell_6t
Xbit_r161_c47 bl[47] br[47] wl[161] vdd gnd cell_6t
Xbit_r162_c47 bl[47] br[47] wl[162] vdd gnd cell_6t
Xbit_r163_c47 bl[47] br[47] wl[163] vdd gnd cell_6t
Xbit_r164_c47 bl[47] br[47] wl[164] vdd gnd cell_6t
Xbit_r165_c47 bl[47] br[47] wl[165] vdd gnd cell_6t
Xbit_r166_c47 bl[47] br[47] wl[166] vdd gnd cell_6t
Xbit_r167_c47 bl[47] br[47] wl[167] vdd gnd cell_6t
Xbit_r168_c47 bl[47] br[47] wl[168] vdd gnd cell_6t
Xbit_r169_c47 bl[47] br[47] wl[169] vdd gnd cell_6t
Xbit_r170_c47 bl[47] br[47] wl[170] vdd gnd cell_6t
Xbit_r171_c47 bl[47] br[47] wl[171] vdd gnd cell_6t
Xbit_r172_c47 bl[47] br[47] wl[172] vdd gnd cell_6t
Xbit_r173_c47 bl[47] br[47] wl[173] vdd gnd cell_6t
Xbit_r174_c47 bl[47] br[47] wl[174] vdd gnd cell_6t
Xbit_r175_c47 bl[47] br[47] wl[175] vdd gnd cell_6t
Xbit_r176_c47 bl[47] br[47] wl[176] vdd gnd cell_6t
Xbit_r177_c47 bl[47] br[47] wl[177] vdd gnd cell_6t
Xbit_r178_c47 bl[47] br[47] wl[178] vdd gnd cell_6t
Xbit_r179_c47 bl[47] br[47] wl[179] vdd gnd cell_6t
Xbit_r180_c47 bl[47] br[47] wl[180] vdd gnd cell_6t
Xbit_r181_c47 bl[47] br[47] wl[181] vdd gnd cell_6t
Xbit_r182_c47 bl[47] br[47] wl[182] vdd gnd cell_6t
Xbit_r183_c47 bl[47] br[47] wl[183] vdd gnd cell_6t
Xbit_r184_c47 bl[47] br[47] wl[184] vdd gnd cell_6t
Xbit_r185_c47 bl[47] br[47] wl[185] vdd gnd cell_6t
Xbit_r186_c47 bl[47] br[47] wl[186] vdd gnd cell_6t
Xbit_r187_c47 bl[47] br[47] wl[187] vdd gnd cell_6t
Xbit_r188_c47 bl[47] br[47] wl[188] vdd gnd cell_6t
Xbit_r189_c47 bl[47] br[47] wl[189] vdd gnd cell_6t
Xbit_r190_c47 bl[47] br[47] wl[190] vdd gnd cell_6t
Xbit_r191_c47 bl[47] br[47] wl[191] vdd gnd cell_6t
Xbit_r192_c47 bl[47] br[47] wl[192] vdd gnd cell_6t
Xbit_r193_c47 bl[47] br[47] wl[193] vdd gnd cell_6t
Xbit_r194_c47 bl[47] br[47] wl[194] vdd gnd cell_6t
Xbit_r195_c47 bl[47] br[47] wl[195] vdd gnd cell_6t
Xbit_r196_c47 bl[47] br[47] wl[196] vdd gnd cell_6t
Xbit_r197_c47 bl[47] br[47] wl[197] vdd gnd cell_6t
Xbit_r198_c47 bl[47] br[47] wl[198] vdd gnd cell_6t
Xbit_r199_c47 bl[47] br[47] wl[199] vdd gnd cell_6t
Xbit_r200_c47 bl[47] br[47] wl[200] vdd gnd cell_6t
Xbit_r201_c47 bl[47] br[47] wl[201] vdd gnd cell_6t
Xbit_r202_c47 bl[47] br[47] wl[202] vdd gnd cell_6t
Xbit_r203_c47 bl[47] br[47] wl[203] vdd gnd cell_6t
Xbit_r204_c47 bl[47] br[47] wl[204] vdd gnd cell_6t
Xbit_r205_c47 bl[47] br[47] wl[205] vdd gnd cell_6t
Xbit_r206_c47 bl[47] br[47] wl[206] vdd gnd cell_6t
Xbit_r207_c47 bl[47] br[47] wl[207] vdd gnd cell_6t
Xbit_r208_c47 bl[47] br[47] wl[208] vdd gnd cell_6t
Xbit_r209_c47 bl[47] br[47] wl[209] vdd gnd cell_6t
Xbit_r210_c47 bl[47] br[47] wl[210] vdd gnd cell_6t
Xbit_r211_c47 bl[47] br[47] wl[211] vdd gnd cell_6t
Xbit_r212_c47 bl[47] br[47] wl[212] vdd gnd cell_6t
Xbit_r213_c47 bl[47] br[47] wl[213] vdd gnd cell_6t
Xbit_r214_c47 bl[47] br[47] wl[214] vdd gnd cell_6t
Xbit_r215_c47 bl[47] br[47] wl[215] vdd gnd cell_6t
Xbit_r216_c47 bl[47] br[47] wl[216] vdd gnd cell_6t
Xbit_r217_c47 bl[47] br[47] wl[217] vdd gnd cell_6t
Xbit_r218_c47 bl[47] br[47] wl[218] vdd gnd cell_6t
Xbit_r219_c47 bl[47] br[47] wl[219] vdd gnd cell_6t
Xbit_r220_c47 bl[47] br[47] wl[220] vdd gnd cell_6t
Xbit_r221_c47 bl[47] br[47] wl[221] vdd gnd cell_6t
Xbit_r222_c47 bl[47] br[47] wl[222] vdd gnd cell_6t
Xbit_r223_c47 bl[47] br[47] wl[223] vdd gnd cell_6t
Xbit_r224_c47 bl[47] br[47] wl[224] vdd gnd cell_6t
Xbit_r225_c47 bl[47] br[47] wl[225] vdd gnd cell_6t
Xbit_r226_c47 bl[47] br[47] wl[226] vdd gnd cell_6t
Xbit_r227_c47 bl[47] br[47] wl[227] vdd gnd cell_6t
Xbit_r228_c47 bl[47] br[47] wl[228] vdd gnd cell_6t
Xbit_r229_c47 bl[47] br[47] wl[229] vdd gnd cell_6t
Xbit_r230_c47 bl[47] br[47] wl[230] vdd gnd cell_6t
Xbit_r231_c47 bl[47] br[47] wl[231] vdd gnd cell_6t
Xbit_r232_c47 bl[47] br[47] wl[232] vdd gnd cell_6t
Xbit_r233_c47 bl[47] br[47] wl[233] vdd gnd cell_6t
Xbit_r234_c47 bl[47] br[47] wl[234] vdd gnd cell_6t
Xbit_r235_c47 bl[47] br[47] wl[235] vdd gnd cell_6t
Xbit_r236_c47 bl[47] br[47] wl[236] vdd gnd cell_6t
Xbit_r237_c47 bl[47] br[47] wl[237] vdd gnd cell_6t
Xbit_r238_c47 bl[47] br[47] wl[238] vdd gnd cell_6t
Xbit_r239_c47 bl[47] br[47] wl[239] vdd gnd cell_6t
Xbit_r240_c47 bl[47] br[47] wl[240] vdd gnd cell_6t
Xbit_r241_c47 bl[47] br[47] wl[241] vdd gnd cell_6t
Xbit_r242_c47 bl[47] br[47] wl[242] vdd gnd cell_6t
Xbit_r243_c47 bl[47] br[47] wl[243] vdd gnd cell_6t
Xbit_r244_c47 bl[47] br[47] wl[244] vdd gnd cell_6t
Xbit_r245_c47 bl[47] br[47] wl[245] vdd gnd cell_6t
Xbit_r246_c47 bl[47] br[47] wl[246] vdd gnd cell_6t
Xbit_r247_c47 bl[47] br[47] wl[247] vdd gnd cell_6t
Xbit_r248_c47 bl[47] br[47] wl[248] vdd gnd cell_6t
Xbit_r249_c47 bl[47] br[47] wl[249] vdd gnd cell_6t
Xbit_r250_c47 bl[47] br[47] wl[250] vdd gnd cell_6t
Xbit_r251_c47 bl[47] br[47] wl[251] vdd gnd cell_6t
Xbit_r252_c47 bl[47] br[47] wl[252] vdd gnd cell_6t
Xbit_r253_c47 bl[47] br[47] wl[253] vdd gnd cell_6t
Xbit_r254_c47 bl[47] br[47] wl[254] vdd gnd cell_6t
Xbit_r255_c47 bl[47] br[47] wl[255] vdd gnd cell_6t
Xbit_r0_c48 bl[48] br[48] wl[0] vdd gnd cell_6t
Xbit_r1_c48 bl[48] br[48] wl[1] vdd gnd cell_6t
Xbit_r2_c48 bl[48] br[48] wl[2] vdd gnd cell_6t
Xbit_r3_c48 bl[48] br[48] wl[3] vdd gnd cell_6t
Xbit_r4_c48 bl[48] br[48] wl[4] vdd gnd cell_6t
Xbit_r5_c48 bl[48] br[48] wl[5] vdd gnd cell_6t
Xbit_r6_c48 bl[48] br[48] wl[6] vdd gnd cell_6t
Xbit_r7_c48 bl[48] br[48] wl[7] vdd gnd cell_6t
Xbit_r8_c48 bl[48] br[48] wl[8] vdd gnd cell_6t
Xbit_r9_c48 bl[48] br[48] wl[9] vdd gnd cell_6t
Xbit_r10_c48 bl[48] br[48] wl[10] vdd gnd cell_6t
Xbit_r11_c48 bl[48] br[48] wl[11] vdd gnd cell_6t
Xbit_r12_c48 bl[48] br[48] wl[12] vdd gnd cell_6t
Xbit_r13_c48 bl[48] br[48] wl[13] vdd gnd cell_6t
Xbit_r14_c48 bl[48] br[48] wl[14] vdd gnd cell_6t
Xbit_r15_c48 bl[48] br[48] wl[15] vdd gnd cell_6t
Xbit_r16_c48 bl[48] br[48] wl[16] vdd gnd cell_6t
Xbit_r17_c48 bl[48] br[48] wl[17] vdd gnd cell_6t
Xbit_r18_c48 bl[48] br[48] wl[18] vdd gnd cell_6t
Xbit_r19_c48 bl[48] br[48] wl[19] vdd gnd cell_6t
Xbit_r20_c48 bl[48] br[48] wl[20] vdd gnd cell_6t
Xbit_r21_c48 bl[48] br[48] wl[21] vdd gnd cell_6t
Xbit_r22_c48 bl[48] br[48] wl[22] vdd gnd cell_6t
Xbit_r23_c48 bl[48] br[48] wl[23] vdd gnd cell_6t
Xbit_r24_c48 bl[48] br[48] wl[24] vdd gnd cell_6t
Xbit_r25_c48 bl[48] br[48] wl[25] vdd gnd cell_6t
Xbit_r26_c48 bl[48] br[48] wl[26] vdd gnd cell_6t
Xbit_r27_c48 bl[48] br[48] wl[27] vdd gnd cell_6t
Xbit_r28_c48 bl[48] br[48] wl[28] vdd gnd cell_6t
Xbit_r29_c48 bl[48] br[48] wl[29] vdd gnd cell_6t
Xbit_r30_c48 bl[48] br[48] wl[30] vdd gnd cell_6t
Xbit_r31_c48 bl[48] br[48] wl[31] vdd gnd cell_6t
Xbit_r32_c48 bl[48] br[48] wl[32] vdd gnd cell_6t
Xbit_r33_c48 bl[48] br[48] wl[33] vdd gnd cell_6t
Xbit_r34_c48 bl[48] br[48] wl[34] vdd gnd cell_6t
Xbit_r35_c48 bl[48] br[48] wl[35] vdd gnd cell_6t
Xbit_r36_c48 bl[48] br[48] wl[36] vdd gnd cell_6t
Xbit_r37_c48 bl[48] br[48] wl[37] vdd gnd cell_6t
Xbit_r38_c48 bl[48] br[48] wl[38] vdd gnd cell_6t
Xbit_r39_c48 bl[48] br[48] wl[39] vdd gnd cell_6t
Xbit_r40_c48 bl[48] br[48] wl[40] vdd gnd cell_6t
Xbit_r41_c48 bl[48] br[48] wl[41] vdd gnd cell_6t
Xbit_r42_c48 bl[48] br[48] wl[42] vdd gnd cell_6t
Xbit_r43_c48 bl[48] br[48] wl[43] vdd gnd cell_6t
Xbit_r44_c48 bl[48] br[48] wl[44] vdd gnd cell_6t
Xbit_r45_c48 bl[48] br[48] wl[45] vdd gnd cell_6t
Xbit_r46_c48 bl[48] br[48] wl[46] vdd gnd cell_6t
Xbit_r47_c48 bl[48] br[48] wl[47] vdd gnd cell_6t
Xbit_r48_c48 bl[48] br[48] wl[48] vdd gnd cell_6t
Xbit_r49_c48 bl[48] br[48] wl[49] vdd gnd cell_6t
Xbit_r50_c48 bl[48] br[48] wl[50] vdd gnd cell_6t
Xbit_r51_c48 bl[48] br[48] wl[51] vdd gnd cell_6t
Xbit_r52_c48 bl[48] br[48] wl[52] vdd gnd cell_6t
Xbit_r53_c48 bl[48] br[48] wl[53] vdd gnd cell_6t
Xbit_r54_c48 bl[48] br[48] wl[54] vdd gnd cell_6t
Xbit_r55_c48 bl[48] br[48] wl[55] vdd gnd cell_6t
Xbit_r56_c48 bl[48] br[48] wl[56] vdd gnd cell_6t
Xbit_r57_c48 bl[48] br[48] wl[57] vdd gnd cell_6t
Xbit_r58_c48 bl[48] br[48] wl[58] vdd gnd cell_6t
Xbit_r59_c48 bl[48] br[48] wl[59] vdd gnd cell_6t
Xbit_r60_c48 bl[48] br[48] wl[60] vdd gnd cell_6t
Xbit_r61_c48 bl[48] br[48] wl[61] vdd gnd cell_6t
Xbit_r62_c48 bl[48] br[48] wl[62] vdd gnd cell_6t
Xbit_r63_c48 bl[48] br[48] wl[63] vdd gnd cell_6t
Xbit_r64_c48 bl[48] br[48] wl[64] vdd gnd cell_6t
Xbit_r65_c48 bl[48] br[48] wl[65] vdd gnd cell_6t
Xbit_r66_c48 bl[48] br[48] wl[66] vdd gnd cell_6t
Xbit_r67_c48 bl[48] br[48] wl[67] vdd gnd cell_6t
Xbit_r68_c48 bl[48] br[48] wl[68] vdd gnd cell_6t
Xbit_r69_c48 bl[48] br[48] wl[69] vdd gnd cell_6t
Xbit_r70_c48 bl[48] br[48] wl[70] vdd gnd cell_6t
Xbit_r71_c48 bl[48] br[48] wl[71] vdd gnd cell_6t
Xbit_r72_c48 bl[48] br[48] wl[72] vdd gnd cell_6t
Xbit_r73_c48 bl[48] br[48] wl[73] vdd gnd cell_6t
Xbit_r74_c48 bl[48] br[48] wl[74] vdd gnd cell_6t
Xbit_r75_c48 bl[48] br[48] wl[75] vdd gnd cell_6t
Xbit_r76_c48 bl[48] br[48] wl[76] vdd gnd cell_6t
Xbit_r77_c48 bl[48] br[48] wl[77] vdd gnd cell_6t
Xbit_r78_c48 bl[48] br[48] wl[78] vdd gnd cell_6t
Xbit_r79_c48 bl[48] br[48] wl[79] vdd gnd cell_6t
Xbit_r80_c48 bl[48] br[48] wl[80] vdd gnd cell_6t
Xbit_r81_c48 bl[48] br[48] wl[81] vdd gnd cell_6t
Xbit_r82_c48 bl[48] br[48] wl[82] vdd gnd cell_6t
Xbit_r83_c48 bl[48] br[48] wl[83] vdd gnd cell_6t
Xbit_r84_c48 bl[48] br[48] wl[84] vdd gnd cell_6t
Xbit_r85_c48 bl[48] br[48] wl[85] vdd gnd cell_6t
Xbit_r86_c48 bl[48] br[48] wl[86] vdd gnd cell_6t
Xbit_r87_c48 bl[48] br[48] wl[87] vdd gnd cell_6t
Xbit_r88_c48 bl[48] br[48] wl[88] vdd gnd cell_6t
Xbit_r89_c48 bl[48] br[48] wl[89] vdd gnd cell_6t
Xbit_r90_c48 bl[48] br[48] wl[90] vdd gnd cell_6t
Xbit_r91_c48 bl[48] br[48] wl[91] vdd gnd cell_6t
Xbit_r92_c48 bl[48] br[48] wl[92] vdd gnd cell_6t
Xbit_r93_c48 bl[48] br[48] wl[93] vdd gnd cell_6t
Xbit_r94_c48 bl[48] br[48] wl[94] vdd gnd cell_6t
Xbit_r95_c48 bl[48] br[48] wl[95] vdd gnd cell_6t
Xbit_r96_c48 bl[48] br[48] wl[96] vdd gnd cell_6t
Xbit_r97_c48 bl[48] br[48] wl[97] vdd gnd cell_6t
Xbit_r98_c48 bl[48] br[48] wl[98] vdd gnd cell_6t
Xbit_r99_c48 bl[48] br[48] wl[99] vdd gnd cell_6t
Xbit_r100_c48 bl[48] br[48] wl[100] vdd gnd cell_6t
Xbit_r101_c48 bl[48] br[48] wl[101] vdd gnd cell_6t
Xbit_r102_c48 bl[48] br[48] wl[102] vdd gnd cell_6t
Xbit_r103_c48 bl[48] br[48] wl[103] vdd gnd cell_6t
Xbit_r104_c48 bl[48] br[48] wl[104] vdd gnd cell_6t
Xbit_r105_c48 bl[48] br[48] wl[105] vdd gnd cell_6t
Xbit_r106_c48 bl[48] br[48] wl[106] vdd gnd cell_6t
Xbit_r107_c48 bl[48] br[48] wl[107] vdd gnd cell_6t
Xbit_r108_c48 bl[48] br[48] wl[108] vdd gnd cell_6t
Xbit_r109_c48 bl[48] br[48] wl[109] vdd gnd cell_6t
Xbit_r110_c48 bl[48] br[48] wl[110] vdd gnd cell_6t
Xbit_r111_c48 bl[48] br[48] wl[111] vdd gnd cell_6t
Xbit_r112_c48 bl[48] br[48] wl[112] vdd gnd cell_6t
Xbit_r113_c48 bl[48] br[48] wl[113] vdd gnd cell_6t
Xbit_r114_c48 bl[48] br[48] wl[114] vdd gnd cell_6t
Xbit_r115_c48 bl[48] br[48] wl[115] vdd gnd cell_6t
Xbit_r116_c48 bl[48] br[48] wl[116] vdd gnd cell_6t
Xbit_r117_c48 bl[48] br[48] wl[117] vdd gnd cell_6t
Xbit_r118_c48 bl[48] br[48] wl[118] vdd gnd cell_6t
Xbit_r119_c48 bl[48] br[48] wl[119] vdd gnd cell_6t
Xbit_r120_c48 bl[48] br[48] wl[120] vdd gnd cell_6t
Xbit_r121_c48 bl[48] br[48] wl[121] vdd gnd cell_6t
Xbit_r122_c48 bl[48] br[48] wl[122] vdd gnd cell_6t
Xbit_r123_c48 bl[48] br[48] wl[123] vdd gnd cell_6t
Xbit_r124_c48 bl[48] br[48] wl[124] vdd gnd cell_6t
Xbit_r125_c48 bl[48] br[48] wl[125] vdd gnd cell_6t
Xbit_r126_c48 bl[48] br[48] wl[126] vdd gnd cell_6t
Xbit_r127_c48 bl[48] br[48] wl[127] vdd gnd cell_6t
Xbit_r128_c48 bl[48] br[48] wl[128] vdd gnd cell_6t
Xbit_r129_c48 bl[48] br[48] wl[129] vdd gnd cell_6t
Xbit_r130_c48 bl[48] br[48] wl[130] vdd gnd cell_6t
Xbit_r131_c48 bl[48] br[48] wl[131] vdd gnd cell_6t
Xbit_r132_c48 bl[48] br[48] wl[132] vdd gnd cell_6t
Xbit_r133_c48 bl[48] br[48] wl[133] vdd gnd cell_6t
Xbit_r134_c48 bl[48] br[48] wl[134] vdd gnd cell_6t
Xbit_r135_c48 bl[48] br[48] wl[135] vdd gnd cell_6t
Xbit_r136_c48 bl[48] br[48] wl[136] vdd gnd cell_6t
Xbit_r137_c48 bl[48] br[48] wl[137] vdd gnd cell_6t
Xbit_r138_c48 bl[48] br[48] wl[138] vdd gnd cell_6t
Xbit_r139_c48 bl[48] br[48] wl[139] vdd gnd cell_6t
Xbit_r140_c48 bl[48] br[48] wl[140] vdd gnd cell_6t
Xbit_r141_c48 bl[48] br[48] wl[141] vdd gnd cell_6t
Xbit_r142_c48 bl[48] br[48] wl[142] vdd gnd cell_6t
Xbit_r143_c48 bl[48] br[48] wl[143] vdd gnd cell_6t
Xbit_r144_c48 bl[48] br[48] wl[144] vdd gnd cell_6t
Xbit_r145_c48 bl[48] br[48] wl[145] vdd gnd cell_6t
Xbit_r146_c48 bl[48] br[48] wl[146] vdd gnd cell_6t
Xbit_r147_c48 bl[48] br[48] wl[147] vdd gnd cell_6t
Xbit_r148_c48 bl[48] br[48] wl[148] vdd gnd cell_6t
Xbit_r149_c48 bl[48] br[48] wl[149] vdd gnd cell_6t
Xbit_r150_c48 bl[48] br[48] wl[150] vdd gnd cell_6t
Xbit_r151_c48 bl[48] br[48] wl[151] vdd gnd cell_6t
Xbit_r152_c48 bl[48] br[48] wl[152] vdd gnd cell_6t
Xbit_r153_c48 bl[48] br[48] wl[153] vdd gnd cell_6t
Xbit_r154_c48 bl[48] br[48] wl[154] vdd gnd cell_6t
Xbit_r155_c48 bl[48] br[48] wl[155] vdd gnd cell_6t
Xbit_r156_c48 bl[48] br[48] wl[156] vdd gnd cell_6t
Xbit_r157_c48 bl[48] br[48] wl[157] vdd gnd cell_6t
Xbit_r158_c48 bl[48] br[48] wl[158] vdd gnd cell_6t
Xbit_r159_c48 bl[48] br[48] wl[159] vdd gnd cell_6t
Xbit_r160_c48 bl[48] br[48] wl[160] vdd gnd cell_6t
Xbit_r161_c48 bl[48] br[48] wl[161] vdd gnd cell_6t
Xbit_r162_c48 bl[48] br[48] wl[162] vdd gnd cell_6t
Xbit_r163_c48 bl[48] br[48] wl[163] vdd gnd cell_6t
Xbit_r164_c48 bl[48] br[48] wl[164] vdd gnd cell_6t
Xbit_r165_c48 bl[48] br[48] wl[165] vdd gnd cell_6t
Xbit_r166_c48 bl[48] br[48] wl[166] vdd gnd cell_6t
Xbit_r167_c48 bl[48] br[48] wl[167] vdd gnd cell_6t
Xbit_r168_c48 bl[48] br[48] wl[168] vdd gnd cell_6t
Xbit_r169_c48 bl[48] br[48] wl[169] vdd gnd cell_6t
Xbit_r170_c48 bl[48] br[48] wl[170] vdd gnd cell_6t
Xbit_r171_c48 bl[48] br[48] wl[171] vdd gnd cell_6t
Xbit_r172_c48 bl[48] br[48] wl[172] vdd gnd cell_6t
Xbit_r173_c48 bl[48] br[48] wl[173] vdd gnd cell_6t
Xbit_r174_c48 bl[48] br[48] wl[174] vdd gnd cell_6t
Xbit_r175_c48 bl[48] br[48] wl[175] vdd gnd cell_6t
Xbit_r176_c48 bl[48] br[48] wl[176] vdd gnd cell_6t
Xbit_r177_c48 bl[48] br[48] wl[177] vdd gnd cell_6t
Xbit_r178_c48 bl[48] br[48] wl[178] vdd gnd cell_6t
Xbit_r179_c48 bl[48] br[48] wl[179] vdd gnd cell_6t
Xbit_r180_c48 bl[48] br[48] wl[180] vdd gnd cell_6t
Xbit_r181_c48 bl[48] br[48] wl[181] vdd gnd cell_6t
Xbit_r182_c48 bl[48] br[48] wl[182] vdd gnd cell_6t
Xbit_r183_c48 bl[48] br[48] wl[183] vdd gnd cell_6t
Xbit_r184_c48 bl[48] br[48] wl[184] vdd gnd cell_6t
Xbit_r185_c48 bl[48] br[48] wl[185] vdd gnd cell_6t
Xbit_r186_c48 bl[48] br[48] wl[186] vdd gnd cell_6t
Xbit_r187_c48 bl[48] br[48] wl[187] vdd gnd cell_6t
Xbit_r188_c48 bl[48] br[48] wl[188] vdd gnd cell_6t
Xbit_r189_c48 bl[48] br[48] wl[189] vdd gnd cell_6t
Xbit_r190_c48 bl[48] br[48] wl[190] vdd gnd cell_6t
Xbit_r191_c48 bl[48] br[48] wl[191] vdd gnd cell_6t
Xbit_r192_c48 bl[48] br[48] wl[192] vdd gnd cell_6t
Xbit_r193_c48 bl[48] br[48] wl[193] vdd gnd cell_6t
Xbit_r194_c48 bl[48] br[48] wl[194] vdd gnd cell_6t
Xbit_r195_c48 bl[48] br[48] wl[195] vdd gnd cell_6t
Xbit_r196_c48 bl[48] br[48] wl[196] vdd gnd cell_6t
Xbit_r197_c48 bl[48] br[48] wl[197] vdd gnd cell_6t
Xbit_r198_c48 bl[48] br[48] wl[198] vdd gnd cell_6t
Xbit_r199_c48 bl[48] br[48] wl[199] vdd gnd cell_6t
Xbit_r200_c48 bl[48] br[48] wl[200] vdd gnd cell_6t
Xbit_r201_c48 bl[48] br[48] wl[201] vdd gnd cell_6t
Xbit_r202_c48 bl[48] br[48] wl[202] vdd gnd cell_6t
Xbit_r203_c48 bl[48] br[48] wl[203] vdd gnd cell_6t
Xbit_r204_c48 bl[48] br[48] wl[204] vdd gnd cell_6t
Xbit_r205_c48 bl[48] br[48] wl[205] vdd gnd cell_6t
Xbit_r206_c48 bl[48] br[48] wl[206] vdd gnd cell_6t
Xbit_r207_c48 bl[48] br[48] wl[207] vdd gnd cell_6t
Xbit_r208_c48 bl[48] br[48] wl[208] vdd gnd cell_6t
Xbit_r209_c48 bl[48] br[48] wl[209] vdd gnd cell_6t
Xbit_r210_c48 bl[48] br[48] wl[210] vdd gnd cell_6t
Xbit_r211_c48 bl[48] br[48] wl[211] vdd gnd cell_6t
Xbit_r212_c48 bl[48] br[48] wl[212] vdd gnd cell_6t
Xbit_r213_c48 bl[48] br[48] wl[213] vdd gnd cell_6t
Xbit_r214_c48 bl[48] br[48] wl[214] vdd gnd cell_6t
Xbit_r215_c48 bl[48] br[48] wl[215] vdd gnd cell_6t
Xbit_r216_c48 bl[48] br[48] wl[216] vdd gnd cell_6t
Xbit_r217_c48 bl[48] br[48] wl[217] vdd gnd cell_6t
Xbit_r218_c48 bl[48] br[48] wl[218] vdd gnd cell_6t
Xbit_r219_c48 bl[48] br[48] wl[219] vdd gnd cell_6t
Xbit_r220_c48 bl[48] br[48] wl[220] vdd gnd cell_6t
Xbit_r221_c48 bl[48] br[48] wl[221] vdd gnd cell_6t
Xbit_r222_c48 bl[48] br[48] wl[222] vdd gnd cell_6t
Xbit_r223_c48 bl[48] br[48] wl[223] vdd gnd cell_6t
Xbit_r224_c48 bl[48] br[48] wl[224] vdd gnd cell_6t
Xbit_r225_c48 bl[48] br[48] wl[225] vdd gnd cell_6t
Xbit_r226_c48 bl[48] br[48] wl[226] vdd gnd cell_6t
Xbit_r227_c48 bl[48] br[48] wl[227] vdd gnd cell_6t
Xbit_r228_c48 bl[48] br[48] wl[228] vdd gnd cell_6t
Xbit_r229_c48 bl[48] br[48] wl[229] vdd gnd cell_6t
Xbit_r230_c48 bl[48] br[48] wl[230] vdd gnd cell_6t
Xbit_r231_c48 bl[48] br[48] wl[231] vdd gnd cell_6t
Xbit_r232_c48 bl[48] br[48] wl[232] vdd gnd cell_6t
Xbit_r233_c48 bl[48] br[48] wl[233] vdd gnd cell_6t
Xbit_r234_c48 bl[48] br[48] wl[234] vdd gnd cell_6t
Xbit_r235_c48 bl[48] br[48] wl[235] vdd gnd cell_6t
Xbit_r236_c48 bl[48] br[48] wl[236] vdd gnd cell_6t
Xbit_r237_c48 bl[48] br[48] wl[237] vdd gnd cell_6t
Xbit_r238_c48 bl[48] br[48] wl[238] vdd gnd cell_6t
Xbit_r239_c48 bl[48] br[48] wl[239] vdd gnd cell_6t
Xbit_r240_c48 bl[48] br[48] wl[240] vdd gnd cell_6t
Xbit_r241_c48 bl[48] br[48] wl[241] vdd gnd cell_6t
Xbit_r242_c48 bl[48] br[48] wl[242] vdd gnd cell_6t
Xbit_r243_c48 bl[48] br[48] wl[243] vdd gnd cell_6t
Xbit_r244_c48 bl[48] br[48] wl[244] vdd gnd cell_6t
Xbit_r245_c48 bl[48] br[48] wl[245] vdd gnd cell_6t
Xbit_r246_c48 bl[48] br[48] wl[246] vdd gnd cell_6t
Xbit_r247_c48 bl[48] br[48] wl[247] vdd gnd cell_6t
Xbit_r248_c48 bl[48] br[48] wl[248] vdd gnd cell_6t
Xbit_r249_c48 bl[48] br[48] wl[249] vdd gnd cell_6t
Xbit_r250_c48 bl[48] br[48] wl[250] vdd gnd cell_6t
Xbit_r251_c48 bl[48] br[48] wl[251] vdd gnd cell_6t
Xbit_r252_c48 bl[48] br[48] wl[252] vdd gnd cell_6t
Xbit_r253_c48 bl[48] br[48] wl[253] vdd gnd cell_6t
Xbit_r254_c48 bl[48] br[48] wl[254] vdd gnd cell_6t
Xbit_r255_c48 bl[48] br[48] wl[255] vdd gnd cell_6t
Xbit_r0_c49 bl[49] br[49] wl[0] vdd gnd cell_6t
Xbit_r1_c49 bl[49] br[49] wl[1] vdd gnd cell_6t
Xbit_r2_c49 bl[49] br[49] wl[2] vdd gnd cell_6t
Xbit_r3_c49 bl[49] br[49] wl[3] vdd gnd cell_6t
Xbit_r4_c49 bl[49] br[49] wl[4] vdd gnd cell_6t
Xbit_r5_c49 bl[49] br[49] wl[5] vdd gnd cell_6t
Xbit_r6_c49 bl[49] br[49] wl[6] vdd gnd cell_6t
Xbit_r7_c49 bl[49] br[49] wl[7] vdd gnd cell_6t
Xbit_r8_c49 bl[49] br[49] wl[8] vdd gnd cell_6t
Xbit_r9_c49 bl[49] br[49] wl[9] vdd gnd cell_6t
Xbit_r10_c49 bl[49] br[49] wl[10] vdd gnd cell_6t
Xbit_r11_c49 bl[49] br[49] wl[11] vdd gnd cell_6t
Xbit_r12_c49 bl[49] br[49] wl[12] vdd gnd cell_6t
Xbit_r13_c49 bl[49] br[49] wl[13] vdd gnd cell_6t
Xbit_r14_c49 bl[49] br[49] wl[14] vdd gnd cell_6t
Xbit_r15_c49 bl[49] br[49] wl[15] vdd gnd cell_6t
Xbit_r16_c49 bl[49] br[49] wl[16] vdd gnd cell_6t
Xbit_r17_c49 bl[49] br[49] wl[17] vdd gnd cell_6t
Xbit_r18_c49 bl[49] br[49] wl[18] vdd gnd cell_6t
Xbit_r19_c49 bl[49] br[49] wl[19] vdd gnd cell_6t
Xbit_r20_c49 bl[49] br[49] wl[20] vdd gnd cell_6t
Xbit_r21_c49 bl[49] br[49] wl[21] vdd gnd cell_6t
Xbit_r22_c49 bl[49] br[49] wl[22] vdd gnd cell_6t
Xbit_r23_c49 bl[49] br[49] wl[23] vdd gnd cell_6t
Xbit_r24_c49 bl[49] br[49] wl[24] vdd gnd cell_6t
Xbit_r25_c49 bl[49] br[49] wl[25] vdd gnd cell_6t
Xbit_r26_c49 bl[49] br[49] wl[26] vdd gnd cell_6t
Xbit_r27_c49 bl[49] br[49] wl[27] vdd gnd cell_6t
Xbit_r28_c49 bl[49] br[49] wl[28] vdd gnd cell_6t
Xbit_r29_c49 bl[49] br[49] wl[29] vdd gnd cell_6t
Xbit_r30_c49 bl[49] br[49] wl[30] vdd gnd cell_6t
Xbit_r31_c49 bl[49] br[49] wl[31] vdd gnd cell_6t
Xbit_r32_c49 bl[49] br[49] wl[32] vdd gnd cell_6t
Xbit_r33_c49 bl[49] br[49] wl[33] vdd gnd cell_6t
Xbit_r34_c49 bl[49] br[49] wl[34] vdd gnd cell_6t
Xbit_r35_c49 bl[49] br[49] wl[35] vdd gnd cell_6t
Xbit_r36_c49 bl[49] br[49] wl[36] vdd gnd cell_6t
Xbit_r37_c49 bl[49] br[49] wl[37] vdd gnd cell_6t
Xbit_r38_c49 bl[49] br[49] wl[38] vdd gnd cell_6t
Xbit_r39_c49 bl[49] br[49] wl[39] vdd gnd cell_6t
Xbit_r40_c49 bl[49] br[49] wl[40] vdd gnd cell_6t
Xbit_r41_c49 bl[49] br[49] wl[41] vdd gnd cell_6t
Xbit_r42_c49 bl[49] br[49] wl[42] vdd gnd cell_6t
Xbit_r43_c49 bl[49] br[49] wl[43] vdd gnd cell_6t
Xbit_r44_c49 bl[49] br[49] wl[44] vdd gnd cell_6t
Xbit_r45_c49 bl[49] br[49] wl[45] vdd gnd cell_6t
Xbit_r46_c49 bl[49] br[49] wl[46] vdd gnd cell_6t
Xbit_r47_c49 bl[49] br[49] wl[47] vdd gnd cell_6t
Xbit_r48_c49 bl[49] br[49] wl[48] vdd gnd cell_6t
Xbit_r49_c49 bl[49] br[49] wl[49] vdd gnd cell_6t
Xbit_r50_c49 bl[49] br[49] wl[50] vdd gnd cell_6t
Xbit_r51_c49 bl[49] br[49] wl[51] vdd gnd cell_6t
Xbit_r52_c49 bl[49] br[49] wl[52] vdd gnd cell_6t
Xbit_r53_c49 bl[49] br[49] wl[53] vdd gnd cell_6t
Xbit_r54_c49 bl[49] br[49] wl[54] vdd gnd cell_6t
Xbit_r55_c49 bl[49] br[49] wl[55] vdd gnd cell_6t
Xbit_r56_c49 bl[49] br[49] wl[56] vdd gnd cell_6t
Xbit_r57_c49 bl[49] br[49] wl[57] vdd gnd cell_6t
Xbit_r58_c49 bl[49] br[49] wl[58] vdd gnd cell_6t
Xbit_r59_c49 bl[49] br[49] wl[59] vdd gnd cell_6t
Xbit_r60_c49 bl[49] br[49] wl[60] vdd gnd cell_6t
Xbit_r61_c49 bl[49] br[49] wl[61] vdd gnd cell_6t
Xbit_r62_c49 bl[49] br[49] wl[62] vdd gnd cell_6t
Xbit_r63_c49 bl[49] br[49] wl[63] vdd gnd cell_6t
Xbit_r64_c49 bl[49] br[49] wl[64] vdd gnd cell_6t
Xbit_r65_c49 bl[49] br[49] wl[65] vdd gnd cell_6t
Xbit_r66_c49 bl[49] br[49] wl[66] vdd gnd cell_6t
Xbit_r67_c49 bl[49] br[49] wl[67] vdd gnd cell_6t
Xbit_r68_c49 bl[49] br[49] wl[68] vdd gnd cell_6t
Xbit_r69_c49 bl[49] br[49] wl[69] vdd gnd cell_6t
Xbit_r70_c49 bl[49] br[49] wl[70] vdd gnd cell_6t
Xbit_r71_c49 bl[49] br[49] wl[71] vdd gnd cell_6t
Xbit_r72_c49 bl[49] br[49] wl[72] vdd gnd cell_6t
Xbit_r73_c49 bl[49] br[49] wl[73] vdd gnd cell_6t
Xbit_r74_c49 bl[49] br[49] wl[74] vdd gnd cell_6t
Xbit_r75_c49 bl[49] br[49] wl[75] vdd gnd cell_6t
Xbit_r76_c49 bl[49] br[49] wl[76] vdd gnd cell_6t
Xbit_r77_c49 bl[49] br[49] wl[77] vdd gnd cell_6t
Xbit_r78_c49 bl[49] br[49] wl[78] vdd gnd cell_6t
Xbit_r79_c49 bl[49] br[49] wl[79] vdd gnd cell_6t
Xbit_r80_c49 bl[49] br[49] wl[80] vdd gnd cell_6t
Xbit_r81_c49 bl[49] br[49] wl[81] vdd gnd cell_6t
Xbit_r82_c49 bl[49] br[49] wl[82] vdd gnd cell_6t
Xbit_r83_c49 bl[49] br[49] wl[83] vdd gnd cell_6t
Xbit_r84_c49 bl[49] br[49] wl[84] vdd gnd cell_6t
Xbit_r85_c49 bl[49] br[49] wl[85] vdd gnd cell_6t
Xbit_r86_c49 bl[49] br[49] wl[86] vdd gnd cell_6t
Xbit_r87_c49 bl[49] br[49] wl[87] vdd gnd cell_6t
Xbit_r88_c49 bl[49] br[49] wl[88] vdd gnd cell_6t
Xbit_r89_c49 bl[49] br[49] wl[89] vdd gnd cell_6t
Xbit_r90_c49 bl[49] br[49] wl[90] vdd gnd cell_6t
Xbit_r91_c49 bl[49] br[49] wl[91] vdd gnd cell_6t
Xbit_r92_c49 bl[49] br[49] wl[92] vdd gnd cell_6t
Xbit_r93_c49 bl[49] br[49] wl[93] vdd gnd cell_6t
Xbit_r94_c49 bl[49] br[49] wl[94] vdd gnd cell_6t
Xbit_r95_c49 bl[49] br[49] wl[95] vdd gnd cell_6t
Xbit_r96_c49 bl[49] br[49] wl[96] vdd gnd cell_6t
Xbit_r97_c49 bl[49] br[49] wl[97] vdd gnd cell_6t
Xbit_r98_c49 bl[49] br[49] wl[98] vdd gnd cell_6t
Xbit_r99_c49 bl[49] br[49] wl[99] vdd gnd cell_6t
Xbit_r100_c49 bl[49] br[49] wl[100] vdd gnd cell_6t
Xbit_r101_c49 bl[49] br[49] wl[101] vdd gnd cell_6t
Xbit_r102_c49 bl[49] br[49] wl[102] vdd gnd cell_6t
Xbit_r103_c49 bl[49] br[49] wl[103] vdd gnd cell_6t
Xbit_r104_c49 bl[49] br[49] wl[104] vdd gnd cell_6t
Xbit_r105_c49 bl[49] br[49] wl[105] vdd gnd cell_6t
Xbit_r106_c49 bl[49] br[49] wl[106] vdd gnd cell_6t
Xbit_r107_c49 bl[49] br[49] wl[107] vdd gnd cell_6t
Xbit_r108_c49 bl[49] br[49] wl[108] vdd gnd cell_6t
Xbit_r109_c49 bl[49] br[49] wl[109] vdd gnd cell_6t
Xbit_r110_c49 bl[49] br[49] wl[110] vdd gnd cell_6t
Xbit_r111_c49 bl[49] br[49] wl[111] vdd gnd cell_6t
Xbit_r112_c49 bl[49] br[49] wl[112] vdd gnd cell_6t
Xbit_r113_c49 bl[49] br[49] wl[113] vdd gnd cell_6t
Xbit_r114_c49 bl[49] br[49] wl[114] vdd gnd cell_6t
Xbit_r115_c49 bl[49] br[49] wl[115] vdd gnd cell_6t
Xbit_r116_c49 bl[49] br[49] wl[116] vdd gnd cell_6t
Xbit_r117_c49 bl[49] br[49] wl[117] vdd gnd cell_6t
Xbit_r118_c49 bl[49] br[49] wl[118] vdd gnd cell_6t
Xbit_r119_c49 bl[49] br[49] wl[119] vdd gnd cell_6t
Xbit_r120_c49 bl[49] br[49] wl[120] vdd gnd cell_6t
Xbit_r121_c49 bl[49] br[49] wl[121] vdd gnd cell_6t
Xbit_r122_c49 bl[49] br[49] wl[122] vdd gnd cell_6t
Xbit_r123_c49 bl[49] br[49] wl[123] vdd gnd cell_6t
Xbit_r124_c49 bl[49] br[49] wl[124] vdd gnd cell_6t
Xbit_r125_c49 bl[49] br[49] wl[125] vdd gnd cell_6t
Xbit_r126_c49 bl[49] br[49] wl[126] vdd gnd cell_6t
Xbit_r127_c49 bl[49] br[49] wl[127] vdd gnd cell_6t
Xbit_r128_c49 bl[49] br[49] wl[128] vdd gnd cell_6t
Xbit_r129_c49 bl[49] br[49] wl[129] vdd gnd cell_6t
Xbit_r130_c49 bl[49] br[49] wl[130] vdd gnd cell_6t
Xbit_r131_c49 bl[49] br[49] wl[131] vdd gnd cell_6t
Xbit_r132_c49 bl[49] br[49] wl[132] vdd gnd cell_6t
Xbit_r133_c49 bl[49] br[49] wl[133] vdd gnd cell_6t
Xbit_r134_c49 bl[49] br[49] wl[134] vdd gnd cell_6t
Xbit_r135_c49 bl[49] br[49] wl[135] vdd gnd cell_6t
Xbit_r136_c49 bl[49] br[49] wl[136] vdd gnd cell_6t
Xbit_r137_c49 bl[49] br[49] wl[137] vdd gnd cell_6t
Xbit_r138_c49 bl[49] br[49] wl[138] vdd gnd cell_6t
Xbit_r139_c49 bl[49] br[49] wl[139] vdd gnd cell_6t
Xbit_r140_c49 bl[49] br[49] wl[140] vdd gnd cell_6t
Xbit_r141_c49 bl[49] br[49] wl[141] vdd gnd cell_6t
Xbit_r142_c49 bl[49] br[49] wl[142] vdd gnd cell_6t
Xbit_r143_c49 bl[49] br[49] wl[143] vdd gnd cell_6t
Xbit_r144_c49 bl[49] br[49] wl[144] vdd gnd cell_6t
Xbit_r145_c49 bl[49] br[49] wl[145] vdd gnd cell_6t
Xbit_r146_c49 bl[49] br[49] wl[146] vdd gnd cell_6t
Xbit_r147_c49 bl[49] br[49] wl[147] vdd gnd cell_6t
Xbit_r148_c49 bl[49] br[49] wl[148] vdd gnd cell_6t
Xbit_r149_c49 bl[49] br[49] wl[149] vdd gnd cell_6t
Xbit_r150_c49 bl[49] br[49] wl[150] vdd gnd cell_6t
Xbit_r151_c49 bl[49] br[49] wl[151] vdd gnd cell_6t
Xbit_r152_c49 bl[49] br[49] wl[152] vdd gnd cell_6t
Xbit_r153_c49 bl[49] br[49] wl[153] vdd gnd cell_6t
Xbit_r154_c49 bl[49] br[49] wl[154] vdd gnd cell_6t
Xbit_r155_c49 bl[49] br[49] wl[155] vdd gnd cell_6t
Xbit_r156_c49 bl[49] br[49] wl[156] vdd gnd cell_6t
Xbit_r157_c49 bl[49] br[49] wl[157] vdd gnd cell_6t
Xbit_r158_c49 bl[49] br[49] wl[158] vdd gnd cell_6t
Xbit_r159_c49 bl[49] br[49] wl[159] vdd gnd cell_6t
Xbit_r160_c49 bl[49] br[49] wl[160] vdd gnd cell_6t
Xbit_r161_c49 bl[49] br[49] wl[161] vdd gnd cell_6t
Xbit_r162_c49 bl[49] br[49] wl[162] vdd gnd cell_6t
Xbit_r163_c49 bl[49] br[49] wl[163] vdd gnd cell_6t
Xbit_r164_c49 bl[49] br[49] wl[164] vdd gnd cell_6t
Xbit_r165_c49 bl[49] br[49] wl[165] vdd gnd cell_6t
Xbit_r166_c49 bl[49] br[49] wl[166] vdd gnd cell_6t
Xbit_r167_c49 bl[49] br[49] wl[167] vdd gnd cell_6t
Xbit_r168_c49 bl[49] br[49] wl[168] vdd gnd cell_6t
Xbit_r169_c49 bl[49] br[49] wl[169] vdd gnd cell_6t
Xbit_r170_c49 bl[49] br[49] wl[170] vdd gnd cell_6t
Xbit_r171_c49 bl[49] br[49] wl[171] vdd gnd cell_6t
Xbit_r172_c49 bl[49] br[49] wl[172] vdd gnd cell_6t
Xbit_r173_c49 bl[49] br[49] wl[173] vdd gnd cell_6t
Xbit_r174_c49 bl[49] br[49] wl[174] vdd gnd cell_6t
Xbit_r175_c49 bl[49] br[49] wl[175] vdd gnd cell_6t
Xbit_r176_c49 bl[49] br[49] wl[176] vdd gnd cell_6t
Xbit_r177_c49 bl[49] br[49] wl[177] vdd gnd cell_6t
Xbit_r178_c49 bl[49] br[49] wl[178] vdd gnd cell_6t
Xbit_r179_c49 bl[49] br[49] wl[179] vdd gnd cell_6t
Xbit_r180_c49 bl[49] br[49] wl[180] vdd gnd cell_6t
Xbit_r181_c49 bl[49] br[49] wl[181] vdd gnd cell_6t
Xbit_r182_c49 bl[49] br[49] wl[182] vdd gnd cell_6t
Xbit_r183_c49 bl[49] br[49] wl[183] vdd gnd cell_6t
Xbit_r184_c49 bl[49] br[49] wl[184] vdd gnd cell_6t
Xbit_r185_c49 bl[49] br[49] wl[185] vdd gnd cell_6t
Xbit_r186_c49 bl[49] br[49] wl[186] vdd gnd cell_6t
Xbit_r187_c49 bl[49] br[49] wl[187] vdd gnd cell_6t
Xbit_r188_c49 bl[49] br[49] wl[188] vdd gnd cell_6t
Xbit_r189_c49 bl[49] br[49] wl[189] vdd gnd cell_6t
Xbit_r190_c49 bl[49] br[49] wl[190] vdd gnd cell_6t
Xbit_r191_c49 bl[49] br[49] wl[191] vdd gnd cell_6t
Xbit_r192_c49 bl[49] br[49] wl[192] vdd gnd cell_6t
Xbit_r193_c49 bl[49] br[49] wl[193] vdd gnd cell_6t
Xbit_r194_c49 bl[49] br[49] wl[194] vdd gnd cell_6t
Xbit_r195_c49 bl[49] br[49] wl[195] vdd gnd cell_6t
Xbit_r196_c49 bl[49] br[49] wl[196] vdd gnd cell_6t
Xbit_r197_c49 bl[49] br[49] wl[197] vdd gnd cell_6t
Xbit_r198_c49 bl[49] br[49] wl[198] vdd gnd cell_6t
Xbit_r199_c49 bl[49] br[49] wl[199] vdd gnd cell_6t
Xbit_r200_c49 bl[49] br[49] wl[200] vdd gnd cell_6t
Xbit_r201_c49 bl[49] br[49] wl[201] vdd gnd cell_6t
Xbit_r202_c49 bl[49] br[49] wl[202] vdd gnd cell_6t
Xbit_r203_c49 bl[49] br[49] wl[203] vdd gnd cell_6t
Xbit_r204_c49 bl[49] br[49] wl[204] vdd gnd cell_6t
Xbit_r205_c49 bl[49] br[49] wl[205] vdd gnd cell_6t
Xbit_r206_c49 bl[49] br[49] wl[206] vdd gnd cell_6t
Xbit_r207_c49 bl[49] br[49] wl[207] vdd gnd cell_6t
Xbit_r208_c49 bl[49] br[49] wl[208] vdd gnd cell_6t
Xbit_r209_c49 bl[49] br[49] wl[209] vdd gnd cell_6t
Xbit_r210_c49 bl[49] br[49] wl[210] vdd gnd cell_6t
Xbit_r211_c49 bl[49] br[49] wl[211] vdd gnd cell_6t
Xbit_r212_c49 bl[49] br[49] wl[212] vdd gnd cell_6t
Xbit_r213_c49 bl[49] br[49] wl[213] vdd gnd cell_6t
Xbit_r214_c49 bl[49] br[49] wl[214] vdd gnd cell_6t
Xbit_r215_c49 bl[49] br[49] wl[215] vdd gnd cell_6t
Xbit_r216_c49 bl[49] br[49] wl[216] vdd gnd cell_6t
Xbit_r217_c49 bl[49] br[49] wl[217] vdd gnd cell_6t
Xbit_r218_c49 bl[49] br[49] wl[218] vdd gnd cell_6t
Xbit_r219_c49 bl[49] br[49] wl[219] vdd gnd cell_6t
Xbit_r220_c49 bl[49] br[49] wl[220] vdd gnd cell_6t
Xbit_r221_c49 bl[49] br[49] wl[221] vdd gnd cell_6t
Xbit_r222_c49 bl[49] br[49] wl[222] vdd gnd cell_6t
Xbit_r223_c49 bl[49] br[49] wl[223] vdd gnd cell_6t
Xbit_r224_c49 bl[49] br[49] wl[224] vdd gnd cell_6t
Xbit_r225_c49 bl[49] br[49] wl[225] vdd gnd cell_6t
Xbit_r226_c49 bl[49] br[49] wl[226] vdd gnd cell_6t
Xbit_r227_c49 bl[49] br[49] wl[227] vdd gnd cell_6t
Xbit_r228_c49 bl[49] br[49] wl[228] vdd gnd cell_6t
Xbit_r229_c49 bl[49] br[49] wl[229] vdd gnd cell_6t
Xbit_r230_c49 bl[49] br[49] wl[230] vdd gnd cell_6t
Xbit_r231_c49 bl[49] br[49] wl[231] vdd gnd cell_6t
Xbit_r232_c49 bl[49] br[49] wl[232] vdd gnd cell_6t
Xbit_r233_c49 bl[49] br[49] wl[233] vdd gnd cell_6t
Xbit_r234_c49 bl[49] br[49] wl[234] vdd gnd cell_6t
Xbit_r235_c49 bl[49] br[49] wl[235] vdd gnd cell_6t
Xbit_r236_c49 bl[49] br[49] wl[236] vdd gnd cell_6t
Xbit_r237_c49 bl[49] br[49] wl[237] vdd gnd cell_6t
Xbit_r238_c49 bl[49] br[49] wl[238] vdd gnd cell_6t
Xbit_r239_c49 bl[49] br[49] wl[239] vdd gnd cell_6t
Xbit_r240_c49 bl[49] br[49] wl[240] vdd gnd cell_6t
Xbit_r241_c49 bl[49] br[49] wl[241] vdd gnd cell_6t
Xbit_r242_c49 bl[49] br[49] wl[242] vdd gnd cell_6t
Xbit_r243_c49 bl[49] br[49] wl[243] vdd gnd cell_6t
Xbit_r244_c49 bl[49] br[49] wl[244] vdd gnd cell_6t
Xbit_r245_c49 bl[49] br[49] wl[245] vdd gnd cell_6t
Xbit_r246_c49 bl[49] br[49] wl[246] vdd gnd cell_6t
Xbit_r247_c49 bl[49] br[49] wl[247] vdd gnd cell_6t
Xbit_r248_c49 bl[49] br[49] wl[248] vdd gnd cell_6t
Xbit_r249_c49 bl[49] br[49] wl[249] vdd gnd cell_6t
Xbit_r250_c49 bl[49] br[49] wl[250] vdd gnd cell_6t
Xbit_r251_c49 bl[49] br[49] wl[251] vdd gnd cell_6t
Xbit_r252_c49 bl[49] br[49] wl[252] vdd gnd cell_6t
Xbit_r253_c49 bl[49] br[49] wl[253] vdd gnd cell_6t
Xbit_r254_c49 bl[49] br[49] wl[254] vdd gnd cell_6t
Xbit_r255_c49 bl[49] br[49] wl[255] vdd gnd cell_6t
Xbit_r0_c50 bl[50] br[50] wl[0] vdd gnd cell_6t
Xbit_r1_c50 bl[50] br[50] wl[1] vdd gnd cell_6t
Xbit_r2_c50 bl[50] br[50] wl[2] vdd gnd cell_6t
Xbit_r3_c50 bl[50] br[50] wl[3] vdd gnd cell_6t
Xbit_r4_c50 bl[50] br[50] wl[4] vdd gnd cell_6t
Xbit_r5_c50 bl[50] br[50] wl[5] vdd gnd cell_6t
Xbit_r6_c50 bl[50] br[50] wl[6] vdd gnd cell_6t
Xbit_r7_c50 bl[50] br[50] wl[7] vdd gnd cell_6t
Xbit_r8_c50 bl[50] br[50] wl[8] vdd gnd cell_6t
Xbit_r9_c50 bl[50] br[50] wl[9] vdd gnd cell_6t
Xbit_r10_c50 bl[50] br[50] wl[10] vdd gnd cell_6t
Xbit_r11_c50 bl[50] br[50] wl[11] vdd gnd cell_6t
Xbit_r12_c50 bl[50] br[50] wl[12] vdd gnd cell_6t
Xbit_r13_c50 bl[50] br[50] wl[13] vdd gnd cell_6t
Xbit_r14_c50 bl[50] br[50] wl[14] vdd gnd cell_6t
Xbit_r15_c50 bl[50] br[50] wl[15] vdd gnd cell_6t
Xbit_r16_c50 bl[50] br[50] wl[16] vdd gnd cell_6t
Xbit_r17_c50 bl[50] br[50] wl[17] vdd gnd cell_6t
Xbit_r18_c50 bl[50] br[50] wl[18] vdd gnd cell_6t
Xbit_r19_c50 bl[50] br[50] wl[19] vdd gnd cell_6t
Xbit_r20_c50 bl[50] br[50] wl[20] vdd gnd cell_6t
Xbit_r21_c50 bl[50] br[50] wl[21] vdd gnd cell_6t
Xbit_r22_c50 bl[50] br[50] wl[22] vdd gnd cell_6t
Xbit_r23_c50 bl[50] br[50] wl[23] vdd gnd cell_6t
Xbit_r24_c50 bl[50] br[50] wl[24] vdd gnd cell_6t
Xbit_r25_c50 bl[50] br[50] wl[25] vdd gnd cell_6t
Xbit_r26_c50 bl[50] br[50] wl[26] vdd gnd cell_6t
Xbit_r27_c50 bl[50] br[50] wl[27] vdd gnd cell_6t
Xbit_r28_c50 bl[50] br[50] wl[28] vdd gnd cell_6t
Xbit_r29_c50 bl[50] br[50] wl[29] vdd gnd cell_6t
Xbit_r30_c50 bl[50] br[50] wl[30] vdd gnd cell_6t
Xbit_r31_c50 bl[50] br[50] wl[31] vdd gnd cell_6t
Xbit_r32_c50 bl[50] br[50] wl[32] vdd gnd cell_6t
Xbit_r33_c50 bl[50] br[50] wl[33] vdd gnd cell_6t
Xbit_r34_c50 bl[50] br[50] wl[34] vdd gnd cell_6t
Xbit_r35_c50 bl[50] br[50] wl[35] vdd gnd cell_6t
Xbit_r36_c50 bl[50] br[50] wl[36] vdd gnd cell_6t
Xbit_r37_c50 bl[50] br[50] wl[37] vdd gnd cell_6t
Xbit_r38_c50 bl[50] br[50] wl[38] vdd gnd cell_6t
Xbit_r39_c50 bl[50] br[50] wl[39] vdd gnd cell_6t
Xbit_r40_c50 bl[50] br[50] wl[40] vdd gnd cell_6t
Xbit_r41_c50 bl[50] br[50] wl[41] vdd gnd cell_6t
Xbit_r42_c50 bl[50] br[50] wl[42] vdd gnd cell_6t
Xbit_r43_c50 bl[50] br[50] wl[43] vdd gnd cell_6t
Xbit_r44_c50 bl[50] br[50] wl[44] vdd gnd cell_6t
Xbit_r45_c50 bl[50] br[50] wl[45] vdd gnd cell_6t
Xbit_r46_c50 bl[50] br[50] wl[46] vdd gnd cell_6t
Xbit_r47_c50 bl[50] br[50] wl[47] vdd gnd cell_6t
Xbit_r48_c50 bl[50] br[50] wl[48] vdd gnd cell_6t
Xbit_r49_c50 bl[50] br[50] wl[49] vdd gnd cell_6t
Xbit_r50_c50 bl[50] br[50] wl[50] vdd gnd cell_6t
Xbit_r51_c50 bl[50] br[50] wl[51] vdd gnd cell_6t
Xbit_r52_c50 bl[50] br[50] wl[52] vdd gnd cell_6t
Xbit_r53_c50 bl[50] br[50] wl[53] vdd gnd cell_6t
Xbit_r54_c50 bl[50] br[50] wl[54] vdd gnd cell_6t
Xbit_r55_c50 bl[50] br[50] wl[55] vdd gnd cell_6t
Xbit_r56_c50 bl[50] br[50] wl[56] vdd gnd cell_6t
Xbit_r57_c50 bl[50] br[50] wl[57] vdd gnd cell_6t
Xbit_r58_c50 bl[50] br[50] wl[58] vdd gnd cell_6t
Xbit_r59_c50 bl[50] br[50] wl[59] vdd gnd cell_6t
Xbit_r60_c50 bl[50] br[50] wl[60] vdd gnd cell_6t
Xbit_r61_c50 bl[50] br[50] wl[61] vdd gnd cell_6t
Xbit_r62_c50 bl[50] br[50] wl[62] vdd gnd cell_6t
Xbit_r63_c50 bl[50] br[50] wl[63] vdd gnd cell_6t
Xbit_r64_c50 bl[50] br[50] wl[64] vdd gnd cell_6t
Xbit_r65_c50 bl[50] br[50] wl[65] vdd gnd cell_6t
Xbit_r66_c50 bl[50] br[50] wl[66] vdd gnd cell_6t
Xbit_r67_c50 bl[50] br[50] wl[67] vdd gnd cell_6t
Xbit_r68_c50 bl[50] br[50] wl[68] vdd gnd cell_6t
Xbit_r69_c50 bl[50] br[50] wl[69] vdd gnd cell_6t
Xbit_r70_c50 bl[50] br[50] wl[70] vdd gnd cell_6t
Xbit_r71_c50 bl[50] br[50] wl[71] vdd gnd cell_6t
Xbit_r72_c50 bl[50] br[50] wl[72] vdd gnd cell_6t
Xbit_r73_c50 bl[50] br[50] wl[73] vdd gnd cell_6t
Xbit_r74_c50 bl[50] br[50] wl[74] vdd gnd cell_6t
Xbit_r75_c50 bl[50] br[50] wl[75] vdd gnd cell_6t
Xbit_r76_c50 bl[50] br[50] wl[76] vdd gnd cell_6t
Xbit_r77_c50 bl[50] br[50] wl[77] vdd gnd cell_6t
Xbit_r78_c50 bl[50] br[50] wl[78] vdd gnd cell_6t
Xbit_r79_c50 bl[50] br[50] wl[79] vdd gnd cell_6t
Xbit_r80_c50 bl[50] br[50] wl[80] vdd gnd cell_6t
Xbit_r81_c50 bl[50] br[50] wl[81] vdd gnd cell_6t
Xbit_r82_c50 bl[50] br[50] wl[82] vdd gnd cell_6t
Xbit_r83_c50 bl[50] br[50] wl[83] vdd gnd cell_6t
Xbit_r84_c50 bl[50] br[50] wl[84] vdd gnd cell_6t
Xbit_r85_c50 bl[50] br[50] wl[85] vdd gnd cell_6t
Xbit_r86_c50 bl[50] br[50] wl[86] vdd gnd cell_6t
Xbit_r87_c50 bl[50] br[50] wl[87] vdd gnd cell_6t
Xbit_r88_c50 bl[50] br[50] wl[88] vdd gnd cell_6t
Xbit_r89_c50 bl[50] br[50] wl[89] vdd gnd cell_6t
Xbit_r90_c50 bl[50] br[50] wl[90] vdd gnd cell_6t
Xbit_r91_c50 bl[50] br[50] wl[91] vdd gnd cell_6t
Xbit_r92_c50 bl[50] br[50] wl[92] vdd gnd cell_6t
Xbit_r93_c50 bl[50] br[50] wl[93] vdd gnd cell_6t
Xbit_r94_c50 bl[50] br[50] wl[94] vdd gnd cell_6t
Xbit_r95_c50 bl[50] br[50] wl[95] vdd gnd cell_6t
Xbit_r96_c50 bl[50] br[50] wl[96] vdd gnd cell_6t
Xbit_r97_c50 bl[50] br[50] wl[97] vdd gnd cell_6t
Xbit_r98_c50 bl[50] br[50] wl[98] vdd gnd cell_6t
Xbit_r99_c50 bl[50] br[50] wl[99] vdd gnd cell_6t
Xbit_r100_c50 bl[50] br[50] wl[100] vdd gnd cell_6t
Xbit_r101_c50 bl[50] br[50] wl[101] vdd gnd cell_6t
Xbit_r102_c50 bl[50] br[50] wl[102] vdd gnd cell_6t
Xbit_r103_c50 bl[50] br[50] wl[103] vdd gnd cell_6t
Xbit_r104_c50 bl[50] br[50] wl[104] vdd gnd cell_6t
Xbit_r105_c50 bl[50] br[50] wl[105] vdd gnd cell_6t
Xbit_r106_c50 bl[50] br[50] wl[106] vdd gnd cell_6t
Xbit_r107_c50 bl[50] br[50] wl[107] vdd gnd cell_6t
Xbit_r108_c50 bl[50] br[50] wl[108] vdd gnd cell_6t
Xbit_r109_c50 bl[50] br[50] wl[109] vdd gnd cell_6t
Xbit_r110_c50 bl[50] br[50] wl[110] vdd gnd cell_6t
Xbit_r111_c50 bl[50] br[50] wl[111] vdd gnd cell_6t
Xbit_r112_c50 bl[50] br[50] wl[112] vdd gnd cell_6t
Xbit_r113_c50 bl[50] br[50] wl[113] vdd gnd cell_6t
Xbit_r114_c50 bl[50] br[50] wl[114] vdd gnd cell_6t
Xbit_r115_c50 bl[50] br[50] wl[115] vdd gnd cell_6t
Xbit_r116_c50 bl[50] br[50] wl[116] vdd gnd cell_6t
Xbit_r117_c50 bl[50] br[50] wl[117] vdd gnd cell_6t
Xbit_r118_c50 bl[50] br[50] wl[118] vdd gnd cell_6t
Xbit_r119_c50 bl[50] br[50] wl[119] vdd gnd cell_6t
Xbit_r120_c50 bl[50] br[50] wl[120] vdd gnd cell_6t
Xbit_r121_c50 bl[50] br[50] wl[121] vdd gnd cell_6t
Xbit_r122_c50 bl[50] br[50] wl[122] vdd gnd cell_6t
Xbit_r123_c50 bl[50] br[50] wl[123] vdd gnd cell_6t
Xbit_r124_c50 bl[50] br[50] wl[124] vdd gnd cell_6t
Xbit_r125_c50 bl[50] br[50] wl[125] vdd gnd cell_6t
Xbit_r126_c50 bl[50] br[50] wl[126] vdd gnd cell_6t
Xbit_r127_c50 bl[50] br[50] wl[127] vdd gnd cell_6t
Xbit_r128_c50 bl[50] br[50] wl[128] vdd gnd cell_6t
Xbit_r129_c50 bl[50] br[50] wl[129] vdd gnd cell_6t
Xbit_r130_c50 bl[50] br[50] wl[130] vdd gnd cell_6t
Xbit_r131_c50 bl[50] br[50] wl[131] vdd gnd cell_6t
Xbit_r132_c50 bl[50] br[50] wl[132] vdd gnd cell_6t
Xbit_r133_c50 bl[50] br[50] wl[133] vdd gnd cell_6t
Xbit_r134_c50 bl[50] br[50] wl[134] vdd gnd cell_6t
Xbit_r135_c50 bl[50] br[50] wl[135] vdd gnd cell_6t
Xbit_r136_c50 bl[50] br[50] wl[136] vdd gnd cell_6t
Xbit_r137_c50 bl[50] br[50] wl[137] vdd gnd cell_6t
Xbit_r138_c50 bl[50] br[50] wl[138] vdd gnd cell_6t
Xbit_r139_c50 bl[50] br[50] wl[139] vdd gnd cell_6t
Xbit_r140_c50 bl[50] br[50] wl[140] vdd gnd cell_6t
Xbit_r141_c50 bl[50] br[50] wl[141] vdd gnd cell_6t
Xbit_r142_c50 bl[50] br[50] wl[142] vdd gnd cell_6t
Xbit_r143_c50 bl[50] br[50] wl[143] vdd gnd cell_6t
Xbit_r144_c50 bl[50] br[50] wl[144] vdd gnd cell_6t
Xbit_r145_c50 bl[50] br[50] wl[145] vdd gnd cell_6t
Xbit_r146_c50 bl[50] br[50] wl[146] vdd gnd cell_6t
Xbit_r147_c50 bl[50] br[50] wl[147] vdd gnd cell_6t
Xbit_r148_c50 bl[50] br[50] wl[148] vdd gnd cell_6t
Xbit_r149_c50 bl[50] br[50] wl[149] vdd gnd cell_6t
Xbit_r150_c50 bl[50] br[50] wl[150] vdd gnd cell_6t
Xbit_r151_c50 bl[50] br[50] wl[151] vdd gnd cell_6t
Xbit_r152_c50 bl[50] br[50] wl[152] vdd gnd cell_6t
Xbit_r153_c50 bl[50] br[50] wl[153] vdd gnd cell_6t
Xbit_r154_c50 bl[50] br[50] wl[154] vdd gnd cell_6t
Xbit_r155_c50 bl[50] br[50] wl[155] vdd gnd cell_6t
Xbit_r156_c50 bl[50] br[50] wl[156] vdd gnd cell_6t
Xbit_r157_c50 bl[50] br[50] wl[157] vdd gnd cell_6t
Xbit_r158_c50 bl[50] br[50] wl[158] vdd gnd cell_6t
Xbit_r159_c50 bl[50] br[50] wl[159] vdd gnd cell_6t
Xbit_r160_c50 bl[50] br[50] wl[160] vdd gnd cell_6t
Xbit_r161_c50 bl[50] br[50] wl[161] vdd gnd cell_6t
Xbit_r162_c50 bl[50] br[50] wl[162] vdd gnd cell_6t
Xbit_r163_c50 bl[50] br[50] wl[163] vdd gnd cell_6t
Xbit_r164_c50 bl[50] br[50] wl[164] vdd gnd cell_6t
Xbit_r165_c50 bl[50] br[50] wl[165] vdd gnd cell_6t
Xbit_r166_c50 bl[50] br[50] wl[166] vdd gnd cell_6t
Xbit_r167_c50 bl[50] br[50] wl[167] vdd gnd cell_6t
Xbit_r168_c50 bl[50] br[50] wl[168] vdd gnd cell_6t
Xbit_r169_c50 bl[50] br[50] wl[169] vdd gnd cell_6t
Xbit_r170_c50 bl[50] br[50] wl[170] vdd gnd cell_6t
Xbit_r171_c50 bl[50] br[50] wl[171] vdd gnd cell_6t
Xbit_r172_c50 bl[50] br[50] wl[172] vdd gnd cell_6t
Xbit_r173_c50 bl[50] br[50] wl[173] vdd gnd cell_6t
Xbit_r174_c50 bl[50] br[50] wl[174] vdd gnd cell_6t
Xbit_r175_c50 bl[50] br[50] wl[175] vdd gnd cell_6t
Xbit_r176_c50 bl[50] br[50] wl[176] vdd gnd cell_6t
Xbit_r177_c50 bl[50] br[50] wl[177] vdd gnd cell_6t
Xbit_r178_c50 bl[50] br[50] wl[178] vdd gnd cell_6t
Xbit_r179_c50 bl[50] br[50] wl[179] vdd gnd cell_6t
Xbit_r180_c50 bl[50] br[50] wl[180] vdd gnd cell_6t
Xbit_r181_c50 bl[50] br[50] wl[181] vdd gnd cell_6t
Xbit_r182_c50 bl[50] br[50] wl[182] vdd gnd cell_6t
Xbit_r183_c50 bl[50] br[50] wl[183] vdd gnd cell_6t
Xbit_r184_c50 bl[50] br[50] wl[184] vdd gnd cell_6t
Xbit_r185_c50 bl[50] br[50] wl[185] vdd gnd cell_6t
Xbit_r186_c50 bl[50] br[50] wl[186] vdd gnd cell_6t
Xbit_r187_c50 bl[50] br[50] wl[187] vdd gnd cell_6t
Xbit_r188_c50 bl[50] br[50] wl[188] vdd gnd cell_6t
Xbit_r189_c50 bl[50] br[50] wl[189] vdd gnd cell_6t
Xbit_r190_c50 bl[50] br[50] wl[190] vdd gnd cell_6t
Xbit_r191_c50 bl[50] br[50] wl[191] vdd gnd cell_6t
Xbit_r192_c50 bl[50] br[50] wl[192] vdd gnd cell_6t
Xbit_r193_c50 bl[50] br[50] wl[193] vdd gnd cell_6t
Xbit_r194_c50 bl[50] br[50] wl[194] vdd gnd cell_6t
Xbit_r195_c50 bl[50] br[50] wl[195] vdd gnd cell_6t
Xbit_r196_c50 bl[50] br[50] wl[196] vdd gnd cell_6t
Xbit_r197_c50 bl[50] br[50] wl[197] vdd gnd cell_6t
Xbit_r198_c50 bl[50] br[50] wl[198] vdd gnd cell_6t
Xbit_r199_c50 bl[50] br[50] wl[199] vdd gnd cell_6t
Xbit_r200_c50 bl[50] br[50] wl[200] vdd gnd cell_6t
Xbit_r201_c50 bl[50] br[50] wl[201] vdd gnd cell_6t
Xbit_r202_c50 bl[50] br[50] wl[202] vdd gnd cell_6t
Xbit_r203_c50 bl[50] br[50] wl[203] vdd gnd cell_6t
Xbit_r204_c50 bl[50] br[50] wl[204] vdd gnd cell_6t
Xbit_r205_c50 bl[50] br[50] wl[205] vdd gnd cell_6t
Xbit_r206_c50 bl[50] br[50] wl[206] vdd gnd cell_6t
Xbit_r207_c50 bl[50] br[50] wl[207] vdd gnd cell_6t
Xbit_r208_c50 bl[50] br[50] wl[208] vdd gnd cell_6t
Xbit_r209_c50 bl[50] br[50] wl[209] vdd gnd cell_6t
Xbit_r210_c50 bl[50] br[50] wl[210] vdd gnd cell_6t
Xbit_r211_c50 bl[50] br[50] wl[211] vdd gnd cell_6t
Xbit_r212_c50 bl[50] br[50] wl[212] vdd gnd cell_6t
Xbit_r213_c50 bl[50] br[50] wl[213] vdd gnd cell_6t
Xbit_r214_c50 bl[50] br[50] wl[214] vdd gnd cell_6t
Xbit_r215_c50 bl[50] br[50] wl[215] vdd gnd cell_6t
Xbit_r216_c50 bl[50] br[50] wl[216] vdd gnd cell_6t
Xbit_r217_c50 bl[50] br[50] wl[217] vdd gnd cell_6t
Xbit_r218_c50 bl[50] br[50] wl[218] vdd gnd cell_6t
Xbit_r219_c50 bl[50] br[50] wl[219] vdd gnd cell_6t
Xbit_r220_c50 bl[50] br[50] wl[220] vdd gnd cell_6t
Xbit_r221_c50 bl[50] br[50] wl[221] vdd gnd cell_6t
Xbit_r222_c50 bl[50] br[50] wl[222] vdd gnd cell_6t
Xbit_r223_c50 bl[50] br[50] wl[223] vdd gnd cell_6t
Xbit_r224_c50 bl[50] br[50] wl[224] vdd gnd cell_6t
Xbit_r225_c50 bl[50] br[50] wl[225] vdd gnd cell_6t
Xbit_r226_c50 bl[50] br[50] wl[226] vdd gnd cell_6t
Xbit_r227_c50 bl[50] br[50] wl[227] vdd gnd cell_6t
Xbit_r228_c50 bl[50] br[50] wl[228] vdd gnd cell_6t
Xbit_r229_c50 bl[50] br[50] wl[229] vdd gnd cell_6t
Xbit_r230_c50 bl[50] br[50] wl[230] vdd gnd cell_6t
Xbit_r231_c50 bl[50] br[50] wl[231] vdd gnd cell_6t
Xbit_r232_c50 bl[50] br[50] wl[232] vdd gnd cell_6t
Xbit_r233_c50 bl[50] br[50] wl[233] vdd gnd cell_6t
Xbit_r234_c50 bl[50] br[50] wl[234] vdd gnd cell_6t
Xbit_r235_c50 bl[50] br[50] wl[235] vdd gnd cell_6t
Xbit_r236_c50 bl[50] br[50] wl[236] vdd gnd cell_6t
Xbit_r237_c50 bl[50] br[50] wl[237] vdd gnd cell_6t
Xbit_r238_c50 bl[50] br[50] wl[238] vdd gnd cell_6t
Xbit_r239_c50 bl[50] br[50] wl[239] vdd gnd cell_6t
Xbit_r240_c50 bl[50] br[50] wl[240] vdd gnd cell_6t
Xbit_r241_c50 bl[50] br[50] wl[241] vdd gnd cell_6t
Xbit_r242_c50 bl[50] br[50] wl[242] vdd gnd cell_6t
Xbit_r243_c50 bl[50] br[50] wl[243] vdd gnd cell_6t
Xbit_r244_c50 bl[50] br[50] wl[244] vdd gnd cell_6t
Xbit_r245_c50 bl[50] br[50] wl[245] vdd gnd cell_6t
Xbit_r246_c50 bl[50] br[50] wl[246] vdd gnd cell_6t
Xbit_r247_c50 bl[50] br[50] wl[247] vdd gnd cell_6t
Xbit_r248_c50 bl[50] br[50] wl[248] vdd gnd cell_6t
Xbit_r249_c50 bl[50] br[50] wl[249] vdd gnd cell_6t
Xbit_r250_c50 bl[50] br[50] wl[250] vdd gnd cell_6t
Xbit_r251_c50 bl[50] br[50] wl[251] vdd gnd cell_6t
Xbit_r252_c50 bl[50] br[50] wl[252] vdd gnd cell_6t
Xbit_r253_c50 bl[50] br[50] wl[253] vdd gnd cell_6t
Xbit_r254_c50 bl[50] br[50] wl[254] vdd gnd cell_6t
Xbit_r255_c50 bl[50] br[50] wl[255] vdd gnd cell_6t
Xbit_r0_c51 bl[51] br[51] wl[0] vdd gnd cell_6t
Xbit_r1_c51 bl[51] br[51] wl[1] vdd gnd cell_6t
Xbit_r2_c51 bl[51] br[51] wl[2] vdd gnd cell_6t
Xbit_r3_c51 bl[51] br[51] wl[3] vdd gnd cell_6t
Xbit_r4_c51 bl[51] br[51] wl[4] vdd gnd cell_6t
Xbit_r5_c51 bl[51] br[51] wl[5] vdd gnd cell_6t
Xbit_r6_c51 bl[51] br[51] wl[6] vdd gnd cell_6t
Xbit_r7_c51 bl[51] br[51] wl[7] vdd gnd cell_6t
Xbit_r8_c51 bl[51] br[51] wl[8] vdd gnd cell_6t
Xbit_r9_c51 bl[51] br[51] wl[9] vdd gnd cell_6t
Xbit_r10_c51 bl[51] br[51] wl[10] vdd gnd cell_6t
Xbit_r11_c51 bl[51] br[51] wl[11] vdd gnd cell_6t
Xbit_r12_c51 bl[51] br[51] wl[12] vdd gnd cell_6t
Xbit_r13_c51 bl[51] br[51] wl[13] vdd gnd cell_6t
Xbit_r14_c51 bl[51] br[51] wl[14] vdd gnd cell_6t
Xbit_r15_c51 bl[51] br[51] wl[15] vdd gnd cell_6t
Xbit_r16_c51 bl[51] br[51] wl[16] vdd gnd cell_6t
Xbit_r17_c51 bl[51] br[51] wl[17] vdd gnd cell_6t
Xbit_r18_c51 bl[51] br[51] wl[18] vdd gnd cell_6t
Xbit_r19_c51 bl[51] br[51] wl[19] vdd gnd cell_6t
Xbit_r20_c51 bl[51] br[51] wl[20] vdd gnd cell_6t
Xbit_r21_c51 bl[51] br[51] wl[21] vdd gnd cell_6t
Xbit_r22_c51 bl[51] br[51] wl[22] vdd gnd cell_6t
Xbit_r23_c51 bl[51] br[51] wl[23] vdd gnd cell_6t
Xbit_r24_c51 bl[51] br[51] wl[24] vdd gnd cell_6t
Xbit_r25_c51 bl[51] br[51] wl[25] vdd gnd cell_6t
Xbit_r26_c51 bl[51] br[51] wl[26] vdd gnd cell_6t
Xbit_r27_c51 bl[51] br[51] wl[27] vdd gnd cell_6t
Xbit_r28_c51 bl[51] br[51] wl[28] vdd gnd cell_6t
Xbit_r29_c51 bl[51] br[51] wl[29] vdd gnd cell_6t
Xbit_r30_c51 bl[51] br[51] wl[30] vdd gnd cell_6t
Xbit_r31_c51 bl[51] br[51] wl[31] vdd gnd cell_6t
Xbit_r32_c51 bl[51] br[51] wl[32] vdd gnd cell_6t
Xbit_r33_c51 bl[51] br[51] wl[33] vdd gnd cell_6t
Xbit_r34_c51 bl[51] br[51] wl[34] vdd gnd cell_6t
Xbit_r35_c51 bl[51] br[51] wl[35] vdd gnd cell_6t
Xbit_r36_c51 bl[51] br[51] wl[36] vdd gnd cell_6t
Xbit_r37_c51 bl[51] br[51] wl[37] vdd gnd cell_6t
Xbit_r38_c51 bl[51] br[51] wl[38] vdd gnd cell_6t
Xbit_r39_c51 bl[51] br[51] wl[39] vdd gnd cell_6t
Xbit_r40_c51 bl[51] br[51] wl[40] vdd gnd cell_6t
Xbit_r41_c51 bl[51] br[51] wl[41] vdd gnd cell_6t
Xbit_r42_c51 bl[51] br[51] wl[42] vdd gnd cell_6t
Xbit_r43_c51 bl[51] br[51] wl[43] vdd gnd cell_6t
Xbit_r44_c51 bl[51] br[51] wl[44] vdd gnd cell_6t
Xbit_r45_c51 bl[51] br[51] wl[45] vdd gnd cell_6t
Xbit_r46_c51 bl[51] br[51] wl[46] vdd gnd cell_6t
Xbit_r47_c51 bl[51] br[51] wl[47] vdd gnd cell_6t
Xbit_r48_c51 bl[51] br[51] wl[48] vdd gnd cell_6t
Xbit_r49_c51 bl[51] br[51] wl[49] vdd gnd cell_6t
Xbit_r50_c51 bl[51] br[51] wl[50] vdd gnd cell_6t
Xbit_r51_c51 bl[51] br[51] wl[51] vdd gnd cell_6t
Xbit_r52_c51 bl[51] br[51] wl[52] vdd gnd cell_6t
Xbit_r53_c51 bl[51] br[51] wl[53] vdd gnd cell_6t
Xbit_r54_c51 bl[51] br[51] wl[54] vdd gnd cell_6t
Xbit_r55_c51 bl[51] br[51] wl[55] vdd gnd cell_6t
Xbit_r56_c51 bl[51] br[51] wl[56] vdd gnd cell_6t
Xbit_r57_c51 bl[51] br[51] wl[57] vdd gnd cell_6t
Xbit_r58_c51 bl[51] br[51] wl[58] vdd gnd cell_6t
Xbit_r59_c51 bl[51] br[51] wl[59] vdd gnd cell_6t
Xbit_r60_c51 bl[51] br[51] wl[60] vdd gnd cell_6t
Xbit_r61_c51 bl[51] br[51] wl[61] vdd gnd cell_6t
Xbit_r62_c51 bl[51] br[51] wl[62] vdd gnd cell_6t
Xbit_r63_c51 bl[51] br[51] wl[63] vdd gnd cell_6t
Xbit_r64_c51 bl[51] br[51] wl[64] vdd gnd cell_6t
Xbit_r65_c51 bl[51] br[51] wl[65] vdd gnd cell_6t
Xbit_r66_c51 bl[51] br[51] wl[66] vdd gnd cell_6t
Xbit_r67_c51 bl[51] br[51] wl[67] vdd gnd cell_6t
Xbit_r68_c51 bl[51] br[51] wl[68] vdd gnd cell_6t
Xbit_r69_c51 bl[51] br[51] wl[69] vdd gnd cell_6t
Xbit_r70_c51 bl[51] br[51] wl[70] vdd gnd cell_6t
Xbit_r71_c51 bl[51] br[51] wl[71] vdd gnd cell_6t
Xbit_r72_c51 bl[51] br[51] wl[72] vdd gnd cell_6t
Xbit_r73_c51 bl[51] br[51] wl[73] vdd gnd cell_6t
Xbit_r74_c51 bl[51] br[51] wl[74] vdd gnd cell_6t
Xbit_r75_c51 bl[51] br[51] wl[75] vdd gnd cell_6t
Xbit_r76_c51 bl[51] br[51] wl[76] vdd gnd cell_6t
Xbit_r77_c51 bl[51] br[51] wl[77] vdd gnd cell_6t
Xbit_r78_c51 bl[51] br[51] wl[78] vdd gnd cell_6t
Xbit_r79_c51 bl[51] br[51] wl[79] vdd gnd cell_6t
Xbit_r80_c51 bl[51] br[51] wl[80] vdd gnd cell_6t
Xbit_r81_c51 bl[51] br[51] wl[81] vdd gnd cell_6t
Xbit_r82_c51 bl[51] br[51] wl[82] vdd gnd cell_6t
Xbit_r83_c51 bl[51] br[51] wl[83] vdd gnd cell_6t
Xbit_r84_c51 bl[51] br[51] wl[84] vdd gnd cell_6t
Xbit_r85_c51 bl[51] br[51] wl[85] vdd gnd cell_6t
Xbit_r86_c51 bl[51] br[51] wl[86] vdd gnd cell_6t
Xbit_r87_c51 bl[51] br[51] wl[87] vdd gnd cell_6t
Xbit_r88_c51 bl[51] br[51] wl[88] vdd gnd cell_6t
Xbit_r89_c51 bl[51] br[51] wl[89] vdd gnd cell_6t
Xbit_r90_c51 bl[51] br[51] wl[90] vdd gnd cell_6t
Xbit_r91_c51 bl[51] br[51] wl[91] vdd gnd cell_6t
Xbit_r92_c51 bl[51] br[51] wl[92] vdd gnd cell_6t
Xbit_r93_c51 bl[51] br[51] wl[93] vdd gnd cell_6t
Xbit_r94_c51 bl[51] br[51] wl[94] vdd gnd cell_6t
Xbit_r95_c51 bl[51] br[51] wl[95] vdd gnd cell_6t
Xbit_r96_c51 bl[51] br[51] wl[96] vdd gnd cell_6t
Xbit_r97_c51 bl[51] br[51] wl[97] vdd gnd cell_6t
Xbit_r98_c51 bl[51] br[51] wl[98] vdd gnd cell_6t
Xbit_r99_c51 bl[51] br[51] wl[99] vdd gnd cell_6t
Xbit_r100_c51 bl[51] br[51] wl[100] vdd gnd cell_6t
Xbit_r101_c51 bl[51] br[51] wl[101] vdd gnd cell_6t
Xbit_r102_c51 bl[51] br[51] wl[102] vdd gnd cell_6t
Xbit_r103_c51 bl[51] br[51] wl[103] vdd gnd cell_6t
Xbit_r104_c51 bl[51] br[51] wl[104] vdd gnd cell_6t
Xbit_r105_c51 bl[51] br[51] wl[105] vdd gnd cell_6t
Xbit_r106_c51 bl[51] br[51] wl[106] vdd gnd cell_6t
Xbit_r107_c51 bl[51] br[51] wl[107] vdd gnd cell_6t
Xbit_r108_c51 bl[51] br[51] wl[108] vdd gnd cell_6t
Xbit_r109_c51 bl[51] br[51] wl[109] vdd gnd cell_6t
Xbit_r110_c51 bl[51] br[51] wl[110] vdd gnd cell_6t
Xbit_r111_c51 bl[51] br[51] wl[111] vdd gnd cell_6t
Xbit_r112_c51 bl[51] br[51] wl[112] vdd gnd cell_6t
Xbit_r113_c51 bl[51] br[51] wl[113] vdd gnd cell_6t
Xbit_r114_c51 bl[51] br[51] wl[114] vdd gnd cell_6t
Xbit_r115_c51 bl[51] br[51] wl[115] vdd gnd cell_6t
Xbit_r116_c51 bl[51] br[51] wl[116] vdd gnd cell_6t
Xbit_r117_c51 bl[51] br[51] wl[117] vdd gnd cell_6t
Xbit_r118_c51 bl[51] br[51] wl[118] vdd gnd cell_6t
Xbit_r119_c51 bl[51] br[51] wl[119] vdd gnd cell_6t
Xbit_r120_c51 bl[51] br[51] wl[120] vdd gnd cell_6t
Xbit_r121_c51 bl[51] br[51] wl[121] vdd gnd cell_6t
Xbit_r122_c51 bl[51] br[51] wl[122] vdd gnd cell_6t
Xbit_r123_c51 bl[51] br[51] wl[123] vdd gnd cell_6t
Xbit_r124_c51 bl[51] br[51] wl[124] vdd gnd cell_6t
Xbit_r125_c51 bl[51] br[51] wl[125] vdd gnd cell_6t
Xbit_r126_c51 bl[51] br[51] wl[126] vdd gnd cell_6t
Xbit_r127_c51 bl[51] br[51] wl[127] vdd gnd cell_6t
Xbit_r128_c51 bl[51] br[51] wl[128] vdd gnd cell_6t
Xbit_r129_c51 bl[51] br[51] wl[129] vdd gnd cell_6t
Xbit_r130_c51 bl[51] br[51] wl[130] vdd gnd cell_6t
Xbit_r131_c51 bl[51] br[51] wl[131] vdd gnd cell_6t
Xbit_r132_c51 bl[51] br[51] wl[132] vdd gnd cell_6t
Xbit_r133_c51 bl[51] br[51] wl[133] vdd gnd cell_6t
Xbit_r134_c51 bl[51] br[51] wl[134] vdd gnd cell_6t
Xbit_r135_c51 bl[51] br[51] wl[135] vdd gnd cell_6t
Xbit_r136_c51 bl[51] br[51] wl[136] vdd gnd cell_6t
Xbit_r137_c51 bl[51] br[51] wl[137] vdd gnd cell_6t
Xbit_r138_c51 bl[51] br[51] wl[138] vdd gnd cell_6t
Xbit_r139_c51 bl[51] br[51] wl[139] vdd gnd cell_6t
Xbit_r140_c51 bl[51] br[51] wl[140] vdd gnd cell_6t
Xbit_r141_c51 bl[51] br[51] wl[141] vdd gnd cell_6t
Xbit_r142_c51 bl[51] br[51] wl[142] vdd gnd cell_6t
Xbit_r143_c51 bl[51] br[51] wl[143] vdd gnd cell_6t
Xbit_r144_c51 bl[51] br[51] wl[144] vdd gnd cell_6t
Xbit_r145_c51 bl[51] br[51] wl[145] vdd gnd cell_6t
Xbit_r146_c51 bl[51] br[51] wl[146] vdd gnd cell_6t
Xbit_r147_c51 bl[51] br[51] wl[147] vdd gnd cell_6t
Xbit_r148_c51 bl[51] br[51] wl[148] vdd gnd cell_6t
Xbit_r149_c51 bl[51] br[51] wl[149] vdd gnd cell_6t
Xbit_r150_c51 bl[51] br[51] wl[150] vdd gnd cell_6t
Xbit_r151_c51 bl[51] br[51] wl[151] vdd gnd cell_6t
Xbit_r152_c51 bl[51] br[51] wl[152] vdd gnd cell_6t
Xbit_r153_c51 bl[51] br[51] wl[153] vdd gnd cell_6t
Xbit_r154_c51 bl[51] br[51] wl[154] vdd gnd cell_6t
Xbit_r155_c51 bl[51] br[51] wl[155] vdd gnd cell_6t
Xbit_r156_c51 bl[51] br[51] wl[156] vdd gnd cell_6t
Xbit_r157_c51 bl[51] br[51] wl[157] vdd gnd cell_6t
Xbit_r158_c51 bl[51] br[51] wl[158] vdd gnd cell_6t
Xbit_r159_c51 bl[51] br[51] wl[159] vdd gnd cell_6t
Xbit_r160_c51 bl[51] br[51] wl[160] vdd gnd cell_6t
Xbit_r161_c51 bl[51] br[51] wl[161] vdd gnd cell_6t
Xbit_r162_c51 bl[51] br[51] wl[162] vdd gnd cell_6t
Xbit_r163_c51 bl[51] br[51] wl[163] vdd gnd cell_6t
Xbit_r164_c51 bl[51] br[51] wl[164] vdd gnd cell_6t
Xbit_r165_c51 bl[51] br[51] wl[165] vdd gnd cell_6t
Xbit_r166_c51 bl[51] br[51] wl[166] vdd gnd cell_6t
Xbit_r167_c51 bl[51] br[51] wl[167] vdd gnd cell_6t
Xbit_r168_c51 bl[51] br[51] wl[168] vdd gnd cell_6t
Xbit_r169_c51 bl[51] br[51] wl[169] vdd gnd cell_6t
Xbit_r170_c51 bl[51] br[51] wl[170] vdd gnd cell_6t
Xbit_r171_c51 bl[51] br[51] wl[171] vdd gnd cell_6t
Xbit_r172_c51 bl[51] br[51] wl[172] vdd gnd cell_6t
Xbit_r173_c51 bl[51] br[51] wl[173] vdd gnd cell_6t
Xbit_r174_c51 bl[51] br[51] wl[174] vdd gnd cell_6t
Xbit_r175_c51 bl[51] br[51] wl[175] vdd gnd cell_6t
Xbit_r176_c51 bl[51] br[51] wl[176] vdd gnd cell_6t
Xbit_r177_c51 bl[51] br[51] wl[177] vdd gnd cell_6t
Xbit_r178_c51 bl[51] br[51] wl[178] vdd gnd cell_6t
Xbit_r179_c51 bl[51] br[51] wl[179] vdd gnd cell_6t
Xbit_r180_c51 bl[51] br[51] wl[180] vdd gnd cell_6t
Xbit_r181_c51 bl[51] br[51] wl[181] vdd gnd cell_6t
Xbit_r182_c51 bl[51] br[51] wl[182] vdd gnd cell_6t
Xbit_r183_c51 bl[51] br[51] wl[183] vdd gnd cell_6t
Xbit_r184_c51 bl[51] br[51] wl[184] vdd gnd cell_6t
Xbit_r185_c51 bl[51] br[51] wl[185] vdd gnd cell_6t
Xbit_r186_c51 bl[51] br[51] wl[186] vdd gnd cell_6t
Xbit_r187_c51 bl[51] br[51] wl[187] vdd gnd cell_6t
Xbit_r188_c51 bl[51] br[51] wl[188] vdd gnd cell_6t
Xbit_r189_c51 bl[51] br[51] wl[189] vdd gnd cell_6t
Xbit_r190_c51 bl[51] br[51] wl[190] vdd gnd cell_6t
Xbit_r191_c51 bl[51] br[51] wl[191] vdd gnd cell_6t
Xbit_r192_c51 bl[51] br[51] wl[192] vdd gnd cell_6t
Xbit_r193_c51 bl[51] br[51] wl[193] vdd gnd cell_6t
Xbit_r194_c51 bl[51] br[51] wl[194] vdd gnd cell_6t
Xbit_r195_c51 bl[51] br[51] wl[195] vdd gnd cell_6t
Xbit_r196_c51 bl[51] br[51] wl[196] vdd gnd cell_6t
Xbit_r197_c51 bl[51] br[51] wl[197] vdd gnd cell_6t
Xbit_r198_c51 bl[51] br[51] wl[198] vdd gnd cell_6t
Xbit_r199_c51 bl[51] br[51] wl[199] vdd gnd cell_6t
Xbit_r200_c51 bl[51] br[51] wl[200] vdd gnd cell_6t
Xbit_r201_c51 bl[51] br[51] wl[201] vdd gnd cell_6t
Xbit_r202_c51 bl[51] br[51] wl[202] vdd gnd cell_6t
Xbit_r203_c51 bl[51] br[51] wl[203] vdd gnd cell_6t
Xbit_r204_c51 bl[51] br[51] wl[204] vdd gnd cell_6t
Xbit_r205_c51 bl[51] br[51] wl[205] vdd gnd cell_6t
Xbit_r206_c51 bl[51] br[51] wl[206] vdd gnd cell_6t
Xbit_r207_c51 bl[51] br[51] wl[207] vdd gnd cell_6t
Xbit_r208_c51 bl[51] br[51] wl[208] vdd gnd cell_6t
Xbit_r209_c51 bl[51] br[51] wl[209] vdd gnd cell_6t
Xbit_r210_c51 bl[51] br[51] wl[210] vdd gnd cell_6t
Xbit_r211_c51 bl[51] br[51] wl[211] vdd gnd cell_6t
Xbit_r212_c51 bl[51] br[51] wl[212] vdd gnd cell_6t
Xbit_r213_c51 bl[51] br[51] wl[213] vdd gnd cell_6t
Xbit_r214_c51 bl[51] br[51] wl[214] vdd gnd cell_6t
Xbit_r215_c51 bl[51] br[51] wl[215] vdd gnd cell_6t
Xbit_r216_c51 bl[51] br[51] wl[216] vdd gnd cell_6t
Xbit_r217_c51 bl[51] br[51] wl[217] vdd gnd cell_6t
Xbit_r218_c51 bl[51] br[51] wl[218] vdd gnd cell_6t
Xbit_r219_c51 bl[51] br[51] wl[219] vdd gnd cell_6t
Xbit_r220_c51 bl[51] br[51] wl[220] vdd gnd cell_6t
Xbit_r221_c51 bl[51] br[51] wl[221] vdd gnd cell_6t
Xbit_r222_c51 bl[51] br[51] wl[222] vdd gnd cell_6t
Xbit_r223_c51 bl[51] br[51] wl[223] vdd gnd cell_6t
Xbit_r224_c51 bl[51] br[51] wl[224] vdd gnd cell_6t
Xbit_r225_c51 bl[51] br[51] wl[225] vdd gnd cell_6t
Xbit_r226_c51 bl[51] br[51] wl[226] vdd gnd cell_6t
Xbit_r227_c51 bl[51] br[51] wl[227] vdd gnd cell_6t
Xbit_r228_c51 bl[51] br[51] wl[228] vdd gnd cell_6t
Xbit_r229_c51 bl[51] br[51] wl[229] vdd gnd cell_6t
Xbit_r230_c51 bl[51] br[51] wl[230] vdd gnd cell_6t
Xbit_r231_c51 bl[51] br[51] wl[231] vdd gnd cell_6t
Xbit_r232_c51 bl[51] br[51] wl[232] vdd gnd cell_6t
Xbit_r233_c51 bl[51] br[51] wl[233] vdd gnd cell_6t
Xbit_r234_c51 bl[51] br[51] wl[234] vdd gnd cell_6t
Xbit_r235_c51 bl[51] br[51] wl[235] vdd gnd cell_6t
Xbit_r236_c51 bl[51] br[51] wl[236] vdd gnd cell_6t
Xbit_r237_c51 bl[51] br[51] wl[237] vdd gnd cell_6t
Xbit_r238_c51 bl[51] br[51] wl[238] vdd gnd cell_6t
Xbit_r239_c51 bl[51] br[51] wl[239] vdd gnd cell_6t
Xbit_r240_c51 bl[51] br[51] wl[240] vdd gnd cell_6t
Xbit_r241_c51 bl[51] br[51] wl[241] vdd gnd cell_6t
Xbit_r242_c51 bl[51] br[51] wl[242] vdd gnd cell_6t
Xbit_r243_c51 bl[51] br[51] wl[243] vdd gnd cell_6t
Xbit_r244_c51 bl[51] br[51] wl[244] vdd gnd cell_6t
Xbit_r245_c51 bl[51] br[51] wl[245] vdd gnd cell_6t
Xbit_r246_c51 bl[51] br[51] wl[246] vdd gnd cell_6t
Xbit_r247_c51 bl[51] br[51] wl[247] vdd gnd cell_6t
Xbit_r248_c51 bl[51] br[51] wl[248] vdd gnd cell_6t
Xbit_r249_c51 bl[51] br[51] wl[249] vdd gnd cell_6t
Xbit_r250_c51 bl[51] br[51] wl[250] vdd gnd cell_6t
Xbit_r251_c51 bl[51] br[51] wl[251] vdd gnd cell_6t
Xbit_r252_c51 bl[51] br[51] wl[252] vdd gnd cell_6t
Xbit_r253_c51 bl[51] br[51] wl[253] vdd gnd cell_6t
Xbit_r254_c51 bl[51] br[51] wl[254] vdd gnd cell_6t
Xbit_r255_c51 bl[51] br[51] wl[255] vdd gnd cell_6t
Xbit_r0_c52 bl[52] br[52] wl[0] vdd gnd cell_6t
Xbit_r1_c52 bl[52] br[52] wl[1] vdd gnd cell_6t
Xbit_r2_c52 bl[52] br[52] wl[2] vdd gnd cell_6t
Xbit_r3_c52 bl[52] br[52] wl[3] vdd gnd cell_6t
Xbit_r4_c52 bl[52] br[52] wl[4] vdd gnd cell_6t
Xbit_r5_c52 bl[52] br[52] wl[5] vdd gnd cell_6t
Xbit_r6_c52 bl[52] br[52] wl[6] vdd gnd cell_6t
Xbit_r7_c52 bl[52] br[52] wl[7] vdd gnd cell_6t
Xbit_r8_c52 bl[52] br[52] wl[8] vdd gnd cell_6t
Xbit_r9_c52 bl[52] br[52] wl[9] vdd gnd cell_6t
Xbit_r10_c52 bl[52] br[52] wl[10] vdd gnd cell_6t
Xbit_r11_c52 bl[52] br[52] wl[11] vdd gnd cell_6t
Xbit_r12_c52 bl[52] br[52] wl[12] vdd gnd cell_6t
Xbit_r13_c52 bl[52] br[52] wl[13] vdd gnd cell_6t
Xbit_r14_c52 bl[52] br[52] wl[14] vdd gnd cell_6t
Xbit_r15_c52 bl[52] br[52] wl[15] vdd gnd cell_6t
Xbit_r16_c52 bl[52] br[52] wl[16] vdd gnd cell_6t
Xbit_r17_c52 bl[52] br[52] wl[17] vdd gnd cell_6t
Xbit_r18_c52 bl[52] br[52] wl[18] vdd gnd cell_6t
Xbit_r19_c52 bl[52] br[52] wl[19] vdd gnd cell_6t
Xbit_r20_c52 bl[52] br[52] wl[20] vdd gnd cell_6t
Xbit_r21_c52 bl[52] br[52] wl[21] vdd gnd cell_6t
Xbit_r22_c52 bl[52] br[52] wl[22] vdd gnd cell_6t
Xbit_r23_c52 bl[52] br[52] wl[23] vdd gnd cell_6t
Xbit_r24_c52 bl[52] br[52] wl[24] vdd gnd cell_6t
Xbit_r25_c52 bl[52] br[52] wl[25] vdd gnd cell_6t
Xbit_r26_c52 bl[52] br[52] wl[26] vdd gnd cell_6t
Xbit_r27_c52 bl[52] br[52] wl[27] vdd gnd cell_6t
Xbit_r28_c52 bl[52] br[52] wl[28] vdd gnd cell_6t
Xbit_r29_c52 bl[52] br[52] wl[29] vdd gnd cell_6t
Xbit_r30_c52 bl[52] br[52] wl[30] vdd gnd cell_6t
Xbit_r31_c52 bl[52] br[52] wl[31] vdd gnd cell_6t
Xbit_r32_c52 bl[52] br[52] wl[32] vdd gnd cell_6t
Xbit_r33_c52 bl[52] br[52] wl[33] vdd gnd cell_6t
Xbit_r34_c52 bl[52] br[52] wl[34] vdd gnd cell_6t
Xbit_r35_c52 bl[52] br[52] wl[35] vdd gnd cell_6t
Xbit_r36_c52 bl[52] br[52] wl[36] vdd gnd cell_6t
Xbit_r37_c52 bl[52] br[52] wl[37] vdd gnd cell_6t
Xbit_r38_c52 bl[52] br[52] wl[38] vdd gnd cell_6t
Xbit_r39_c52 bl[52] br[52] wl[39] vdd gnd cell_6t
Xbit_r40_c52 bl[52] br[52] wl[40] vdd gnd cell_6t
Xbit_r41_c52 bl[52] br[52] wl[41] vdd gnd cell_6t
Xbit_r42_c52 bl[52] br[52] wl[42] vdd gnd cell_6t
Xbit_r43_c52 bl[52] br[52] wl[43] vdd gnd cell_6t
Xbit_r44_c52 bl[52] br[52] wl[44] vdd gnd cell_6t
Xbit_r45_c52 bl[52] br[52] wl[45] vdd gnd cell_6t
Xbit_r46_c52 bl[52] br[52] wl[46] vdd gnd cell_6t
Xbit_r47_c52 bl[52] br[52] wl[47] vdd gnd cell_6t
Xbit_r48_c52 bl[52] br[52] wl[48] vdd gnd cell_6t
Xbit_r49_c52 bl[52] br[52] wl[49] vdd gnd cell_6t
Xbit_r50_c52 bl[52] br[52] wl[50] vdd gnd cell_6t
Xbit_r51_c52 bl[52] br[52] wl[51] vdd gnd cell_6t
Xbit_r52_c52 bl[52] br[52] wl[52] vdd gnd cell_6t
Xbit_r53_c52 bl[52] br[52] wl[53] vdd gnd cell_6t
Xbit_r54_c52 bl[52] br[52] wl[54] vdd gnd cell_6t
Xbit_r55_c52 bl[52] br[52] wl[55] vdd gnd cell_6t
Xbit_r56_c52 bl[52] br[52] wl[56] vdd gnd cell_6t
Xbit_r57_c52 bl[52] br[52] wl[57] vdd gnd cell_6t
Xbit_r58_c52 bl[52] br[52] wl[58] vdd gnd cell_6t
Xbit_r59_c52 bl[52] br[52] wl[59] vdd gnd cell_6t
Xbit_r60_c52 bl[52] br[52] wl[60] vdd gnd cell_6t
Xbit_r61_c52 bl[52] br[52] wl[61] vdd gnd cell_6t
Xbit_r62_c52 bl[52] br[52] wl[62] vdd gnd cell_6t
Xbit_r63_c52 bl[52] br[52] wl[63] vdd gnd cell_6t
Xbit_r64_c52 bl[52] br[52] wl[64] vdd gnd cell_6t
Xbit_r65_c52 bl[52] br[52] wl[65] vdd gnd cell_6t
Xbit_r66_c52 bl[52] br[52] wl[66] vdd gnd cell_6t
Xbit_r67_c52 bl[52] br[52] wl[67] vdd gnd cell_6t
Xbit_r68_c52 bl[52] br[52] wl[68] vdd gnd cell_6t
Xbit_r69_c52 bl[52] br[52] wl[69] vdd gnd cell_6t
Xbit_r70_c52 bl[52] br[52] wl[70] vdd gnd cell_6t
Xbit_r71_c52 bl[52] br[52] wl[71] vdd gnd cell_6t
Xbit_r72_c52 bl[52] br[52] wl[72] vdd gnd cell_6t
Xbit_r73_c52 bl[52] br[52] wl[73] vdd gnd cell_6t
Xbit_r74_c52 bl[52] br[52] wl[74] vdd gnd cell_6t
Xbit_r75_c52 bl[52] br[52] wl[75] vdd gnd cell_6t
Xbit_r76_c52 bl[52] br[52] wl[76] vdd gnd cell_6t
Xbit_r77_c52 bl[52] br[52] wl[77] vdd gnd cell_6t
Xbit_r78_c52 bl[52] br[52] wl[78] vdd gnd cell_6t
Xbit_r79_c52 bl[52] br[52] wl[79] vdd gnd cell_6t
Xbit_r80_c52 bl[52] br[52] wl[80] vdd gnd cell_6t
Xbit_r81_c52 bl[52] br[52] wl[81] vdd gnd cell_6t
Xbit_r82_c52 bl[52] br[52] wl[82] vdd gnd cell_6t
Xbit_r83_c52 bl[52] br[52] wl[83] vdd gnd cell_6t
Xbit_r84_c52 bl[52] br[52] wl[84] vdd gnd cell_6t
Xbit_r85_c52 bl[52] br[52] wl[85] vdd gnd cell_6t
Xbit_r86_c52 bl[52] br[52] wl[86] vdd gnd cell_6t
Xbit_r87_c52 bl[52] br[52] wl[87] vdd gnd cell_6t
Xbit_r88_c52 bl[52] br[52] wl[88] vdd gnd cell_6t
Xbit_r89_c52 bl[52] br[52] wl[89] vdd gnd cell_6t
Xbit_r90_c52 bl[52] br[52] wl[90] vdd gnd cell_6t
Xbit_r91_c52 bl[52] br[52] wl[91] vdd gnd cell_6t
Xbit_r92_c52 bl[52] br[52] wl[92] vdd gnd cell_6t
Xbit_r93_c52 bl[52] br[52] wl[93] vdd gnd cell_6t
Xbit_r94_c52 bl[52] br[52] wl[94] vdd gnd cell_6t
Xbit_r95_c52 bl[52] br[52] wl[95] vdd gnd cell_6t
Xbit_r96_c52 bl[52] br[52] wl[96] vdd gnd cell_6t
Xbit_r97_c52 bl[52] br[52] wl[97] vdd gnd cell_6t
Xbit_r98_c52 bl[52] br[52] wl[98] vdd gnd cell_6t
Xbit_r99_c52 bl[52] br[52] wl[99] vdd gnd cell_6t
Xbit_r100_c52 bl[52] br[52] wl[100] vdd gnd cell_6t
Xbit_r101_c52 bl[52] br[52] wl[101] vdd gnd cell_6t
Xbit_r102_c52 bl[52] br[52] wl[102] vdd gnd cell_6t
Xbit_r103_c52 bl[52] br[52] wl[103] vdd gnd cell_6t
Xbit_r104_c52 bl[52] br[52] wl[104] vdd gnd cell_6t
Xbit_r105_c52 bl[52] br[52] wl[105] vdd gnd cell_6t
Xbit_r106_c52 bl[52] br[52] wl[106] vdd gnd cell_6t
Xbit_r107_c52 bl[52] br[52] wl[107] vdd gnd cell_6t
Xbit_r108_c52 bl[52] br[52] wl[108] vdd gnd cell_6t
Xbit_r109_c52 bl[52] br[52] wl[109] vdd gnd cell_6t
Xbit_r110_c52 bl[52] br[52] wl[110] vdd gnd cell_6t
Xbit_r111_c52 bl[52] br[52] wl[111] vdd gnd cell_6t
Xbit_r112_c52 bl[52] br[52] wl[112] vdd gnd cell_6t
Xbit_r113_c52 bl[52] br[52] wl[113] vdd gnd cell_6t
Xbit_r114_c52 bl[52] br[52] wl[114] vdd gnd cell_6t
Xbit_r115_c52 bl[52] br[52] wl[115] vdd gnd cell_6t
Xbit_r116_c52 bl[52] br[52] wl[116] vdd gnd cell_6t
Xbit_r117_c52 bl[52] br[52] wl[117] vdd gnd cell_6t
Xbit_r118_c52 bl[52] br[52] wl[118] vdd gnd cell_6t
Xbit_r119_c52 bl[52] br[52] wl[119] vdd gnd cell_6t
Xbit_r120_c52 bl[52] br[52] wl[120] vdd gnd cell_6t
Xbit_r121_c52 bl[52] br[52] wl[121] vdd gnd cell_6t
Xbit_r122_c52 bl[52] br[52] wl[122] vdd gnd cell_6t
Xbit_r123_c52 bl[52] br[52] wl[123] vdd gnd cell_6t
Xbit_r124_c52 bl[52] br[52] wl[124] vdd gnd cell_6t
Xbit_r125_c52 bl[52] br[52] wl[125] vdd gnd cell_6t
Xbit_r126_c52 bl[52] br[52] wl[126] vdd gnd cell_6t
Xbit_r127_c52 bl[52] br[52] wl[127] vdd gnd cell_6t
Xbit_r128_c52 bl[52] br[52] wl[128] vdd gnd cell_6t
Xbit_r129_c52 bl[52] br[52] wl[129] vdd gnd cell_6t
Xbit_r130_c52 bl[52] br[52] wl[130] vdd gnd cell_6t
Xbit_r131_c52 bl[52] br[52] wl[131] vdd gnd cell_6t
Xbit_r132_c52 bl[52] br[52] wl[132] vdd gnd cell_6t
Xbit_r133_c52 bl[52] br[52] wl[133] vdd gnd cell_6t
Xbit_r134_c52 bl[52] br[52] wl[134] vdd gnd cell_6t
Xbit_r135_c52 bl[52] br[52] wl[135] vdd gnd cell_6t
Xbit_r136_c52 bl[52] br[52] wl[136] vdd gnd cell_6t
Xbit_r137_c52 bl[52] br[52] wl[137] vdd gnd cell_6t
Xbit_r138_c52 bl[52] br[52] wl[138] vdd gnd cell_6t
Xbit_r139_c52 bl[52] br[52] wl[139] vdd gnd cell_6t
Xbit_r140_c52 bl[52] br[52] wl[140] vdd gnd cell_6t
Xbit_r141_c52 bl[52] br[52] wl[141] vdd gnd cell_6t
Xbit_r142_c52 bl[52] br[52] wl[142] vdd gnd cell_6t
Xbit_r143_c52 bl[52] br[52] wl[143] vdd gnd cell_6t
Xbit_r144_c52 bl[52] br[52] wl[144] vdd gnd cell_6t
Xbit_r145_c52 bl[52] br[52] wl[145] vdd gnd cell_6t
Xbit_r146_c52 bl[52] br[52] wl[146] vdd gnd cell_6t
Xbit_r147_c52 bl[52] br[52] wl[147] vdd gnd cell_6t
Xbit_r148_c52 bl[52] br[52] wl[148] vdd gnd cell_6t
Xbit_r149_c52 bl[52] br[52] wl[149] vdd gnd cell_6t
Xbit_r150_c52 bl[52] br[52] wl[150] vdd gnd cell_6t
Xbit_r151_c52 bl[52] br[52] wl[151] vdd gnd cell_6t
Xbit_r152_c52 bl[52] br[52] wl[152] vdd gnd cell_6t
Xbit_r153_c52 bl[52] br[52] wl[153] vdd gnd cell_6t
Xbit_r154_c52 bl[52] br[52] wl[154] vdd gnd cell_6t
Xbit_r155_c52 bl[52] br[52] wl[155] vdd gnd cell_6t
Xbit_r156_c52 bl[52] br[52] wl[156] vdd gnd cell_6t
Xbit_r157_c52 bl[52] br[52] wl[157] vdd gnd cell_6t
Xbit_r158_c52 bl[52] br[52] wl[158] vdd gnd cell_6t
Xbit_r159_c52 bl[52] br[52] wl[159] vdd gnd cell_6t
Xbit_r160_c52 bl[52] br[52] wl[160] vdd gnd cell_6t
Xbit_r161_c52 bl[52] br[52] wl[161] vdd gnd cell_6t
Xbit_r162_c52 bl[52] br[52] wl[162] vdd gnd cell_6t
Xbit_r163_c52 bl[52] br[52] wl[163] vdd gnd cell_6t
Xbit_r164_c52 bl[52] br[52] wl[164] vdd gnd cell_6t
Xbit_r165_c52 bl[52] br[52] wl[165] vdd gnd cell_6t
Xbit_r166_c52 bl[52] br[52] wl[166] vdd gnd cell_6t
Xbit_r167_c52 bl[52] br[52] wl[167] vdd gnd cell_6t
Xbit_r168_c52 bl[52] br[52] wl[168] vdd gnd cell_6t
Xbit_r169_c52 bl[52] br[52] wl[169] vdd gnd cell_6t
Xbit_r170_c52 bl[52] br[52] wl[170] vdd gnd cell_6t
Xbit_r171_c52 bl[52] br[52] wl[171] vdd gnd cell_6t
Xbit_r172_c52 bl[52] br[52] wl[172] vdd gnd cell_6t
Xbit_r173_c52 bl[52] br[52] wl[173] vdd gnd cell_6t
Xbit_r174_c52 bl[52] br[52] wl[174] vdd gnd cell_6t
Xbit_r175_c52 bl[52] br[52] wl[175] vdd gnd cell_6t
Xbit_r176_c52 bl[52] br[52] wl[176] vdd gnd cell_6t
Xbit_r177_c52 bl[52] br[52] wl[177] vdd gnd cell_6t
Xbit_r178_c52 bl[52] br[52] wl[178] vdd gnd cell_6t
Xbit_r179_c52 bl[52] br[52] wl[179] vdd gnd cell_6t
Xbit_r180_c52 bl[52] br[52] wl[180] vdd gnd cell_6t
Xbit_r181_c52 bl[52] br[52] wl[181] vdd gnd cell_6t
Xbit_r182_c52 bl[52] br[52] wl[182] vdd gnd cell_6t
Xbit_r183_c52 bl[52] br[52] wl[183] vdd gnd cell_6t
Xbit_r184_c52 bl[52] br[52] wl[184] vdd gnd cell_6t
Xbit_r185_c52 bl[52] br[52] wl[185] vdd gnd cell_6t
Xbit_r186_c52 bl[52] br[52] wl[186] vdd gnd cell_6t
Xbit_r187_c52 bl[52] br[52] wl[187] vdd gnd cell_6t
Xbit_r188_c52 bl[52] br[52] wl[188] vdd gnd cell_6t
Xbit_r189_c52 bl[52] br[52] wl[189] vdd gnd cell_6t
Xbit_r190_c52 bl[52] br[52] wl[190] vdd gnd cell_6t
Xbit_r191_c52 bl[52] br[52] wl[191] vdd gnd cell_6t
Xbit_r192_c52 bl[52] br[52] wl[192] vdd gnd cell_6t
Xbit_r193_c52 bl[52] br[52] wl[193] vdd gnd cell_6t
Xbit_r194_c52 bl[52] br[52] wl[194] vdd gnd cell_6t
Xbit_r195_c52 bl[52] br[52] wl[195] vdd gnd cell_6t
Xbit_r196_c52 bl[52] br[52] wl[196] vdd gnd cell_6t
Xbit_r197_c52 bl[52] br[52] wl[197] vdd gnd cell_6t
Xbit_r198_c52 bl[52] br[52] wl[198] vdd gnd cell_6t
Xbit_r199_c52 bl[52] br[52] wl[199] vdd gnd cell_6t
Xbit_r200_c52 bl[52] br[52] wl[200] vdd gnd cell_6t
Xbit_r201_c52 bl[52] br[52] wl[201] vdd gnd cell_6t
Xbit_r202_c52 bl[52] br[52] wl[202] vdd gnd cell_6t
Xbit_r203_c52 bl[52] br[52] wl[203] vdd gnd cell_6t
Xbit_r204_c52 bl[52] br[52] wl[204] vdd gnd cell_6t
Xbit_r205_c52 bl[52] br[52] wl[205] vdd gnd cell_6t
Xbit_r206_c52 bl[52] br[52] wl[206] vdd gnd cell_6t
Xbit_r207_c52 bl[52] br[52] wl[207] vdd gnd cell_6t
Xbit_r208_c52 bl[52] br[52] wl[208] vdd gnd cell_6t
Xbit_r209_c52 bl[52] br[52] wl[209] vdd gnd cell_6t
Xbit_r210_c52 bl[52] br[52] wl[210] vdd gnd cell_6t
Xbit_r211_c52 bl[52] br[52] wl[211] vdd gnd cell_6t
Xbit_r212_c52 bl[52] br[52] wl[212] vdd gnd cell_6t
Xbit_r213_c52 bl[52] br[52] wl[213] vdd gnd cell_6t
Xbit_r214_c52 bl[52] br[52] wl[214] vdd gnd cell_6t
Xbit_r215_c52 bl[52] br[52] wl[215] vdd gnd cell_6t
Xbit_r216_c52 bl[52] br[52] wl[216] vdd gnd cell_6t
Xbit_r217_c52 bl[52] br[52] wl[217] vdd gnd cell_6t
Xbit_r218_c52 bl[52] br[52] wl[218] vdd gnd cell_6t
Xbit_r219_c52 bl[52] br[52] wl[219] vdd gnd cell_6t
Xbit_r220_c52 bl[52] br[52] wl[220] vdd gnd cell_6t
Xbit_r221_c52 bl[52] br[52] wl[221] vdd gnd cell_6t
Xbit_r222_c52 bl[52] br[52] wl[222] vdd gnd cell_6t
Xbit_r223_c52 bl[52] br[52] wl[223] vdd gnd cell_6t
Xbit_r224_c52 bl[52] br[52] wl[224] vdd gnd cell_6t
Xbit_r225_c52 bl[52] br[52] wl[225] vdd gnd cell_6t
Xbit_r226_c52 bl[52] br[52] wl[226] vdd gnd cell_6t
Xbit_r227_c52 bl[52] br[52] wl[227] vdd gnd cell_6t
Xbit_r228_c52 bl[52] br[52] wl[228] vdd gnd cell_6t
Xbit_r229_c52 bl[52] br[52] wl[229] vdd gnd cell_6t
Xbit_r230_c52 bl[52] br[52] wl[230] vdd gnd cell_6t
Xbit_r231_c52 bl[52] br[52] wl[231] vdd gnd cell_6t
Xbit_r232_c52 bl[52] br[52] wl[232] vdd gnd cell_6t
Xbit_r233_c52 bl[52] br[52] wl[233] vdd gnd cell_6t
Xbit_r234_c52 bl[52] br[52] wl[234] vdd gnd cell_6t
Xbit_r235_c52 bl[52] br[52] wl[235] vdd gnd cell_6t
Xbit_r236_c52 bl[52] br[52] wl[236] vdd gnd cell_6t
Xbit_r237_c52 bl[52] br[52] wl[237] vdd gnd cell_6t
Xbit_r238_c52 bl[52] br[52] wl[238] vdd gnd cell_6t
Xbit_r239_c52 bl[52] br[52] wl[239] vdd gnd cell_6t
Xbit_r240_c52 bl[52] br[52] wl[240] vdd gnd cell_6t
Xbit_r241_c52 bl[52] br[52] wl[241] vdd gnd cell_6t
Xbit_r242_c52 bl[52] br[52] wl[242] vdd gnd cell_6t
Xbit_r243_c52 bl[52] br[52] wl[243] vdd gnd cell_6t
Xbit_r244_c52 bl[52] br[52] wl[244] vdd gnd cell_6t
Xbit_r245_c52 bl[52] br[52] wl[245] vdd gnd cell_6t
Xbit_r246_c52 bl[52] br[52] wl[246] vdd gnd cell_6t
Xbit_r247_c52 bl[52] br[52] wl[247] vdd gnd cell_6t
Xbit_r248_c52 bl[52] br[52] wl[248] vdd gnd cell_6t
Xbit_r249_c52 bl[52] br[52] wl[249] vdd gnd cell_6t
Xbit_r250_c52 bl[52] br[52] wl[250] vdd gnd cell_6t
Xbit_r251_c52 bl[52] br[52] wl[251] vdd gnd cell_6t
Xbit_r252_c52 bl[52] br[52] wl[252] vdd gnd cell_6t
Xbit_r253_c52 bl[52] br[52] wl[253] vdd gnd cell_6t
Xbit_r254_c52 bl[52] br[52] wl[254] vdd gnd cell_6t
Xbit_r255_c52 bl[52] br[52] wl[255] vdd gnd cell_6t
Xbit_r0_c53 bl[53] br[53] wl[0] vdd gnd cell_6t
Xbit_r1_c53 bl[53] br[53] wl[1] vdd gnd cell_6t
Xbit_r2_c53 bl[53] br[53] wl[2] vdd gnd cell_6t
Xbit_r3_c53 bl[53] br[53] wl[3] vdd gnd cell_6t
Xbit_r4_c53 bl[53] br[53] wl[4] vdd gnd cell_6t
Xbit_r5_c53 bl[53] br[53] wl[5] vdd gnd cell_6t
Xbit_r6_c53 bl[53] br[53] wl[6] vdd gnd cell_6t
Xbit_r7_c53 bl[53] br[53] wl[7] vdd gnd cell_6t
Xbit_r8_c53 bl[53] br[53] wl[8] vdd gnd cell_6t
Xbit_r9_c53 bl[53] br[53] wl[9] vdd gnd cell_6t
Xbit_r10_c53 bl[53] br[53] wl[10] vdd gnd cell_6t
Xbit_r11_c53 bl[53] br[53] wl[11] vdd gnd cell_6t
Xbit_r12_c53 bl[53] br[53] wl[12] vdd gnd cell_6t
Xbit_r13_c53 bl[53] br[53] wl[13] vdd gnd cell_6t
Xbit_r14_c53 bl[53] br[53] wl[14] vdd gnd cell_6t
Xbit_r15_c53 bl[53] br[53] wl[15] vdd gnd cell_6t
Xbit_r16_c53 bl[53] br[53] wl[16] vdd gnd cell_6t
Xbit_r17_c53 bl[53] br[53] wl[17] vdd gnd cell_6t
Xbit_r18_c53 bl[53] br[53] wl[18] vdd gnd cell_6t
Xbit_r19_c53 bl[53] br[53] wl[19] vdd gnd cell_6t
Xbit_r20_c53 bl[53] br[53] wl[20] vdd gnd cell_6t
Xbit_r21_c53 bl[53] br[53] wl[21] vdd gnd cell_6t
Xbit_r22_c53 bl[53] br[53] wl[22] vdd gnd cell_6t
Xbit_r23_c53 bl[53] br[53] wl[23] vdd gnd cell_6t
Xbit_r24_c53 bl[53] br[53] wl[24] vdd gnd cell_6t
Xbit_r25_c53 bl[53] br[53] wl[25] vdd gnd cell_6t
Xbit_r26_c53 bl[53] br[53] wl[26] vdd gnd cell_6t
Xbit_r27_c53 bl[53] br[53] wl[27] vdd gnd cell_6t
Xbit_r28_c53 bl[53] br[53] wl[28] vdd gnd cell_6t
Xbit_r29_c53 bl[53] br[53] wl[29] vdd gnd cell_6t
Xbit_r30_c53 bl[53] br[53] wl[30] vdd gnd cell_6t
Xbit_r31_c53 bl[53] br[53] wl[31] vdd gnd cell_6t
Xbit_r32_c53 bl[53] br[53] wl[32] vdd gnd cell_6t
Xbit_r33_c53 bl[53] br[53] wl[33] vdd gnd cell_6t
Xbit_r34_c53 bl[53] br[53] wl[34] vdd gnd cell_6t
Xbit_r35_c53 bl[53] br[53] wl[35] vdd gnd cell_6t
Xbit_r36_c53 bl[53] br[53] wl[36] vdd gnd cell_6t
Xbit_r37_c53 bl[53] br[53] wl[37] vdd gnd cell_6t
Xbit_r38_c53 bl[53] br[53] wl[38] vdd gnd cell_6t
Xbit_r39_c53 bl[53] br[53] wl[39] vdd gnd cell_6t
Xbit_r40_c53 bl[53] br[53] wl[40] vdd gnd cell_6t
Xbit_r41_c53 bl[53] br[53] wl[41] vdd gnd cell_6t
Xbit_r42_c53 bl[53] br[53] wl[42] vdd gnd cell_6t
Xbit_r43_c53 bl[53] br[53] wl[43] vdd gnd cell_6t
Xbit_r44_c53 bl[53] br[53] wl[44] vdd gnd cell_6t
Xbit_r45_c53 bl[53] br[53] wl[45] vdd gnd cell_6t
Xbit_r46_c53 bl[53] br[53] wl[46] vdd gnd cell_6t
Xbit_r47_c53 bl[53] br[53] wl[47] vdd gnd cell_6t
Xbit_r48_c53 bl[53] br[53] wl[48] vdd gnd cell_6t
Xbit_r49_c53 bl[53] br[53] wl[49] vdd gnd cell_6t
Xbit_r50_c53 bl[53] br[53] wl[50] vdd gnd cell_6t
Xbit_r51_c53 bl[53] br[53] wl[51] vdd gnd cell_6t
Xbit_r52_c53 bl[53] br[53] wl[52] vdd gnd cell_6t
Xbit_r53_c53 bl[53] br[53] wl[53] vdd gnd cell_6t
Xbit_r54_c53 bl[53] br[53] wl[54] vdd gnd cell_6t
Xbit_r55_c53 bl[53] br[53] wl[55] vdd gnd cell_6t
Xbit_r56_c53 bl[53] br[53] wl[56] vdd gnd cell_6t
Xbit_r57_c53 bl[53] br[53] wl[57] vdd gnd cell_6t
Xbit_r58_c53 bl[53] br[53] wl[58] vdd gnd cell_6t
Xbit_r59_c53 bl[53] br[53] wl[59] vdd gnd cell_6t
Xbit_r60_c53 bl[53] br[53] wl[60] vdd gnd cell_6t
Xbit_r61_c53 bl[53] br[53] wl[61] vdd gnd cell_6t
Xbit_r62_c53 bl[53] br[53] wl[62] vdd gnd cell_6t
Xbit_r63_c53 bl[53] br[53] wl[63] vdd gnd cell_6t
Xbit_r64_c53 bl[53] br[53] wl[64] vdd gnd cell_6t
Xbit_r65_c53 bl[53] br[53] wl[65] vdd gnd cell_6t
Xbit_r66_c53 bl[53] br[53] wl[66] vdd gnd cell_6t
Xbit_r67_c53 bl[53] br[53] wl[67] vdd gnd cell_6t
Xbit_r68_c53 bl[53] br[53] wl[68] vdd gnd cell_6t
Xbit_r69_c53 bl[53] br[53] wl[69] vdd gnd cell_6t
Xbit_r70_c53 bl[53] br[53] wl[70] vdd gnd cell_6t
Xbit_r71_c53 bl[53] br[53] wl[71] vdd gnd cell_6t
Xbit_r72_c53 bl[53] br[53] wl[72] vdd gnd cell_6t
Xbit_r73_c53 bl[53] br[53] wl[73] vdd gnd cell_6t
Xbit_r74_c53 bl[53] br[53] wl[74] vdd gnd cell_6t
Xbit_r75_c53 bl[53] br[53] wl[75] vdd gnd cell_6t
Xbit_r76_c53 bl[53] br[53] wl[76] vdd gnd cell_6t
Xbit_r77_c53 bl[53] br[53] wl[77] vdd gnd cell_6t
Xbit_r78_c53 bl[53] br[53] wl[78] vdd gnd cell_6t
Xbit_r79_c53 bl[53] br[53] wl[79] vdd gnd cell_6t
Xbit_r80_c53 bl[53] br[53] wl[80] vdd gnd cell_6t
Xbit_r81_c53 bl[53] br[53] wl[81] vdd gnd cell_6t
Xbit_r82_c53 bl[53] br[53] wl[82] vdd gnd cell_6t
Xbit_r83_c53 bl[53] br[53] wl[83] vdd gnd cell_6t
Xbit_r84_c53 bl[53] br[53] wl[84] vdd gnd cell_6t
Xbit_r85_c53 bl[53] br[53] wl[85] vdd gnd cell_6t
Xbit_r86_c53 bl[53] br[53] wl[86] vdd gnd cell_6t
Xbit_r87_c53 bl[53] br[53] wl[87] vdd gnd cell_6t
Xbit_r88_c53 bl[53] br[53] wl[88] vdd gnd cell_6t
Xbit_r89_c53 bl[53] br[53] wl[89] vdd gnd cell_6t
Xbit_r90_c53 bl[53] br[53] wl[90] vdd gnd cell_6t
Xbit_r91_c53 bl[53] br[53] wl[91] vdd gnd cell_6t
Xbit_r92_c53 bl[53] br[53] wl[92] vdd gnd cell_6t
Xbit_r93_c53 bl[53] br[53] wl[93] vdd gnd cell_6t
Xbit_r94_c53 bl[53] br[53] wl[94] vdd gnd cell_6t
Xbit_r95_c53 bl[53] br[53] wl[95] vdd gnd cell_6t
Xbit_r96_c53 bl[53] br[53] wl[96] vdd gnd cell_6t
Xbit_r97_c53 bl[53] br[53] wl[97] vdd gnd cell_6t
Xbit_r98_c53 bl[53] br[53] wl[98] vdd gnd cell_6t
Xbit_r99_c53 bl[53] br[53] wl[99] vdd gnd cell_6t
Xbit_r100_c53 bl[53] br[53] wl[100] vdd gnd cell_6t
Xbit_r101_c53 bl[53] br[53] wl[101] vdd gnd cell_6t
Xbit_r102_c53 bl[53] br[53] wl[102] vdd gnd cell_6t
Xbit_r103_c53 bl[53] br[53] wl[103] vdd gnd cell_6t
Xbit_r104_c53 bl[53] br[53] wl[104] vdd gnd cell_6t
Xbit_r105_c53 bl[53] br[53] wl[105] vdd gnd cell_6t
Xbit_r106_c53 bl[53] br[53] wl[106] vdd gnd cell_6t
Xbit_r107_c53 bl[53] br[53] wl[107] vdd gnd cell_6t
Xbit_r108_c53 bl[53] br[53] wl[108] vdd gnd cell_6t
Xbit_r109_c53 bl[53] br[53] wl[109] vdd gnd cell_6t
Xbit_r110_c53 bl[53] br[53] wl[110] vdd gnd cell_6t
Xbit_r111_c53 bl[53] br[53] wl[111] vdd gnd cell_6t
Xbit_r112_c53 bl[53] br[53] wl[112] vdd gnd cell_6t
Xbit_r113_c53 bl[53] br[53] wl[113] vdd gnd cell_6t
Xbit_r114_c53 bl[53] br[53] wl[114] vdd gnd cell_6t
Xbit_r115_c53 bl[53] br[53] wl[115] vdd gnd cell_6t
Xbit_r116_c53 bl[53] br[53] wl[116] vdd gnd cell_6t
Xbit_r117_c53 bl[53] br[53] wl[117] vdd gnd cell_6t
Xbit_r118_c53 bl[53] br[53] wl[118] vdd gnd cell_6t
Xbit_r119_c53 bl[53] br[53] wl[119] vdd gnd cell_6t
Xbit_r120_c53 bl[53] br[53] wl[120] vdd gnd cell_6t
Xbit_r121_c53 bl[53] br[53] wl[121] vdd gnd cell_6t
Xbit_r122_c53 bl[53] br[53] wl[122] vdd gnd cell_6t
Xbit_r123_c53 bl[53] br[53] wl[123] vdd gnd cell_6t
Xbit_r124_c53 bl[53] br[53] wl[124] vdd gnd cell_6t
Xbit_r125_c53 bl[53] br[53] wl[125] vdd gnd cell_6t
Xbit_r126_c53 bl[53] br[53] wl[126] vdd gnd cell_6t
Xbit_r127_c53 bl[53] br[53] wl[127] vdd gnd cell_6t
Xbit_r128_c53 bl[53] br[53] wl[128] vdd gnd cell_6t
Xbit_r129_c53 bl[53] br[53] wl[129] vdd gnd cell_6t
Xbit_r130_c53 bl[53] br[53] wl[130] vdd gnd cell_6t
Xbit_r131_c53 bl[53] br[53] wl[131] vdd gnd cell_6t
Xbit_r132_c53 bl[53] br[53] wl[132] vdd gnd cell_6t
Xbit_r133_c53 bl[53] br[53] wl[133] vdd gnd cell_6t
Xbit_r134_c53 bl[53] br[53] wl[134] vdd gnd cell_6t
Xbit_r135_c53 bl[53] br[53] wl[135] vdd gnd cell_6t
Xbit_r136_c53 bl[53] br[53] wl[136] vdd gnd cell_6t
Xbit_r137_c53 bl[53] br[53] wl[137] vdd gnd cell_6t
Xbit_r138_c53 bl[53] br[53] wl[138] vdd gnd cell_6t
Xbit_r139_c53 bl[53] br[53] wl[139] vdd gnd cell_6t
Xbit_r140_c53 bl[53] br[53] wl[140] vdd gnd cell_6t
Xbit_r141_c53 bl[53] br[53] wl[141] vdd gnd cell_6t
Xbit_r142_c53 bl[53] br[53] wl[142] vdd gnd cell_6t
Xbit_r143_c53 bl[53] br[53] wl[143] vdd gnd cell_6t
Xbit_r144_c53 bl[53] br[53] wl[144] vdd gnd cell_6t
Xbit_r145_c53 bl[53] br[53] wl[145] vdd gnd cell_6t
Xbit_r146_c53 bl[53] br[53] wl[146] vdd gnd cell_6t
Xbit_r147_c53 bl[53] br[53] wl[147] vdd gnd cell_6t
Xbit_r148_c53 bl[53] br[53] wl[148] vdd gnd cell_6t
Xbit_r149_c53 bl[53] br[53] wl[149] vdd gnd cell_6t
Xbit_r150_c53 bl[53] br[53] wl[150] vdd gnd cell_6t
Xbit_r151_c53 bl[53] br[53] wl[151] vdd gnd cell_6t
Xbit_r152_c53 bl[53] br[53] wl[152] vdd gnd cell_6t
Xbit_r153_c53 bl[53] br[53] wl[153] vdd gnd cell_6t
Xbit_r154_c53 bl[53] br[53] wl[154] vdd gnd cell_6t
Xbit_r155_c53 bl[53] br[53] wl[155] vdd gnd cell_6t
Xbit_r156_c53 bl[53] br[53] wl[156] vdd gnd cell_6t
Xbit_r157_c53 bl[53] br[53] wl[157] vdd gnd cell_6t
Xbit_r158_c53 bl[53] br[53] wl[158] vdd gnd cell_6t
Xbit_r159_c53 bl[53] br[53] wl[159] vdd gnd cell_6t
Xbit_r160_c53 bl[53] br[53] wl[160] vdd gnd cell_6t
Xbit_r161_c53 bl[53] br[53] wl[161] vdd gnd cell_6t
Xbit_r162_c53 bl[53] br[53] wl[162] vdd gnd cell_6t
Xbit_r163_c53 bl[53] br[53] wl[163] vdd gnd cell_6t
Xbit_r164_c53 bl[53] br[53] wl[164] vdd gnd cell_6t
Xbit_r165_c53 bl[53] br[53] wl[165] vdd gnd cell_6t
Xbit_r166_c53 bl[53] br[53] wl[166] vdd gnd cell_6t
Xbit_r167_c53 bl[53] br[53] wl[167] vdd gnd cell_6t
Xbit_r168_c53 bl[53] br[53] wl[168] vdd gnd cell_6t
Xbit_r169_c53 bl[53] br[53] wl[169] vdd gnd cell_6t
Xbit_r170_c53 bl[53] br[53] wl[170] vdd gnd cell_6t
Xbit_r171_c53 bl[53] br[53] wl[171] vdd gnd cell_6t
Xbit_r172_c53 bl[53] br[53] wl[172] vdd gnd cell_6t
Xbit_r173_c53 bl[53] br[53] wl[173] vdd gnd cell_6t
Xbit_r174_c53 bl[53] br[53] wl[174] vdd gnd cell_6t
Xbit_r175_c53 bl[53] br[53] wl[175] vdd gnd cell_6t
Xbit_r176_c53 bl[53] br[53] wl[176] vdd gnd cell_6t
Xbit_r177_c53 bl[53] br[53] wl[177] vdd gnd cell_6t
Xbit_r178_c53 bl[53] br[53] wl[178] vdd gnd cell_6t
Xbit_r179_c53 bl[53] br[53] wl[179] vdd gnd cell_6t
Xbit_r180_c53 bl[53] br[53] wl[180] vdd gnd cell_6t
Xbit_r181_c53 bl[53] br[53] wl[181] vdd gnd cell_6t
Xbit_r182_c53 bl[53] br[53] wl[182] vdd gnd cell_6t
Xbit_r183_c53 bl[53] br[53] wl[183] vdd gnd cell_6t
Xbit_r184_c53 bl[53] br[53] wl[184] vdd gnd cell_6t
Xbit_r185_c53 bl[53] br[53] wl[185] vdd gnd cell_6t
Xbit_r186_c53 bl[53] br[53] wl[186] vdd gnd cell_6t
Xbit_r187_c53 bl[53] br[53] wl[187] vdd gnd cell_6t
Xbit_r188_c53 bl[53] br[53] wl[188] vdd gnd cell_6t
Xbit_r189_c53 bl[53] br[53] wl[189] vdd gnd cell_6t
Xbit_r190_c53 bl[53] br[53] wl[190] vdd gnd cell_6t
Xbit_r191_c53 bl[53] br[53] wl[191] vdd gnd cell_6t
Xbit_r192_c53 bl[53] br[53] wl[192] vdd gnd cell_6t
Xbit_r193_c53 bl[53] br[53] wl[193] vdd gnd cell_6t
Xbit_r194_c53 bl[53] br[53] wl[194] vdd gnd cell_6t
Xbit_r195_c53 bl[53] br[53] wl[195] vdd gnd cell_6t
Xbit_r196_c53 bl[53] br[53] wl[196] vdd gnd cell_6t
Xbit_r197_c53 bl[53] br[53] wl[197] vdd gnd cell_6t
Xbit_r198_c53 bl[53] br[53] wl[198] vdd gnd cell_6t
Xbit_r199_c53 bl[53] br[53] wl[199] vdd gnd cell_6t
Xbit_r200_c53 bl[53] br[53] wl[200] vdd gnd cell_6t
Xbit_r201_c53 bl[53] br[53] wl[201] vdd gnd cell_6t
Xbit_r202_c53 bl[53] br[53] wl[202] vdd gnd cell_6t
Xbit_r203_c53 bl[53] br[53] wl[203] vdd gnd cell_6t
Xbit_r204_c53 bl[53] br[53] wl[204] vdd gnd cell_6t
Xbit_r205_c53 bl[53] br[53] wl[205] vdd gnd cell_6t
Xbit_r206_c53 bl[53] br[53] wl[206] vdd gnd cell_6t
Xbit_r207_c53 bl[53] br[53] wl[207] vdd gnd cell_6t
Xbit_r208_c53 bl[53] br[53] wl[208] vdd gnd cell_6t
Xbit_r209_c53 bl[53] br[53] wl[209] vdd gnd cell_6t
Xbit_r210_c53 bl[53] br[53] wl[210] vdd gnd cell_6t
Xbit_r211_c53 bl[53] br[53] wl[211] vdd gnd cell_6t
Xbit_r212_c53 bl[53] br[53] wl[212] vdd gnd cell_6t
Xbit_r213_c53 bl[53] br[53] wl[213] vdd gnd cell_6t
Xbit_r214_c53 bl[53] br[53] wl[214] vdd gnd cell_6t
Xbit_r215_c53 bl[53] br[53] wl[215] vdd gnd cell_6t
Xbit_r216_c53 bl[53] br[53] wl[216] vdd gnd cell_6t
Xbit_r217_c53 bl[53] br[53] wl[217] vdd gnd cell_6t
Xbit_r218_c53 bl[53] br[53] wl[218] vdd gnd cell_6t
Xbit_r219_c53 bl[53] br[53] wl[219] vdd gnd cell_6t
Xbit_r220_c53 bl[53] br[53] wl[220] vdd gnd cell_6t
Xbit_r221_c53 bl[53] br[53] wl[221] vdd gnd cell_6t
Xbit_r222_c53 bl[53] br[53] wl[222] vdd gnd cell_6t
Xbit_r223_c53 bl[53] br[53] wl[223] vdd gnd cell_6t
Xbit_r224_c53 bl[53] br[53] wl[224] vdd gnd cell_6t
Xbit_r225_c53 bl[53] br[53] wl[225] vdd gnd cell_6t
Xbit_r226_c53 bl[53] br[53] wl[226] vdd gnd cell_6t
Xbit_r227_c53 bl[53] br[53] wl[227] vdd gnd cell_6t
Xbit_r228_c53 bl[53] br[53] wl[228] vdd gnd cell_6t
Xbit_r229_c53 bl[53] br[53] wl[229] vdd gnd cell_6t
Xbit_r230_c53 bl[53] br[53] wl[230] vdd gnd cell_6t
Xbit_r231_c53 bl[53] br[53] wl[231] vdd gnd cell_6t
Xbit_r232_c53 bl[53] br[53] wl[232] vdd gnd cell_6t
Xbit_r233_c53 bl[53] br[53] wl[233] vdd gnd cell_6t
Xbit_r234_c53 bl[53] br[53] wl[234] vdd gnd cell_6t
Xbit_r235_c53 bl[53] br[53] wl[235] vdd gnd cell_6t
Xbit_r236_c53 bl[53] br[53] wl[236] vdd gnd cell_6t
Xbit_r237_c53 bl[53] br[53] wl[237] vdd gnd cell_6t
Xbit_r238_c53 bl[53] br[53] wl[238] vdd gnd cell_6t
Xbit_r239_c53 bl[53] br[53] wl[239] vdd gnd cell_6t
Xbit_r240_c53 bl[53] br[53] wl[240] vdd gnd cell_6t
Xbit_r241_c53 bl[53] br[53] wl[241] vdd gnd cell_6t
Xbit_r242_c53 bl[53] br[53] wl[242] vdd gnd cell_6t
Xbit_r243_c53 bl[53] br[53] wl[243] vdd gnd cell_6t
Xbit_r244_c53 bl[53] br[53] wl[244] vdd gnd cell_6t
Xbit_r245_c53 bl[53] br[53] wl[245] vdd gnd cell_6t
Xbit_r246_c53 bl[53] br[53] wl[246] vdd gnd cell_6t
Xbit_r247_c53 bl[53] br[53] wl[247] vdd gnd cell_6t
Xbit_r248_c53 bl[53] br[53] wl[248] vdd gnd cell_6t
Xbit_r249_c53 bl[53] br[53] wl[249] vdd gnd cell_6t
Xbit_r250_c53 bl[53] br[53] wl[250] vdd gnd cell_6t
Xbit_r251_c53 bl[53] br[53] wl[251] vdd gnd cell_6t
Xbit_r252_c53 bl[53] br[53] wl[252] vdd gnd cell_6t
Xbit_r253_c53 bl[53] br[53] wl[253] vdd gnd cell_6t
Xbit_r254_c53 bl[53] br[53] wl[254] vdd gnd cell_6t
Xbit_r255_c53 bl[53] br[53] wl[255] vdd gnd cell_6t
Xbit_r0_c54 bl[54] br[54] wl[0] vdd gnd cell_6t
Xbit_r1_c54 bl[54] br[54] wl[1] vdd gnd cell_6t
Xbit_r2_c54 bl[54] br[54] wl[2] vdd gnd cell_6t
Xbit_r3_c54 bl[54] br[54] wl[3] vdd gnd cell_6t
Xbit_r4_c54 bl[54] br[54] wl[4] vdd gnd cell_6t
Xbit_r5_c54 bl[54] br[54] wl[5] vdd gnd cell_6t
Xbit_r6_c54 bl[54] br[54] wl[6] vdd gnd cell_6t
Xbit_r7_c54 bl[54] br[54] wl[7] vdd gnd cell_6t
Xbit_r8_c54 bl[54] br[54] wl[8] vdd gnd cell_6t
Xbit_r9_c54 bl[54] br[54] wl[9] vdd gnd cell_6t
Xbit_r10_c54 bl[54] br[54] wl[10] vdd gnd cell_6t
Xbit_r11_c54 bl[54] br[54] wl[11] vdd gnd cell_6t
Xbit_r12_c54 bl[54] br[54] wl[12] vdd gnd cell_6t
Xbit_r13_c54 bl[54] br[54] wl[13] vdd gnd cell_6t
Xbit_r14_c54 bl[54] br[54] wl[14] vdd gnd cell_6t
Xbit_r15_c54 bl[54] br[54] wl[15] vdd gnd cell_6t
Xbit_r16_c54 bl[54] br[54] wl[16] vdd gnd cell_6t
Xbit_r17_c54 bl[54] br[54] wl[17] vdd gnd cell_6t
Xbit_r18_c54 bl[54] br[54] wl[18] vdd gnd cell_6t
Xbit_r19_c54 bl[54] br[54] wl[19] vdd gnd cell_6t
Xbit_r20_c54 bl[54] br[54] wl[20] vdd gnd cell_6t
Xbit_r21_c54 bl[54] br[54] wl[21] vdd gnd cell_6t
Xbit_r22_c54 bl[54] br[54] wl[22] vdd gnd cell_6t
Xbit_r23_c54 bl[54] br[54] wl[23] vdd gnd cell_6t
Xbit_r24_c54 bl[54] br[54] wl[24] vdd gnd cell_6t
Xbit_r25_c54 bl[54] br[54] wl[25] vdd gnd cell_6t
Xbit_r26_c54 bl[54] br[54] wl[26] vdd gnd cell_6t
Xbit_r27_c54 bl[54] br[54] wl[27] vdd gnd cell_6t
Xbit_r28_c54 bl[54] br[54] wl[28] vdd gnd cell_6t
Xbit_r29_c54 bl[54] br[54] wl[29] vdd gnd cell_6t
Xbit_r30_c54 bl[54] br[54] wl[30] vdd gnd cell_6t
Xbit_r31_c54 bl[54] br[54] wl[31] vdd gnd cell_6t
Xbit_r32_c54 bl[54] br[54] wl[32] vdd gnd cell_6t
Xbit_r33_c54 bl[54] br[54] wl[33] vdd gnd cell_6t
Xbit_r34_c54 bl[54] br[54] wl[34] vdd gnd cell_6t
Xbit_r35_c54 bl[54] br[54] wl[35] vdd gnd cell_6t
Xbit_r36_c54 bl[54] br[54] wl[36] vdd gnd cell_6t
Xbit_r37_c54 bl[54] br[54] wl[37] vdd gnd cell_6t
Xbit_r38_c54 bl[54] br[54] wl[38] vdd gnd cell_6t
Xbit_r39_c54 bl[54] br[54] wl[39] vdd gnd cell_6t
Xbit_r40_c54 bl[54] br[54] wl[40] vdd gnd cell_6t
Xbit_r41_c54 bl[54] br[54] wl[41] vdd gnd cell_6t
Xbit_r42_c54 bl[54] br[54] wl[42] vdd gnd cell_6t
Xbit_r43_c54 bl[54] br[54] wl[43] vdd gnd cell_6t
Xbit_r44_c54 bl[54] br[54] wl[44] vdd gnd cell_6t
Xbit_r45_c54 bl[54] br[54] wl[45] vdd gnd cell_6t
Xbit_r46_c54 bl[54] br[54] wl[46] vdd gnd cell_6t
Xbit_r47_c54 bl[54] br[54] wl[47] vdd gnd cell_6t
Xbit_r48_c54 bl[54] br[54] wl[48] vdd gnd cell_6t
Xbit_r49_c54 bl[54] br[54] wl[49] vdd gnd cell_6t
Xbit_r50_c54 bl[54] br[54] wl[50] vdd gnd cell_6t
Xbit_r51_c54 bl[54] br[54] wl[51] vdd gnd cell_6t
Xbit_r52_c54 bl[54] br[54] wl[52] vdd gnd cell_6t
Xbit_r53_c54 bl[54] br[54] wl[53] vdd gnd cell_6t
Xbit_r54_c54 bl[54] br[54] wl[54] vdd gnd cell_6t
Xbit_r55_c54 bl[54] br[54] wl[55] vdd gnd cell_6t
Xbit_r56_c54 bl[54] br[54] wl[56] vdd gnd cell_6t
Xbit_r57_c54 bl[54] br[54] wl[57] vdd gnd cell_6t
Xbit_r58_c54 bl[54] br[54] wl[58] vdd gnd cell_6t
Xbit_r59_c54 bl[54] br[54] wl[59] vdd gnd cell_6t
Xbit_r60_c54 bl[54] br[54] wl[60] vdd gnd cell_6t
Xbit_r61_c54 bl[54] br[54] wl[61] vdd gnd cell_6t
Xbit_r62_c54 bl[54] br[54] wl[62] vdd gnd cell_6t
Xbit_r63_c54 bl[54] br[54] wl[63] vdd gnd cell_6t
Xbit_r64_c54 bl[54] br[54] wl[64] vdd gnd cell_6t
Xbit_r65_c54 bl[54] br[54] wl[65] vdd gnd cell_6t
Xbit_r66_c54 bl[54] br[54] wl[66] vdd gnd cell_6t
Xbit_r67_c54 bl[54] br[54] wl[67] vdd gnd cell_6t
Xbit_r68_c54 bl[54] br[54] wl[68] vdd gnd cell_6t
Xbit_r69_c54 bl[54] br[54] wl[69] vdd gnd cell_6t
Xbit_r70_c54 bl[54] br[54] wl[70] vdd gnd cell_6t
Xbit_r71_c54 bl[54] br[54] wl[71] vdd gnd cell_6t
Xbit_r72_c54 bl[54] br[54] wl[72] vdd gnd cell_6t
Xbit_r73_c54 bl[54] br[54] wl[73] vdd gnd cell_6t
Xbit_r74_c54 bl[54] br[54] wl[74] vdd gnd cell_6t
Xbit_r75_c54 bl[54] br[54] wl[75] vdd gnd cell_6t
Xbit_r76_c54 bl[54] br[54] wl[76] vdd gnd cell_6t
Xbit_r77_c54 bl[54] br[54] wl[77] vdd gnd cell_6t
Xbit_r78_c54 bl[54] br[54] wl[78] vdd gnd cell_6t
Xbit_r79_c54 bl[54] br[54] wl[79] vdd gnd cell_6t
Xbit_r80_c54 bl[54] br[54] wl[80] vdd gnd cell_6t
Xbit_r81_c54 bl[54] br[54] wl[81] vdd gnd cell_6t
Xbit_r82_c54 bl[54] br[54] wl[82] vdd gnd cell_6t
Xbit_r83_c54 bl[54] br[54] wl[83] vdd gnd cell_6t
Xbit_r84_c54 bl[54] br[54] wl[84] vdd gnd cell_6t
Xbit_r85_c54 bl[54] br[54] wl[85] vdd gnd cell_6t
Xbit_r86_c54 bl[54] br[54] wl[86] vdd gnd cell_6t
Xbit_r87_c54 bl[54] br[54] wl[87] vdd gnd cell_6t
Xbit_r88_c54 bl[54] br[54] wl[88] vdd gnd cell_6t
Xbit_r89_c54 bl[54] br[54] wl[89] vdd gnd cell_6t
Xbit_r90_c54 bl[54] br[54] wl[90] vdd gnd cell_6t
Xbit_r91_c54 bl[54] br[54] wl[91] vdd gnd cell_6t
Xbit_r92_c54 bl[54] br[54] wl[92] vdd gnd cell_6t
Xbit_r93_c54 bl[54] br[54] wl[93] vdd gnd cell_6t
Xbit_r94_c54 bl[54] br[54] wl[94] vdd gnd cell_6t
Xbit_r95_c54 bl[54] br[54] wl[95] vdd gnd cell_6t
Xbit_r96_c54 bl[54] br[54] wl[96] vdd gnd cell_6t
Xbit_r97_c54 bl[54] br[54] wl[97] vdd gnd cell_6t
Xbit_r98_c54 bl[54] br[54] wl[98] vdd gnd cell_6t
Xbit_r99_c54 bl[54] br[54] wl[99] vdd gnd cell_6t
Xbit_r100_c54 bl[54] br[54] wl[100] vdd gnd cell_6t
Xbit_r101_c54 bl[54] br[54] wl[101] vdd gnd cell_6t
Xbit_r102_c54 bl[54] br[54] wl[102] vdd gnd cell_6t
Xbit_r103_c54 bl[54] br[54] wl[103] vdd gnd cell_6t
Xbit_r104_c54 bl[54] br[54] wl[104] vdd gnd cell_6t
Xbit_r105_c54 bl[54] br[54] wl[105] vdd gnd cell_6t
Xbit_r106_c54 bl[54] br[54] wl[106] vdd gnd cell_6t
Xbit_r107_c54 bl[54] br[54] wl[107] vdd gnd cell_6t
Xbit_r108_c54 bl[54] br[54] wl[108] vdd gnd cell_6t
Xbit_r109_c54 bl[54] br[54] wl[109] vdd gnd cell_6t
Xbit_r110_c54 bl[54] br[54] wl[110] vdd gnd cell_6t
Xbit_r111_c54 bl[54] br[54] wl[111] vdd gnd cell_6t
Xbit_r112_c54 bl[54] br[54] wl[112] vdd gnd cell_6t
Xbit_r113_c54 bl[54] br[54] wl[113] vdd gnd cell_6t
Xbit_r114_c54 bl[54] br[54] wl[114] vdd gnd cell_6t
Xbit_r115_c54 bl[54] br[54] wl[115] vdd gnd cell_6t
Xbit_r116_c54 bl[54] br[54] wl[116] vdd gnd cell_6t
Xbit_r117_c54 bl[54] br[54] wl[117] vdd gnd cell_6t
Xbit_r118_c54 bl[54] br[54] wl[118] vdd gnd cell_6t
Xbit_r119_c54 bl[54] br[54] wl[119] vdd gnd cell_6t
Xbit_r120_c54 bl[54] br[54] wl[120] vdd gnd cell_6t
Xbit_r121_c54 bl[54] br[54] wl[121] vdd gnd cell_6t
Xbit_r122_c54 bl[54] br[54] wl[122] vdd gnd cell_6t
Xbit_r123_c54 bl[54] br[54] wl[123] vdd gnd cell_6t
Xbit_r124_c54 bl[54] br[54] wl[124] vdd gnd cell_6t
Xbit_r125_c54 bl[54] br[54] wl[125] vdd gnd cell_6t
Xbit_r126_c54 bl[54] br[54] wl[126] vdd gnd cell_6t
Xbit_r127_c54 bl[54] br[54] wl[127] vdd gnd cell_6t
Xbit_r128_c54 bl[54] br[54] wl[128] vdd gnd cell_6t
Xbit_r129_c54 bl[54] br[54] wl[129] vdd gnd cell_6t
Xbit_r130_c54 bl[54] br[54] wl[130] vdd gnd cell_6t
Xbit_r131_c54 bl[54] br[54] wl[131] vdd gnd cell_6t
Xbit_r132_c54 bl[54] br[54] wl[132] vdd gnd cell_6t
Xbit_r133_c54 bl[54] br[54] wl[133] vdd gnd cell_6t
Xbit_r134_c54 bl[54] br[54] wl[134] vdd gnd cell_6t
Xbit_r135_c54 bl[54] br[54] wl[135] vdd gnd cell_6t
Xbit_r136_c54 bl[54] br[54] wl[136] vdd gnd cell_6t
Xbit_r137_c54 bl[54] br[54] wl[137] vdd gnd cell_6t
Xbit_r138_c54 bl[54] br[54] wl[138] vdd gnd cell_6t
Xbit_r139_c54 bl[54] br[54] wl[139] vdd gnd cell_6t
Xbit_r140_c54 bl[54] br[54] wl[140] vdd gnd cell_6t
Xbit_r141_c54 bl[54] br[54] wl[141] vdd gnd cell_6t
Xbit_r142_c54 bl[54] br[54] wl[142] vdd gnd cell_6t
Xbit_r143_c54 bl[54] br[54] wl[143] vdd gnd cell_6t
Xbit_r144_c54 bl[54] br[54] wl[144] vdd gnd cell_6t
Xbit_r145_c54 bl[54] br[54] wl[145] vdd gnd cell_6t
Xbit_r146_c54 bl[54] br[54] wl[146] vdd gnd cell_6t
Xbit_r147_c54 bl[54] br[54] wl[147] vdd gnd cell_6t
Xbit_r148_c54 bl[54] br[54] wl[148] vdd gnd cell_6t
Xbit_r149_c54 bl[54] br[54] wl[149] vdd gnd cell_6t
Xbit_r150_c54 bl[54] br[54] wl[150] vdd gnd cell_6t
Xbit_r151_c54 bl[54] br[54] wl[151] vdd gnd cell_6t
Xbit_r152_c54 bl[54] br[54] wl[152] vdd gnd cell_6t
Xbit_r153_c54 bl[54] br[54] wl[153] vdd gnd cell_6t
Xbit_r154_c54 bl[54] br[54] wl[154] vdd gnd cell_6t
Xbit_r155_c54 bl[54] br[54] wl[155] vdd gnd cell_6t
Xbit_r156_c54 bl[54] br[54] wl[156] vdd gnd cell_6t
Xbit_r157_c54 bl[54] br[54] wl[157] vdd gnd cell_6t
Xbit_r158_c54 bl[54] br[54] wl[158] vdd gnd cell_6t
Xbit_r159_c54 bl[54] br[54] wl[159] vdd gnd cell_6t
Xbit_r160_c54 bl[54] br[54] wl[160] vdd gnd cell_6t
Xbit_r161_c54 bl[54] br[54] wl[161] vdd gnd cell_6t
Xbit_r162_c54 bl[54] br[54] wl[162] vdd gnd cell_6t
Xbit_r163_c54 bl[54] br[54] wl[163] vdd gnd cell_6t
Xbit_r164_c54 bl[54] br[54] wl[164] vdd gnd cell_6t
Xbit_r165_c54 bl[54] br[54] wl[165] vdd gnd cell_6t
Xbit_r166_c54 bl[54] br[54] wl[166] vdd gnd cell_6t
Xbit_r167_c54 bl[54] br[54] wl[167] vdd gnd cell_6t
Xbit_r168_c54 bl[54] br[54] wl[168] vdd gnd cell_6t
Xbit_r169_c54 bl[54] br[54] wl[169] vdd gnd cell_6t
Xbit_r170_c54 bl[54] br[54] wl[170] vdd gnd cell_6t
Xbit_r171_c54 bl[54] br[54] wl[171] vdd gnd cell_6t
Xbit_r172_c54 bl[54] br[54] wl[172] vdd gnd cell_6t
Xbit_r173_c54 bl[54] br[54] wl[173] vdd gnd cell_6t
Xbit_r174_c54 bl[54] br[54] wl[174] vdd gnd cell_6t
Xbit_r175_c54 bl[54] br[54] wl[175] vdd gnd cell_6t
Xbit_r176_c54 bl[54] br[54] wl[176] vdd gnd cell_6t
Xbit_r177_c54 bl[54] br[54] wl[177] vdd gnd cell_6t
Xbit_r178_c54 bl[54] br[54] wl[178] vdd gnd cell_6t
Xbit_r179_c54 bl[54] br[54] wl[179] vdd gnd cell_6t
Xbit_r180_c54 bl[54] br[54] wl[180] vdd gnd cell_6t
Xbit_r181_c54 bl[54] br[54] wl[181] vdd gnd cell_6t
Xbit_r182_c54 bl[54] br[54] wl[182] vdd gnd cell_6t
Xbit_r183_c54 bl[54] br[54] wl[183] vdd gnd cell_6t
Xbit_r184_c54 bl[54] br[54] wl[184] vdd gnd cell_6t
Xbit_r185_c54 bl[54] br[54] wl[185] vdd gnd cell_6t
Xbit_r186_c54 bl[54] br[54] wl[186] vdd gnd cell_6t
Xbit_r187_c54 bl[54] br[54] wl[187] vdd gnd cell_6t
Xbit_r188_c54 bl[54] br[54] wl[188] vdd gnd cell_6t
Xbit_r189_c54 bl[54] br[54] wl[189] vdd gnd cell_6t
Xbit_r190_c54 bl[54] br[54] wl[190] vdd gnd cell_6t
Xbit_r191_c54 bl[54] br[54] wl[191] vdd gnd cell_6t
Xbit_r192_c54 bl[54] br[54] wl[192] vdd gnd cell_6t
Xbit_r193_c54 bl[54] br[54] wl[193] vdd gnd cell_6t
Xbit_r194_c54 bl[54] br[54] wl[194] vdd gnd cell_6t
Xbit_r195_c54 bl[54] br[54] wl[195] vdd gnd cell_6t
Xbit_r196_c54 bl[54] br[54] wl[196] vdd gnd cell_6t
Xbit_r197_c54 bl[54] br[54] wl[197] vdd gnd cell_6t
Xbit_r198_c54 bl[54] br[54] wl[198] vdd gnd cell_6t
Xbit_r199_c54 bl[54] br[54] wl[199] vdd gnd cell_6t
Xbit_r200_c54 bl[54] br[54] wl[200] vdd gnd cell_6t
Xbit_r201_c54 bl[54] br[54] wl[201] vdd gnd cell_6t
Xbit_r202_c54 bl[54] br[54] wl[202] vdd gnd cell_6t
Xbit_r203_c54 bl[54] br[54] wl[203] vdd gnd cell_6t
Xbit_r204_c54 bl[54] br[54] wl[204] vdd gnd cell_6t
Xbit_r205_c54 bl[54] br[54] wl[205] vdd gnd cell_6t
Xbit_r206_c54 bl[54] br[54] wl[206] vdd gnd cell_6t
Xbit_r207_c54 bl[54] br[54] wl[207] vdd gnd cell_6t
Xbit_r208_c54 bl[54] br[54] wl[208] vdd gnd cell_6t
Xbit_r209_c54 bl[54] br[54] wl[209] vdd gnd cell_6t
Xbit_r210_c54 bl[54] br[54] wl[210] vdd gnd cell_6t
Xbit_r211_c54 bl[54] br[54] wl[211] vdd gnd cell_6t
Xbit_r212_c54 bl[54] br[54] wl[212] vdd gnd cell_6t
Xbit_r213_c54 bl[54] br[54] wl[213] vdd gnd cell_6t
Xbit_r214_c54 bl[54] br[54] wl[214] vdd gnd cell_6t
Xbit_r215_c54 bl[54] br[54] wl[215] vdd gnd cell_6t
Xbit_r216_c54 bl[54] br[54] wl[216] vdd gnd cell_6t
Xbit_r217_c54 bl[54] br[54] wl[217] vdd gnd cell_6t
Xbit_r218_c54 bl[54] br[54] wl[218] vdd gnd cell_6t
Xbit_r219_c54 bl[54] br[54] wl[219] vdd gnd cell_6t
Xbit_r220_c54 bl[54] br[54] wl[220] vdd gnd cell_6t
Xbit_r221_c54 bl[54] br[54] wl[221] vdd gnd cell_6t
Xbit_r222_c54 bl[54] br[54] wl[222] vdd gnd cell_6t
Xbit_r223_c54 bl[54] br[54] wl[223] vdd gnd cell_6t
Xbit_r224_c54 bl[54] br[54] wl[224] vdd gnd cell_6t
Xbit_r225_c54 bl[54] br[54] wl[225] vdd gnd cell_6t
Xbit_r226_c54 bl[54] br[54] wl[226] vdd gnd cell_6t
Xbit_r227_c54 bl[54] br[54] wl[227] vdd gnd cell_6t
Xbit_r228_c54 bl[54] br[54] wl[228] vdd gnd cell_6t
Xbit_r229_c54 bl[54] br[54] wl[229] vdd gnd cell_6t
Xbit_r230_c54 bl[54] br[54] wl[230] vdd gnd cell_6t
Xbit_r231_c54 bl[54] br[54] wl[231] vdd gnd cell_6t
Xbit_r232_c54 bl[54] br[54] wl[232] vdd gnd cell_6t
Xbit_r233_c54 bl[54] br[54] wl[233] vdd gnd cell_6t
Xbit_r234_c54 bl[54] br[54] wl[234] vdd gnd cell_6t
Xbit_r235_c54 bl[54] br[54] wl[235] vdd gnd cell_6t
Xbit_r236_c54 bl[54] br[54] wl[236] vdd gnd cell_6t
Xbit_r237_c54 bl[54] br[54] wl[237] vdd gnd cell_6t
Xbit_r238_c54 bl[54] br[54] wl[238] vdd gnd cell_6t
Xbit_r239_c54 bl[54] br[54] wl[239] vdd gnd cell_6t
Xbit_r240_c54 bl[54] br[54] wl[240] vdd gnd cell_6t
Xbit_r241_c54 bl[54] br[54] wl[241] vdd gnd cell_6t
Xbit_r242_c54 bl[54] br[54] wl[242] vdd gnd cell_6t
Xbit_r243_c54 bl[54] br[54] wl[243] vdd gnd cell_6t
Xbit_r244_c54 bl[54] br[54] wl[244] vdd gnd cell_6t
Xbit_r245_c54 bl[54] br[54] wl[245] vdd gnd cell_6t
Xbit_r246_c54 bl[54] br[54] wl[246] vdd gnd cell_6t
Xbit_r247_c54 bl[54] br[54] wl[247] vdd gnd cell_6t
Xbit_r248_c54 bl[54] br[54] wl[248] vdd gnd cell_6t
Xbit_r249_c54 bl[54] br[54] wl[249] vdd gnd cell_6t
Xbit_r250_c54 bl[54] br[54] wl[250] vdd gnd cell_6t
Xbit_r251_c54 bl[54] br[54] wl[251] vdd gnd cell_6t
Xbit_r252_c54 bl[54] br[54] wl[252] vdd gnd cell_6t
Xbit_r253_c54 bl[54] br[54] wl[253] vdd gnd cell_6t
Xbit_r254_c54 bl[54] br[54] wl[254] vdd gnd cell_6t
Xbit_r255_c54 bl[54] br[54] wl[255] vdd gnd cell_6t
Xbit_r0_c55 bl[55] br[55] wl[0] vdd gnd cell_6t
Xbit_r1_c55 bl[55] br[55] wl[1] vdd gnd cell_6t
Xbit_r2_c55 bl[55] br[55] wl[2] vdd gnd cell_6t
Xbit_r3_c55 bl[55] br[55] wl[3] vdd gnd cell_6t
Xbit_r4_c55 bl[55] br[55] wl[4] vdd gnd cell_6t
Xbit_r5_c55 bl[55] br[55] wl[5] vdd gnd cell_6t
Xbit_r6_c55 bl[55] br[55] wl[6] vdd gnd cell_6t
Xbit_r7_c55 bl[55] br[55] wl[7] vdd gnd cell_6t
Xbit_r8_c55 bl[55] br[55] wl[8] vdd gnd cell_6t
Xbit_r9_c55 bl[55] br[55] wl[9] vdd gnd cell_6t
Xbit_r10_c55 bl[55] br[55] wl[10] vdd gnd cell_6t
Xbit_r11_c55 bl[55] br[55] wl[11] vdd gnd cell_6t
Xbit_r12_c55 bl[55] br[55] wl[12] vdd gnd cell_6t
Xbit_r13_c55 bl[55] br[55] wl[13] vdd gnd cell_6t
Xbit_r14_c55 bl[55] br[55] wl[14] vdd gnd cell_6t
Xbit_r15_c55 bl[55] br[55] wl[15] vdd gnd cell_6t
Xbit_r16_c55 bl[55] br[55] wl[16] vdd gnd cell_6t
Xbit_r17_c55 bl[55] br[55] wl[17] vdd gnd cell_6t
Xbit_r18_c55 bl[55] br[55] wl[18] vdd gnd cell_6t
Xbit_r19_c55 bl[55] br[55] wl[19] vdd gnd cell_6t
Xbit_r20_c55 bl[55] br[55] wl[20] vdd gnd cell_6t
Xbit_r21_c55 bl[55] br[55] wl[21] vdd gnd cell_6t
Xbit_r22_c55 bl[55] br[55] wl[22] vdd gnd cell_6t
Xbit_r23_c55 bl[55] br[55] wl[23] vdd gnd cell_6t
Xbit_r24_c55 bl[55] br[55] wl[24] vdd gnd cell_6t
Xbit_r25_c55 bl[55] br[55] wl[25] vdd gnd cell_6t
Xbit_r26_c55 bl[55] br[55] wl[26] vdd gnd cell_6t
Xbit_r27_c55 bl[55] br[55] wl[27] vdd gnd cell_6t
Xbit_r28_c55 bl[55] br[55] wl[28] vdd gnd cell_6t
Xbit_r29_c55 bl[55] br[55] wl[29] vdd gnd cell_6t
Xbit_r30_c55 bl[55] br[55] wl[30] vdd gnd cell_6t
Xbit_r31_c55 bl[55] br[55] wl[31] vdd gnd cell_6t
Xbit_r32_c55 bl[55] br[55] wl[32] vdd gnd cell_6t
Xbit_r33_c55 bl[55] br[55] wl[33] vdd gnd cell_6t
Xbit_r34_c55 bl[55] br[55] wl[34] vdd gnd cell_6t
Xbit_r35_c55 bl[55] br[55] wl[35] vdd gnd cell_6t
Xbit_r36_c55 bl[55] br[55] wl[36] vdd gnd cell_6t
Xbit_r37_c55 bl[55] br[55] wl[37] vdd gnd cell_6t
Xbit_r38_c55 bl[55] br[55] wl[38] vdd gnd cell_6t
Xbit_r39_c55 bl[55] br[55] wl[39] vdd gnd cell_6t
Xbit_r40_c55 bl[55] br[55] wl[40] vdd gnd cell_6t
Xbit_r41_c55 bl[55] br[55] wl[41] vdd gnd cell_6t
Xbit_r42_c55 bl[55] br[55] wl[42] vdd gnd cell_6t
Xbit_r43_c55 bl[55] br[55] wl[43] vdd gnd cell_6t
Xbit_r44_c55 bl[55] br[55] wl[44] vdd gnd cell_6t
Xbit_r45_c55 bl[55] br[55] wl[45] vdd gnd cell_6t
Xbit_r46_c55 bl[55] br[55] wl[46] vdd gnd cell_6t
Xbit_r47_c55 bl[55] br[55] wl[47] vdd gnd cell_6t
Xbit_r48_c55 bl[55] br[55] wl[48] vdd gnd cell_6t
Xbit_r49_c55 bl[55] br[55] wl[49] vdd gnd cell_6t
Xbit_r50_c55 bl[55] br[55] wl[50] vdd gnd cell_6t
Xbit_r51_c55 bl[55] br[55] wl[51] vdd gnd cell_6t
Xbit_r52_c55 bl[55] br[55] wl[52] vdd gnd cell_6t
Xbit_r53_c55 bl[55] br[55] wl[53] vdd gnd cell_6t
Xbit_r54_c55 bl[55] br[55] wl[54] vdd gnd cell_6t
Xbit_r55_c55 bl[55] br[55] wl[55] vdd gnd cell_6t
Xbit_r56_c55 bl[55] br[55] wl[56] vdd gnd cell_6t
Xbit_r57_c55 bl[55] br[55] wl[57] vdd gnd cell_6t
Xbit_r58_c55 bl[55] br[55] wl[58] vdd gnd cell_6t
Xbit_r59_c55 bl[55] br[55] wl[59] vdd gnd cell_6t
Xbit_r60_c55 bl[55] br[55] wl[60] vdd gnd cell_6t
Xbit_r61_c55 bl[55] br[55] wl[61] vdd gnd cell_6t
Xbit_r62_c55 bl[55] br[55] wl[62] vdd gnd cell_6t
Xbit_r63_c55 bl[55] br[55] wl[63] vdd gnd cell_6t
Xbit_r64_c55 bl[55] br[55] wl[64] vdd gnd cell_6t
Xbit_r65_c55 bl[55] br[55] wl[65] vdd gnd cell_6t
Xbit_r66_c55 bl[55] br[55] wl[66] vdd gnd cell_6t
Xbit_r67_c55 bl[55] br[55] wl[67] vdd gnd cell_6t
Xbit_r68_c55 bl[55] br[55] wl[68] vdd gnd cell_6t
Xbit_r69_c55 bl[55] br[55] wl[69] vdd gnd cell_6t
Xbit_r70_c55 bl[55] br[55] wl[70] vdd gnd cell_6t
Xbit_r71_c55 bl[55] br[55] wl[71] vdd gnd cell_6t
Xbit_r72_c55 bl[55] br[55] wl[72] vdd gnd cell_6t
Xbit_r73_c55 bl[55] br[55] wl[73] vdd gnd cell_6t
Xbit_r74_c55 bl[55] br[55] wl[74] vdd gnd cell_6t
Xbit_r75_c55 bl[55] br[55] wl[75] vdd gnd cell_6t
Xbit_r76_c55 bl[55] br[55] wl[76] vdd gnd cell_6t
Xbit_r77_c55 bl[55] br[55] wl[77] vdd gnd cell_6t
Xbit_r78_c55 bl[55] br[55] wl[78] vdd gnd cell_6t
Xbit_r79_c55 bl[55] br[55] wl[79] vdd gnd cell_6t
Xbit_r80_c55 bl[55] br[55] wl[80] vdd gnd cell_6t
Xbit_r81_c55 bl[55] br[55] wl[81] vdd gnd cell_6t
Xbit_r82_c55 bl[55] br[55] wl[82] vdd gnd cell_6t
Xbit_r83_c55 bl[55] br[55] wl[83] vdd gnd cell_6t
Xbit_r84_c55 bl[55] br[55] wl[84] vdd gnd cell_6t
Xbit_r85_c55 bl[55] br[55] wl[85] vdd gnd cell_6t
Xbit_r86_c55 bl[55] br[55] wl[86] vdd gnd cell_6t
Xbit_r87_c55 bl[55] br[55] wl[87] vdd gnd cell_6t
Xbit_r88_c55 bl[55] br[55] wl[88] vdd gnd cell_6t
Xbit_r89_c55 bl[55] br[55] wl[89] vdd gnd cell_6t
Xbit_r90_c55 bl[55] br[55] wl[90] vdd gnd cell_6t
Xbit_r91_c55 bl[55] br[55] wl[91] vdd gnd cell_6t
Xbit_r92_c55 bl[55] br[55] wl[92] vdd gnd cell_6t
Xbit_r93_c55 bl[55] br[55] wl[93] vdd gnd cell_6t
Xbit_r94_c55 bl[55] br[55] wl[94] vdd gnd cell_6t
Xbit_r95_c55 bl[55] br[55] wl[95] vdd gnd cell_6t
Xbit_r96_c55 bl[55] br[55] wl[96] vdd gnd cell_6t
Xbit_r97_c55 bl[55] br[55] wl[97] vdd gnd cell_6t
Xbit_r98_c55 bl[55] br[55] wl[98] vdd gnd cell_6t
Xbit_r99_c55 bl[55] br[55] wl[99] vdd gnd cell_6t
Xbit_r100_c55 bl[55] br[55] wl[100] vdd gnd cell_6t
Xbit_r101_c55 bl[55] br[55] wl[101] vdd gnd cell_6t
Xbit_r102_c55 bl[55] br[55] wl[102] vdd gnd cell_6t
Xbit_r103_c55 bl[55] br[55] wl[103] vdd gnd cell_6t
Xbit_r104_c55 bl[55] br[55] wl[104] vdd gnd cell_6t
Xbit_r105_c55 bl[55] br[55] wl[105] vdd gnd cell_6t
Xbit_r106_c55 bl[55] br[55] wl[106] vdd gnd cell_6t
Xbit_r107_c55 bl[55] br[55] wl[107] vdd gnd cell_6t
Xbit_r108_c55 bl[55] br[55] wl[108] vdd gnd cell_6t
Xbit_r109_c55 bl[55] br[55] wl[109] vdd gnd cell_6t
Xbit_r110_c55 bl[55] br[55] wl[110] vdd gnd cell_6t
Xbit_r111_c55 bl[55] br[55] wl[111] vdd gnd cell_6t
Xbit_r112_c55 bl[55] br[55] wl[112] vdd gnd cell_6t
Xbit_r113_c55 bl[55] br[55] wl[113] vdd gnd cell_6t
Xbit_r114_c55 bl[55] br[55] wl[114] vdd gnd cell_6t
Xbit_r115_c55 bl[55] br[55] wl[115] vdd gnd cell_6t
Xbit_r116_c55 bl[55] br[55] wl[116] vdd gnd cell_6t
Xbit_r117_c55 bl[55] br[55] wl[117] vdd gnd cell_6t
Xbit_r118_c55 bl[55] br[55] wl[118] vdd gnd cell_6t
Xbit_r119_c55 bl[55] br[55] wl[119] vdd gnd cell_6t
Xbit_r120_c55 bl[55] br[55] wl[120] vdd gnd cell_6t
Xbit_r121_c55 bl[55] br[55] wl[121] vdd gnd cell_6t
Xbit_r122_c55 bl[55] br[55] wl[122] vdd gnd cell_6t
Xbit_r123_c55 bl[55] br[55] wl[123] vdd gnd cell_6t
Xbit_r124_c55 bl[55] br[55] wl[124] vdd gnd cell_6t
Xbit_r125_c55 bl[55] br[55] wl[125] vdd gnd cell_6t
Xbit_r126_c55 bl[55] br[55] wl[126] vdd gnd cell_6t
Xbit_r127_c55 bl[55] br[55] wl[127] vdd gnd cell_6t
Xbit_r128_c55 bl[55] br[55] wl[128] vdd gnd cell_6t
Xbit_r129_c55 bl[55] br[55] wl[129] vdd gnd cell_6t
Xbit_r130_c55 bl[55] br[55] wl[130] vdd gnd cell_6t
Xbit_r131_c55 bl[55] br[55] wl[131] vdd gnd cell_6t
Xbit_r132_c55 bl[55] br[55] wl[132] vdd gnd cell_6t
Xbit_r133_c55 bl[55] br[55] wl[133] vdd gnd cell_6t
Xbit_r134_c55 bl[55] br[55] wl[134] vdd gnd cell_6t
Xbit_r135_c55 bl[55] br[55] wl[135] vdd gnd cell_6t
Xbit_r136_c55 bl[55] br[55] wl[136] vdd gnd cell_6t
Xbit_r137_c55 bl[55] br[55] wl[137] vdd gnd cell_6t
Xbit_r138_c55 bl[55] br[55] wl[138] vdd gnd cell_6t
Xbit_r139_c55 bl[55] br[55] wl[139] vdd gnd cell_6t
Xbit_r140_c55 bl[55] br[55] wl[140] vdd gnd cell_6t
Xbit_r141_c55 bl[55] br[55] wl[141] vdd gnd cell_6t
Xbit_r142_c55 bl[55] br[55] wl[142] vdd gnd cell_6t
Xbit_r143_c55 bl[55] br[55] wl[143] vdd gnd cell_6t
Xbit_r144_c55 bl[55] br[55] wl[144] vdd gnd cell_6t
Xbit_r145_c55 bl[55] br[55] wl[145] vdd gnd cell_6t
Xbit_r146_c55 bl[55] br[55] wl[146] vdd gnd cell_6t
Xbit_r147_c55 bl[55] br[55] wl[147] vdd gnd cell_6t
Xbit_r148_c55 bl[55] br[55] wl[148] vdd gnd cell_6t
Xbit_r149_c55 bl[55] br[55] wl[149] vdd gnd cell_6t
Xbit_r150_c55 bl[55] br[55] wl[150] vdd gnd cell_6t
Xbit_r151_c55 bl[55] br[55] wl[151] vdd gnd cell_6t
Xbit_r152_c55 bl[55] br[55] wl[152] vdd gnd cell_6t
Xbit_r153_c55 bl[55] br[55] wl[153] vdd gnd cell_6t
Xbit_r154_c55 bl[55] br[55] wl[154] vdd gnd cell_6t
Xbit_r155_c55 bl[55] br[55] wl[155] vdd gnd cell_6t
Xbit_r156_c55 bl[55] br[55] wl[156] vdd gnd cell_6t
Xbit_r157_c55 bl[55] br[55] wl[157] vdd gnd cell_6t
Xbit_r158_c55 bl[55] br[55] wl[158] vdd gnd cell_6t
Xbit_r159_c55 bl[55] br[55] wl[159] vdd gnd cell_6t
Xbit_r160_c55 bl[55] br[55] wl[160] vdd gnd cell_6t
Xbit_r161_c55 bl[55] br[55] wl[161] vdd gnd cell_6t
Xbit_r162_c55 bl[55] br[55] wl[162] vdd gnd cell_6t
Xbit_r163_c55 bl[55] br[55] wl[163] vdd gnd cell_6t
Xbit_r164_c55 bl[55] br[55] wl[164] vdd gnd cell_6t
Xbit_r165_c55 bl[55] br[55] wl[165] vdd gnd cell_6t
Xbit_r166_c55 bl[55] br[55] wl[166] vdd gnd cell_6t
Xbit_r167_c55 bl[55] br[55] wl[167] vdd gnd cell_6t
Xbit_r168_c55 bl[55] br[55] wl[168] vdd gnd cell_6t
Xbit_r169_c55 bl[55] br[55] wl[169] vdd gnd cell_6t
Xbit_r170_c55 bl[55] br[55] wl[170] vdd gnd cell_6t
Xbit_r171_c55 bl[55] br[55] wl[171] vdd gnd cell_6t
Xbit_r172_c55 bl[55] br[55] wl[172] vdd gnd cell_6t
Xbit_r173_c55 bl[55] br[55] wl[173] vdd gnd cell_6t
Xbit_r174_c55 bl[55] br[55] wl[174] vdd gnd cell_6t
Xbit_r175_c55 bl[55] br[55] wl[175] vdd gnd cell_6t
Xbit_r176_c55 bl[55] br[55] wl[176] vdd gnd cell_6t
Xbit_r177_c55 bl[55] br[55] wl[177] vdd gnd cell_6t
Xbit_r178_c55 bl[55] br[55] wl[178] vdd gnd cell_6t
Xbit_r179_c55 bl[55] br[55] wl[179] vdd gnd cell_6t
Xbit_r180_c55 bl[55] br[55] wl[180] vdd gnd cell_6t
Xbit_r181_c55 bl[55] br[55] wl[181] vdd gnd cell_6t
Xbit_r182_c55 bl[55] br[55] wl[182] vdd gnd cell_6t
Xbit_r183_c55 bl[55] br[55] wl[183] vdd gnd cell_6t
Xbit_r184_c55 bl[55] br[55] wl[184] vdd gnd cell_6t
Xbit_r185_c55 bl[55] br[55] wl[185] vdd gnd cell_6t
Xbit_r186_c55 bl[55] br[55] wl[186] vdd gnd cell_6t
Xbit_r187_c55 bl[55] br[55] wl[187] vdd gnd cell_6t
Xbit_r188_c55 bl[55] br[55] wl[188] vdd gnd cell_6t
Xbit_r189_c55 bl[55] br[55] wl[189] vdd gnd cell_6t
Xbit_r190_c55 bl[55] br[55] wl[190] vdd gnd cell_6t
Xbit_r191_c55 bl[55] br[55] wl[191] vdd gnd cell_6t
Xbit_r192_c55 bl[55] br[55] wl[192] vdd gnd cell_6t
Xbit_r193_c55 bl[55] br[55] wl[193] vdd gnd cell_6t
Xbit_r194_c55 bl[55] br[55] wl[194] vdd gnd cell_6t
Xbit_r195_c55 bl[55] br[55] wl[195] vdd gnd cell_6t
Xbit_r196_c55 bl[55] br[55] wl[196] vdd gnd cell_6t
Xbit_r197_c55 bl[55] br[55] wl[197] vdd gnd cell_6t
Xbit_r198_c55 bl[55] br[55] wl[198] vdd gnd cell_6t
Xbit_r199_c55 bl[55] br[55] wl[199] vdd gnd cell_6t
Xbit_r200_c55 bl[55] br[55] wl[200] vdd gnd cell_6t
Xbit_r201_c55 bl[55] br[55] wl[201] vdd gnd cell_6t
Xbit_r202_c55 bl[55] br[55] wl[202] vdd gnd cell_6t
Xbit_r203_c55 bl[55] br[55] wl[203] vdd gnd cell_6t
Xbit_r204_c55 bl[55] br[55] wl[204] vdd gnd cell_6t
Xbit_r205_c55 bl[55] br[55] wl[205] vdd gnd cell_6t
Xbit_r206_c55 bl[55] br[55] wl[206] vdd gnd cell_6t
Xbit_r207_c55 bl[55] br[55] wl[207] vdd gnd cell_6t
Xbit_r208_c55 bl[55] br[55] wl[208] vdd gnd cell_6t
Xbit_r209_c55 bl[55] br[55] wl[209] vdd gnd cell_6t
Xbit_r210_c55 bl[55] br[55] wl[210] vdd gnd cell_6t
Xbit_r211_c55 bl[55] br[55] wl[211] vdd gnd cell_6t
Xbit_r212_c55 bl[55] br[55] wl[212] vdd gnd cell_6t
Xbit_r213_c55 bl[55] br[55] wl[213] vdd gnd cell_6t
Xbit_r214_c55 bl[55] br[55] wl[214] vdd gnd cell_6t
Xbit_r215_c55 bl[55] br[55] wl[215] vdd gnd cell_6t
Xbit_r216_c55 bl[55] br[55] wl[216] vdd gnd cell_6t
Xbit_r217_c55 bl[55] br[55] wl[217] vdd gnd cell_6t
Xbit_r218_c55 bl[55] br[55] wl[218] vdd gnd cell_6t
Xbit_r219_c55 bl[55] br[55] wl[219] vdd gnd cell_6t
Xbit_r220_c55 bl[55] br[55] wl[220] vdd gnd cell_6t
Xbit_r221_c55 bl[55] br[55] wl[221] vdd gnd cell_6t
Xbit_r222_c55 bl[55] br[55] wl[222] vdd gnd cell_6t
Xbit_r223_c55 bl[55] br[55] wl[223] vdd gnd cell_6t
Xbit_r224_c55 bl[55] br[55] wl[224] vdd gnd cell_6t
Xbit_r225_c55 bl[55] br[55] wl[225] vdd gnd cell_6t
Xbit_r226_c55 bl[55] br[55] wl[226] vdd gnd cell_6t
Xbit_r227_c55 bl[55] br[55] wl[227] vdd gnd cell_6t
Xbit_r228_c55 bl[55] br[55] wl[228] vdd gnd cell_6t
Xbit_r229_c55 bl[55] br[55] wl[229] vdd gnd cell_6t
Xbit_r230_c55 bl[55] br[55] wl[230] vdd gnd cell_6t
Xbit_r231_c55 bl[55] br[55] wl[231] vdd gnd cell_6t
Xbit_r232_c55 bl[55] br[55] wl[232] vdd gnd cell_6t
Xbit_r233_c55 bl[55] br[55] wl[233] vdd gnd cell_6t
Xbit_r234_c55 bl[55] br[55] wl[234] vdd gnd cell_6t
Xbit_r235_c55 bl[55] br[55] wl[235] vdd gnd cell_6t
Xbit_r236_c55 bl[55] br[55] wl[236] vdd gnd cell_6t
Xbit_r237_c55 bl[55] br[55] wl[237] vdd gnd cell_6t
Xbit_r238_c55 bl[55] br[55] wl[238] vdd gnd cell_6t
Xbit_r239_c55 bl[55] br[55] wl[239] vdd gnd cell_6t
Xbit_r240_c55 bl[55] br[55] wl[240] vdd gnd cell_6t
Xbit_r241_c55 bl[55] br[55] wl[241] vdd gnd cell_6t
Xbit_r242_c55 bl[55] br[55] wl[242] vdd gnd cell_6t
Xbit_r243_c55 bl[55] br[55] wl[243] vdd gnd cell_6t
Xbit_r244_c55 bl[55] br[55] wl[244] vdd gnd cell_6t
Xbit_r245_c55 bl[55] br[55] wl[245] vdd gnd cell_6t
Xbit_r246_c55 bl[55] br[55] wl[246] vdd gnd cell_6t
Xbit_r247_c55 bl[55] br[55] wl[247] vdd gnd cell_6t
Xbit_r248_c55 bl[55] br[55] wl[248] vdd gnd cell_6t
Xbit_r249_c55 bl[55] br[55] wl[249] vdd gnd cell_6t
Xbit_r250_c55 bl[55] br[55] wl[250] vdd gnd cell_6t
Xbit_r251_c55 bl[55] br[55] wl[251] vdd gnd cell_6t
Xbit_r252_c55 bl[55] br[55] wl[252] vdd gnd cell_6t
Xbit_r253_c55 bl[55] br[55] wl[253] vdd gnd cell_6t
Xbit_r254_c55 bl[55] br[55] wl[254] vdd gnd cell_6t
Xbit_r255_c55 bl[55] br[55] wl[255] vdd gnd cell_6t
Xbit_r0_c56 bl[56] br[56] wl[0] vdd gnd cell_6t
Xbit_r1_c56 bl[56] br[56] wl[1] vdd gnd cell_6t
Xbit_r2_c56 bl[56] br[56] wl[2] vdd gnd cell_6t
Xbit_r3_c56 bl[56] br[56] wl[3] vdd gnd cell_6t
Xbit_r4_c56 bl[56] br[56] wl[4] vdd gnd cell_6t
Xbit_r5_c56 bl[56] br[56] wl[5] vdd gnd cell_6t
Xbit_r6_c56 bl[56] br[56] wl[6] vdd gnd cell_6t
Xbit_r7_c56 bl[56] br[56] wl[7] vdd gnd cell_6t
Xbit_r8_c56 bl[56] br[56] wl[8] vdd gnd cell_6t
Xbit_r9_c56 bl[56] br[56] wl[9] vdd gnd cell_6t
Xbit_r10_c56 bl[56] br[56] wl[10] vdd gnd cell_6t
Xbit_r11_c56 bl[56] br[56] wl[11] vdd gnd cell_6t
Xbit_r12_c56 bl[56] br[56] wl[12] vdd gnd cell_6t
Xbit_r13_c56 bl[56] br[56] wl[13] vdd gnd cell_6t
Xbit_r14_c56 bl[56] br[56] wl[14] vdd gnd cell_6t
Xbit_r15_c56 bl[56] br[56] wl[15] vdd gnd cell_6t
Xbit_r16_c56 bl[56] br[56] wl[16] vdd gnd cell_6t
Xbit_r17_c56 bl[56] br[56] wl[17] vdd gnd cell_6t
Xbit_r18_c56 bl[56] br[56] wl[18] vdd gnd cell_6t
Xbit_r19_c56 bl[56] br[56] wl[19] vdd gnd cell_6t
Xbit_r20_c56 bl[56] br[56] wl[20] vdd gnd cell_6t
Xbit_r21_c56 bl[56] br[56] wl[21] vdd gnd cell_6t
Xbit_r22_c56 bl[56] br[56] wl[22] vdd gnd cell_6t
Xbit_r23_c56 bl[56] br[56] wl[23] vdd gnd cell_6t
Xbit_r24_c56 bl[56] br[56] wl[24] vdd gnd cell_6t
Xbit_r25_c56 bl[56] br[56] wl[25] vdd gnd cell_6t
Xbit_r26_c56 bl[56] br[56] wl[26] vdd gnd cell_6t
Xbit_r27_c56 bl[56] br[56] wl[27] vdd gnd cell_6t
Xbit_r28_c56 bl[56] br[56] wl[28] vdd gnd cell_6t
Xbit_r29_c56 bl[56] br[56] wl[29] vdd gnd cell_6t
Xbit_r30_c56 bl[56] br[56] wl[30] vdd gnd cell_6t
Xbit_r31_c56 bl[56] br[56] wl[31] vdd gnd cell_6t
Xbit_r32_c56 bl[56] br[56] wl[32] vdd gnd cell_6t
Xbit_r33_c56 bl[56] br[56] wl[33] vdd gnd cell_6t
Xbit_r34_c56 bl[56] br[56] wl[34] vdd gnd cell_6t
Xbit_r35_c56 bl[56] br[56] wl[35] vdd gnd cell_6t
Xbit_r36_c56 bl[56] br[56] wl[36] vdd gnd cell_6t
Xbit_r37_c56 bl[56] br[56] wl[37] vdd gnd cell_6t
Xbit_r38_c56 bl[56] br[56] wl[38] vdd gnd cell_6t
Xbit_r39_c56 bl[56] br[56] wl[39] vdd gnd cell_6t
Xbit_r40_c56 bl[56] br[56] wl[40] vdd gnd cell_6t
Xbit_r41_c56 bl[56] br[56] wl[41] vdd gnd cell_6t
Xbit_r42_c56 bl[56] br[56] wl[42] vdd gnd cell_6t
Xbit_r43_c56 bl[56] br[56] wl[43] vdd gnd cell_6t
Xbit_r44_c56 bl[56] br[56] wl[44] vdd gnd cell_6t
Xbit_r45_c56 bl[56] br[56] wl[45] vdd gnd cell_6t
Xbit_r46_c56 bl[56] br[56] wl[46] vdd gnd cell_6t
Xbit_r47_c56 bl[56] br[56] wl[47] vdd gnd cell_6t
Xbit_r48_c56 bl[56] br[56] wl[48] vdd gnd cell_6t
Xbit_r49_c56 bl[56] br[56] wl[49] vdd gnd cell_6t
Xbit_r50_c56 bl[56] br[56] wl[50] vdd gnd cell_6t
Xbit_r51_c56 bl[56] br[56] wl[51] vdd gnd cell_6t
Xbit_r52_c56 bl[56] br[56] wl[52] vdd gnd cell_6t
Xbit_r53_c56 bl[56] br[56] wl[53] vdd gnd cell_6t
Xbit_r54_c56 bl[56] br[56] wl[54] vdd gnd cell_6t
Xbit_r55_c56 bl[56] br[56] wl[55] vdd gnd cell_6t
Xbit_r56_c56 bl[56] br[56] wl[56] vdd gnd cell_6t
Xbit_r57_c56 bl[56] br[56] wl[57] vdd gnd cell_6t
Xbit_r58_c56 bl[56] br[56] wl[58] vdd gnd cell_6t
Xbit_r59_c56 bl[56] br[56] wl[59] vdd gnd cell_6t
Xbit_r60_c56 bl[56] br[56] wl[60] vdd gnd cell_6t
Xbit_r61_c56 bl[56] br[56] wl[61] vdd gnd cell_6t
Xbit_r62_c56 bl[56] br[56] wl[62] vdd gnd cell_6t
Xbit_r63_c56 bl[56] br[56] wl[63] vdd gnd cell_6t
Xbit_r64_c56 bl[56] br[56] wl[64] vdd gnd cell_6t
Xbit_r65_c56 bl[56] br[56] wl[65] vdd gnd cell_6t
Xbit_r66_c56 bl[56] br[56] wl[66] vdd gnd cell_6t
Xbit_r67_c56 bl[56] br[56] wl[67] vdd gnd cell_6t
Xbit_r68_c56 bl[56] br[56] wl[68] vdd gnd cell_6t
Xbit_r69_c56 bl[56] br[56] wl[69] vdd gnd cell_6t
Xbit_r70_c56 bl[56] br[56] wl[70] vdd gnd cell_6t
Xbit_r71_c56 bl[56] br[56] wl[71] vdd gnd cell_6t
Xbit_r72_c56 bl[56] br[56] wl[72] vdd gnd cell_6t
Xbit_r73_c56 bl[56] br[56] wl[73] vdd gnd cell_6t
Xbit_r74_c56 bl[56] br[56] wl[74] vdd gnd cell_6t
Xbit_r75_c56 bl[56] br[56] wl[75] vdd gnd cell_6t
Xbit_r76_c56 bl[56] br[56] wl[76] vdd gnd cell_6t
Xbit_r77_c56 bl[56] br[56] wl[77] vdd gnd cell_6t
Xbit_r78_c56 bl[56] br[56] wl[78] vdd gnd cell_6t
Xbit_r79_c56 bl[56] br[56] wl[79] vdd gnd cell_6t
Xbit_r80_c56 bl[56] br[56] wl[80] vdd gnd cell_6t
Xbit_r81_c56 bl[56] br[56] wl[81] vdd gnd cell_6t
Xbit_r82_c56 bl[56] br[56] wl[82] vdd gnd cell_6t
Xbit_r83_c56 bl[56] br[56] wl[83] vdd gnd cell_6t
Xbit_r84_c56 bl[56] br[56] wl[84] vdd gnd cell_6t
Xbit_r85_c56 bl[56] br[56] wl[85] vdd gnd cell_6t
Xbit_r86_c56 bl[56] br[56] wl[86] vdd gnd cell_6t
Xbit_r87_c56 bl[56] br[56] wl[87] vdd gnd cell_6t
Xbit_r88_c56 bl[56] br[56] wl[88] vdd gnd cell_6t
Xbit_r89_c56 bl[56] br[56] wl[89] vdd gnd cell_6t
Xbit_r90_c56 bl[56] br[56] wl[90] vdd gnd cell_6t
Xbit_r91_c56 bl[56] br[56] wl[91] vdd gnd cell_6t
Xbit_r92_c56 bl[56] br[56] wl[92] vdd gnd cell_6t
Xbit_r93_c56 bl[56] br[56] wl[93] vdd gnd cell_6t
Xbit_r94_c56 bl[56] br[56] wl[94] vdd gnd cell_6t
Xbit_r95_c56 bl[56] br[56] wl[95] vdd gnd cell_6t
Xbit_r96_c56 bl[56] br[56] wl[96] vdd gnd cell_6t
Xbit_r97_c56 bl[56] br[56] wl[97] vdd gnd cell_6t
Xbit_r98_c56 bl[56] br[56] wl[98] vdd gnd cell_6t
Xbit_r99_c56 bl[56] br[56] wl[99] vdd gnd cell_6t
Xbit_r100_c56 bl[56] br[56] wl[100] vdd gnd cell_6t
Xbit_r101_c56 bl[56] br[56] wl[101] vdd gnd cell_6t
Xbit_r102_c56 bl[56] br[56] wl[102] vdd gnd cell_6t
Xbit_r103_c56 bl[56] br[56] wl[103] vdd gnd cell_6t
Xbit_r104_c56 bl[56] br[56] wl[104] vdd gnd cell_6t
Xbit_r105_c56 bl[56] br[56] wl[105] vdd gnd cell_6t
Xbit_r106_c56 bl[56] br[56] wl[106] vdd gnd cell_6t
Xbit_r107_c56 bl[56] br[56] wl[107] vdd gnd cell_6t
Xbit_r108_c56 bl[56] br[56] wl[108] vdd gnd cell_6t
Xbit_r109_c56 bl[56] br[56] wl[109] vdd gnd cell_6t
Xbit_r110_c56 bl[56] br[56] wl[110] vdd gnd cell_6t
Xbit_r111_c56 bl[56] br[56] wl[111] vdd gnd cell_6t
Xbit_r112_c56 bl[56] br[56] wl[112] vdd gnd cell_6t
Xbit_r113_c56 bl[56] br[56] wl[113] vdd gnd cell_6t
Xbit_r114_c56 bl[56] br[56] wl[114] vdd gnd cell_6t
Xbit_r115_c56 bl[56] br[56] wl[115] vdd gnd cell_6t
Xbit_r116_c56 bl[56] br[56] wl[116] vdd gnd cell_6t
Xbit_r117_c56 bl[56] br[56] wl[117] vdd gnd cell_6t
Xbit_r118_c56 bl[56] br[56] wl[118] vdd gnd cell_6t
Xbit_r119_c56 bl[56] br[56] wl[119] vdd gnd cell_6t
Xbit_r120_c56 bl[56] br[56] wl[120] vdd gnd cell_6t
Xbit_r121_c56 bl[56] br[56] wl[121] vdd gnd cell_6t
Xbit_r122_c56 bl[56] br[56] wl[122] vdd gnd cell_6t
Xbit_r123_c56 bl[56] br[56] wl[123] vdd gnd cell_6t
Xbit_r124_c56 bl[56] br[56] wl[124] vdd gnd cell_6t
Xbit_r125_c56 bl[56] br[56] wl[125] vdd gnd cell_6t
Xbit_r126_c56 bl[56] br[56] wl[126] vdd gnd cell_6t
Xbit_r127_c56 bl[56] br[56] wl[127] vdd gnd cell_6t
Xbit_r128_c56 bl[56] br[56] wl[128] vdd gnd cell_6t
Xbit_r129_c56 bl[56] br[56] wl[129] vdd gnd cell_6t
Xbit_r130_c56 bl[56] br[56] wl[130] vdd gnd cell_6t
Xbit_r131_c56 bl[56] br[56] wl[131] vdd gnd cell_6t
Xbit_r132_c56 bl[56] br[56] wl[132] vdd gnd cell_6t
Xbit_r133_c56 bl[56] br[56] wl[133] vdd gnd cell_6t
Xbit_r134_c56 bl[56] br[56] wl[134] vdd gnd cell_6t
Xbit_r135_c56 bl[56] br[56] wl[135] vdd gnd cell_6t
Xbit_r136_c56 bl[56] br[56] wl[136] vdd gnd cell_6t
Xbit_r137_c56 bl[56] br[56] wl[137] vdd gnd cell_6t
Xbit_r138_c56 bl[56] br[56] wl[138] vdd gnd cell_6t
Xbit_r139_c56 bl[56] br[56] wl[139] vdd gnd cell_6t
Xbit_r140_c56 bl[56] br[56] wl[140] vdd gnd cell_6t
Xbit_r141_c56 bl[56] br[56] wl[141] vdd gnd cell_6t
Xbit_r142_c56 bl[56] br[56] wl[142] vdd gnd cell_6t
Xbit_r143_c56 bl[56] br[56] wl[143] vdd gnd cell_6t
Xbit_r144_c56 bl[56] br[56] wl[144] vdd gnd cell_6t
Xbit_r145_c56 bl[56] br[56] wl[145] vdd gnd cell_6t
Xbit_r146_c56 bl[56] br[56] wl[146] vdd gnd cell_6t
Xbit_r147_c56 bl[56] br[56] wl[147] vdd gnd cell_6t
Xbit_r148_c56 bl[56] br[56] wl[148] vdd gnd cell_6t
Xbit_r149_c56 bl[56] br[56] wl[149] vdd gnd cell_6t
Xbit_r150_c56 bl[56] br[56] wl[150] vdd gnd cell_6t
Xbit_r151_c56 bl[56] br[56] wl[151] vdd gnd cell_6t
Xbit_r152_c56 bl[56] br[56] wl[152] vdd gnd cell_6t
Xbit_r153_c56 bl[56] br[56] wl[153] vdd gnd cell_6t
Xbit_r154_c56 bl[56] br[56] wl[154] vdd gnd cell_6t
Xbit_r155_c56 bl[56] br[56] wl[155] vdd gnd cell_6t
Xbit_r156_c56 bl[56] br[56] wl[156] vdd gnd cell_6t
Xbit_r157_c56 bl[56] br[56] wl[157] vdd gnd cell_6t
Xbit_r158_c56 bl[56] br[56] wl[158] vdd gnd cell_6t
Xbit_r159_c56 bl[56] br[56] wl[159] vdd gnd cell_6t
Xbit_r160_c56 bl[56] br[56] wl[160] vdd gnd cell_6t
Xbit_r161_c56 bl[56] br[56] wl[161] vdd gnd cell_6t
Xbit_r162_c56 bl[56] br[56] wl[162] vdd gnd cell_6t
Xbit_r163_c56 bl[56] br[56] wl[163] vdd gnd cell_6t
Xbit_r164_c56 bl[56] br[56] wl[164] vdd gnd cell_6t
Xbit_r165_c56 bl[56] br[56] wl[165] vdd gnd cell_6t
Xbit_r166_c56 bl[56] br[56] wl[166] vdd gnd cell_6t
Xbit_r167_c56 bl[56] br[56] wl[167] vdd gnd cell_6t
Xbit_r168_c56 bl[56] br[56] wl[168] vdd gnd cell_6t
Xbit_r169_c56 bl[56] br[56] wl[169] vdd gnd cell_6t
Xbit_r170_c56 bl[56] br[56] wl[170] vdd gnd cell_6t
Xbit_r171_c56 bl[56] br[56] wl[171] vdd gnd cell_6t
Xbit_r172_c56 bl[56] br[56] wl[172] vdd gnd cell_6t
Xbit_r173_c56 bl[56] br[56] wl[173] vdd gnd cell_6t
Xbit_r174_c56 bl[56] br[56] wl[174] vdd gnd cell_6t
Xbit_r175_c56 bl[56] br[56] wl[175] vdd gnd cell_6t
Xbit_r176_c56 bl[56] br[56] wl[176] vdd gnd cell_6t
Xbit_r177_c56 bl[56] br[56] wl[177] vdd gnd cell_6t
Xbit_r178_c56 bl[56] br[56] wl[178] vdd gnd cell_6t
Xbit_r179_c56 bl[56] br[56] wl[179] vdd gnd cell_6t
Xbit_r180_c56 bl[56] br[56] wl[180] vdd gnd cell_6t
Xbit_r181_c56 bl[56] br[56] wl[181] vdd gnd cell_6t
Xbit_r182_c56 bl[56] br[56] wl[182] vdd gnd cell_6t
Xbit_r183_c56 bl[56] br[56] wl[183] vdd gnd cell_6t
Xbit_r184_c56 bl[56] br[56] wl[184] vdd gnd cell_6t
Xbit_r185_c56 bl[56] br[56] wl[185] vdd gnd cell_6t
Xbit_r186_c56 bl[56] br[56] wl[186] vdd gnd cell_6t
Xbit_r187_c56 bl[56] br[56] wl[187] vdd gnd cell_6t
Xbit_r188_c56 bl[56] br[56] wl[188] vdd gnd cell_6t
Xbit_r189_c56 bl[56] br[56] wl[189] vdd gnd cell_6t
Xbit_r190_c56 bl[56] br[56] wl[190] vdd gnd cell_6t
Xbit_r191_c56 bl[56] br[56] wl[191] vdd gnd cell_6t
Xbit_r192_c56 bl[56] br[56] wl[192] vdd gnd cell_6t
Xbit_r193_c56 bl[56] br[56] wl[193] vdd gnd cell_6t
Xbit_r194_c56 bl[56] br[56] wl[194] vdd gnd cell_6t
Xbit_r195_c56 bl[56] br[56] wl[195] vdd gnd cell_6t
Xbit_r196_c56 bl[56] br[56] wl[196] vdd gnd cell_6t
Xbit_r197_c56 bl[56] br[56] wl[197] vdd gnd cell_6t
Xbit_r198_c56 bl[56] br[56] wl[198] vdd gnd cell_6t
Xbit_r199_c56 bl[56] br[56] wl[199] vdd gnd cell_6t
Xbit_r200_c56 bl[56] br[56] wl[200] vdd gnd cell_6t
Xbit_r201_c56 bl[56] br[56] wl[201] vdd gnd cell_6t
Xbit_r202_c56 bl[56] br[56] wl[202] vdd gnd cell_6t
Xbit_r203_c56 bl[56] br[56] wl[203] vdd gnd cell_6t
Xbit_r204_c56 bl[56] br[56] wl[204] vdd gnd cell_6t
Xbit_r205_c56 bl[56] br[56] wl[205] vdd gnd cell_6t
Xbit_r206_c56 bl[56] br[56] wl[206] vdd gnd cell_6t
Xbit_r207_c56 bl[56] br[56] wl[207] vdd gnd cell_6t
Xbit_r208_c56 bl[56] br[56] wl[208] vdd gnd cell_6t
Xbit_r209_c56 bl[56] br[56] wl[209] vdd gnd cell_6t
Xbit_r210_c56 bl[56] br[56] wl[210] vdd gnd cell_6t
Xbit_r211_c56 bl[56] br[56] wl[211] vdd gnd cell_6t
Xbit_r212_c56 bl[56] br[56] wl[212] vdd gnd cell_6t
Xbit_r213_c56 bl[56] br[56] wl[213] vdd gnd cell_6t
Xbit_r214_c56 bl[56] br[56] wl[214] vdd gnd cell_6t
Xbit_r215_c56 bl[56] br[56] wl[215] vdd gnd cell_6t
Xbit_r216_c56 bl[56] br[56] wl[216] vdd gnd cell_6t
Xbit_r217_c56 bl[56] br[56] wl[217] vdd gnd cell_6t
Xbit_r218_c56 bl[56] br[56] wl[218] vdd gnd cell_6t
Xbit_r219_c56 bl[56] br[56] wl[219] vdd gnd cell_6t
Xbit_r220_c56 bl[56] br[56] wl[220] vdd gnd cell_6t
Xbit_r221_c56 bl[56] br[56] wl[221] vdd gnd cell_6t
Xbit_r222_c56 bl[56] br[56] wl[222] vdd gnd cell_6t
Xbit_r223_c56 bl[56] br[56] wl[223] vdd gnd cell_6t
Xbit_r224_c56 bl[56] br[56] wl[224] vdd gnd cell_6t
Xbit_r225_c56 bl[56] br[56] wl[225] vdd gnd cell_6t
Xbit_r226_c56 bl[56] br[56] wl[226] vdd gnd cell_6t
Xbit_r227_c56 bl[56] br[56] wl[227] vdd gnd cell_6t
Xbit_r228_c56 bl[56] br[56] wl[228] vdd gnd cell_6t
Xbit_r229_c56 bl[56] br[56] wl[229] vdd gnd cell_6t
Xbit_r230_c56 bl[56] br[56] wl[230] vdd gnd cell_6t
Xbit_r231_c56 bl[56] br[56] wl[231] vdd gnd cell_6t
Xbit_r232_c56 bl[56] br[56] wl[232] vdd gnd cell_6t
Xbit_r233_c56 bl[56] br[56] wl[233] vdd gnd cell_6t
Xbit_r234_c56 bl[56] br[56] wl[234] vdd gnd cell_6t
Xbit_r235_c56 bl[56] br[56] wl[235] vdd gnd cell_6t
Xbit_r236_c56 bl[56] br[56] wl[236] vdd gnd cell_6t
Xbit_r237_c56 bl[56] br[56] wl[237] vdd gnd cell_6t
Xbit_r238_c56 bl[56] br[56] wl[238] vdd gnd cell_6t
Xbit_r239_c56 bl[56] br[56] wl[239] vdd gnd cell_6t
Xbit_r240_c56 bl[56] br[56] wl[240] vdd gnd cell_6t
Xbit_r241_c56 bl[56] br[56] wl[241] vdd gnd cell_6t
Xbit_r242_c56 bl[56] br[56] wl[242] vdd gnd cell_6t
Xbit_r243_c56 bl[56] br[56] wl[243] vdd gnd cell_6t
Xbit_r244_c56 bl[56] br[56] wl[244] vdd gnd cell_6t
Xbit_r245_c56 bl[56] br[56] wl[245] vdd gnd cell_6t
Xbit_r246_c56 bl[56] br[56] wl[246] vdd gnd cell_6t
Xbit_r247_c56 bl[56] br[56] wl[247] vdd gnd cell_6t
Xbit_r248_c56 bl[56] br[56] wl[248] vdd gnd cell_6t
Xbit_r249_c56 bl[56] br[56] wl[249] vdd gnd cell_6t
Xbit_r250_c56 bl[56] br[56] wl[250] vdd gnd cell_6t
Xbit_r251_c56 bl[56] br[56] wl[251] vdd gnd cell_6t
Xbit_r252_c56 bl[56] br[56] wl[252] vdd gnd cell_6t
Xbit_r253_c56 bl[56] br[56] wl[253] vdd gnd cell_6t
Xbit_r254_c56 bl[56] br[56] wl[254] vdd gnd cell_6t
Xbit_r255_c56 bl[56] br[56] wl[255] vdd gnd cell_6t
Xbit_r0_c57 bl[57] br[57] wl[0] vdd gnd cell_6t
Xbit_r1_c57 bl[57] br[57] wl[1] vdd gnd cell_6t
Xbit_r2_c57 bl[57] br[57] wl[2] vdd gnd cell_6t
Xbit_r3_c57 bl[57] br[57] wl[3] vdd gnd cell_6t
Xbit_r4_c57 bl[57] br[57] wl[4] vdd gnd cell_6t
Xbit_r5_c57 bl[57] br[57] wl[5] vdd gnd cell_6t
Xbit_r6_c57 bl[57] br[57] wl[6] vdd gnd cell_6t
Xbit_r7_c57 bl[57] br[57] wl[7] vdd gnd cell_6t
Xbit_r8_c57 bl[57] br[57] wl[8] vdd gnd cell_6t
Xbit_r9_c57 bl[57] br[57] wl[9] vdd gnd cell_6t
Xbit_r10_c57 bl[57] br[57] wl[10] vdd gnd cell_6t
Xbit_r11_c57 bl[57] br[57] wl[11] vdd gnd cell_6t
Xbit_r12_c57 bl[57] br[57] wl[12] vdd gnd cell_6t
Xbit_r13_c57 bl[57] br[57] wl[13] vdd gnd cell_6t
Xbit_r14_c57 bl[57] br[57] wl[14] vdd gnd cell_6t
Xbit_r15_c57 bl[57] br[57] wl[15] vdd gnd cell_6t
Xbit_r16_c57 bl[57] br[57] wl[16] vdd gnd cell_6t
Xbit_r17_c57 bl[57] br[57] wl[17] vdd gnd cell_6t
Xbit_r18_c57 bl[57] br[57] wl[18] vdd gnd cell_6t
Xbit_r19_c57 bl[57] br[57] wl[19] vdd gnd cell_6t
Xbit_r20_c57 bl[57] br[57] wl[20] vdd gnd cell_6t
Xbit_r21_c57 bl[57] br[57] wl[21] vdd gnd cell_6t
Xbit_r22_c57 bl[57] br[57] wl[22] vdd gnd cell_6t
Xbit_r23_c57 bl[57] br[57] wl[23] vdd gnd cell_6t
Xbit_r24_c57 bl[57] br[57] wl[24] vdd gnd cell_6t
Xbit_r25_c57 bl[57] br[57] wl[25] vdd gnd cell_6t
Xbit_r26_c57 bl[57] br[57] wl[26] vdd gnd cell_6t
Xbit_r27_c57 bl[57] br[57] wl[27] vdd gnd cell_6t
Xbit_r28_c57 bl[57] br[57] wl[28] vdd gnd cell_6t
Xbit_r29_c57 bl[57] br[57] wl[29] vdd gnd cell_6t
Xbit_r30_c57 bl[57] br[57] wl[30] vdd gnd cell_6t
Xbit_r31_c57 bl[57] br[57] wl[31] vdd gnd cell_6t
Xbit_r32_c57 bl[57] br[57] wl[32] vdd gnd cell_6t
Xbit_r33_c57 bl[57] br[57] wl[33] vdd gnd cell_6t
Xbit_r34_c57 bl[57] br[57] wl[34] vdd gnd cell_6t
Xbit_r35_c57 bl[57] br[57] wl[35] vdd gnd cell_6t
Xbit_r36_c57 bl[57] br[57] wl[36] vdd gnd cell_6t
Xbit_r37_c57 bl[57] br[57] wl[37] vdd gnd cell_6t
Xbit_r38_c57 bl[57] br[57] wl[38] vdd gnd cell_6t
Xbit_r39_c57 bl[57] br[57] wl[39] vdd gnd cell_6t
Xbit_r40_c57 bl[57] br[57] wl[40] vdd gnd cell_6t
Xbit_r41_c57 bl[57] br[57] wl[41] vdd gnd cell_6t
Xbit_r42_c57 bl[57] br[57] wl[42] vdd gnd cell_6t
Xbit_r43_c57 bl[57] br[57] wl[43] vdd gnd cell_6t
Xbit_r44_c57 bl[57] br[57] wl[44] vdd gnd cell_6t
Xbit_r45_c57 bl[57] br[57] wl[45] vdd gnd cell_6t
Xbit_r46_c57 bl[57] br[57] wl[46] vdd gnd cell_6t
Xbit_r47_c57 bl[57] br[57] wl[47] vdd gnd cell_6t
Xbit_r48_c57 bl[57] br[57] wl[48] vdd gnd cell_6t
Xbit_r49_c57 bl[57] br[57] wl[49] vdd gnd cell_6t
Xbit_r50_c57 bl[57] br[57] wl[50] vdd gnd cell_6t
Xbit_r51_c57 bl[57] br[57] wl[51] vdd gnd cell_6t
Xbit_r52_c57 bl[57] br[57] wl[52] vdd gnd cell_6t
Xbit_r53_c57 bl[57] br[57] wl[53] vdd gnd cell_6t
Xbit_r54_c57 bl[57] br[57] wl[54] vdd gnd cell_6t
Xbit_r55_c57 bl[57] br[57] wl[55] vdd gnd cell_6t
Xbit_r56_c57 bl[57] br[57] wl[56] vdd gnd cell_6t
Xbit_r57_c57 bl[57] br[57] wl[57] vdd gnd cell_6t
Xbit_r58_c57 bl[57] br[57] wl[58] vdd gnd cell_6t
Xbit_r59_c57 bl[57] br[57] wl[59] vdd gnd cell_6t
Xbit_r60_c57 bl[57] br[57] wl[60] vdd gnd cell_6t
Xbit_r61_c57 bl[57] br[57] wl[61] vdd gnd cell_6t
Xbit_r62_c57 bl[57] br[57] wl[62] vdd gnd cell_6t
Xbit_r63_c57 bl[57] br[57] wl[63] vdd gnd cell_6t
Xbit_r64_c57 bl[57] br[57] wl[64] vdd gnd cell_6t
Xbit_r65_c57 bl[57] br[57] wl[65] vdd gnd cell_6t
Xbit_r66_c57 bl[57] br[57] wl[66] vdd gnd cell_6t
Xbit_r67_c57 bl[57] br[57] wl[67] vdd gnd cell_6t
Xbit_r68_c57 bl[57] br[57] wl[68] vdd gnd cell_6t
Xbit_r69_c57 bl[57] br[57] wl[69] vdd gnd cell_6t
Xbit_r70_c57 bl[57] br[57] wl[70] vdd gnd cell_6t
Xbit_r71_c57 bl[57] br[57] wl[71] vdd gnd cell_6t
Xbit_r72_c57 bl[57] br[57] wl[72] vdd gnd cell_6t
Xbit_r73_c57 bl[57] br[57] wl[73] vdd gnd cell_6t
Xbit_r74_c57 bl[57] br[57] wl[74] vdd gnd cell_6t
Xbit_r75_c57 bl[57] br[57] wl[75] vdd gnd cell_6t
Xbit_r76_c57 bl[57] br[57] wl[76] vdd gnd cell_6t
Xbit_r77_c57 bl[57] br[57] wl[77] vdd gnd cell_6t
Xbit_r78_c57 bl[57] br[57] wl[78] vdd gnd cell_6t
Xbit_r79_c57 bl[57] br[57] wl[79] vdd gnd cell_6t
Xbit_r80_c57 bl[57] br[57] wl[80] vdd gnd cell_6t
Xbit_r81_c57 bl[57] br[57] wl[81] vdd gnd cell_6t
Xbit_r82_c57 bl[57] br[57] wl[82] vdd gnd cell_6t
Xbit_r83_c57 bl[57] br[57] wl[83] vdd gnd cell_6t
Xbit_r84_c57 bl[57] br[57] wl[84] vdd gnd cell_6t
Xbit_r85_c57 bl[57] br[57] wl[85] vdd gnd cell_6t
Xbit_r86_c57 bl[57] br[57] wl[86] vdd gnd cell_6t
Xbit_r87_c57 bl[57] br[57] wl[87] vdd gnd cell_6t
Xbit_r88_c57 bl[57] br[57] wl[88] vdd gnd cell_6t
Xbit_r89_c57 bl[57] br[57] wl[89] vdd gnd cell_6t
Xbit_r90_c57 bl[57] br[57] wl[90] vdd gnd cell_6t
Xbit_r91_c57 bl[57] br[57] wl[91] vdd gnd cell_6t
Xbit_r92_c57 bl[57] br[57] wl[92] vdd gnd cell_6t
Xbit_r93_c57 bl[57] br[57] wl[93] vdd gnd cell_6t
Xbit_r94_c57 bl[57] br[57] wl[94] vdd gnd cell_6t
Xbit_r95_c57 bl[57] br[57] wl[95] vdd gnd cell_6t
Xbit_r96_c57 bl[57] br[57] wl[96] vdd gnd cell_6t
Xbit_r97_c57 bl[57] br[57] wl[97] vdd gnd cell_6t
Xbit_r98_c57 bl[57] br[57] wl[98] vdd gnd cell_6t
Xbit_r99_c57 bl[57] br[57] wl[99] vdd gnd cell_6t
Xbit_r100_c57 bl[57] br[57] wl[100] vdd gnd cell_6t
Xbit_r101_c57 bl[57] br[57] wl[101] vdd gnd cell_6t
Xbit_r102_c57 bl[57] br[57] wl[102] vdd gnd cell_6t
Xbit_r103_c57 bl[57] br[57] wl[103] vdd gnd cell_6t
Xbit_r104_c57 bl[57] br[57] wl[104] vdd gnd cell_6t
Xbit_r105_c57 bl[57] br[57] wl[105] vdd gnd cell_6t
Xbit_r106_c57 bl[57] br[57] wl[106] vdd gnd cell_6t
Xbit_r107_c57 bl[57] br[57] wl[107] vdd gnd cell_6t
Xbit_r108_c57 bl[57] br[57] wl[108] vdd gnd cell_6t
Xbit_r109_c57 bl[57] br[57] wl[109] vdd gnd cell_6t
Xbit_r110_c57 bl[57] br[57] wl[110] vdd gnd cell_6t
Xbit_r111_c57 bl[57] br[57] wl[111] vdd gnd cell_6t
Xbit_r112_c57 bl[57] br[57] wl[112] vdd gnd cell_6t
Xbit_r113_c57 bl[57] br[57] wl[113] vdd gnd cell_6t
Xbit_r114_c57 bl[57] br[57] wl[114] vdd gnd cell_6t
Xbit_r115_c57 bl[57] br[57] wl[115] vdd gnd cell_6t
Xbit_r116_c57 bl[57] br[57] wl[116] vdd gnd cell_6t
Xbit_r117_c57 bl[57] br[57] wl[117] vdd gnd cell_6t
Xbit_r118_c57 bl[57] br[57] wl[118] vdd gnd cell_6t
Xbit_r119_c57 bl[57] br[57] wl[119] vdd gnd cell_6t
Xbit_r120_c57 bl[57] br[57] wl[120] vdd gnd cell_6t
Xbit_r121_c57 bl[57] br[57] wl[121] vdd gnd cell_6t
Xbit_r122_c57 bl[57] br[57] wl[122] vdd gnd cell_6t
Xbit_r123_c57 bl[57] br[57] wl[123] vdd gnd cell_6t
Xbit_r124_c57 bl[57] br[57] wl[124] vdd gnd cell_6t
Xbit_r125_c57 bl[57] br[57] wl[125] vdd gnd cell_6t
Xbit_r126_c57 bl[57] br[57] wl[126] vdd gnd cell_6t
Xbit_r127_c57 bl[57] br[57] wl[127] vdd gnd cell_6t
Xbit_r128_c57 bl[57] br[57] wl[128] vdd gnd cell_6t
Xbit_r129_c57 bl[57] br[57] wl[129] vdd gnd cell_6t
Xbit_r130_c57 bl[57] br[57] wl[130] vdd gnd cell_6t
Xbit_r131_c57 bl[57] br[57] wl[131] vdd gnd cell_6t
Xbit_r132_c57 bl[57] br[57] wl[132] vdd gnd cell_6t
Xbit_r133_c57 bl[57] br[57] wl[133] vdd gnd cell_6t
Xbit_r134_c57 bl[57] br[57] wl[134] vdd gnd cell_6t
Xbit_r135_c57 bl[57] br[57] wl[135] vdd gnd cell_6t
Xbit_r136_c57 bl[57] br[57] wl[136] vdd gnd cell_6t
Xbit_r137_c57 bl[57] br[57] wl[137] vdd gnd cell_6t
Xbit_r138_c57 bl[57] br[57] wl[138] vdd gnd cell_6t
Xbit_r139_c57 bl[57] br[57] wl[139] vdd gnd cell_6t
Xbit_r140_c57 bl[57] br[57] wl[140] vdd gnd cell_6t
Xbit_r141_c57 bl[57] br[57] wl[141] vdd gnd cell_6t
Xbit_r142_c57 bl[57] br[57] wl[142] vdd gnd cell_6t
Xbit_r143_c57 bl[57] br[57] wl[143] vdd gnd cell_6t
Xbit_r144_c57 bl[57] br[57] wl[144] vdd gnd cell_6t
Xbit_r145_c57 bl[57] br[57] wl[145] vdd gnd cell_6t
Xbit_r146_c57 bl[57] br[57] wl[146] vdd gnd cell_6t
Xbit_r147_c57 bl[57] br[57] wl[147] vdd gnd cell_6t
Xbit_r148_c57 bl[57] br[57] wl[148] vdd gnd cell_6t
Xbit_r149_c57 bl[57] br[57] wl[149] vdd gnd cell_6t
Xbit_r150_c57 bl[57] br[57] wl[150] vdd gnd cell_6t
Xbit_r151_c57 bl[57] br[57] wl[151] vdd gnd cell_6t
Xbit_r152_c57 bl[57] br[57] wl[152] vdd gnd cell_6t
Xbit_r153_c57 bl[57] br[57] wl[153] vdd gnd cell_6t
Xbit_r154_c57 bl[57] br[57] wl[154] vdd gnd cell_6t
Xbit_r155_c57 bl[57] br[57] wl[155] vdd gnd cell_6t
Xbit_r156_c57 bl[57] br[57] wl[156] vdd gnd cell_6t
Xbit_r157_c57 bl[57] br[57] wl[157] vdd gnd cell_6t
Xbit_r158_c57 bl[57] br[57] wl[158] vdd gnd cell_6t
Xbit_r159_c57 bl[57] br[57] wl[159] vdd gnd cell_6t
Xbit_r160_c57 bl[57] br[57] wl[160] vdd gnd cell_6t
Xbit_r161_c57 bl[57] br[57] wl[161] vdd gnd cell_6t
Xbit_r162_c57 bl[57] br[57] wl[162] vdd gnd cell_6t
Xbit_r163_c57 bl[57] br[57] wl[163] vdd gnd cell_6t
Xbit_r164_c57 bl[57] br[57] wl[164] vdd gnd cell_6t
Xbit_r165_c57 bl[57] br[57] wl[165] vdd gnd cell_6t
Xbit_r166_c57 bl[57] br[57] wl[166] vdd gnd cell_6t
Xbit_r167_c57 bl[57] br[57] wl[167] vdd gnd cell_6t
Xbit_r168_c57 bl[57] br[57] wl[168] vdd gnd cell_6t
Xbit_r169_c57 bl[57] br[57] wl[169] vdd gnd cell_6t
Xbit_r170_c57 bl[57] br[57] wl[170] vdd gnd cell_6t
Xbit_r171_c57 bl[57] br[57] wl[171] vdd gnd cell_6t
Xbit_r172_c57 bl[57] br[57] wl[172] vdd gnd cell_6t
Xbit_r173_c57 bl[57] br[57] wl[173] vdd gnd cell_6t
Xbit_r174_c57 bl[57] br[57] wl[174] vdd gnd cell_6t
Xbit_r175_c57 bl[57] br[57] wl[175] vdd gnd cell_6t
Xbit_r176_c57 bl[57] br[57] wl[176] vdd gnd cell_6t
Xbit_r177_c57 bl[57] br[57] wl[177] vdd gnd cell_6t
Xbit_r178_c57 bl[57] br[57] wl[178] vdd gnd cell_6t
Xbit_r179_c57 bl[57] br[57] wl[179] vdd gnd cell_6t
Xbit_r180_c57 bl[57] br[57] wl[180] vdd gnd cell_6t
Xbit_r181_c57 bl[57] br[57] wl[181] vdd gnd cell_6t
Xbit_r182_c57 bl[57] br[57] wl[182] vdd gnd cell_6t
Xbit_r183_c57 bl[57] br[57] wl[183] vdd gnd cell_6t
Xbit_r184_c57 bl[57] br[57] wl[184] vdd gnd cell_6t
Xbit_r185_c57 bl[57] br[57] wl[185] vdd gnd cell_6t
Xbit_r186_c57 bl[57] br[57] wl[186] vdd gnd cell_6t
Xbit_r187_c57 bl[57] br[57] wl[187] vdd gnd cell_6t
Xbit_r188_c57 bl[57] br[57] wl[188] vdd gnd cell_6t
Xbit_r189_c57 bl[57] br[57] wl[189] vdd gnd cell_6t
Xbit_r190_c57 bl[57] br[57] wl[190] vdd gnd cell_6t
Xbit_r191_c57 bl[57] br[57] wl[191] vdd gnd cell_6t
Xbit_r192_c57 bl[57] br[57] wl[192] vdd gnd cell_6t
Xbit_r193_c57 bl[57] br[57] wl[193] vdd gnd cell_6t
Xbit_r194_c57 bl[57] br[57] wl[194] vdd gnd cell_6t
Xbit_r195_c57 bl[57] br[57] wl[195] vdd gnd cell_6t
Xbit_r196_c57 bl[57] br[57] wl[196] vdd gnd cell_6t
Xbit_r197_c57 bl[57] br[57] wl[197] vdd gnd cell_6t
Xbit_r198_c57 bl[57] br[57] wl[198] vdd gnd cell_6t
Xbit_r199_c57 bl[57] br[57] wl[199] vdd gnd cell_6t
Xbit_r200_c57 bl[57] br[57] wl[200] vdd gnd cell_6t
Xbit_r201_c57 bl[57] br[57] wl[201] vdd gnd cell_6t
Xbit_r202_c57 bl[57] br[57] wl[202] vdd gnd cell_6t
Xbit_r203_c57 bl[57] br[57] wl[203] vdd gnd cell_6t
Xbit_r204_c57 bl[57] br[57] wl[204] vdd gnd cell_6t
Xbit_r205_c57 bl[57] br[57] wl[205] vdd gnd cell_6t
Xbit_r206_c57 bl[57] br[57] wl[206] vdd gnd cell_6t
Xbit_r207_c57 bl[57] br[57] wl[207] vdd gnd cell_6t
Xbit_r208_c57 bl[57] br[57] wl[208] vdd gnd cell_6t
Xbit_r209_c57 bl[57] br[57] wl[209] vdd gnd cell_6t
Xbit_r210_c57 bl[57] br[57] wl[210] vdd gnd cell_6t
Xbit_r211_c57 bl[57] br[57] wl[211] vdd gnd cell_6t
Xbit_r212_c57 bl[57] br[57] wl[212] vdd gnd cell_6t
Xbit_r213_c57 bl[57] br[57] wl[213] vdd gnd cell_6t
Xbit_r214_c57 bl[57] br[57] wl[214] vdd gnd cell_6t
Xbit_r215_c57 bl[57] br[57] wl[215] vdd gnd cell_6t
Xbit_r216_c57 bl[57] br[57] wl[216] vdd gnd cell_6t
Xbit_r217_c57 bl[57] br[57] wl[217] vdd gnd cell_6t
Xbit_r218_c57 bl[57] br[57] wl[218] vdd gnd cell_6t
Xbit_r219_c57 bl[57] br[57] wl[219] vdd gnd cell_6t
Xbit_r220_c57 bl[57] br[57] wl[220] vdd gnd cell_6t
Xbit_r221_c57 bl[57] br[57] wl[221] vdd gnd cell_6t
Xbit_r222_c57 bl[57] br[57] wl[222] vdd gnd cell_6t
Xbit_r223_c57 bl[57] br[57] wl[223] vdd gnd cell_6t
Xbit_r224_c57 bl[57] br[57] wl[224] vdd gnd cell_6t
Xbit_r225_c57 bl[57] br[57] wl[225] vdd gnd cell_6t
Xbit_r226_c57 bl[57] br[57] wl[226] vdd gnd cell_6t
Xbit_r227_c57 bl[57] br[57] wl[227] vdd gnd cell_6t
Xbit_r228_c57 bl[57] br[57] wl[228] vdd gnd cell_6t
Xbit_r229_c57 bl[57] br[57] wl[229] vdd gnd cell_6t
Xbit_r230_c57 bl[57] br[57] wl[230] vdd gnd cell_6t
Xbit_r231_c57 bl[57] br[57] wl[231] vdd gnd cell_6t
Xbit_r232_c57 bl[57] br[57] wl[232] vdd gnd cell_6t
Xbit_r233_c57 bl[57] br[57] wl[233] vdd gnd cell_6t
Xbit_r234_c57 bl[57] br[57] wl[234] vdd gnd cell_6t
Xbit_r235_c57 bl[57] br[57] wl[235] vdd gnd cell_6t
Xbit_r236_c57 bl[57] br[57] wl[236] vdd gnd cell_6t
Xbit_r237_c57 bl[57] br[57] wl[237] vdd gnd cell_6t
Xbit_r238_c57 bl[57] br[57] wl[238] vdd gnd cell_6t
Xbit_r239_c57 bl[57] br[57] wl[239] vdd gnd cell_6t
Xbit_r240_c57 bl[57] br[57] wl[240] vdd gnd cell_6t
Xbit_r241_c57 bl[57] br[57] wl[241] vdd gnd cell_6t
Xbit_r242_c57 bl[57] br[57] wl[242] vdd gnd cell_6t
Xbit_r243_c57 bl[57] br[57] wl[243] vdd gnd cell_6t
Xbit_r244_c57 bl[57] br[57] wl[244] vdd gnd cell_6t
Xbit_r245_c57 bl[57] br[57] wl[245] vdd gnd cell_6t
Xbit_r246_c57 bl[57] br[57] wl[246] vdd gnd cell_6t
Xbit_r247_c57 bl[57] br[57] wl[247] vdd gnd cell_6t
Xbit_r248_c57 bl[57] br[57] wl[248] vdd gnd cell_6t
Xbit_r249_c57 bl[57] br[57] wl[249] vdd gnd cell_6t
Xbit_r250_c57 bl[57] br[57] wl[250] vdd gnd cell_6t
Xbit_r251_c57 bl[57] br[57] wl[251] vdd gnd cell_6t
Xbit_r252_c57 bl[57] br[57] wl[252] vdd gnd cell_6t
Xbit_r253_c57 bl[57] br[57] wl[253] vdd gnd cell_6t
Xbit_r254_c57 bl[57] br[57] wl[254] vdd gnd cell_6t
Xbit_r255_c57 bl[57] br[57] wl[255] vdd gnd cell_6t
Xbit_r0_c58 bl[58] br[58] wl[0] vdd gnd cell_6t
Xbit_r1_c58 bl[58] br[58] wl[1] vdd gnd cell_6t
Xbit_r2_c58 bl[58] br[58] wl[2] vdd gnd cell_6t
Xbit_r3_c58 bl[58] br[58] wl[3] vdd gnd cell_6t
Xbit_r4_c58 bl[58] br[58] wl[4] vdd gnd cell_6t
Xbit_r5_c58 bl[58] br[58] wl[5] vdd gnd cell_6t
Xbit_r6_c58 bl[58] br[58] wl[6] vdd gnd cell_6t
Xbit_r7_c58 bl[58] br[58] wl[7] vdd gnd cell_6t
Xbit_r8_c58 bl[58] br[58] wl[8] vdd gnd cell_6t
Xbit_r9_c58 bl[58] br[58] wl[9] vdd gnd cell_6t
Xbit_r10_c58 bl[58] br[58] wl[10] vdd gnd cell_6t
Xbit_r11_c58 bl[58] br[58] wl[11] vdd gnd cell_6t
Xbit_r12_c58 bl[58] br[58] wl[12] vdd gnd cell_6t
Xbit_r13_c58 bl[58] br[58] wl[13] vdd gnd cell_6t
Xbit_r14_c58 bl[58] br[58] wl[14] vdd gnd cell_6t
Xbit_r15_c58 bl[58] br[58] wl[15] vdd gnd cell_6t
Xbit_r16_c58 bl[58] br[58] wl[16] vdd gnd cell_6t
Xbit_r17_c58 bl[58] br[58] wl[17] vdd gnd cell_6t
Xbit_r18_c58 bl[58] br[58] wl[18] vdd gnd cell_6t
Xbit_r19_c58 bl[58] br[58] wl[19] vdd gnd cell_6t
Xbit_r20_c58 bl[58] br[58] wl[20] vdd gnd cell_6t
Xbit_r21_c58 bl[58] br[58] wl[21] vdd gnd cell_6t
Xbit_r22_c58 bl[58] br[58] wl[22] vdd gnd cell_6t
Xbit_r23_c58 bl[58] br[58] wl[23] vdd gnd cell_6t
Xbit_r24_c58 bl[58] br[58] wl[24] vdd gnd cell_6t
Xbit_r25_c58 bl[58] br[58] wl[25] vdd gnd cell_6t
Xbit_r26_c58 bl[58] br[58] wl[26] vdd gnd cell_6t
Xbit_r27_c58 bl[58] br[58] wl[27] vdd gnd cell_6t
Xbit_r28_c58 bl[58] br[58] wl[28] vdd gnd cell_6t
Xbit_r29_c58 bl[58] br[58] wl[29] vdd gnd cell_6t
Xbit_r30_c58 bl[58] br[58] wl[30] vdd gnd cell_6t
Xbit_r31_c58 bl[58] br[58] wl[31] vdd gnd cell_6t
Xbit_r32_c58 bl[58] br[58] wl[32] vdd gnd cell_6t
Xbit_r33_c58 bl[58] br[58] wl[33] vdd gnd cell_6t
Xbit_r34_c58 bl[58] br[58] wl[34] vdd gnd cell_6t
Xbit_r35_c58 bl[58] br[58] wl[35] vdd gnd cell_6t
Xbit_r36_c58 bl[58] br[58] wl[36] vdd gnd cell_6t
Xbit_r37_c58 bl[58] br[58] wl[37] vdd gnd cell_6t
Xbit_r38_c58 bl[58] br[58] wl[38] vdd gnd cell_6t
Xbit_r39_c58 bl[58] br[58] wl[39] vdd gnd cell_6t
Xbit_r40_c58 bl[58] br[58] wl[40] vdd gnd cell_6t
Xbit_r41_c58 bl[58] br[58] wl[41] vdd gnd cell_6t
Xbit_r42_c58 bl[58] br[58] wl[42] vdd gnd cell_6t
Xbit_r43_c58 bl[58] br[58] wl[43] vdd gnd cell_6t
Xbit_r44_c58 bl[58] br[58] wl[44] vdd gnd cell_6t
Xbit_r45_c58 bl[58] br[58] wl[45] vdd gnd cell_6t
Xbit_r46_c58 bl[58] br[58] wl[46] vdd gnd cell_6t
Xbit_r47_c58 bl[58] br[58] wl[47] vdd gnd cell_6t
Xbit_r48_c58 bl[58] br[58] wl[48] vdd gnd cell_6t
Xbit_r49_c58 bl[58] br[58] wl[49] vdd gnd cell_6t
Xbit_r50_c58 bl[58] br[58] wl[50] vdd gnd cell_6t
Xbit_r51_c58 bl[58] br[58] wl[51] vdd gnd cell_6t
Xbit_r52_c58 bl[58] br[58] wl[52] vdd gnd cell_6t
Xbit_r53_c58 bl[58] br[58] wl[53] vdd gnd cell_6t
Xbit_r54_c58 bl[58] br[58] wl[54] vdd gnd cell_6t
Xbit_r55_c58 bl[58] br[58] wl[55] vdd gnd cell_6t
Xbit_r56_c58 bl[58] br[58] wl[56] vdd gnd cell_6t
Xbit_r57_c58 bl[58] br[58] wl[57] vdd gnd cell_6t
Xbit_r58_c58 bl[58] br[58] wl[58] vdd gnd cell_6t
Xbit_r59_c58 bl[58] br[58] wl[59] vdd gnd cell_6t
Xbit_r60_c58 bl[58] br[58] wl[60] vdd gnd cell_6t
Xbit_r61_c58 bl[58] br[58] wl[61] vdd gnd cell_6t
Xbit_r62_c58 bl[58] br[58] wl[62] vdd gnd cell_6t
Xbit_r63_c58 bl[58] br[58] wl[63] vdd gnd cell_6t
Xbit_r64_c58 bl[58] br[58] wl[64] vdd gnd cell_6t
Xbit_r65_c58 bl[58] br[58] wl[65] vdd gnd cell_6t
Xbit_r66_c58 bl[58] br[58] wl[66] vdd gnd cell_6t
Xbit_r67_c58 bl[58] br[58] wl[67] vdd gnd cell_6t
Xbit_r68_c58 bl[58] br[58] wl[68] vdd gnd cell_6t
Xbit_r69_c58 bl[58] br[58] wl[69] vdd gnd cell_6t
Xbit_r70_c58 bl[58] br[58] wl[70] vdd gnd cell_6t
Xbit_r71_c58 bl[58] br[58] wl[71] vdd gnd cell_6t
Xbit_r72_c58 bl[58] br[58] wl[72] vdd gnd cell_6t
Xbit_r73_c58 bl[58] br[58] wl[73] vdd gnd cell_6t
Xbit_r74_c58 bl[58] br[58] wl[74] vdd gnd cell_6t
Xbit_r75_c58 bl[58] br[58] wl[75] vdd gnd cell_6t
Xbit_r76_c58 bl[58] br[58] wl[76] vdd gnd cell_6t
Xbit_r77_c58 bl[58] br[58] wl[77] vdd gnd cell_6t
Xbit_r78_c58 bl[58] br[58] wl[78] vdd gnd cell_6t
Xbit_r79_c58 bl[58] br[58] wl[79] vdd gnd cell_6t
Xbit_r80_c58 bl[58] br[58] wl[80] vdd gnd cell_6t
Xbit_r81_c58 bl[58] br[58] wl[81] vdd gnd cell_6t
Xbit_r82_c58 bl[58] br[58] wl[82] vdd gnd cell_6t
Xbit_r83_c58 bl[58] br[58] wl[83] vdd gnd cell_6t
Xbit_r84_c58 bl[58] br[58] wl[84] vdd gnd cell_6t
Xbit_r85_c58 bl[58] br[58] wl[85] vdd gnd cell_6t
Xbit_r86_c58 bl[58] br[58] wl[86] vdd gnd cell_6t
Xbit_r87_c58 bl[58] br[58] wl[87] vdd gnd cell_6t
Xbit_r88_c58 bl[58] br[58] wl[88] vdd gnd cell_6t
Xbit_r89_c58 bl[58] br[58] wl[89] vdd gnd cell_6t
Xbit_r90_c58 bl[58] br[58] wl[90] vdd gnd cell_6t
Xbit_r91_c58 bl[58] br[58] wl[91] vdd gnd cell_6t
Xbit_r92_c58 bl[58] br[58] wl[92] vdd gnd cell_6t
Xbit_r93_c58 bl[58] br[58] wl[93] vdd gnd cell_6t
Xbit_r94_c58 bl[58] br[58] wl[94] vdd gnd cell_6t
Xbit_r95_c58 bl[58] br[58] wl[95] vdd gnd cell_6t
Xbit_r96_c58 bl[58] br[58] wl[96] vdd gnd cell_6t
Xbit_r97_c58 bl[58] br[58] wl[97] vdd gnd cell_6t
Xbit_r98_c58 bl[58] br[58] wl[98] vdd gnd cell_6t
Xbit_r99_c58 bl[58] br[58] wl[99] vdd gnd cell_6t
Xbit_r100_c58 bl[58] br[58] wl[100] vdd gnd cell_6t
Xbit_r101_c58 bl[58] br[58] wl[101] vdd gnd cell_6t
Xbit_r102_c58 bl[58] br[58] wl[102] vdd gnd cell_6t
Xbit_r103_c58 bl[58] br[58] wl[103] vdd gnd cell_6t
Xbit_r104_c58 bl[58] br[58] wl[104] vdd gnd cell_6t
Xbit_r105_c58 bl[58] br[58] wl[105] vdd gnd cell_6t
Xbit_r106_c58 bl[58] br[58] wl[106] vdd gnd cell_6t
Xbit_r107_c58 bl[58] br[58] wl[107] vdd gnd cell_6t
Xbit_r108_c58 bl[58] br[58] wl[108] vdd gnd cell_6t
Xbit_r109_c58 bl[58] br[58] wl[109] vdd gnd cell_6t
Xbit_r110_c58 bl[58] br[58] wl[110] vdd gnd cell_6t
Xbit_r111_c58 bl[58] br[58] wl[111] vdd gnd cell_6t
Xbit_r112_c58 bl[58] br[58] wl[112] vdd gnd cell_6t
Xbit_r113_c58 bl[58] br[58] wl[113] vdd gnd cell_6t
Xbit_r114_c58 bl[58] br[58] wl[114] vdd gnd cell_6t
Xbit_r115_c58 bl[58] br[58] wl[115] vdd gnd cell_6t
Xbit_r116_c58 bl[58] br[58] wl[116] vdd gnd cell_6t
Xbit_r117_c58 bl[58] br[58] wl[117] vdd gnd cell_6t
Xbit_r118_c58 bl[58] br[58] wl[118] vdd gnd cell_6t
Xbit_r119_c58 bl[58] br[58] wl[119] vdd gnd cell_6t
Xbit_r120_c58 bl[58] br[58] wl[120] vdd gnd cell_6t
Xbit_r121_c58 bl[58] br[58] wl[121] vdd gnd cell_6t
Xbit_r122_c58 bl[58] br[58] wl[122] vdd gnd cell_6t
Xbit_r123_c58 bl[58] br[58] wl[123] vdd gnd cell_6t
Xbit_r124_c58 bl[58] br[58] wl[124] vdd gnd cell_6t
Xbit_r125_c58 bl[58] br[58] wl[125] vdd gnd cell_6t
Xbit_r126_c58 bl[58] br[58] wl[126] vdd gnd cell_6t
Xbit_r127_c58 bl[58] br[58] wl[127] vdd gnd cell_6t
Xbit_r128_c58 bl[58] br[58] wl[128] vdd gnd cell_6t
Xbit_r129_c58 bl[58] br[58] wl[129] vdd gnd cell_6t
Xbit_r130_c58 bl[58] br[58] wl[130] vdd gnd cell_6t
Xbit_r131_c58 bl[58] br[58] wl[131] vdd gnd cell_6t
Xbit_r132_c58 bl[58] br[58] wl[132] vdd gnd cell_6t
Xbit_r133_c58 bl[58] br[58] wl[133] vdd gnd cell_6t
Xbit_r134_c58 bl[58] br[58] wl[134] vdd gnd cell_6t
Xbit_r135_c58 bl[58] br[58] wl[135] vdd gnd cell_6t
Xbit_r136_c58 bl[58] br[58] wl[136] vdd gnd cell_6t
Xbit_r137_c58 bl[58] br[58] wl[137] vdd gnd cell_6t
Xbit_r138_c58 bl[58] br[58] wl[138] vdd gnd cell_6t
Xbit_r139_c58 bl[58] br[58] wl[139] vdd gnd cell_6t
Xbit_r140_c58 bl[58] br[58] wl[140] vdd gnd cell_6t
Xbit_r141_c58 bl[58] br[58] wl[141] vdd gnd cell_6t
Xbit_r142_c58 bl[58] br[58] wl[142] vdd gnd cell_6t
Xbit_r143_c58 bl[58] br[58] wl[143] vdd gnd cell_6t
Xbit_r144_c58 bl[58] br[58] wl[144] vdd gnd cell_6t
Xbit_r145_c58 bl[58] br[58] wl[145] vdd gnd cell_6t
Xbit_r146_c58 bl[58] br[58] wl[146] vdd gnd cell_6t
Xbit_r147_c58 bl[58] br[58] wl[147] vdd gnd cell_6t
Xbit_r148_c58 bl[58] br[58] wl[148] vdd gnd cell_6t
Xbit_r149_c58 bl[58] br[58] wl[149] vdd gnd cell_6t
Xbit_r150_c58 bl[58] br[58] wl[150] vdd gnd cell_6t
Xbit_r151_c58 bl[58] br[58] wl[151] vdd gnd cell_6t
Xbit_r152_c58 bl[58] br[58] wl[152] vdd gnd cell_6t
Xbit_r153_c58 bl[58] br[58] wl[153] vdd gnd cell_6t
Xbit_r154_c58 bl[58] br[58] wl[154] vdd gnd cell_6t
Xbit_r155_c58 bl[58] br[58] wl[155] vdd gnd cell_6t
Xbit_r156_c58 bl[58] br[58] wl[156] vdd gnd cell_6t
Xbit_r157_c58 bl[58] br[58] wl[157] vdd gnd cell_6t
Xbit_r158_c58 bl[58] br[58] wl[158] vdd gnd cell_6t
Xbit_r159_c58 bl[58] br[58] wl[159] vdd gnd cell_6t
Xbit_r160_c58 bl[58] br[58] wl[160] vdd gnd cell_6t
Xbit_r161_c58 bl[58] br[58] wl[161] vdd gnd cell_6t
Xbit_r162_c58 bl[58] br[58] wl[162] vdd gnd cell_6t
Xbit_r163_c58 bl[58] br[58] wl[163] vdd gnd cell_6t
Xbit_r164_c58 bl[58] br[58] wl[164] vdd gnd cell_6t
Xbit_r165_c58 bl[58] br[58] wl[165] vdd gnd cell_6t
Xbit_r166_c58 bl[58] br[58] wl[166] vdd gnd cell_6t
Xbit_r167_c58 bl[58] br[58] wl[167] vdd gnd cell_6t
Xbit_r168_c58 bl[58] br[58] wl[168] vdd gnd cell_6t
Xbit_r169_c58 bl[58] br[58] wl[169] vdd gnd cell_6t
Xbit_r170_c58 bl[58] br[58] wl[170] vdd gnd cell_6t
Xbit_r171_c58 bl[58] br[58] wl[171] vdd gnd cell_6t
Xbit_r172_c58 bl[58] br[58] wl[172] vdd gnd cell_6t
Xbit_r173_c58 bl[58] br[58] wl[173] vdd gnd cell_6t
Xbit_r174_c58 bl[58] br[58] wl[174] vdd gnd cell_6t
Xbit_r175_c58 bl[58] br[58] wl[175] vdd gnd cell_6t
Xbit_r176_c58 bl[58] br[58] wl[176] vdd gnd cell_6t
Xbit_r177_c58 bl[58] br[58] wl[177] vdd gnd cell_6t
Xbit_r178_c58 bl[58] br[58] wl[178] vdd gnd cell_6t
Xbit_r179_c58 bl[58] br[58] wl[179] vdd gnd cell_6t
Xbit_r180_c58 bl[58] br[58] wl[180] vdd gnd cell_6t
Xbit_r181_c58 bl[58] br[58] wl[181] vdd gnd cell_6t
Xbit_r182_c58 bl[58] br[58] wl[182] vdd gnd cell_6t
Xbit_r183_c58 bl[58] br[58] wl[183] vdd gnd cell_6t
Xbit_r184_c58 bl[58] br[58] wl[184] vdd gnd cell_6t
Xbit_r185_c58 bl[58] br[58] wl[185] vdd gnd cell_6t
Xbit_r186_c58 bl[58] br[58] wl[186] vdd gnd cell_6t
Xbit_r187_c58 bl[58] br[58] wl[187] vdd gnd cell_6t
Xbit_r188_c58 bl[58] br[58] wl[188] vdd gnd cell_6t
Xbit_r189_c58 bl[58] br[58] wl[189] vdd gnd cell_6t
Xbit_r190_c58 bl[58] br[58] wl[190] vdd gnd cell_6t
Xbit_r191_c58 bl[58] br[58] wl[191] vdd gnd cell_6t
Xbit_r192_c58 bl[58] br[58] wl[192] vdd gnd cell_6t
Xbit_r193_c58 bl[58] br[58] wl[193] vdd gnd cell_6t
Xbit_r194_c58 bl[58] br[58] wl[194] vdd gnd cell_6t
Xbit_r195_c58 bl[58] br[58] wl[195] vdd gnd cell_6t
Xbit_r196_c58 bl[58] br[58] wl[196] vdd gnd cell_6t
Xbit_r197_c58 bl[58] br[58] wl[197] vdd gnd cell_6t
Xbit_r198_c58 bl[58] br[58] wl[198] vdd gnd cell_6t
Xbit_r199_c58 bl[58] br[58] wl[199] vdd gnd cell_6t
Xbit_r200_c58 bl[58] br[58] wl[200] vdd gnd cell_6t
Xbit_r201_c58 bl[58] br[58] wl[201] vdd gnd cell_6t
Xbit_r202_c58 bl[58] br[58] wl[202] vdd gnd cell_6t
Xbit_r203_c58 bl[58] br[58] wl[203] vdd gnd cell_6t
Xbit_r204_c58 bl[58] br[58] wl[204] vdd gnd cell_6t
Xbit_r205_c58 bl[58] br[58] wl[205] vdd gnd cell_6t
Xbit_r206_c58 bl[58] br[58] wl[206] vdd gnd cell_6t
Xbit_r207_c58 bl[58] br[58] wl[207] vdd gnd cell_6t
Xbit_r208_c58 bl[58] br[58] wl[208] vdd gnd cell_6t
Xbit_r209_c58 bl[58] br[58] wl[209] vdd gnd cell_6t
Xbit_r210_c58 bl[58] br[58] wl[210] vdd gnd cell_6t
Xbit_r211_c58 bl[58] br[58] wl[211] vdd gnd cell_6t
Xbit_r212_c58 bl[58] br[58] wl[212] vdd gnd cell_6t
Xbit_r213_c58 bl[58] br[58] wl[213] vdd gnd cell_6t
Xbit_r214_c58 bl[58] br[58] wl[214] vdd gnd cell_6t
Xbit_r215_c58 bl[58] br[58] wl[215] vdd gnd cell_6t
Xbit_r216_c58 bl[58] br[58] wl[216] vdd gnd cell_6t
Xbit_r217_c58 bl[58] br[58] wl[217] vdd gnd cell_6t
Xbit_r218_c58 bl[58] br[58] wl[218] vdd gnd cell_6t
Xbit_r219_c58 bl[58] br[58] wl[219] vdd gnd cell_6t
Xbit_r220_c58 bl[58] br[58] wl[220] vdd gnd cell_6t
Xbit_r221_c58 bl[58] br[58] wl[221] vdd gnd cell_6t
Xbit_r222_c58 bl[58] br[58] wl[222] vdd gnd cell_6t
Xbit_r223_c58 bl[58] br[58] wl[223] vdd gnd cell_6t
Xbit_r224_c58 bl[58] br[58] wl[224] vdd gnd cell_6t
Xbit_r225_c58 bl[58] br[58] wl[225] vdd gnd cell_6t
Xbit_r226_c58 bl[58] br[58] wl[226] vdd gnd cell_6t
Xbit_r227_c58 bl[58] br[58] wl[227] vdd gnd cell_6t
Xbit_r228_c58 bl[58] br[58] wl[228] vdd gnd cell_6t
Xbit_r229_c58 bl[58] br[58] wl[229] vdd gnd cell_6t
Xbit_r230_c58 bl[58] br[58] wl[230] vdd gnd cell_6t
Xbit_r231_c58 bl[58] br[58] wl[231] vdd gnd cell_6t
Xbit_r232_c58 bl[58] br[58] wl[232] vdd gnd cell_6t
Xbit_r233_c58 bl[58] br[58] wl[233] vdd gnd cell_6t
Xbit_r234_c58 bl[58] br[58] wl[234] vdd gnd cell_6t
Xbit_r235_c58 bl[58] br[58] wl[235] vdd gnd cell_6t
Xbit_r236_c58 bl[58] br[58] wl[236] vdd gnd cell_6t
Xbit_r237_c58 bl[58] br[58] wl[237] vdd gnd cell_6t
Xbit_r238_c58 bl[58] br[58] wl[238] vdd gnd cell_6t
Xbit_r239_c58 bl[58] br[58] wl[239] vdd gnd cell_6t
Xbit_r240_c58 bl[58] br[58] wl[240] vdd gnd cell_6t
Xbit_r241_c58 bl[58] br[58] wl[241] vdd gnd cell_6t
Xbit_r242_c58 bl[58] br[58] wl[242] vdd gnd cell_6t
Xbit_r243_c58 bl[58] br[58] wl[243] vdd gnd cell_6t
Xbit_r244_c58 bl[58] br[58] wl[244] vdd gnd cell_6t
Xbit_r245_c58 bl[58] br[58] wl[245] vdd gnd cell_6t
Xbit_r246_c58 bl[58] br[58] wl[246] vdd gnd cell_6t
Xbit_r247_c58 bl[58] br[58] wl[247] vdd gnd cell_6t
Xbit_r248_c58 bl[58] br[58] wl[248] vdd gnd cell_6t
Xbit_r249_c58 bl[58] br[58] wl[249] vdd gnd cell_6t
Xbit_r250_c58 bl[58] br[58] wl[250] vdd gnd cell_6t
Xbit_r251_c58 bl[58] br[58] wl[251] vdd gnd cell_6t
Xbit_r252_c58 bl[58] br[58] wl[252] vdd gnd cell_6t
Xbit_r253_c58 bl[58] br[58] wl[253] vdd gnd cell_6t
Xbit_r254_c58 bl[58] br[58] wl[254] vdd gnd cell_6t
Xbit_r255_c58 bl[58] br[58] wl[255] vdd gnd cell_6t
Xbit_r0_c59 bl[59] br[59] wl[0] vdd gnd cell_6t
Xbit_r1_c59 bl[59] br[59] wl[1] vdd gnd cell_6t
Xbit_r2_c59 bl[59] br[59] wl[2] vdd gnd cell_6t
Xbit_r3_c59 bl[59] br[59] wl[3] vdd gnd cell_6t
Xbit_r4_c59 bl[59] br[59] wl[4] vdd gnd cell_6t
Xbit_r5_c59 bl[59] br[59] wl[5] vdd gnd cell_6t
Xbit_r6_c59 bl[59] br[59] wl[6] vdd gnd cell_6t
Xbit_r7_c59 bl[59] br[59] wl[7] vdd gnd cell_6t
Xbit_r8_c59 bl[59] br[59] wl[8] vdd gnd cell_6t
Xbit_r9_c59 bl[59] br[59] wl[9] vdd gnd cell_6t
Xbit_r10_c59 bl[59] br[59] wl[10] vdd gnd cell_6t
Xbit_r11_c59 bl[59] br[59] wl[11] vdd gnd cell_6t
Xbit_r12_c59 bl[59] br[59] wl[12] vdd gnd cell_6t
Xbit_r13_c59 bl[59] br[59] wl[13] vdd gnd cell_6t
Xbit_r14_c59 bl[59] br[59] wl[14] vdd gnd cell_6t
Xbit_r15_c59 bl[59] br[59] wl[15] vdd gnd cell_6t
Xbit_r16_c59 bl[59] br[59] wl[16] vdd gnd cell_6t
Xbit_r17_c59 bl[59] br[59] wl[17] vdd gnd cell_6t
Xbit_r18_c59 bl[59] br[59] wl[18] vdd gnd cell_6t
Xbit_r19_c59 bl[59] br[59] wl[19] vdd gnd cell_6t
Xbit_r20_c59 bl[59] br[59] wl[20] vdd gnd cell_6t
Xbit_r21_c59 bl[59] br[59] wl[21] vdd gnd cell_6t
Xbit_r22_c59 bl[59] br[59] wl[22] vdd gnd cell_6t
Xbit_r23_c59 bl[59] br[59] wl[23] vdd gnd cell_6t
Xbit_r24_c59 bl[59] br[59] wl[24] vdd gnd cell_6t
Xbit_r25_c59 bl[59] br[59] wl[25] vdd gnd cell_6t
Xbit_r26_c59 bl[59] br[59] wl[26] vdd gnd cell_6t
Xbit_r27_c59 bl[59] br[59] wl[27] vdd gnd cell_6t
Xbit_r28_c59 bl[59] br[59] wl[28] vdd gnd cell_6t
Xbit_r29_c59 bl[59] br[59] wl[29] vdd gnd cell_6t
Xbit_r30_c59 bl[59] br[59] wl[30] vdd gnd cell_6t
Xbit_r31_c59 bl[59] br[59] wl[31] vdd gnd cell_6t
Xbit_r32_c59 bl[59] br[59] wl[32] vdd gnd cell_6t
Xbit_r33_c59 bl[59] br[59] wl[33] vdd gnd cell_6t
Xbit_r34_c59 bl[59] br[59] wl[34] vdd gnd cell_6t
Xbit_r35_c59 bl[59] br[59] wl[35] vdd gnd cell_6t
Xbit_r36_c59 bl[59] br[59] wl[36] vdd gnd cell_6t
Xbit_r37_c59 bl[59] br[59] wl[37] vdd gnd cell_6t
Xbit_r38_c59 bl[59] br[59] wl[38] vdd gnd cell_6t
Xbit_r39_c59 bl[59] br[59] wl[39] vdd gnd cell_6t
Xbit_r40_c59 bl[59] br[59] wl[40] vdd gnd cell_6t
Xbit_r41_c59 bl[59] br[59] wl[41] vdd gnd cell_6t
Xbit_r42_c59 bl[59] br[59] wl[42] vdd gnd cell_6t
Xbit_r43_c59 bl[59] br[59] wl[43] vdd gnd cell_6t
Xbit_r44_c59 bl[59] br[59] wl[44] vdd gnd cell_6t
Xbit_r45_c59 bl[59] br[59] wl[45] vdd gnd cell_6t
Xbit_r46_c59 bl[59] br[59] wl[46] vdd gnd cell_6t
Xbit_r47_c59 bl[59] br[59] wl[47] vdd gnd cell_6t
Xbit_r48_c59 bl[59] br[59] wl[48] vdd gnd cell_6t
Xbit_r49_c59 bl[59] br[59] wl[49] vdd gnd cell_6t
Xbit_r50_c59 bl[59] br[59] wl[50] vdd gnd cell_6t
Xbit_r51_c59 bl[59] br[59] wl[51] vdd gnd cell_6t
Xbit_r52_c59 bl[59] br[59] wl[52] vdd gnd cell_6t
Xbit_r53_c59 bl[59] br[59] wl[53] vdd gnd cell_6t
Xbit_r54_c59 bl[59] br[59] wl[54] vdd gnd cell_6t
Xbit_r55_c59 bl[59] br[59] wl[55] vdd gnd cell_6t
Xbit_r56_c59 bl[59] br[59] wl[56] vdd gnd cell_6t
Xbit_r57_c59 bl[59] br[59] wl[57] vdd gnd cell_6t
Xbit_r58_c59 bl[59] br[59] wl[58] vdd gnd cell_6t
Xbit_r59_c59 bl[59] br[59] wl[59] vdd gnd cell_6t
Xbit_r60_c59 bl[59] br[59] wl[60] vdd gnd cell_6t
Xbit_r61_c59 bl[59] br[59] wl[61] vdd gnd cell_6t
Xbit_r62_c59 bl[59] br[59] wl[62] vdd gnd cell_6t
Xbit_r63_c59 bl[59] br[59] wl[63] vdd gnd cell_6t
Xbit_r64_c59 bl[59] br[59] wl[64] vdd gnd cell_6t
Xbit_r65_c59 bl[59] br[59] wl[65] vdd gnd cell_6t
Xbit_r66_c59 bl[59] br[59] wl[66] vdd gnd cell_6t
Xbit_r67_c59 bl[59] br[59] wl[67] vdd gnd cell_6t
Xbit_r68_c59 bl[59] br[59] wl[68] vdd gnd cell_6t
Xbit_r69_c59 bl[59] br[59] wl[69] vdd gnd cell_6t
Xbit_r70_c59 bl[59] br[59] wl[70] vdd gnd cell_6t
Xbit_r71_c59 bl[59] br[59] wl[71] vdd gnd cell_6t
Xbit_r72_c59 bl[59] br[59] wl[72] vdd gnd cell_6t
Xbit_r73_c59 bl[59] br[59] wl[73] vdd gnd cell_6t
Xbit_r74_c59 bl[59] br[59] wl[74] vdd gnd cell_6t
Xbit_r75_c59 bl[59] br[59] wl[75] vdd gnd cell_6t
Xbit_r76_c59 bl[59] br[59] wl[76] vdd gnd cell_6t
Xbit_r77_c59 bl[59] br[59] wl[77] vdd gnd cell_6t
Xbit_r78_c59 bl[59] br[59] wl[78] vdd gnd cell_6t
Xbit_r79_c59 bl[59] br[59] wl[79] vdd gnd cell_6t
Xbit_r80_c59 bl[59] br[59] wl[80] vdd gnd cell_6t
Xbit_r81_c59 bl[59] br[59] wl[81] vdd gnd cell_6t
Xbit_r82_c59 bl[59] br[59] wl[82] vdd gnd cell_6t
Xbit_r83_c59 bl[59] br[59] wl[83] vdd gnd cell_6t
Xbit_r84_c59 bl[59] br[59] wl[84] vdd gnd cell_6t
Xbit_r85_c59 bl[59] br[59] wl[85] vdd gnd cell_6t
Xbit_r86_c59 bl[59] br[59] wl[86] vdd gnd cell_6t
Xbit_r87_c59 bl[59] br[59] wl[87] vdd gnd cell_6t
Xbit_r88_c59 bl[59] br[59] wl[88] vdd gnd cell_6t
Xbit_r89_c59 bl[59] br[59] wl[89] vdd gnd cell_6t
Xbit_r90_c59 bl[59] br[59] wl[90] vdd gnd cell_6t
Xbit_r91_c59 bl[59] br[59] wl[91] vdd gnd cell_6t
Xbit_r92_c59 bl[59] br[59] wl[92] vdd gnd cell_6t
Xbit_r93_c59 bl[59] br[59] wl[93] vdd gnd cell_6t
Xbit_r94_c59 bl[59] br[59] wl[94] vdd gnd cell_6t
Xbit_r95_c59 bl[59] br[59] wl[95] vdd gnd cell_6t
Xbit_r96_c59 bl[59] br[59] wl[96] vdd gnd cell_6t
Xbit_r97_c59 bl[59] br[59] wl[97] vdd gnd cell_6t
Xbit_r98_c59 bl[59] br[59] wl[98] vdd gnd cell_6t
Xbit_r99_c59 bl[59] br[59] wl[99] vdd gnd cell_6t
Xbit_r100_c59 bl[59] br[59] wl[100] vdd gnd cell_6t
Xbit_r101_c59 bl[59] br[59] wl[101] vdd gnd cell_6t
Xbit_r102_c59 bl[59] br[59] wl[102] vdd gnd cell_6t
Xbit_r103_c59 bl[59] br[59] wl[103] vdd gnd cell_6t
Xbit_r104_c59 bl[59] br[59] wl[104] vdd gnd cell_6t
Xbit_r105_c59 bl[59] br[59] wl[105] vdd gnd cell_6t
Xbit_r106_c59 bl[59] br[59] wl[106] vdd gnd cell_6t
Xbit_r107_c59 bl[59] br[59] wl[107] vdd gnd cell_6t
Xbit_r108_c59 bl[59] br[59] wl[108] vdd gnd cell_6t
Xbit_r109_c59 bl[59] br[59] wl[109] vdd gnd cell_6t
Xbit_r110_c59 bl[59] br[59] wl[110] vdd gnd cell_6t
Xbit_r111_c59 bl[59] br[59] wl[111] vdd gnd cell_6t
Xbit_r112_c59 bl[59] br[59] wl[112] vdd gnd cell_6t
Xbit_r113_c59 bl[59] br[59] wl[113] vdd gnd cell_6t
Xbit_r114_c59 bl[59] br[59] wl[114] vdd gnd cell_6t
Xbit_r115_c59 bl[59] br[59] wl[115] vdd gnd cell_6t
Xbit_r116_c59 bl[59] br[59] wl[116] vdd gnd cell_6t
Xbit_r117_c59 bl[59] br[59] wl[117] vdd gnd cell_6t
Xbit_r118_c59 bl[59] br[59] wl[118] vdd gnd cell_6t
Xbit_r119_c59 bl[59] br[59] wl[119] vdd gnd cell_6t
Xbit_r120_c59 bl[59] br[59] wl[120] vdd gnd cell_6t
Xbit_r121_c59 bl[59] br[59] wl[121] vdd gnd cell_6t
Xbit_r122_c59 bl[59] br[59] wl[122] vdd gnd cell_6t
Xbit_r123_c59 bl[59] br[59] wl[123] vdd gnd cell_6t
Xbit_r124_c59 bl[59] br[59] wl[124] vdd gnd cell_6t
Xbit_r125_c59 bl[59] br[59] wl[125] vdd gnd cell_6t
Xbit_r126_c59 bl[59] br[59] wl[126] vdd gnd cell_6t
Xbit_r127_c59 bl[59] br[59] wl[127] vdd gnd cell_6t
Xbit_r128_c59 bl[59] br[59] wl[128] vdd gnd cell_6t
Xbit_r129_c59 bl[59] br[59] wl[129] vdd gnd cell_6t
Xbit_r130_c59 bl[59] br[59] wl[130] vdd gnd cell_6t
Xbit_r131_c59 bl[59] br[59] wl[131] vdd gnd cell_6t
Xbit_r132_c59 bl[59] br[59] wl[132] vdd gnd cell_6t
Xbit_r133_c59 bl[59] br[59] wl[133] vdd gnd cell_6t
Xbit_r134_c59 bl[59] br[59] wl[134] vdd gnd cell_6t
Xbit_r135_c59 bl[59] br[59] wl[135] vdd gnd cell_6t
Xbit_r136_c59 bl[59] br[59] wl[136] vdd gnd cell_6t
Xbit_r137_c59 bl[59] br[59] wl[137] vdd gnd cell_6t
Xbit_r138_c59 bl[59] br[59] wl[138] vdd gnd cell_6t
Xbit_r139_c59 bl[59] br[59] wl[139] vdd gnd cell_6t
Xbit_r140_c59 bl[59] br[59] wl[140] vdd gnd cell_6t
Xbit_r141_c59 bl[59] br[59] wl[141] vdd gnd cell_6t
Xbit_r142_c59 bl[59] br[59] wl[142] vdd gnd cell_6t
Xbit_r143_c59 bl[59] br[59] wl[143] vdd gnd cell_6t
Xbit_r144_c59 bl[59] br[59] wl[144] vdd gnd cell_6t
Xbit_r145_c59 bl[59] br[59] wl[145] vdd gnd cell_6t
Xbit_r146_c59 bl[59] br[59] wl[146] vdd gnd cell_6t
Xbit_r147_c59 bl[59] br[59] wl[147] vdd gnd cell_6t
Xbit_r148_c59 bl[59] br[59] wl[148] vdd gnd cell_6t
Xbit_r149_c59 bl[59] br[59] wl[149] vdd gnd cell_6t
Xbit_r150_c59 bl[59] br[59] wl[150] vdd gnd cell_6t
Xbit_r151_c59 bl[59] br[59] wl[151] vdd gnd cell_6t
Xbit_r152_c59 bl[59] br[59] wl[152] vdd gnd cell_6t
Xbit_r153_c59 bl[59] br[59] wl[153] vdd gnd cell_6t
Xbit_r154_c59 bl[59] br[59] wl[154] vdd gnd cell_6t
Xbit_r155_c59 bl[59] br[59] wl[155] vdd gnd cell_6t
Xbit_r156_c59 bl[59] br[59] wl[156] vdd gnd cell_6t
Xbit_r157_c59 bl[59] br[59] wl[157] vdd gnd cell_6t
Xbit_r158_c59 bl[59] br[59] wl[158] vdd gnd cell_6t
Xbit_r159_c59 bl[59] br[59] wl[159] vdd gnd cell_6t
Xbit_r160_c59 bl[59] br[59] wl[160] vdd gnd cell_6t
Xbit_r161_c59 bl[59] br[59] wl[161] vdd gnd cell_6t
Xbit_r162_c59 bl[59] br[59] wl[162] vdd gnd cell_6t
Xbit_r163_c59 bl[59] br[59] wl[163] vdd gnd cell_6t
Xbit_r164_c59 bl[59] br[59] wl[164] vdd gnd cell_6t
Xbit_r165_c59 bl[59] br[59] wl[165] vdd gnd cell_6t
Xbit_r166_c59 bl[59] br[59] wl[166] vdd gnd cell_6t
Xbit_r167_c59 bl[59] br[59] wl[167] vdd gnd cell_6t
Xbit_r168_c59 bl[59] br[59] wl[168] vdd gnd cell_6t
Xbit_r169_c59 bl[59] br[59] wl[169] vdd gnd cell_6t
Xbit_r170_c59 bl[59] br[59] wl[170] vdd gnd cell_6t
Xbit_r171_c59 bl[59] br[59] wl[171] vdd gnd cell_6t
Xbit_r172_c59 bl[59] br[59] wl[172] vdd gnd cell_6t
Xbit_r173_c59 bl[59] br[59] wl[173] vdd gnd cell_6t
Xbit_r174_c59 bl[59] br[59] wl[174] vdd gnd cell_6t
Xbit_r175_c59 bl[59] br[59] wl[175] vdd gnd cell_6t
Xbit_r176_c59 bl[59] br[59] wl[176] vdd gnd cell_6t
Xbit_r177_c59 bl[59] br[59] wl[177] vdd gnd cell_6t
Xbit_r178_c59 bl[59] br[59] wl[178] vdd gnd cell_6t
Xbit_r179_c59 bl[59] br[59] wl[179] vdd gnd cell_6t
Xbit_r180_c59 bl[59] br[59] wl[180] vdd gnd cell_6t
Xbit_r181_c59 bl[59] br[59] wl[181] vdd gnd cell_6t
Xbit_r182_c59 bl[59] br[59] wl[182] vdd gnd cell_6t
Xbit_r183_c59 bl[59] br[59] wl[183] vdd gnd cell_6t
Xbit_r184_c59 bl[59] br[59] wl[184] vdd gnd cell_6t
Xbit_r185_c59 bl[59] br[59] wl[185] vdd gnd cell_6t
Xbit_r186_c59 bl[59] br[59] wl[186] vdd gnd cell_6t
Xbit_r187_c59 bl[59] br[59] wl[187] vdd gnd cell_6t
Xbit_r188_c59 bl[59] br[59] wl[188] vdd gnd cell_6t
Xbit_r189_c59 bl[59] br[59] wl[189] vdd gnd cell_6t
Xbit_r190_c59 bl[59] br[59] wl[190] vdd gnd cell_6t
Xbit_r191_c59 bl[59] br[59] wl[191] vdd gnd cell_6t
Xbit_r192_c59 bl[59] br[59] wl[192] vdd gnd cell_6t
Xbit_r193_c59 bl[59] br[59] wl[193] vdd gnd cell_6t
Xbit_r194_c59 bl[59] br[59] wl[194] vdd gnd cell_6t
Xbit_r195_c59 bl[59] br[59] wl[195] vdd gnd cell_6t
Xbit_r196_c59 bl[59] br[59] wl[196] vdd gnd cell_6t
Xbit_r197_c59 bl[59] br[59] wl[197] vdd gnd cell_6t
Xbit_r198_c59 bl[59] br[59] wl[198] vdd gnd cell_6t
Xbit_r199_c59 bl[59] br[59] wl[199] vdd gnd cell_6t
Xbit_r200_c59 bl[59] br[59] wl[200] vdd gnd cell_6t
Xbit_r201_c59 bl[59] br[59] wl[201] vdd gnd cell_6t
Xbit_r202_c59 bl[59] br[59] wl[202] vdd gnd cell_6t
Xbit_r203_c59 bl[59] br[59] wl[203] vdd gnd cell_6t
Xbit_r204_c59 bl[59] br[59] wl[204] vdd gnd cell_6t
Xbit_r205_c59 bl[59] br[59] wl[205] vdd gnd cell_6t
Xbit_r206_c59 bl[59] br[59] wl[206] vdd gnd cell_6t
Xbit_r207_c59 bl[59] br[59] wl[207] vdd gnd cell_6t
Xbit_r208_c59 bl[59] br[59] wl[208] vdd gnd cell_6t
Xbit_r209_c59 bl[59] br[59] wl[209] vdd gnd cell_6t
Xbit_r210_c59 bl[59] br[59] wl[210] vdd gnd cell_6t
Xbit_r211_c59 bl[59] br[59] wl[211] vdd gnd cell_6t
Xbit_r212_c59 bl[59] br[59] wl[212] vdd gnd cell_6t
Xbit_r213_c59 bl[59] br[59] wl[213] vdd gnd cell_6t
Xbit_r214_c59 bl[59] br[59] wl[214] vdd gnd cell_6t
Xbit_r215_c59 bl[59] br[59] wl[215] vdd gnd cell_6t
Xbit_r216_c59 bl[59] br[59] wl[216] vdd gnd cell_6t
Xbit_r217_c59 bl[59] br[59] wl[217] vdd gnd cell_6t
Xbit_r218_c59 bl[59] br[59] wl[218] vdd gnd cell_6t
Xbit_r219_c59 bl[59] br[59] wl[219] vdd gnd cell_6t
Xbit_r220_c59 bl[59] br[59] wl[220] vdd gnd cell_6t
Xbit_r221_c59 bl[59] br[59] wl[221] vdd gnd cell_6t
Xbit_r222_c59 bl[59] br[59] wl[222] vdd gnd cell_6t
Xbit_r223_c59 bl[59] br[59] wl[223] vdd gnd cell_6t
Xbit_r224_c59 bl[59] br[59] wl[224] vdd gnd cell_6t
Xbit_r225_c59 bl[59] br[59] wl[225] vdd gnd cell_6t
Xbit_r226_c59 bl[59] br[59] wl[226] vdd gnd cell_6t
Xbit_r227_c59 bl[59] br[59] wl[227] vdd gnd cell_6t
Xbit_r228_c59 bl[59] br[59] wl[228] vdd gnd cell_6t
Xbit_r229_c59 bl[59] br[59] wl[229] vdd gnd cell_6t
Xbit_r230_c59 bl[59] br[59] wl[230] vdd gnd cell_6t
Xbit_r231_c59 bl[59] br[59] wl[231] vdd gnd cell_6t
Xbit_r232_c59 bl[59] br[59] wl[232] vdd gnd cell_6t
Xbit_r233_c59 bl[59] br[59] wl[233] vdd gnd cell_6t
Xbit_r234_c59 bl[59] br[59] wl[234] vdd gnd cell_6t
Xbit_r235_c59 bl[59] br[59] wl[235] vdd gnd cell_6t
Xbit_r236_c59 bl[59] br[59] wl[236] vdd gnd cell_6t
Xbit_r237_c59 bl[59] br[59] wl[237] vdd gnd cell_6t
Xbit_r238_c59 bl[59] br[59] wl[238] vdd gnd cell_6t
Xbit_r239_c59 bl[59] br[59] wl[239] vdd gnd cell_6t
Xbit_r240_c59 bl[59] br[59] wl[240] vdd gnd cell_6t
Xbit_r241_c59 bl[59] br[59] wl[241] vdd gnd cell_6t
Xbit_r242_c59 bl[59] br[59] wl[242] vdd gnd cell_6t
Xbit_r243_c59 bl[59] br[59] wl[243] vdd gnd cell_6t
Xbit_r244_c59 bl[59] br[59] wl[244] vdd gnd cell_6t
Xbit_r245_c59 bl[59] br[59] wl[245] vdd gnd cell_6t
Xbit_r246_c59 bl[59] br[59] wl[246] vdd gnd cell_6t
Xbit_r247_c59 bl[59] br[59] wl[247] vdd gnd cell_6t
Xbit_r248_c59 bl[59] br[59] wl[248] vdd gnd cell_6t
Xbit_r249_c59 bl[59] br[59] wl[249] vdd gnd cell_6t
Xbit_r250_c59 bl[59] br[59] wl[250] vdd gnd cell_6t
Xbit_r251_c59 bl[59] br[59] wl[251] vdd gnd cell_6t
Xbit_r252_c59 bl[59] br[59] wl[252] vdd gnd cell_6t
Xbit_r253_c59 bl[59] br[59] wl[253] vdd gnd cell_6t
Xbit_r254_c59 bl[59] br[59] wl[254] vdd gnd cell_6t
Xbit_r255_c59 bl[59] br[59] wl[255] vdd gnd cell_6t
Xbit_r0_c60 bl[60] br[60] wl[0] vdd gnd cell_6t
Xbit_r1_c60 bl[60] br[60] wl[1] vdd gnd cell_6t
Xbit_r2_c60 bl[60] br[60] wl[2] vdd gnd cell_6t
Xbit_r3_c60 bl[60] br[60] wl[3] vdd gnd cell_6t
Xbit_r4_c60 bl[60] br[60] wl[4] vdd gnd cell_6t
Xbit_r5_c60 bl[60] br[60] wl[5] vdd gnd cell_6t
Xbit_r6_c60 bl[60] br[60] wl[6] vdd gnd cell_6t
Xbit_r7_c60 bl[60] br[60] wl[7] vdd gnd cell_6t
Xbit_r8_c60 bl[60] br[60] wl[8] vdd gnd cell_6t
Xbit_r9_c60 bl[60] br[60] wl[9] vdd gnd cell_6t
Xbit_r10_c60 bl[60] br[60] wl[10] vdd gnd cell_6t
Xbit_r11_c60 bl[60] br[60] wl[11] vdd gnd cell_6t
Xbit_r12_c60 bl[60] br[60] wl[12] vdd gnd cell_6t
Xbit_r13_c60 bl[60] br[60] wl[13] vdd gnd cell_6t
Xbit_r14_c60 bl[60] br[60] wl[14] vdd gnd cell_6t
Xbit_r15_c60 bl[60] br[60] wl[15] vdd gnd cell_6t
Xbit_r16_c60 bl[60] br[60] wl[16] vdd gnd cell_6t
Xbit_r17_c60 bl[60] br[60] wl[17] vdd gnd cell_6t
Xbit_r18_c60 bl[60] br[60] wl[18] vdd gnd cell_6t
Xbit_r19_c60 bl[60] br[60] wl[19] vdd gnd cell_6t
Xbit_r20_c60 bl[60] br[60] wl[20] vdd gnd cell_6t
Xbit_r21_c60 bl[60] br[60] wl[21] vdd gnd cell_6t
Xbit_r22_c60 bl[60] br[60] wl[22] vdd gnd cell_6t
Xbit_r23_c60 bl[60] br[60] wl[23] vdd gnd cell_6t
Xbit_r24_c60 bl[60] br[60] wl[24] vdd gnd cell_6t
Xbit_r25_c60 bl[60] br[60] wl[25] vdd gnd cell_6t
Xbit_r26_c60 bl[60] br[60] wl[26] vdd gnd cell_6t
Xbit_r27_c60 bl[60] br[60] wl[27] vdd gnd cell_6t
Xbit_r28_c60 bl[60] br[60] wl[28] vdd gnd cell_6t
Xbit_r29_c60 bl[60] br[60] wl[29] vdd gnd cell_6t
Xbit_r30_c60 bl[60] br[60] wl[30] vdd gnd cell_6t
Xbit_r31_c60 bl[60] br[60] wl[31] vdd gnd cell_6t
Xbit_r32_c60 bl[60] br[60] wl[32] vdd gnd cell_6t
Xbit_r33_c60 bl[60] br[60] wl[33] vdd gnd cell_6t
Xbit_r34_c60 bl[60] br[60] wl[34] vdd gnd cell_6t
Xbit_r35_c60 bl[60] br[60] wl[35] vdd gnd cell_6t
Xbit_r36_c60 bl[60] br[60] wl[36] vdd gnd cell_6t
Xbit_r37_c60 bl[60] br[60] wl[37] vdd gnd cell_6t
Xbit_r38_c60 bl[60] br[60] wl[38] vdd gnd cell_6t
Xbit_r39_c60 bl[60] br[60] wl[39] vdd gnd cell_6t
Xbit_r40_c60 bl[60] br[60] wl[40] vdd gnd cell_6t
Xbit_r41_c60 bl[60] br[60] wl[41] vdd gnd cell_6t
Xbit_r42_c60 bl[60] br[60] wl[42] vdd gnd cell_6t
Xbit_r43_c60 bl[60] br[60] wl[43] vdd gnd cell_6t
Xbit_r44_c60 bl[60] br[60] wl[44] vdd gnd cell_6t
Xbit_r45_c60 bl[60] br[60] wl[45] vdd gnd cell_6t
Xbit_r46_c60 bl[60] br[60] wl[46] vdd gnd cell_6t
Xbit_r47_c60 bl[60] br[60] wl[47] vdd gnd cell_6t
Xbit_r48_c60 bl[60] br[60] wl[48] vdd gnd cell_6t
Xbit_r49_c60 bl[60] br[60] wl[49] vdd gnd cell_6t
Xbit_r50_c60 bl[60] br[60] wl[50] vdd gnd cell_6t
Xbit_r51_c60 bl[60] br[60] wl[51] vdd gnd cell_6t
Xbit_r52_c60 bl[60] br[60] wl[52] vdd gnd cell_6t
Xbit_r53_c60 bl[60] br[60] wl[53] vdd gnd cell_6t
Xbit_r54_c60 bl[60] br[60] wl[54] vdd gnd cell_6t
Xbit_r55_c60 bl[60] br[60] wl[55] vdd gnd cell_6t
Xbit_r56_c60 bl[60] br[60] wl[56] vdd gnd cell_6t
Xbit_r57_c60 bl[60] br[60] wl[57] vdd gnd cell_6t
Xbit_r58_c60 bl[60] br[60] wl[58] vdd gnd cell_6t
Xbit_r59_c60 bl[60] br[60] wl[59] vdd gnd cell_6t
Xbit_r60_c60 bl[60] br[60] wl[60] vdd gnd cell_6t
Xbit_r61_c60 bl[60] br[60] wl[61] vdd gnd cell_6t
Xbit_r62_c60 bl[60] br[60] wl[62] vdd gnd cell_6t
Xbit_r63_c60 bl[60] br[60] wl[63] vdd gnd cell_6t
Xbit_r64_c60 bl[60] br[60] wl[64] vdd gnd cell_6t
Xbit_r65_c60 bl[60] br[60] wl[65] vdd gnd cell_6t
Xbit_r66_c60 bl[60] br[60] wl[66] vdd gnd cell_6t
Xbit_r67_c60 bl[60] br[60] wl[67] vdd gnd cell_6t
Xbit_r68_c60 bl[60] br[60] wl[68] vdd gnd cell_6t
Xbit_r69_c60 bl[60] br[60] wl[69] vdd gnd cell_6t
Xbit_r70_c60 bl[60] br[60] wl[70] vdd gnd cell_6t
Xbit_r71_c60 bl[60] br[60] wl[71] vdd gnd cell_6t
Xbit_r72_c60 bl[60] br[60] wl[72] vdd gnd cell_6t
Xbit_r73_c60 bl[60] br[60] wl[73] vdd gnd cell_6t
Xbit_r74_c60 bl[60] br[60] wl[74] vdd gnd cell_6t
Xbit_r75_c60 bl[60] br[60] wl[75] vdd gnd cell_6t
Xbit_r76_c60 bl[60] br[60] wl[76] vdd gnd cell_6t
Xbit_r77_c60 bl[60] br[60] wl[77] vdd gnd cell_6t
Xbit_r78_c60 bl[60] br[60] wl[78] vdd gnd cell_6t
Xbit_r79_c60 bl[60] br[60] wl[79] vdd gnd cell_6t
Xbit_r80_c60 bl[60] br[60] wl[80] vdd gnd cell_6t
Xbit_r81_c60 bl[60] br[60] wl[81] vdd gnd cell_6t
Xbit_r82_c60 bl[60] br[60] wl[82] vdd gnd cell_6t
Xbit_r83_c60 bl[60] br[60] wl[83] vdd gnd cell_6t
Xbit_r84_c60 bl[60] br[60] wl[84] vdd gnd cell_6t
Xbit_r85_c60 bl[60] br[60] wl[85] vdd gnd cell_6t
Xbit_r86_c60 bl[60] br[60] wl[86] vdd gnd cell_6t
Xbit_r87_c60 bl[60] br[60] wl[87] vdd gnd cell_6t
Xbit_r88_c60 bl[60] br[60] wl[88] vdd gnd cell_6t
Xbit_r89_c60 bl[60] br[60] wl[89] vdd gnd cell_6t
Xbit_r90_c60 bl[60] br[60] wl[90] vdd gnd cell_6t
Xbit_r91_c60 bl[60] br[60] wl[91] vdd gnd cell_6t
Xbit_r92_c60 bl[60] br[60] wl[92] vdd gnd cell_6t
Xbit_r93_c60 bl[60] br[60] wl[93] vdd gnd cell_6t
Xbit_r94_c60 bl[60] br[60] wl[94] vdd gnd cell_6t
Xbit_r95_c60 bl[60] br[60] wl[95] vdd gnd cell_6t
Xbit_r96_c60 bl[60] br[60] wl[96] vdd gnd cell_6t
Xbit_r97_c60 bl[60] br[60] wl[97] vdd gnd cell_6t
Xbit_r98_c60 bl[60] br[60] wl[98] vdd gnd cell_6t
Xbit_r99_c60 bl[60] br[60] wl[99] vdd gnd cell_6t
Xbit_r100_c60 bl[60] br[60] wl[100] vdd gnd cell_6t
Xbit_r101_c60 bl[60] br[60] wl[101] vdd gnd cell_6t
Xbit_r102_c60 bl[60] br[60] wl[102] vdd gnd cell_6t
Xbit_r103_c60 bl[60] br[60] wl[103] vdd gnd cell_6t
Xbit_r104_c60 bl[60] br[60] wl[104] vdd gnd cell_6t
Xbit_r105_c60 bl[60] br[60] wl[105] vdd gnd cell_6t
Xbit_r106_c60 bl[60] br[60] wl[106] vdd gnd cell_6t
Xbit_r107_c60 bl[60] br[60] wl[107] vdd gnd cell_6t
Xbit_r108_c60 bl[60] br[60] wl[108] vdd gnd cell_6t
Xbit_r109_c60 bl[60] br[60] wl[109] vdd gnd cell_6t
Xbit_r110_c60 bl[60] br[60] wl[110] vdd gnd cell_6t
Xbit_r111_c60 bl[60] br[60] wl[111] vdd gnd cell_6t
Xbit_r112_c60 bl[60] br[60] wl[112] vdd gnd cell_6t
Xbit_r113_c60 bl[60] br[60] wl[113] vdd gnd cell_6t
Xbit_r114_c60 bl[60] br[60] wl[114] vdd gnd cell_6t
Xbit_r115_c60 bl[60] br[60] wl[115] vdd gnd cell_6t
Xbit_r116_c60 bl[60] br[60] wl[116] vdd gnd cell_6t
Xbit_r117_c60 bl[60] br[60] wl[117] vdd gnd cell_6t
Xbit_r118_c60 bl[60] br[60] wl[118] vdd gnd cell_6t
Xbit_r119_c60 bl[60] br[60] wl[119] vdd gnd cell_6t
Xbit_r120_c60 bl[60] br[60] wl[120] vdd gnd cell_6t
Xbit_r121_c60 bl[60] br[60] wl[121] vdd gnd cell_6t
Xbit_r122_c60 bl[60] br[60] wl[122] vdd gnd cell_6t
Xbit_r123_c60 bl[60] br[60] wl[123] vdd gnd cell_6t
Xbit_r124_c60 bl[60] br[60] wl[124] vdd gnd cell_6t
Xbit_r125_c60 bl[60] br[60] wl[125] vdd gnd cell_6t
Xbit_r126_c60 bl[60] br[60] wl[126] vdd gnd cell_6t
Xbit_r127_c60 bl[60] br[60] wl[127] vdd gnd cell_6t
Xbit_r128_c60 bl[60] br[60] wl[128] vdd gnd cell_6t
Xbit_r129_c60 bl[60] br[60] wl[129] vdd gnd cell_6t
Xbit_r130_c60 bl[60] br[60] wl[130] vdd gnd cell_6t
Xbit_r131_c60 bl[60] br[60] wl[131] vdd gnd cell_6t
Xbit_r132_c60 bl[60] br[60] wl[132] vdd gnd cell_6t
Xbit_r133_c60 bl[60] br[60] wl[133] vdd gnd cell_6t
Xbit_r134_c60 bl[60] br[60] wl[134] vdd gnd cell_6t
Xbit_r135_c60 bl[60] br[60] wl[135] vdd gnd cell_6t
Xbit_r136_c60 bl[60] br[60] wl[136] vdd gnd cell_6t
Xbit_r137_c60 bl[60] br[60] wl[137] vdd gnd cell_6t
Xbit_r138_c60 bl[60] br[60] wl[138] vdd gnd cell_6t
Xbit_r139_c60 bl[60] br[60] wl[139] vdd gnd cell_6t
Xbit_r140_c60 bl[60] br[60] wl[140] vdd gnd cell_6t
Xbit_r141_c60 bl[60] br[60] wl[141] vdd gnd cell_6t
Xbit_r142_c60 bl[60] br[60] wl[142] vdd gnd cell_6t
Xbit_r143_c60 bl[60] br[60] wl[143] vdd gnd cell_6t
Xbit_r144_c60 bl[60] br[60] wl[144] vdd gnd cell_6t
Xbit_r145_c60 bl[60] br[60] wl[145] vdd gnd cell_6t
Xbit_r146_c60 bl[60] br[60] wl[146] vdd gnd cell_6t
Xbit_r147_c60 bl[60] br[60] wl[147] vdd gnd cell_6t
Xbit_r148_c60 bl[60] br[60] wl[148] vdd gnd cell_6t
Xbit_r149_c60 bl[60] br[60] wl[149] vdd gnd cell_6t
Xbit_r150_c60 bl[60] br[60] wl[150] vdd gnd cell_6t
Xbit_r151_c60 bl[60] br[60] wl[151] vdd gnd cell_6t
Xbit_r152_c60 bl[60] br[60] wl[152] vdd gnd cell_6t
Xbit_r153_c60 bl[60] br[60] wl[153] vdd gnd cell_6t
Xbit_r154_c60 bl[60] br[60] wl[154] vdd gnd cell_6t
Xbit_r155_c60 bl[60] br[60] wl[155] vdd gnd cell_6t
Xbit_r156_c60 bl[60] br[60] wl[156] vdd gnd cell_6t
Xbit_r157_c60 bl[60] br[60] wl[157] vdd gnd cell_6t
Xbit_r158_c60 bl[60] br[60] wl[158] vdd gnd cell_6t
Xbit_r159_c60 bl[60] br[60] wl[159] vdd gnd cell_6t
Xbit_r160_c60 bl[60] br[60] wl[160] vdd gnd cell_6t
Xbit_r161_c60 bl[60] br[60] wl[161] vdd gnd cell_6t
Xbit_r162_c60 bl[60] br[60] wl[162] vdd gnd cell_6t
Xbit_r163_c60 bl[60] br[60] wl[163] vdd gnd cell_6t
Xbit_r164_c60 bl[60] br[60] wl[164] vdd gnd cell_6t
Xbit_r165_c60 bl[60] br[60] wl[165] vdd gnd cell_6t
Xbit_r166_c60 bl[60] br[60] wl[166] vdd gnd cell_6t
Xbit_r167_c60 bl[60] br[60] wl[167] vdd gnd cell_6t
Xbit_r168_c60 bl[60] br[60] wl[168] vdd gnd cell_6t
Xbit_r169_c60 bl[60] br[60] wl[169] vdd gnd cell_6t
Xbit_r170_c60 bl[60] br[60] wl[170] vdd gnd cell_6t
Xbit_r171_c60 bl[60] br[60] wl[171] vdd gnd cell_6t
Xbit_r172_c60 bl[60] br[60] wl[172] vdd gnd cell_6t
Xbit_r173_c60 bl[60] br[60] wl[173] vdd gnd cell_6t
Xbit_r174_c60 bl[60] br[60] wl[174] vdd gnd cell_6t
Xbit_r175_c60 bl[60] br[60] wl[175] vdd gnd cell_6t
Xbit_r176_c60 bl[60] br[60] wl[176] vdd gnd cell_6t
Xbit_r177_c60 bl[60] br[60] wl[177] vdd gnd cell_6t
Xbit_r178_c60 bl[60] br[60] wl[178] vdd gnd cell_6t
Xbit_r179_c60 bl[60] br[60] wl[179] vdd gnd cell_6t
Xbit_r180_c60 bl[60] br[60] wl[180] vdd gnd cell_6t
Xbit_r181_c60 bl[60] br[60] wl[181] vdd gnd cell_6t
Xbit_r182_c60 bl[60] br[60] wl[182] vdd gnd cell_6t
Xbit_r183_c60 bl[60] br[60] wl[183] vdd gnd cell_6t
Xbit_r184_c60 bl[60] br[60] wl[184] vdd gnd cell_6t
Xbit_r185_c60 bl[60] br[60] wl[185] vdd gnd cell_6t
Xbit_r186_c60 bl[60] br[60] wl[186] vdd gnd cell_6t
Xbit_r187_c60 bl[60] br[60] wl[187] vdd gnd cell_6t
Xbit_r188_c60 bl[60] br[60] wl[188] vdd gnd cell_6t
Xbit_r189_c60 bl[60] br[60] wl[189] vdd gnd cell_6t
Xbit_r190_c60 bl[60] br[60] wl[190] vdd gnd cell_6t
Xbit_r191_c60 bl[60] br[60] wl[191] vdd gnd cell_6t
Xbit_r192_c60 bl[60] br[60] wl[192] vdd gnd cell_6t
Xbit_r193_c60 bl[60] br[60] wl[193] vdd gnd cell_6t
Xbit_r194_c60 bl[60] br[60] wl[194] vdd gnd cell_6t
Xbit_r195_c60 bl[60] br[60] wl[195] vdd gnd cell_6t
Xbit_r196_c60 bl[60] br[60] wl[196] vdd gnd cell_6t
Xbit_r197_c60 bl[60] br[60] wl[197] vdd gnd cell_6t
Xbit_r198_c60 bl[60] br[60] wl[198] vdd gnd cell_6t
Xbit_r199_c60 bl[60] br[60] wl[199] vdd gnd cell_6t
Xbit_r200_c60 bl[60] br[60] wl[200] vdd gnd cell_6t
Xbit_r201_c60 bl[60] br[60] wl[201] vdd gnd cell_6t
Xbit_r202_c60 bl[60] br[60] wl[202] vdd gnd cell_6t
Xbit_r203_c60 bl[60] br[60] wl[203] vdd gnd cell_6t
Xbit_r204_c60 bl[60] br[60] wl[204] vdd gnd cell_6t
Xbit_r205_c60 bl[60] br[60] wl[205] vdd gnd cell_6t
Xbit_r206_c60 bl[60] br[60] wl[206] vdd gnd cell_6t
Xbit_r207_c60 bl[60] br[60] wl[207] vdd gnd cell_6t
Xbit_r208_c60 bl[60] br[60] wl[208] vdd gnd cell_6t
Xbit_r209_c60 bl[60] br[60] wl[209] vdd gnd cell_6t
Xbit_r210_c60 bl[60] br[60] wl[210] vdd gnd cell_6t
Xbit_r211_c60 bl[60] br[60] wl[211] vdd gnd cell_6t
Xbit_r212_c60 bl[60] br[60] wl[212] vdd gnd cell_6t
Xbit_r213_c60 bl[60] br[60] wl[213] vdd gnd cell_6t
Xbit_r214_c60 bl[60] br[60] wl[214] vdd gnd cell_6t
Xbit_r215_c60 bl[60] br[60] wl[215] vdd gnd cell_6t
Xbit_r216_c60 bl[60] br[60] wl[216] vdd gnd cell_6t
Xbit_r217_c60 bl[60] br[60] wl[217] vdd gnd cell_6t
Xbit_r218_c60 bl[60] br[60] wl[218] vdd gnd cell_6t
Xbit_r219_c60 bl[60] br[60] wl[219] vdd gnd cell_6t
Xbit_r220_c60 bl[60] br[60] wl[220] vdd gnd cell_6t
Xbit_r221_c60 bl[60] br[60] wl[221] vdd gnd cell_6t
Xbit_r222_c60 bl[60] br[60] wl[222] vdd gnd cell_6t
Xbit_r223_c60 bl[60] br[60] wl[223] vdd gnd cell_6t
Xbit_r224_c60 bl[60] br[60] wl[224] vdd gnd cell_6t
Xbit_r225_c60 bl[60] br[60] wl[225] vdd gnd cell_6t
Xbit_r226_c60 bl[60] br[60] wl[226] vdd gnd cell_6t
Xbit_r227_c60 bl[60] br[60] wl[227] vdd gnd cell_6t
Xbit_r228_c60 bl[60] br[60] wl[228] vdd gnd cell_6t
Xbit_r229_c60 bl[60] br[60] wl[229] vdd gnd cell_6t
Xbit_r230_c60 bl[60] br[60] wl[230] vdd gnd cell_6t
Xbit_r231_c60 bl[60] br[60] wl[231] vdd gnd cell_6t
Xbit_r232_c60 bl[60] br[60] wl[232] vdd gnd cell_6t
Xbit_r233_c60 bl[60] br[60] wl[233] vdd gnd cell_6t
Xbit_r234_c60 bl[60] br[60] wl[234] vdd gnd cell_6t
Xbit_r235_c60 bl[60] br[60] wl[235] vdd gnd cell_6t
Xbit_r236_c60 bl[60] br[60] wl[236] vdd gnd cell_6t
Xbit_r237_c60 bl[60] br[60] wl[237] vdd gnd cell_6t
Xbit_r238_c60 bl[60] br[60] wl[238] vdd gnd cell_6t
Xbit_r239_c60 bl[60] br[60] wl[239] vdd gnd cell_6t
Xbit_r240_c60 bl[60] br[60] wl[240] vdd gnd cell_6t
Xbit_r241_c60 bl[60] br[60] wl[241] vdd gnd cell_6t
Xbit_r242_c60 bl[60] br[60] wl[242] vdd gnd cell_6t
Xbit_r243_c60 bl[60] br[60] wl[243] vdd gnd cell_6t
Xbit_r244_c60 bl[60] br[60] wl[244] vdd gnd cell_6t
Xbit_r245_c60 bl[60] br[60] wl[245] vdd gnd cell_6t
Xbit_r246_c60 bl[60] br[60] wl[246] vdd gnd cell_6t
Xbit_r247_c60 bl[60] br[60] wl[247] vdd gnd cell_6t
Xbit_r248_c60 bl[60] br[60] wl[248] vdd gnd cell_6t
Xbit_r249_c60 bl[60] br[60] wl[249] vdd gnd cell_6t
Xbit_r250_c60 bl[60] br[60] wl[250] vdd gnd cell_6t
Xbit_r251_c60 bl[60] br[60] wl[251] vdd gnd cell_6t
Xbit_r252_c60 bl[60] br[60] wl[252] vdd gnd cell_6t
Xbit_r253_c60 bl[60] br[60] wl[253] vdd gnd cell_6t
Xbit_r254_c60 bl[60] br[60] wl[254] vdd gnd cell_6t
Xbit_r255_c60 bl[60] br[60] wl[255] vdd gnd cell_6t
Xbit_r0_c61 bl[61] br[61] wl[0] vdd gnd cell_6t
Xbit_r1_c61 bl[61] br[61] wl[1] vdd gnd cell_6t
Xbit_r2_c61 bl[61] br[61] wl[2] vdd gnd cell_6t
Xbit_r3_c61 bl[61] br[61] wl[3] vdd gnd cell_6t
Xbit_r4_c61 bl[61] br[61] wl[4] vdd gnd cell_6t
Xbit_r5_c61 bl[61] br[61] wl[5] vdd gnd cell_6t
Xbit_r6_c61 bl[61] br[61] wl[6] vdd gnd cell_6t
Xbit_r7_c61 bl[61] br[61] wl[7] vdd gnd cell_6t
Xbit_r8_c61 bl[61] br[61] wl[8] vdd gnd cell_6t
Xbit_r9_c61 bl[61] br[61] wl[9] vdd gnd cell_6t
Xbit_r10_c61 bl[61] br[61] wl[10] vdd gnd cell_6t
Xbit_r11_c61 bl[61] br[61] wl[11] vdd gnd cell_6t
Xbit_r12_c61 bl[61] br[61] wl[12] vdd gnd cell_6t
Xbit_r13_c61 bl[61] br[61] wl[13] vdd gnd cell_6t
Xbit_r14_c61 bl[61] br[61] wl[14] vdd gnd cell_6t
Xbit_r15_c61 bl[61] br[61] wl[15] vdd gnd cell_6t
Xbit_r16_c61 bl[61] br[61] wl[16] vdd gnd cell_6t
Xbit_r17_c61 bl[61] br[61] wl[17] vdd gnd cell_6t
Xbit_r18_c61 bl[61] br[61] wl[18] vdd gnd cell_6t
Xbit_r19_c61 bl[61] br[61] wl[19] vdd gnd cell_6t
Xbit_r20_c61 bl[61] br[61] wl[20] vdd gnd cell_6t
Xbit_r21_c61 bl[61] br[61] wl[21] vdd gnd cell_6t
Xbit_r22_c61 bl[61] br[61] wl[22] vdd gnd cell_6t
Xbit_r23_c61 bl[61] br[61] wl[23] vdd gnd cell_6t
Xbit_r24_c61 bl[61] br[61] wl[24] vdd gnd cell_6t
Xbit_r25_c61 bl[61] br[61] wl[25] vdd gnd cell_6t
Xbit_r26_c61 bl[61] br[61] wl[26] vdd gnd cell_6t
Xbit_r27_c61 bl[61] br[61] wl[27] vdd gnd cell_6t
Xbit_r28_c61 bl[61] br[61] wl[28] vdd gnd cell_6t
Xbit_r29_c61 bl[61] br[61] wl[29] vdd gnd cell_6t
Xbit_r30_c61 bl[61] br[61] wl[30] vdd gnd cell_6t
Xbit_r31_c61 bl[61] br[61] wl[31] vdd gnd cell_6t
Xbit_r32_c61 bl[61] br[61] wl[32] vdd gnd cell_6t
Xbit_r33_c61 bl[61] br[61] wl[33] vdd gnd cell_6t
Xbit_r34_c61 bl[61] br[61] wl[34] vdd gnd cell_6t
Xbit_r35_c61 bl[61] br[61] wl[35] vdd gnd cell_6t
Xbit_r36_c61 bl[61] br[61] wl[36] vdd gnd cell_6t
Xbit_r37_c61 bl[61] br[61] wl[37] vdd gnd cell_6t
Xbit_r38_c61 bl[61] br[61] wl[38] vdd gnd cell_6t
Xbit_r39_c61 bl[61] br[61] wl[39] vdd gnd cell_6t
Xbit_r40_c61 bl[61] br[61] wl[40] vdd gnd cell_6t
Xbit_r41_c61 bl[61] br[61] wl[41] vdd gnd cell_6t
Xbit_r42_c61 bl[61] br[61] wl[42] vdd gnd cell_6t
Xbit_r43_c61 bl[61] br[61] wl[43] vdd gnd cell_6t
Xbit_r44_c61 bl[61] br[61] wl[44] vdd gnd cell_6t
Xbit_r45_c61 bl[61] br[61] wl[45] vdd gnd cell_6t
Xbit_r46_c61 bl[61] br[61] wl[46] vdd gnd cell_6t
Xbit_r47_c61 bl[61] br[61] wl[47] vdd gnd cell_6t
Xbit_r48_c61 bl[61] br[61] wl[48] vdd gnd cell_6t
Xbit_r49_c61 bl[61] br[61] wl[49] vdd gnd cell_6t
Xbit_r50_c61 bl[61] br[61] wl[50] vdd gnd cell_6t
Xbit_r51_c61 bl[61] br[61] wl[51] vdd gnd cell_6t
Xbit_r52_c61 bl[61] br[61] wl[52] vdd gnd cell_6t
Xbit_r53_c61 bl[61] br[61] wl[53] vdd gnd cell_6t
Xbit_r54_c61 bl[61] br[61] wl[54] vdd gnd cell_6t
Xbit_r55_c61 bl[61] br[61] wl[55] vdd gnd cell_6t
Xbit_r56_c61 bl[61] br[61] wl[56] vdd gnd cell_6t
Xbit_r57_c61 bl[61] br[61] wl[57] vdd gnd cell_6t
Xbit_r58_c61 bl[61] br[61] wl[58] vdd gnd cell_6t
Xbit_r59_c61 bl[61] br[61] wl[59] vdd gnd cell_6t
Xbit_r60_c61 bl[61] br[61] wl[60] vdd gnd cell_6t
Xbit_r61_c61 bl[61] br[61] wl[61] vdd gnd cell_6t
Xbit_r62_c61 bl[61] br[61] wl[62] vdd gnd cell_6t
Xbit_r63_c61 bl[61] br[61] wl[63] vdd gnd cell_6t
Xbit_r64_c61 bl[61] br[61] wl[64] vdd gnd cell_6t
Xbit_r65_c61 bl[61] br[61] wl[65] vdd gnd cell_6t
Xbit_r66_c61 bl[61] br[61] wl[66] vdd gnd cell_6t
Xbit_r67_c61 bl[61] br[61] wl[67] vdd gnd cell_6t
Xbit_r68_c61 bl[61] br[61] wl[68] vdd gnd cell_6t
Xbit_r69_c61 bl[61] br[61] wl[69] vdd gnd cell_6t
Xbit_r70_c61 bl[61] br[61] wl[70] vdd gnd cell_6t
Xbit_r71_c61 bl[61] br[61] wl[71] vdd gnd cell_6t
Xbit_r72_c61 bl[61] br[61] wl[72] vdd gnd cell_6t
Xbit_r73_c61 bl[61] br[61] wl[73] vdd gnd cell_6t
Xbit_r74_c61 bl[61] br[61] wl[74] vdd gnd cell_6t
Xbit_r75_c61 bl[61] br[61] wl[75] vdd gnd cell_6t
Xbit_r76_c61 bl[61] br[61] wl[76] vdd gnd cell_6t
Xbit_r77_c61 bl[61] br[61] wl[77] vdd gnd cell_6t
Xbit_r78_c61 bl[61] br[61] wl[78] vdd gnd cell_6t
Xbit_r79_c61 bl[61] br[61] wl[79] vdd gnd cell_6t
Xbit_r80_c61 bl[61] br[61] wl[80] vdd gnd cell_6t
Xbit_r81_c61 bl[61] br[61] wl[81] vdd gnd cell_6t
Xbit_r82_c61 bl[61] br[61] wl[82] vdd gnd cell_6t
Xbit_r83_c61 bl[61] br[61] wl[83] vdd gnd cell_6t
Xbit_r84_c61 bl[61] br[61] wl[84] vdd gnd cell_6t
Xbit_r85_c61 bl[61] br[61] wl[85] vdd gnd cell_6t
Xbit_r86_c61 bl[61] br[61] wl[86] vdd gnd cell_6t
Xbit_r87_c61 bl[61] br[61] wl[87] vdd gnd cell_6t
Xbit_r88_c61 bl[61] br[61] wl[88] vdd gnd cell_6t
Xbit_r89_c61 bl[61] br[61] wl[89] vdd gnd cell_6t
Xbit_r90_c61 bl[61] br[61] wl[90] vdd gnd cell_6t
Xbit_r91_c61 bl[61] br[61] wl[91] vdd gnd cell_6t
Xbit_r92_c61 bl[61] br[61] wl[92] vdd gnd cell_6t
Xbit_r93_c61 bl[61] br[61] wl[93] vdd gnd cell_6t
Xbit_r94_c61 bl[61] br[61] wl[94] vdd gnd cell_6t
Xbit_r95_c61 bl[61] br[61] wl[95] vdd gnd cell_6t
Xbit_r96_c61 bl[61] br[61] wl[96] vdd gnd cell_6t
Xbit_r97_c61 bl[61] br[61] wl[97] vdd gnd cell_6t
Xbit_r98_c61 bl[61] br[61] wl[98] vdd gnd cell_6t
Xbit_r99_c61 bl[61] br[61] wl[99] vdd gnd cell_6t
Xbit_r100_c61 bl[61] br[61] wl[100] vdd gnd cell_6t
Xbit_r101_c61 bl[61] br[61] wl[101] vdd gnd cell_6t
Xbit_r102_c61 bl[61] br[61] wl[102] vdd gnd cell_6t
Xbit_r103_c61 bl[61] br[61] wl[103] vdd gnd cell_6t
Xbit_r104_c61 bl[61] br[61] wl[104] vdd gnd cell_6t
Xbit_r105_c61 bl[61] br[61] wl[105] vdd gnd cell_6t
Xbit_r106_c61 bl[61] br[61] wl[106] vdd gnd cell_6t
Xbit_r107_c61 bl[61] br[61] wl[107] vdd gnd cell_6t
Xbit_r108_c61 bl[61] br[61] wl[108] vdd gnd cell_6t
Xbit_r109_c61 bl[61] br[61] wl[109] vdd gnd cell_6t
Xbit_r110_c61 bl[61] br[61] wl[110] vdd gnd cell_6t
Xbit_r111_c61 bl[61] br[61] wl[111] vdd gnd cell_6t
Xbit_r112_c61 bl[61] br[61] wl[112] vdd gnd cell_6t
Xbit_r113_c61 bl[61] br[61] wl[113] vdd gnd cell_6t
Xbit_r114_c61 bl[61] br[61] wl[114] vdd gnd cell_6t
Xbit_r115_c61 bl[61] br[61] wl[115] vdd gnd cell_6t
Xbit_r116_c61 bl[61] br[61] wl[116] vdd gnd cell_6t
Xbit_r117_c61 bl[61] br[61] wl[117] vdd gnd cell_6t
Xbit_r118_c61 bl[61] br[61] wl[118] vdd gnd cell_6t
Xbit_r119_c61 bl[61] br[61] wl[119] vdd gnd cell_6t
Xbit_r120_c61 bl[61] br[61] wl[120] vdd gnd cell_6t
Xbit_r121_c61 bl[61] br[61] wl[121] vdd gnd cell_6t
Xbit_r122_c61 bl[61] br[61] wl[122] vdd gnd cell_6t
Xbit_r123_c61 bl[61] br[61] wl[123] vdd gnd cell_6t
Xbit_r124_c61 bl[61] br[61] wl[124] vdd gnd cell_6t
Xbit_r125_c61 bl[61] br[61] wl[125] vdd gnd cell_6t
Xbit_r126_c61 bl[61] br[61] wl[126] vdd gnd cell_6t
Xbit_r127_c61 bl[61] br[61] wl[127] vdd gnd cell_6t
Xbit_r128_c61 bl[61] br[61] wl[128] vdd gnd cell_6t
Xbit_r129_c61 bl[61] br[61] wl[129] vdd gnd cell_6t
Xbit_r130_c61 bl[61] br[61] wl[130] vdd gnd cell_6t
Xbit_r131_c61 bl[61] br[61] wl[131] vdd gnd cell_6t
Xbit_r132_c61 bl[61] br[61] wl[132] vdd gnd cell_6t
Xbit_r133_c61 bl[61] br[61] wl[133] vdd gnd cell_6t
Xbit_r134_c61 bl[61] br[61] wl[134] vdd gnd cell_6t
Xbit_r135_c61 bl[61] br[61] wl[135] vdd gnd cell_6t
Xbit_r136_c61 bl[61] br[61] wl[136] vdd gnd cell_6t
Xbit_r137_c61 bl[61] br[61] wl[137] vdd gnd cell_6t
Xbit_r138_c61 bl[61] br[61] wl[138] vdd gnd cell_6t
Xbit_r139_c61 bl[61] br[61] wl[139] vdd gnd cell_6t
Xbit_r140_c61 bl[61] br[61] wl[140] vdd gnd cell_6t
Xbit_r141_c61 bl[61] br[61] wl[141] vdd gnd cell_6t
Xbit_r142_c61 bl[61] br[61] wl[142] vdd gnd cell_6t
Xbit_r143_c61 bl[61] br[61] wl[143] vdd gnd cell_6t
Xbit_r144_c61 bl[61] br[61] wl[144] vdd gnd cell_6t
Xbit_r145_c61 bl[61] br[61] wl[145] vdd gnd cell_6t
Xbit_r146_c61 bl[61] br[61] wl[146] vdd gnd cell_6t
Xbit_r147_c61 bl[61] br[61] wl[147] vdd gnd cell_6t
Xbit_r148_c61 bl[61] br[61] wl[148] vdd gnd cell_6t
Xbit_r149_c61 bl[61] br[61] wl[149] vdd gnd cell_6t
Xbit_r150_c61 bl[61] br[61] wl[150] vdd gnd cell_6t
Xbit_r151_c61 bl[61] br[61] wl[151] vdd gnd cell_6t
Xbit_r152_c61 bl[61] br[61] wl[152] vdd gnd cell_6t
Xbit_r153_c61 bl[61] br[61] wl[153] vdd gnd cell_6t
Xbit_r154_c61 bl[61] br[61] wl[154] vdd gnd cell_6t
Xbit_r155_c61 bl[61] br[61] wl[155] vdd gnd cell_6t
Xbit_r156_c61 bl[61] br[61] wl[156] vdd gnd cell_6t
Xbit_r157_c61 bl[61] br[61] wl[157] vdd gnd cell_6t
Xbit_r158_c61 bl[61] br[61] wl[158] vdd gnd cell_6t
Xbit_r159_c61 bl[61] br[61] wl[159] vdd gnd cell_6t
Xbit_r160_c61 bl[61] br[61] wl[160] vdd gnd cell_6t
Xbit_r161_c61 bl[61] br[61] wl[161] vdd gnd cell_6t
Xbit_r162_c61 bl[61] br[61] wl[162] vdd gnd cell_6t
Xbit_r163_c61 bl[61] br[61] wl[163] vdd gnd cell_6t
Xbit_r164_c61 bl[61] br[61] wl[164] vdd gnd cell_6t
Xbit_r165_c61 bl[61] br[61] wl[165] vdd gnd cell_6t
Xbit_r166_c61 bl[61] br[61] wl[166] vdd gnd cell_6t
Xbit_r167_c61 bl[61] br[61] wl[167] vdd gnd cell_6t
Xbit_r168_c61 bl[61] br[61] wl[168] vdd gnd cell_6t
Xbit_r169_c61 bl[61] br[61] wl[169] vdd gnd cell_6t
Xbit_r170_c61 bl[61] br[61] wl[170] vdd gnd cell_6t
Xbit_r171_c61 bl[61] br[61] wl[171] vdd gnd cell_6t
Xbit_r172_c61 bl[61] br[61] wl[172] vdd gnd cell_6t
Xbit_r173_c61 bl[61] br[61] wl[173] vdd gnd cell_6t
Xbit_r174_c61 bl[61] br[61] wl[174] vdd gnd cell_6t
Xbit_r175_c61 bl[61] br[61] wl[175] vdd gnd cell_6t
Xbit_r176_c61 bl[61] br[61] wl[176] vdd gnd cell_6t
Xbit_r177_c61 bl[61] br[61] wl[177] vdd gnd cell_6t
Xbit_r178_c61 bl[61] br[61] wl[178] vdd gnd cell_6t
Xbit_r179_c61 bl[61] br[61] wl[179] vdd gnd cell_6t
Xbit_r180_c61 bl[61] br[61] wl[180] vdd gnd cell_6t
Xbit_r181_c61 bl[61] br[61] wl[181] vdd gnd cell_6t
Xbit_r182_c61 bl[61] br[61] wl[182] vdd gnd cell_6t
Xbit_r183_c61 bl[61] br[61] wl[183] vdd gnd cell_6t
Xbit_r184_c61 bl[61] br[61] wl[184] vdd gnd cell_6t
Xbit_r185_c61 bl[61] br[61] wl[185] vdd gnd cell_6t
Xbit_r186_c61 bl[61] br[61] wl[186] vdd gnd cell_6t
Xbit_r187_c61 bl[61] br[61] wl[187] vdd gnd cell_6t
Xbit_r188_c61 bl[61] br[61] wl[188] vdd gnd cell_6t
Xbit_r189_c61 bl[61] br[61] wl[189] vdd gnd cell_6t
Xbit_r190_c61 bl[61] br[61] wl[190] vdd gnd cell_6t
Xbit_r191_c61 bl[61] br[61] wl[191] vdd gnd cell_6t
Xbit_r192_c61 bl[61] br[61] wl[192] vdd gnd cell_6t
Xbit_r193_c61 bl[61] br[61] wl[193] vdd gnd cell_6t
Xbit_r194_c61 bl[61] br[61] wl[194] vdd gnd cell_6t
Xbit_r195_c61 bl[61] br[61] wl[195] vdd gnd cell_6t
Xbit_r196_c61 bl[61] br[61] wl[196] vdd gnd cell_6t
Xbit_r197_c61 bl[61] br[61] wl[197] vdd gnd cell_6t
Xbit_r198_c61 bl[61] br[61] wl[198] vdd gnd cell_6t
Xbit_r199_c61 bl[61] br[61] wl[199] vdd gnd cell_6t
Xbit_r200_c61 bl[61] br[61] wl[200] vdd gnd cell_6t
Xbit_r201_c61 bl[61] br[61] wl[201] vdd gnd cell_6t
Xbit_r202_c61 bl[61] br[61] wl[202] vdd gnd cell_6t
Xbit_r203_c61 bl[61] br[61] wl[203] vdd gnd cell_6t
Xbit_r204_c61 bl[61] br[61] wl[204] vdd gnd cell_6t
Xbit_r205_c61 bl[61] br[61] wl[205] vdd gnd cell_6t
Xbit_r206_c61 bl[61] br[61] wl[206] vdd gnd cell_6t
Xbit_r207_c61 bl[61] br[61] wl[207] vdd gnd cell_6t
Xbit_r208_c61 bl[61] br[61] wl[208] vdd gnd cell_6t
Xbit_r209_c61 bl[61] br[61] wl[209] vdd gnd cell_6t
Xbit_r210_c61 bl[61] br[61] wl[210] vdd gnd cell_6t
Xbit_r211_c61 bl[61] br[61] wl[211] vdd gnd cell_6t
Xbit_r212_c61 bl[61] br[61] wl[212] vdd gnd cell_6t
Xbit_r213_c61 bl[61] br[61] wl[213] vdd gnd cell_6t
Xbit_r214_c61 bl[61] br[61] wl[214] vdd gnd cell_6t
Xbit_r215_c61 bl[61] br[61] wl[215] vdd gnd cell_6t
Xbit_r216_c61 bl[61] br[61] wl[216] vdd gnd cell_6t
Xbit_r217_c61 bl[61] br[61] wl[217] vdd gnd cell_6t
Xbit_r218_c61 bl[61] br[61] wl[218] vdd gnd cell_6t
Xbit_r219_c61 bl[61] br[61] wl[219] vdd gnd cell_6t
Xbit_r220_c61 bl[61] br[61] wl[220] vdd gnd cell_6t
Xbit_r221_c61 bl[61] br[61] wl[221] vdd gnd cell_6t
Xbit_r222_c61 bl[61] br[61] wl[222] vdd gnd cell_6t
Xbit_r223_c61 bl[61] br[61] wl[223] vdd gnd cell_6t
Xbit_r224_c61 bl[61] br[61] wl[224] vdd gnd cell_6t
Xbit_r225_c61 bl[61] br[61] wl[225] vdd gnd cell_6t
Xbit_r226_c61 bl[61] br[61] wl[226] vdd gnd cell_6t
Xbit_r227_c61 bl[61] br[61] wl[227] vdd gnd cell_6t
Xbit_r228_c61 bl[61] br[61] wl[228] vdd gnd cell_6t
Xbit_r229_c61 bl[61] br[61] wl[229] vdd gnd cell_6t
Xbit_r230_c61 bl[61] br[61] wl[230] vdd gnd cell_6t
Xbit_r231_c61 bl[61] br[61] wl[231] vdd gnd cell_6t
Xbit_r232_c61 bl[61] br[61] wl[232] vdd gnd cell_6t
Xbit_r233_c61 bl[61] br[61] wl[233] vdd gnd cell_6t
Xbit_r234_c61 bl[61] br[61] wl[234] vdd gnd cell_6t
Xbit_r235_c61 bl[61] br[61] wl[235] vdd gnd cell_6t
Xbit_r236_c61 bl[61] br[61] wl[236] vdd gnd cell_6t
Xbit_r237_c61 bl[61] br[61] wl[237] vdd gnd cell_6t
Xbit_r238_c61 bl[61] br[61] wl[238] vdd gnd cell_6t
Xbit_r239_c61 bl[61] br[61] wl[239] vdd gnd cell_6t
Xbit_r240_c61 bl[61] br[61] wl[240] vdd gnd cell_6t
Xbit_r241_c61 bl[61] br[61] wl[241] vdd gnd cell_6t
Xbit_r242_c61 bl[61] br[61] wl[242] vdd gnd cell_6t
Xbit_r243_c61 bl[61] br[61] wl[243] vdd gnd cell_6t
Xbit_r244_c61 bl[61] br[61] wl[244] vdd gnd cell_6t
Xbit_r245_c61 bl[61] br[61] wl[245] vdd gnd cell_6t
Xbit_r246_c61 bl[61] br[61] wl[246] vdd gnd cell_6t
Xbit_r247_c61 bl[61] br[61] wl[247] vdd gnd cell_6t
Xbit_r248_c61 bl[61] br[61] wl[248] vdd gnd cell_6t
Xbit_r249_c61 bl[61] br[61] wl[249] vdd gnd cell_6t
Xbit_r250_c61 bl[61] br[61] wl[250] vdd gnd cell_6t
Xbit_r251_c61 bl[61] br[61] wl[251] vdd gnd cell_6t
Xbit_r252_c61 bl[61] br[61] wl[252] vdd gnd cell_6t
Xbit_r253_c61 bl[61] br[61] wl[253] vdd gnd cell_6t
Xbit_r254_c61 bl[61] br[61] wl[254] vdd gnd cell_6t
Xbit_r255_c61 bl[61] br[61] wl[255] vdd gnd cell_6t
Xbit_r0_c62 bl[62] br[62] wl[0] vdd gnd cell_6t
Xbit_r1_c62 bl[62] br[62] wl[1] vdd gnd cell_6t
Xbit_r2_c62 bl[62] br[62] wl[2] vdd gnd cell_6t
Xbit_r3_c62 bl[62] br[62] wl[3] vdd gnd cell_6t
Xbit_r4_c62 bl[62] br[62] wl[4] vdd gnd cell_6t
Xbit_r5_c62 bl[62] br[62] wl[5] vdd gnd cell_6t
Xbit_r6_c62 bl[62] br[62] wl[6] vdd gnd cell_6t
Xbit_r7_c62 bl[62] br[62] wl[7] vdd gnd cell_6t
Xbit_r8_c62 bl[62] br[62] wl[8] vdd gnd cell_6t
Xbit_r9_c62 bl[62] br[62] wl[9] vdd gnd cell_6t
Xbit_r10_c62 bl[62] br[62] wl[10] vdd gnd cell_6t
Xbit_r11_c62 bl[62] br[62] wl[11] vdd gnd cell_6t
Xbit_r12_c62 bl[62] br[62] wl[12] vdd gnd cell_6t
Xbit_r13_c62 bl[62] br[62] wl[13] vdd gnd cell_6t
Xbit_r14_c62 bl[62] br[62] wl[14] vdd gnd cell_6t
Xbit_r15_c62 bl[62] br[62] wl[15] vdd gnd cell_6t
Xbit_r16_c62 bl[62] br[62] wl[16] vdd gnd cell_6t
Xbit_r17_c62 bl[62] br[62] wl[17] vdd gnd cell_6t
Xbit_r18_c62 bl[62] br[62] wl[18] vdd gnd cell_6t
Xbit_r19_c62 bl[62] br[62] wl[19] vdd gnd cell_6t
Xbit_r20_c62 bl[62] br[62] wl[20] vdd gnd cell_6t
Xbit_r21_c62 bl[62] br[62] wl[21] vdd gnd cell_6t
Xbit_r22_c62 bl[62] br[62] wl[22] vdd gnd cell_6t
Xbit_r23_c62 bl[62] br[62] wl[23] vdd gnd cell_6t
Xbit_r24_c62 bl[62] br[62] wl[24] vdd gnd cell_6t
Xbit_r25_c62 bl[62] br[62] wl[25] vdd gnd cell_6t
Xbit_r26_c62 bl[62] br[62] wl[26] vdd gnd cell_6t
Xbit_r27_c62 bl[62] br[62] wl[27] vdd gnd cell_6t
Xbit_r28_c62 bl[62] br[62] wl[28] vdd gnd cell_6t
Xbit_r29_c62 bl[62] br[62] wl[29] vdd gnd cell_6t
Xbit_r30_c62 bl[62] br[62] wl[30] vdd gnd cell_6t
Xbit_r31_c62 bl[62] br[62] wl[31] vdd gnd cell_6t
Xbit_r32_c62 bl[62] br[62] wl[32] vdd gnd cell_6t
Xbit_r33_c62 bl[62] br[62] wl[33] vdd gnd cell_6t
Xbit_r34_c62 bl[62] br[62] wl[34] vdd gnd cell_6t
Xbit_r35_c62 bl[62] br[62] wl[35] vdd gnd cell_6t
Xbit_r36_c62 bl[62] br[62] wl[36] vdd gnd cell_6t
Xbit_r37_c62 bl[62] br[62] wl[37] vdd gnd cell_6t
Xbit_r38_c62 bl[62] br[62] wl[38] vdd gnd cell_6t
Xbit_r39_c62 bl[62] br[62] wl[39] vdd gnd cell_6t
Xbit_r40_c62 bl[62] br[62] wl[40] vdd gnd cell_6t
Xbit_r41_c62 bl[62] br[62] wl[41] vdd gnd cell_6t
Xbit_r42_c62 bl[62] br[62] wl[42] vdd gnd cell_6t
Xbit_r43_c62 bl[62] br[62] wl[43] vdd gnd cell_6t
Xbit_r44_c62 bl[62] br[62] wl[44] vdd gnd cell_6t
Xbit_r45_c62 bl[62] br[62] wl[45] vdd gnd cell_6t
Xbit_r46_c62 bl[62] br[62] wl[46] vdd gnd cell_6t
Xbit_r47_c62 bl[62] br[62] wl[47] vdd gnd cell_6t
Xbit_r48_c62 bl[62] br[62] wl[48] vdd gnd cell_6t
Xbit_r49_c62 bl[62] br[62] wl[49] vdd gnd cell_6t
Xbit_r50_c62 bl[62] br[62] wl[50] vdd gnd cell_6t
Xbit_r51_c62 bl[62] br[62] wl[51] vdd gnd cell_6t
Xbit_r52_c62 bl[62] br[62] wl[52] vdd gnd cell_6t
Xbit_r53_c62 bl[62] br[62] wl[53] vdd gnd cell_6t
Xbit_r54_c62 bl[62] br[62] wl[54] vdd gnd cell_6t
Xbit_r55_c62 bl[62] br[62] wl[55] vdd gnd cell_6t
Xbit_r56_c62 bl[62] br[62] wl[56] vdd gnd cell_6t
Xbit_r57_c62 bl[62] br[62] wl[57] vdd gnd cell_6t
Xbit_r58_c62 bl[62] br[62] wl[58] vdd gnd cell_6t
Xbit_r59_c62 bl[62] br[62] wl[59] vdd gnd cell_6t
Xbit_r60_c62 bl[62] br[62] wl[60] vdd gnd cell_6t
Xbit_r61_c62 bl[62] br[62] wl[61] vdd gnd cell_6t
Xbit_r62_c62 bl[62] br[62] wl[62] vdd gnd cell_6t
Xbit_r63_c62 bl[62] br[62] wl[63] vdd gnd cell_6t
Xbit_r64_c62 bl[62] br[62] wl[64] vdd gnd cell_6t
Xbit_r65_c62 bl[62] br[62] wl[65] vdd gnd cell_6t
Xbit_r66_c62 bl[62] br[62] wl[66] vdd gnd cell_6t
Xbit_r67_c62 bl[62] br[62] wl[67] vdd gnd cell_6t
Xbit_r68_c62 bl[62] br[62] wl[68] vdd gnd cell_6t
Xbit_r69_c62 bl[62] br[62] wl[69] vdd gnd cell_6t
Xbit_r70_c62 bl[62] br[62] wl[70] vdd gnd cell_6t
Xbit_r71_c62 bl[62] br[62] wl[71] vdd gnd cell_6t
Xbit_r72_c62 bl[62] br[62] wl[72] vdd gnd cell_6t
Xbit_r73_c62 bl[62] br[62] wl[73] vdd gnd cell_6t
Xbit_r74_c62 bl[62] br[62] wl[74] vdd gnd cell_6t
Xbit_r75_c62 bl[62] br[62] wl[75] vdd gnd cell_6t
Xbit_r76_c62 bl[62] br[62] wl[76] vdd gnd cell_6t
Xbit_r77_c62 bl[62] br[62] wl[77] vdd gnd cell_6t
Xbit_r78_c62 bl[62] br[62] wl[78] vdd gnd cell_6t
Xbit_r79_c62 bl[62] br[62] wl[79] vdd gnd cell_6t
Xbit_r80_c62 bl[62] br[62] wl[80] vdd gnd cell_6t
Xbit_r81_c62 bl[62] br[62] wl[81] vdd gnd cell_6t
Xbit_r82_c62 bl[62] br[62] wl[82] vdd gnd cell_6t
Xbit_r83_c62 bl[62] br[62] wl[83] vdd gnd cell_6t
Xbit_r84_c62 bl[62] br[62] wl[84] vdd gnd cell_6t
Xbit_r85_c62 bl[62] br[62] wl[85] vdd gnd cell_6t
Xbit_r86_c62 bl[62] br[62] wl[86] vdd gnd cell_6t
Xbit_r87_c62 bl[62] br[62] wl[87] vdd gnd cell_6t
Xbit_r88_c62 bl[62] br[62] wl[88] vdd gnd cell_6t
Xbit_r89_c62 bl[62] br[62] wl[89] vdd gnd cell_6t
Xbit_r90_c62 bl[62] br[62] wl[90] vdd gnd cell_6t
Xbit_r91_c62 bl[62] br[62] wl[91] vdd gnd cell_6t
Xbit_r92_c62 bl[62] br[62] wl[92] vdd gnd cell_6t
Xbit_r93_c62 bl[62] br[62] wl[93] vdd gnd cell_6t
Xbit_r94_c62 bl[62] br[62] wl[94] vdd gnd cell_6t
Xbit_r95_c62 bl[62] br[62] wl[95] vdd gnd cell_6t
Xbit_r96_c62 bl[62] br[62] wl[96] vdd gnd cell_6t
Xbit_r97_c62 bl[62] br[62] wl[97] vdd gnd cell_6t
Xbit_r98_c62 bl[62] br[62] wl[98] vdd gnd cell_6t
Xbit_r99_c62 bl[62] br[62] wl[99] vdd gnd cell_6t
Xbit_r100_c62 bl[62] br[62] wl[100] vdd gnd cell_6t
Xbit_r101_c62 bl[62] br[62] wl[101] vdd gnd cell_6t
Xbit_r102_c62 bl[62] br[62] wl[102] vdd gnd cell_6t
Xbit_r103_c62 bl[62] br[62] wl[103] vdd gnd cell_6t
Xbit_r104_c62 bl[62] br[62] wl[104] vdd gnd cell_6t
Xbit_r105_c62 bl[62] br[62] wl[105] vdd gnd cell_6t
Xbit_r106_c62 bl[62] br[62] wl[106] vdd gnd cell_6t
Xbit_r107_c62 bl[62] br[62] wl[107] vdd gnd cell_6t
Xbit_r108_c62 bl[62] br[62] wl[108] vdd gnd cell_6t
Xbit_r109_c62 bl[62] br[62] wl[109] vdd gnd cell_6t
Xbit_r110_c62 bl[62] br[62] wl[110] vdd gnd cell_6t
Xbit_r111_c62 bl[62] br[62] wl[111] vdd gnd cell_6t
Xbit_r112_c62 bl[62] br[62] wl[112] vdd gnd cell_6t
Xbit_r113_c62 bl[62] br[62] wl[113] vdd gnd cell_6t
Xbit_r114_c62 bl[62] br[62] wl[114] vdd gnd cell_6t
Xbit_r115_c62 bl[62] br[62] wl[115] vdd gnd cell_6t
Xbit_r116_c62 bl[62] br[62] wl[116] vdd gnd cell_6t
Xbit_r117_c62 bl[62] br[62] wl[117] vdd gnd cell_6t
Xbit_r118_c62 bl[62] br[62] wl[118] vdd gnd cell_6t
Xbit_r119_c62 bl[62] br[62] wl[119] vdd gnd cell_6t
Xbit_r120_c62 bl[62] br[62] wl[120] vdd gnd cell_6t
Xbit_r121_c62 bl[62] br[62] wl[121] vdd gnd cell_6t
Xbit_r122_c62 bl[62] br[62] wl[122] vdd gnd cell_6t
Xbit_r123_c62 bl[62] br[62] wl[123] vdd gnd cell_6t
Xbit_r124_c62 bl[62] br[62] wl[124] vdd gnd cell_6t
Xbit_r125_c62 bl[62] br[62] wl[125] vdd gnd cell_6t
Xbit_r126_c62 bl[62] br[62] wl[126] vdd gnd cell_6t
Xbit_r127_c62 bl[62] br[62] wl[127] vdd gnd cell_6t
Xbit_r128_c62 bl[62] br[62] wl[128] vdd gnd cell_6t
Xbit_r129_c62 bl[62] br[62] wl[129] vdd gnd cell_6t
Xbit_r130_c62 bl[62] br[62] wl[130] vdd gnd cell_6t
Xbit_r131_c62 bl[62] br[62] wl[131] vdd gnd cell_6t
Xbit_r132_c62 bl[62] br[62] wl[132] vdd gnd cell_6t
Xbit_r133_c62 bl[62] br[62] wl[133] vdd gnd cell_6t
Xbit_r134_c62 bl[62] br[62] wl[134] vdd gnd cell_6t
Xbit_r135_c62 bl[62] br[62] wl[135] vdd gnd cell_6t
Xbit_r136_c62 bl[62] br[62] wl[136] vdd gnd cell_6t
Xbit_r137_c62 bl[62] br[62] wl[137] vdd gnd cell_6t
Xbit_r138_c62 bl[62] br[62] wl[138] vdd gnd cell_6t
Xbit_r139_c62 bl[62] br[62] wl[139] vdd gnd cell_6t
Xbit_r140_c62 bl[62] br[62] wl[140] vdd gnd cell_6t
Xbit_r141_c62 bl[62] br[62] wl[141] vdd gnd cell_6t
Xbit_r142_c62 bl[62] br[62] wl[142] vdd gnd cell_6t
Xbit_r143_c62 bl[62] br[62] wl[143] vdd gnd cell_6t
Xbit_r144_c62 bl[62] br[62] wl[144] vdd gnd cell_6t
Xbit_r145_c62 bl[62] br[62] wl[145] vdd gnd cell_6t
Xbit_r146_c62 bl[62] br[62] wl[146] vdd gnd cell_6t
Xbit_r147_c62 bl[62] br[62] wl[147] vdd gnd cell_6t
Xbit_r148_c62 bl[62] br[62] wl[148] vdd gnd cell_6t
Xbit_r149_c62 bl[62] br[62] wl[149] vdd gnd cell_6t
Xbit_r150_c62 bl[62] br[62] wl[150] vdd gnd cell_6t
Xbit_r151_c62 bl[62] br[62] wl[151] vdd gnd cell_6t
Xbit_r152_c62 bl[62] br[62] wl[152] vdd gnd cell_6t
Xbit_r153_c62 bl[62] br[62] wl[153] vdd gnd cell_6t
Xbit_r154_c62 bl[62] br[62] wl[154] vdd gnd cell_6t
Xbit_r155_c62 bl[62] br[62] wl[155] vdd gnd cell_6t
Xbit_r156_c62 bl[62] br[62] wl[156] vdd gnd cell_6t
Xbit_r157_c62 bl[62] br[62] wl[157] vdd gnd cell_6t
Xbit_r158_c62 bl[62] br[62] wl[158] vdd gnd cell_6t
Xbit_r159_c62 bl[62] br[62] wl[159] vdd gnd cell_6t
Xbit_r160_c62 bl[62] br[62] wl[160] vdd gnd cell_6t
Xbit_r161_c62 bl[62] br[62] wl[161] vdd gnd cell_6t
Xbit_r162_c62 bl[62] br[62] wl[162] vdd gnd cell_6t
Xbit_r163_c62 bl[62] br[62] wl[163] vdd gnd cell_6t
Xbit_r164_c62 bl[62] br[62] wl[164] vdd gnd cell_6t
Xbit_r165_c62 bl[62] br[62] wl[165] vdd gnd cell_6t
Xbit_r166_c62 bl[62] br[62] wl[166] vdd gnd cell_6t
Xbit_r167_c62 bl[62] br[62] wl[167] vdd gnd cell_6t
Xbit_r168_c62 bl[62] br[62] wl[168] vdd gnd cell_6t
Xbit_r169_c62 bl[62] br[62] wl[169] vdd gnd cell_6t
Xbit_r170_c62 bl[62] br[62] wl[170] vdd gnd cell_6t
Xbit_r171_c62 bl[62] br[62] wl[171] vdd gnd cell_6t
Xbit_r172_c62 bl[62] br[62] wl[172] vdd gnd cell_6t
Xbit_r173_c62 bl[62] br[62] wl[173] vdd gnd cell_6t
Xbit_r174_c62 bl[62] br[62] wl[174] vdd gnd cell_6t
Xbit_r175_c62 bl[62] br[62] wl[175] vdd gnd cell_6t
Xbit_r176_c62 bl[62] br[62] wl[176] vdd gnd cell_6t
Xbit_r177_c62 bl[62] br[62] wl[177] vdd gnd cell_6t
Xbit_r178_c62 bl[62] br[62] wl[178] vdd gnd cell_6t
Xbit_r179_c62 bl[62] br[62] wl[179] vdd gnd cell_6t
Xbit_r180_c62 bl[62] br[62] wl[180] vdd gnd cell_6t
Xbit_r181_c62 bl[62] br[62] wl[181] vdd gnd cell_6t
Xbit_r182_c62 bl[62] br[62] wl[182] vdd gnd cell_6t
Xbit_r183_c62 bl[62] br[62] wl[183] vdd gnd cell_6t
Xbit_r184_c62 bl[62] br[62] wl[184] vdd gnd cell_6t
Xbit_r185_c62 bl[62] br[62] wl[185] vdd gnd cell_6t
Xbit_r186_c62 bl[62] br[62] wl[186] vdd gnd cell_6t
Xbit_r187_c62 bl[62] br[62] wl[187] vdd gnd cell_6t
Xbit_r188_c62 bl[62] br[62] wl[188] vdd gnd cell_6t
Xbit_r189_c62 bl[62] br[62] wl[189] vdd gnd cell_6t
Xbit_r190_c62 bl[62] br[62] wl[190] vdd gnd cell_6t
Xbit_r191_c62 bl[62] br[62] wl[191] vdd gnd cell_6t
Xbit_r192_c62 bl[62] br[62] wl[192] vdd gnd cell_6t
Xbit_r193_c62 bl[62] br[62] wl[193] vdd gnd cell_6t
Xbit_r194_c62 bl[62] br[62] wl[194] vdd gnd cell_6t
Xbit_r195_c62 bl[62] br[62] wl[195] vdd gnd cell_6t
Xbit_r196_c62 bl[62] br[62] wl[196] vdd gnd cell_6t
Xbit_r197_c62 bl[62] br[62] wl[197] vdd gnd cell_6t
Xbit_r198_c62 bl[62] br[62] wl[198] vdd gnd cell_6t
Xbit_r199_c62 bl[62] br[62] wl[199] vdd gnd cell_6t
Xbit_r200_c62 bl[62] br[62] wl[200] vdd gnd cell_6t
Xbit_r201_c62 bl[62] br[62] wl[201] vdd gnd cell_6t
Xbit_r202_c62 bl[62] br[62] wl[202] vdd gnd cell_6t
Xbit_r203_c62 bl[62] br[62] wl[203] vdd gnd cell_6t
Xbit_r204_c62 bl[62] br[62] wl[204] vdd gnd cell_6t
Xbit_r205_c62 bl[62] br[62] wl[205] vdd gnd cell_6t
Xbit_r206_c62 bl[62] br[62] wl[206] vdd gnd cell_6t
Xbit_r207_c62 bl[62] br[62] wl[207] vdd gnd cell_6t
Xbit_r208_c62 bl[62] br[62] wl[208] vdd gnd cell_6t
Xbit_r209_c62 bl[62] br[62] wl[209] vdd gnd cell_6t
Xbit_r210_c62 bl[62] br[62] wl[210] vdd gnd cell_6t
Xbit_r211_c62 bl[62] br[62] wl[211] vdd gnd cell_6t
Xbit_r212_c62 bl[62] br[62] wl[212] vdd gnd cell_6t
Xbit_r213_c62 bl[62] br[62] wl[213] vdd gnd cell_6t
Xbit_r214_c62 bl[62] br[62] wl[214] vdd gnd cell_6t
Xbit_r215_c62 bl[62] br[62] wl[215] vdd gnd cell_6t
Xbit_r216_c62 bl[62] br[62] wl[216] vdd gnd cell_6t
Xbit_r217_c62 bl[62] br[62] wl[217] vdd gnd cell_6t
Xbit_r218_c62 bl[62] br[62] wl[218] vdd gnd cell_6t
Xbit_r219_c62 bl[62] br[62] wl[219] vdd gnd cell_6t
Xbit_r220_c62 bl[62] br[62] wl[220] vdd gnd cell_6t
Xbit_r221_c62 bl[62] br[62] wl[221] vdd gnd cell_6t
Xbit_r222_c62 bl[62] br[62] wl[222] vdd gnd cell_6t
Xbit_r223_c62 bl[62] br[62] wl[223] vdd gnd cell_6t
Xbit_r224_c62 bl[62] br[62] wl[224] vdd gnd cell_6t
Xbit_r225_c62 bl[62] br[62] wl[225] vdd gnd cell_6t
Xbit_r226_c62 bl[62] br[62] wl[226] vdd gnd cell_6t
Xbit_r227_c62 bl[62] br[62] wl[227] vdd gnd cell_6t
Xbit_r228_c62 bl[62] br[62] wl[228] vdd gnd cell_6t
Xbit_r229_c62 bl[62] br[62] wl[229] vdd gnd cell_6t
Xbit_r230_c62 bl[62] br[62] wl[230] vdd gnd cell_6t
Xbit_r231_c62 bl[62] br[62] wl[231] vdd gnd cell_6t
Xbit_r232_c62 bl[62] br[62] wl[232] vdd gnd cell_6t
Xbit_r233_c62 bl[62] br[62] wl[233] vdd gnd cell_6t
Xbit_r234_c62 bl[62] br[62] wl[234] vdd gnd cell_6t
Xbit_r235_c62 bl[62] br[62] wl[235] vdd gnd cell_6t
Xbit_r236_c62 bl[62] br[62] wl[236] vdd gnd cell_6t
Xbit_r237_c62 bl[62] br[62] wl[237] vdd gnd cell_6t
Xbit_r238_c62 bl[62] br[62] wl[238] vdd gnd cell_6t
Xbit_r239_c62 bl[62] br[62] wl[239] vdd gnd cell_6t
Xbit_r240_c62 bl[62] br[62] wl[240] vdd gnd cell_6t
Xbit_r241_c62 bl[62] br[62] wl[241] vdd gnd cell_6t
Xbit_r242_c62 bl[62] br[62] wl[242] vdd gnd cell_6t
Xbit_r243_c62 bl[62] br[62] wl[243] vdd gnd cell_6t
Xbit_r244_c62 bl[62] br[62] wl[244] vdd gnd cell_6t
Xbit_r245_c62 bl[62] br[62] wl[245] vdd gnd cell_6t
Xbit_r246_c62 bl[62] br[62] wl[246] vdd gnd cell_6t
Xbit_r247_c62 bl[62] br[62] wl[247] vdd gnd cell_6t
Xbit_r248_c62 bl[62] br[62] wl[248] vdd gnd cell_6t
Xbit_r249_c62 bl[62] br[62] wl[249] vdd gnd cell_6t
Xbit_r250_c62 bl[62] br[62] wl[250] vdd gnd cell_6t
Xbit_r251_c62 bl[62] br[62] wl[251] vdd gnd cell_6t
Xbit_r252_c62 bl[62] br[62] wl[252] vdd gnd cell_6t
Xbit_r253_c62 bl[62] br[62] wl[253] vdd gnd cell_6t
Xbit_r254_c62 bl[62] br[62] wl[254] vdd gnd cell_6t
Xbit_r255_c62 bl[62] br[62] wl[255] vdd gnd cell_6t
Xbit_r0_c63 bl[63] br[63] wl[0] vdd gnd cell_6t
Xbit_r1_c63 bl[63] br[63] wl[1] vdd gnd cell_6t
Xbit_r2_c63 bl[63] br[63] wl[2] vdd gnd cell_6t
Xbit_r3_c63 bl[63] br[63] wl[3] vdd gnd cell_6t
Xbit_r4_c63 bl[63] br[63] wl[4] vdd gnd cell_6t
Xbit_r5_c63 bl[63] br[63] wl[5] vdd gnd cell_6t
Xbit_r6_c63 bl[63] br[63] wl[6] vdd gnd cell_6t
Xbit_r7_c63 bl[63] br[63] wl[7] vdd gnd cell_6t
Xbit_r8_c63 bl[63] br[63] wl[8] vdd gnd cell_6t
Xbit_r9_c63 bl[63] br[63] wl[9] vdd gnd cell_6t
Xbit_r10_c63 bl[63] br[63] wl[10] vdd gnd cell_6t
Xbit_r11_c63 bl[63] br[63] wl[11] vdd gnd cell_6t
Xbit_r12_c63 bl[63] br[63] wl[12] vdd gnd cell_6t
Xbit_r13_c63 bl[63] br[63] wl[13] vdd gnd cell_6t
Xbit_r14_c63 bl[63] br[63] wl[14] vdd gnd cell_6t
Xbit_r15_c63 bl[63] br[63] wl[15] vdd gnd cell_6t
Xbit_r16_c63 bl[63] br[63] wl[16] vdd gnd cell_6t
Xbit_r17_c63 bl[63] br[63] wl[17] vdd gnd cell_6t
Xbit_r18_c63 bl[63] br[63] wl[18] vdd gnd cell_6t
Xbit_r19_c63 bl[63] br[63] wl[19] vdd gnd cell_6t
Xbit_r20_c63 bl[63] br[63] wl[20] vdd gnd cell_6t
Xbit_r21_c63 bl[63] br[63] wl[21] vdd gnd cell_6t
Xbit_r22_c63 bl[63] br[63] wl[22] vdd gnd cell_6t
Xbit_r23_c63 bl[63] br[63] wl[23] vdd gnd cell_6t
Xbit_r24_c63 bl[63] br[63] wl[24] vdd gnd cell_6t
Xbit_r25_c63 bl[63] br[63] wl[25] vdd gnd cell_6t
Xbit_r26_c63 bl[63] br[63] wl[26] vdd gnd cell_6t
Xbit_r27_c63 bl[63] br[63] wl[27] vdd gnd cell_6t
Xbit_r28_c63 bl[63] br[63] wl[28] vdd gnd cell_6t
Xbit_r29_c63 bl[63] br[63] wl[29] vdd gnd cell_6t
Xbit_r30_c63 bl[63] br[63] wl[30] vdd gnd cell_6t
Xbit_r31_c63 bl[63] br[63] wl[31] vdd gnd cell_6t
Xbit_r32_c63 bl[63] br[63] wl[32] vdd gnd cell_6t
Xbit_r33_c63 bl[63] br[63] wl[33] vdd gnd cell_6t
Xbit_r34_c63 bl[63] br[63] wl[34] vdd gnd cell_6t
Xbit_r35_c63 bl[63] br[63] wl[35] vdd gnd cell_6t
Xbit_r36_c63 bl[63] br[63] wl[36] vdd gnd cell_6t
Xbit_r37_c63 bl[63] br[63] wl[37] vdd gnd cell_6t
Xbit_r38_c63 bl[63] br[63] wl[38] vdd gnd cell_6t
Xbit_r39_c63 bl[63] br[63] wl[39] vdd gnd cell_6t
Xbit_r40_c63 bl[63] br[63] wl[40] vdd gnd cell_6t
Xbit_r41_c63 bl[63] br[63] wl[41] vdd gnd cell_6t
Xbit_r42_c63 bl[63] br[63] wl[42] vdd gnd cell_6t
Xbit_r43_c63 bl[63] br[63] wl[43] vdd gnd cell_6t
Xbit_r44_c63 bl[63] br[63] wl[44] vdd gnd cell_6t
Xbit_r45_c63 bl[63] br[63] wl[45] vdd gnd cell_6t
Xbit_r46_c63 bl[63] br[63] wl[46] vdd gnd cell_6t
Xbit_r47_c63 bl[63] br[63] wl[47] vdd gnd cell_6t
Xbit_r48_c63 bl[63] br[63] wl[48] vdd gnd cell_6t
Xbit_r49_c63 bl[63] br[63] wl[49] vdd gnd cell_6t
Xbit_r50_c63 bl[63] br[63] wl[50] vdd gnd cell_6t
Xbit_r51_c63 bl[63] br[63] wl[51] vdd gnd cell_6t
Xbit_r52_c63 bl[63] br[63] wl[52] vdd gnd cell_6t
Xbit_r53_c63 bl[63] br[63] wl[53] vdd gnd cell_6t
Xbit_r54_c63 bl[63] br[63] wl[54] vdd gnd cell_6t
Xbit_r55_c63 bl[63] br[63] wl[55] vdd gnd cell_6t
Xbit_r56_c63 bl[63] br[63] wl[56] vdd gnd cell_6t
Xbit_r57_c63 bl[63] br[63] wl[57] vdd gnd cell_6t
Xbit_r58_c63 bl[63] br[63] wl[58] vdd gnd cell_6t
Xbit_r59_c63 bl[63] br[63] wl[59] vdd gnd cell_6t
Xbit_r60_c63 bl[63] br[63] wl[60] vdd gnd cell_6t
Xbit_r61_c63 bl[63] br[63] wl[61] vdd gnd cell_6t
Xbit_r62_c63 bl[63] br[63] wl[62] vdd gnd cell_6t
Xbit_r63_c63 bl[63] br[63] wl[63] vdd gnd cell_6t
Xbit_r64_c63 bl[63] br[63] wl[64] vdd gnd cell_6t
Xbit_r65_c63 bl[63] br[63] wl[65] vdd gnd cell_6t
Xbit_r66_c63 bl[63] br[63] wl[66] vdd gnd cell_6t
Xbit_r67_c63 bl[63] br[63] wl[67] vdd gnd cell_6t
Xbit_r68_c63 bl[63] br[63] wl[68] vdd gnd cell_6t
Xbit_r69_c63 bl[63] br[63] wl[69] vdd gnd cell_6t
Xbit_r70_c63 bl[63] br[63] wl[70] vdd gnd cell_6t
Xbit_r71_c63 bl[63] br[63] wl[71] vdd gnd cell_6t
Xbit_r72_c63 bl[63] br[63] wl[72] vdd gnd cell_6t
Xbit_r73_c63 bl[63] br[63] wl[73] vdd gnd cell_6t
Xbit_r74_c63 bl[63] br[63] wl[74] vdd gnd cell_6t
Xbit_r75_c63 bl[63] br[63] wl[75] vdd gnd cell_6t
Xbit_r76_c63 bl[63] br[63] wl[76] vdd gnd cell_6t
Xbit_r77_c63 bl[63] br[63] wl[77] vdd gnd cell_6t
Xbit_r78_c63 bl[63] br[63] wl[78] vdd gnd cell_6t
Xbit_r79_c63 bl[63] br[63] wl[79] vdd gnd cell_6t
Xbit_r80_c63 bl[63] br[63] wl[80] vdd gnd cell_6t
Xbit_r81_c63 bl[63] br[63] wl[81] vdd gnd cell_6t
Xbit_r82_c63 bl[63] br[63] wl[82] vdd gnd cell_6t
Xbit_r83_c63 bl[63] br[63] wl[83] vdd gnd cell_6t
Xbit_r84_c63 bl[63] br[63] wl[84] vdd gnd cell_6t
Xbit_r85_c63 bl[63] br[63] wl[85] vdd gnd cell_6t
Xbit_r86_c63 bl[63] br[63] wl[86] vdd gnd cell_6t
Xbit_r87_c63 bl[63] br[63] wl[87] vdd gnd cell_6t
Xbit_r88_c63 bl[63] br[63] wl[88] vdd gnd cell_6t
Xbit_r89_c63 bl[63] br[63] wl[89] vdd gnd cell_6t
Xbit_r90_c63 bl[63] br[63] wl[90] vdd gnd cell_6t
Xbit_r91_c63 bl[63] br[63] wl[91] vdd gnd cell_6t
Xbit_r92_c63 bl[63] br[63] wl[92] vdd gnd cell_6t
Xbit_r93_c63 bl[63] br[63] wl[93] vdd gnd cell_6t
Xbit_r94_c63 bl[63] br[63] wl[94] vdd gnd cell_6t
Xbit_r95_c63 bl[63] br[63] wl[95] vdd gnd cell_6t
Xbit_r96_c63 bl[63] br[63] wl[96] vdd gnd cell_6t
Xbit_r97_c63 bl[63] br[63] wl[97] vdd gnd cell_6t
Xbit_r98_c63 bl[63] br[63] wl[98] vdd gnd cell_6t
Xbit_r99_c63 bl[63] br[63] wl[99] vdd gnd cell_6t
Xbit_r100_c63 bl[63] br[63] wl[100] vdd gnd cell_6t
Xbit_r101_c63 bl[63] br[63] wl[101] vdd gnd cell_6t
Xbit_r102_c63 bl[63] br[63] wl[102] vdd gnd cell_6t
Xbit_r103_c63 bl[63] br[63] wl[103] vdd gnd cell_6t
Xbit_r104_c63 bl[63] br[63] wl[104] vdd gnd cell_6t
Xbit_r105_c63 bl[63] br[63] wl[105] vdd gnd cell_6t
Xbit_r106_c63 bl[63] br[63] wl[106] vdd gnd cell_6t
Xbit_r107_c63 bl[63] br[63] wl[107] vdd gnd cell_6t
Xbit_r108_c63 bl[63] br[63] wl[108] vdd gnd cell_6t
Xbit_r109_c63 bl[63] br[63] wl[109] vdd gnd cell_6t
Xbit_r110_c63 bl[63] br[63] wl[110] vdd gnd cell_6t
Xbit_r111_c63 bl[63] br[63] wl[111] vdd gnd cell_6t
Xbit_r112_c63 bl[63] br[63] wl[112] vdd gnd cell_6t
Xbit_r113_c63 bl[63] br[63] wl[113] vdd gnd cell_6t
Xbit_r114_c63 bl[63] br[63] wl[114] vdd gnd cell_6t
Xbit_r115_c63 bl[63] br[63] wl[115] vdd gnd cell_6t
Xbit_r116_c63 bl[63] br[63] wl[116] vdd gnd cell_6t
Xbit_r117_c63 bl[63] br[63] wl[117] vdd gnd cell_6t
Xbit_r118_c63 bl[63] br[63] wl[118] vdd gnd cell_6t
Xbit_r119_c63 bl[63] br[63] wl[119] vdd gnd cell_6t
Xbit_r120_c63 bl[63] br[63] wl[120] vdd gnd cell_6t
Xbit_r121_c63 bl[63] br[63] wl[121] vdd gnd cell_6t
Xbit_r122_c63 bl[63] br[63] wl[122] vdd gnd cell_6t
Xbit_r123_c63 bl[63] br[63] wl[123] vdd gnd cell_6t
Xbit_r124_c63 bl[63] br[63] wl[124] vdd gnd cell_6t
Xbit_r125_c63 bl[63] br[63] wl[125] vdd gnd cell_6t
Xbit_r126_c63 bl[63] br[63] wl[126] vdd gnd cell_6t
Xbit_r127_c63 bl[63] br[63] wl[127] vdd gnd cell_6t
Xbit_r128_c63 bl[63] br[63] wl[128] vdd gnd cell_6t
Xbit_r129_c63 bl[63] br[63] wl[129] vdd gnd cell_6t
Xbit_r130_c63 bl[63] br[63] wl[130] vdd gnd cell_6t
Xbit_r131_c63 bl[63] br[63] wl[131] vdd gnd cell_6t
Xbit_r132_c63 bl[63] br[63] wl[132] vdd gnd cell_6t
Xbit_r133_c63 bl[63] br[63] wl[133] vdd gnd cell_6t
Xbit_r134_c63 bl[63] br[63] wl[134] vdd gnd cell_6t
Xbit_r135_c63 bl[63] br[63] wl[135] vdd gnd cell_6t
Xbit_r136_c63 bl[63] br[63] wl[136] vdd gnd cell_6t
Xbit_r137_c63 bl[63] br[63] wl[137] vdd gnd cell_6t
Xbit_r138_c63 bl[63] br[63] wl[138] vdd gnd cell_6t
Xbit_r139_c63 bl[63] br[63] wl[139] vdd gnd cell_6t
Xbit_r140_c63 bl[63] br[63] wl[140] vdd gnd cell_6t
Xbit_r141_c63 bl[63] br[63] wl[141] vdd gnd cell_6t
Xbit_r142_c63 bl[63] br[63] wl[142] vdd gnd cell_6t
Xbit_r143_c63 bl[63] br[63] wl[143] vdd gnd cell_6t
Xbit_r144_c63 bl[63] br[63] wl[144] vdd gnd cell_6t
Xbit_r145_c63 bl[63] br[63] wl[145] vdd gnd cell_6t
Xbit_r146_c63 bl[63] br[63] wl[146] vdd gnd cell_6t
Xbit_r147_c63 bl[63] br[63] wl[147] vdd gnd cell_6t
Xbit_r148_c63 bl[63] br[63] wl[148] vdd gnd cell_6t
Xbit_r149_c63 bl[63] br[63] wl[149] vdd gnd cell_6t
Xbit_r150_c63 bl[63] br[63] wl[150] vdd gnd cell_6t
Xbit_r151_c63 bl[63] br[63] wl[151] vdd gnd cell_6t
Xbit_r152_c63 bl[63] br[63] wl[152] vdd gnd cell_6t
Xbit_r153_c63 bl[63] br[63] wl[153] vdd gnd cell_6t
Xbit_r154_c63 bl[63] br[63] wl[154] vdd gnd cell_6t
Xbit_r155_c63 bl[63] br[63] wl[155] vdd gnd cell_6t
Xbit_r156_c63 bl[63] br[63] wl[156] vdd gnd cell_6t
Xbit_r157_c63 bl[63] br[63] wl[157] vdd gnd cell_6t
Xbit_r158_c63 bl[63] br[63] wl[158] vdd gnd cell_6t
Xbit_r159_c63 bl[63] br[63] wl[159] vdd gnd cell_6t
Xbit_r160_c63 bl[63] br[63] wl[160] vdd gnd cell_6t
Xbit_r161_c63 bl[63] br[63] wl[161] vdd gnd cell_6t
Xbit_r162_c63 bl[63] br[63] wl[162] vdd gnd cell_6t
Xbit_r163_c63 bl[63] br[63] wl[163] vdd gnd cell_6t
Xbit_r164_c63 bl[63] br[63] wl[164] vdd gnd cell_6t
Xbit_r165_c63 bl[63] br[63] wl[165] vdd gnd cell_6t
Xbit_r166_c63 bl[63] br[63] wl[166] vdd gnd cell_6t
Xbit_r167_c63 bl[63] br[63] wl[167] vdd gnd cell_6t
Xbit_r168_c63 bl[63] br[63] wl[168] vdd gnd cell_6t
Xbit_r169_c63 bl[63] br[63] wl[169] vdd gnd cell_6t
Xbit_r170_c63 bl[63] br[63] wl[170] vdd gnd cell_6t
Xbit_r171_c63 bl[63] br[63] wl[171] vdd gnd cell_6t
Xbit_r172_c63 bl[63] br[63] wl[172] vdd gnd cell_6t
Xbit_r173_c63 bl[63] br[63] wl[173] vdd gnd cell_6t
Xbit_r174_c63 bl[63] br[63] wl[174] vdd gnd cell_6t
Xbit_r175_c63 bl[63] br[63] wl[175] vdd gnd cell_6t
Xbit_r176_c63 bl[63] br[63] wl[176] vdd gnd cell_6t
Xbit_r177_c63 bl[63] br[63] wl[177] vdd gnd cell_6t
Xbit_r178_c63 bl[63] br[63] wl[178] vdd gnd cell_6t
Xbit_r179_c63 bl[63] br[63] wl[179] vdd gnd cell_6t
Xbit_r180_c63 bl[63] br[63] wl[180] vdd gnd cell_6t
Xbit_r181_c63 bl[63] br[63] wl[181] vdd gnd cell_6t
Xbit_r182_c63 bl[63] br[63] wl[182] vdd gnd cell_6t
Xbit_r183_c63 bl[63] br[63] wl[183] vdd gnd cell_6t
Xbit_r184_c63 bl[63] br[63] wl[184] vdd gnd cell_6t
Xbit_r185_c63 bl[63] br[63] wl[185] vdd gnd cell_6t
Xbit_r186_c63 bl[63] br[63] wl[186] vdd gnd cell_6t
Xbit_r187_c63 bl[63] br[63] wl[187] vdd gnd cell_6t
Xbit_r188_c63 bl[63] br[63] wl[188] vdd gnd cell_6t
Xbit_r189_c63 bl[63] br[63] wl[189] vdd gnd cell_6t
Xbit_r190_c63 bl[63] br[63] wl[190] vdd gnd cell_6t
Xbit_r191_c63 bl[63] br[63] wl[191] vdd gnd cell_6t
Xbit_r192_c63 bl[63] br[63] wl[192] vdd gnd cell_6t
Xbit_r193_c63 bl[63] br[63] wl[193] vdd gnd cell_6t
Xbit_r194_c63 bl[63] br[63] wl[194] vdd gnd cell_6t
Xbit_r195_c63 bl[63] br[63] wl[195] vdd gnd cell_6t
Xbit_r196_c63 bl[63] br[63] wl[196] vdd gnd cell_6t
Xbit_r197_c63 bl[63] br[63] wl[197] vdd gnd cell_6t
Xbit_r198_c63 bl[63] br[63] wl[198] vdd gnd cell_6t
Xbit_r199_c63 bl[63] br[63] wl[199] vdd gnd cell_6t
Xbit_r200_c63 bl[63] br[63] wl[200] vdd gnd cell_6t
Xbit_r201_c63 bl[63] br[63] wl[201] vdd gnd cell_6t
Xbit_r202_c63 bl[63] br[63] wl[202] vdd gnd cell_6t
Xbit_r203_c63 bl[63] br[63] wl[203] vdd gnd cell_6t
Xbit_r204_c63 bl[63] br[63] wl[204] vdd gnd cell_6t
Xbit_r205_c63 bl[63] br[63] wl[205] vdd gnd cell_6t
Xbit_r206_c63 bl[63] br[63] wl[206] vdd gnd cell_6t
Xbit_r207_c63 bl[63] br[63] wl[207] vdd gnd cell_6t
Xbit_r208_c63 bl[63] br[63] wl[208] vdd gnd cell_6t
Xbit_r209_c63 bl[63] br[63] wl[209] vdd gnd cell_6t
Xbit_r210_c63 bl[63] br[63] wl[210] vdd gnd cell_6t
Xbit_r211_c63 bl[63] br[63] wl[211] vdd gnd cell_6t
Xbit_r212_c63 bl[63] br[63] wl[212] vdd gnd cell_6t
Xbit_r213_c63 bl[63] br[63] wl[213] vdd gnd cell_6t
Xbit_r214_c63 bl[63] br[63] wl[214] vdd gnd cell_6t
Xbit_r215_c63 bl[63] br[63] wl[215] vdd gnd cell_6t
Xbit_r216_c63 bl[63] br[63] wl[216] vdd gnd cell_6t
Xbit_r217_c63 bl[63] br[63] wl[217] vdd gnd cell_6t
Xbit_r218_c63 bl[63] br[63] wl[218] vdd gnd cell_6t
Xbit_r219_c63 bl[63] br[63] wl[219] vdd gnd cell_6t
Xbit_r220_c63 bl[63] br[63] wl[220] vdd gnd cell_6t
Xbit_r221_c63 bl[63] br[63] wl[221] vdd gnd cell_6t
Xbit_r222_c63 bl[63] br[63] wl[222] vdd gnd cell_6t
Xbit_r223_c63 bl[63] br[63] wl[223] vdd gnd cell_6t
Xbit_r224_c63 bl[63] br[63] wl[224] vdd gnd cell_6t
Xbit_r225_c63 bl[63] br[63] wl[225] vdd gnd cell_6t
Xbit_r226_c63 bl[63] br[63] wl[226] vdd gnd cell_6t
Xbit_r227_c63 bl[63] br[63] wl[227] vdd gnd cell_6t
Xbit_r228_c63 bl[63] br[63] wl[228] vdd gnd cell_6t
Xbit_r229_c63 bl[63] br[63] wl[229] vdd gnd cell_6t
Xbit_r230_c63 bl[63] br[63] wl[230] vdd gnd cell_6t
Xbit_r231_c63 bl[63] br[63] wl[231] vdd gnd cell_6t
Xbit_r232_c63 bl[63] br[63] wl[232] vdd gnd cell_6t
Xbit_r233_c63 bl[63] br[63] wl[233] vdd gnd cell_6t
Xbit_r234_c63 bl[63] br[63] wl[234] vdd gnd cell_6t
Xbit_r235_c63 bl[63] br[63] wl[235] vdd gnd cell_6t
Xbit_r236_c63 bl[63] br[63] wl[236] vdd gnd cell_6t
Xbit_r237_c63 bl[63] br[63] wl[237] vdd gnd cell_6t
Xbit_r238_c63 bl[63] br[63] wl[238] vdd gnd cell_6t
Xbit_r239_c63 bl[63] br[63] wl[239] vdd gnd cell_6t
Xbit_r240_c63 bl[63] br[63] wl[240] vdd gnd cell_6t
Xbit_r241_c63 bl[63] br[63] wl[241] vdd gnd cell_6t
Xbit_r242_c63 bl[63] br[63] wl[242] vdd gnd cell_6t
Xbit_r243_c63 bl[63] br[63] wl[243] vdd gnd cell_6t
Xbit_r244_c63 bl[63] br[63] wl[244] vdd gnd cell_6t
Xbit_r245_c63 bl[63] br[63] wl[245] vdd gnd cell_6t
Xbit_r246_c63 bl[63] br[63] wl[246] vdd gnd cell_6t
Xbit_r247_c63 bl[63] br[63] wl[247] vdd gnd cell_6t
Xbit_r248_c63 bl[63] br[63] wl[248] vdd gnd cell_6t
Xbit_r249_c63 bl[63] br[63] wl[249] vdd gnd cell_6t
Xbit_r250_c63 bl[63] br[63] wl[250] vdd gnd cell_6t
Xbit_r251_c63 bl[63] br[63] wl[251] vdd gnd cell_6t
Xbit_r252_c63 bl[63] br[63] wl[252] vdd gnd cell_6t
Xbit_r253_c63 bl[63] br[63] wl[253] vdd gnd cell_6t
Xbit_r254_c63 bl[63] br[63] wl[254] vdd gnd cell_6t
Xbit_r255_c63 bl[63] br[63] wl[255] vdd gnd cell_6t
Xbit_r0_c64 bl[64] br[64] wl[0] vdd gnd cell_6t
Xbit_r1_c64 bl[64] br[64] wl[1] vdd gnd cell_6t
Xbit_r2_c64 bl[64] br[64] wl[2] vdd gnd cell_6t
Xbit_r3_c64 bl[64] br[64] wl[3] vdd gnd cell_6t
Xbit_r4_c64 bl[64] br[64] wl[4] vdd gnd cell_6t
Xbit_r5_c64 bl[64] br[64] wl[5] vdd gnd cell_6t
Xbit_r6_c64 bl[64] br[64] wl[6] vdd gnd cell_6t
Xbit_r7_c64 bl[64] br[64] wl[7] vdd gnd cell_6t
Xbit_r8_c64 bl[64] br[64] wl[8] vdd gnd cell_6t
Xbit_r9_c64 bl[64] br[64] wl[9] vdd gnd cell_6t
Xbit_r10_c64 bl[64] br[64] wl[10] vdd gnd cell_6t
Xbit_r11_c64 bl[64] br[64] wl[11] vdd gnd cell_6t
Xbit_r12_c64 bl[64] br[64] wl[12] vdd gnd cell_6t
Xbit_r13_c64 bl[64] br[64] wl[13] vdd gnd cell_6t
Xbit_r14_c64 bl[64] br[64] wl[14] vdd gnd cell_6t
Xbit_r15_c64 bl[64] br[64] wl[15] vdd gnd cell_6t
Xbit_r16_c64 bl[64] br[64] wl[16] vdd gnd cell_6t
Xbit_r17_c64 bl[64] br[64] wl[17] vdd gnd cell_6t
Xbit_r18_c64 bl[64] br[64] wl[18] vdd gnd cell_6t
Xbit_r19_c64 bl[64] br[64] wl[19] vdd gnd cell_6t
Xbit_r20_c64 bl[64] br[64] wl[20] vdd gnd cell_6t
Xbit_r21_c64 bl[64] br[64] wl[21] vdd gnd cell_6t
Xbit_r22_c64 bl[64] br[64] wl[22] vdd gnd cell_6t
Xbit_r23_c64 bl[64] br[64] wl[23] vdd gnd cell_6t
Xbit_r24_c64 bl[64] br[64] wl[24] vdd gnd cell_6t
Xbit_r25_c64 bl[64] br[64] wl[25] vdd gnd cell_6t
Xbit_r26_c64 bl[64] br[64] wl[26] vdd gnd cell_6t
Xbit_r27_c64 bl[64] br[64] wl[27] vdd gnd cell_6t
Xbit_r28_c64 bl[64] br[64] wl[28] vdd gnd cell_6t
Xbit_r29_c64 bl[64] br[64] wl[29] vdd gnd cell_6t
Xbit_r30_c64 bl[64] br[64] wl[30] vdd gnd cell_6t
Xbit_r31_c64 bl[64] br[64] wl[31] vdd gnd cell_6t
Xbit_r32_c64 bl[64] br[64] wl[32] vdd gnd cell_6t
Xbit_r33_c64 bl[64] br[64] wl[33] vdd gnd cell_6t
Xbit_r34_c64 bl[64] br[64] wl[34] vdd gnd cell_6t
Xbit_r35_c64 bl[64] br[64] wl[35] vdd gnd cell_6t
Xbit_r36_c64 bl[64] br[64] wl[36] vdd gnd cell_6t
Xbit_r37_c64 bl[64] br[64] wl[37] vdd gnd cell_6t
Xbit_r38_c64 bl[64] br[64] wl[38] vdd gnd cell_6t
Xbit_r39_c64 bl[64] br[64] wl[39] vdd gnd cell_6t
Xbit_r40_c64 bl[64] br[64] wl[40] vdd gnd cell_6t
Xbit_r41_c64 bl[64] br[64] wl[41] vdd gnd cell_6t
Xbit_r42_c64 bl[64] br[64] wl[42] vdd gnd cell_6t
Xbit_r43_c64 bl[64] br[64] wl[43] vdd gnd cell_6t
Xbit_r44_c64 bl[64] br[64] wl[44] vdd gnd cell_6t
Xbit_r45_c64 bl[64] br[64] wl[45] vdd gnd cell_6t
Xbit_r46_c64 bl[64] br[64] wl[46] vdd gnd cell_6t
Xbit_r47_c64 bl[64] br[64] wl[47] vdd gnd cell_6t
Xbit_r48_c64 bl[64] br[64] wl[48] vdd gnd cell_6t
Xbit_r49_c64 bl[64] br[64] wl[49] vdd gnd cell_6t
Xbit_r50_c64 bl[64] br[64] wl[50] vdd gnd cell_6t
Xbit_r51_c64 bl[64] br[64] wl[51] vdd gnd cell_6t
Xbit_r52_c64 bl[64] br[64] wl[52] vdd gnd cell_6t
Xbit_r53_c64 bl[64] br[64] wl[53] vdd gnd cell_6t
Xbit_r54_c64 bl[64] br[64] wl[54] vdd gnd cell_6t
Xbit_r55_c64 bl[64] br[64] wl[55] vdd gnd cell_6t
Xbit_r56_c64 bl[64] br[64] wl[56] vdd gnd cell_6t
Xbit_r57_c64 bl[64] br[64] wl[57] vdd gnd cell_6t
Xbit_r58_c64 bl[64] br[64] wl[58] vdd gnd cell_6t
Xbit_r59_c64 bl[64] br[64] wl[59] vdd gnd cell_6t
Xbit_r60_c64 bl[64] br[64] wl[60] vdd gnd cell_6t
Xbit_r61_c64 bl[64] br[64] wl[61] vdd gnd cell_6t
Xbit_r62_c64 bl[64] br[64] wl[62] vdd gnd cell_6t
Xbit_r63_c64 bl[64] br[64] wl[63] vdd gnd cell_6t
Xbit_r64_c64 bl[64] br[64] wl[64] vdd gnd cell_6t
Xbit_r65_c64 bl[64] br[64] wl[65] vdd gnd cell_6t
Xbit_r66_c64 bl[64] br[64] wl[66] vdd gnd cell_6t
Xbit_r67_c64 bl[64] br[64] wl[67] vdd gnd cell_6t
Xbit_r68_c64 bl[64] br[64] wl[68] vdd gnd cell_6t
Xbit_r69_c64 bl[64] br[64] wl[69] vdd gnd cell_6t
Xbit_r70_c64 bl[64] br[64] wl[70] vdd gnd cell_6t
Xbit_r71_c64 bl[64] br[64] wl[71] vdd gnd cell_6t
Xbit_r72_c64 bl[64] br[64] wl[72] vdd gnd cell_6t
Xbit_r73_c64 bl[64] br[64] wl[73] vdd gnd cell_6t
Xbit_r74_c64 bl[64] br[64] wl[74] vdd gnd cell_6t
Xbit_r75_c64 bl[64] br[64] wl[75] vdd gnd cell_6t
Xbit_r76_c64 bl[64] br[64] wl[76] vdd gnd cell_6t
Xbit_r77_c64 bl[64] br[64] wl[77] vdd gnd cell_6t
Xbit_r78_c64 bl[64] br[64] wl[78] vdd gnd cell_6t
Xbit_r79_c64 bl[64] br[64] wl[79] vdd gnd cell_6t
Xbit_r80_c64 bl[64] br[64] wl[80] vdd gnd cell_6t
Xbit_r81_c64 bl[64] br[64] wl[81] vdd gnd cell_6t
Xbit_r82_c64 bl[64] br[64] wl[82] vdd gnd cell_6t
Xbit_r83_c64 bl[64] br[64] wl[83] vdd gnd cell_6t
Xbit_r84_c64 bl[64] br[64] wl[84] vdd gnd cell_6t
Xbit_r85_c64 bl[64] br[64] wl[85] vdd gnd cell_6t
Xbit_r86_c64 bl[64] br[64] wl[86] vdd gnd cell_6t
Xbit_r87_c64 bl[64] br[64] wl[87] vdd gnd cell_6t
Xbit_r88_c64 bl[64] br[64] wl[88] vdd gnd cell_6t
Xbit_r89_c64 bl[64] br[64] wl[89] vdd gnd cell_6t
Xbit_r90_c64 bl[64] br[64] wl[90] vdd gnd cell_6t
Xbit_r91_c64 bl[64] br[64] wl[91] vdd gnd cell_6t
Xbit_r92_c64 bl[64] br[64] wl[92] vdd gnd cell_6t
Xbit_r93_c64 bl[64] br[64] wl[93] vdd gnd cell_6t
Xbit_r94_c64 bl[64] br[64] wl[94] vdd gnd cell_6t
Xbit_r95_c64 bl[64] br[64] wl[95] vdd gnd cell_6t
Xbit_r96_c64 bl[64] br[64] wl[96] vdd gnd cell_6t
Xbit_r97_c64 bl[64] br[64] wl[97] vdd gnd cell_6t
Xbit_r98_c64 bl[64] br[64] wl[98] vdd gnd cell_6t
Xbit_r99_c64 bl[64] br[64] wl[99] vdd gnd cell_6t
Xbit_r100_c64 bl[64] br[64] wl[100] vdd gnd cell_6t
Xbit_r101_c64 bl[64] br[64] wl[101] vdd gnd cell_6t
Xbit_r102_c64 bl[64] br[64] wl[102] vdd gnd cell_6t
Xbit_r103_c64 bl[64] br[64] wl[103] vdd gnd cell_6t
Xbit_r104_c64 bl[64] br[64] wl[104] vdd gnd cell_6t
Xbit_r105_c64 bl[64] br[64] wl[105] vdd gnd cell_6t
Xbit_r106_c64 bl[64] br[64] wl[106] vdd gnd cell_6t
Xbit_r107_c64 bl[64] br[64] wl[107] vdd gnd cell_6t
Xbit_r108_c64 bl[64] br[64] wl[108] vdd gnd cell_6t
Xbit_r109_c64 bl[64] br[64] wl[109] vdd gnd cell_6t
Xbit_r110_c64 bl[64] br[64] wl[110] vdd gnd cell_6t
Xbit_r111_c64 bl[64] br[64] wl[111] vdd gnd cell_6t
Xbit_r112_c64 bl[64] br[64] wl[112] vdd gnd cell_6t
Xbit_r113_c64 bl[64] br[64] wl[113] vdd gnd cell_6t
Xbit_r114_c64 bl[64] br[64] wl[114] vdd gnd cell_6t
Xbit_r115_c64 bl[64] br[64] wl[115] vdd gnd cell_6t
Xbit_r116_c64 bl[64] br[64] wl[116] vdd gnd cell_6t
Xbit_r117_c64 bl[64] br[64] wl[117] vdd gnd cell_6t
Xbit_r118_c64 bl[64] br[64] wl[118] vdd gnd cell_6t
Xbit_r119_c64 bl[64] br[64] wl[119] vdd gnd cell_6t
Xbit_r120_c64 bl[64] br[64] wl[120] vdd gnd cell_6t
Xbit_r121_c64 bl[64] br[64] wl[121] vdd gnd cell_6t
Xbit_r122_c64 bl[64] br[64] wl[122] vdd gnd cell_6t
Xbit_r123_c64 bl[64] br[64] wl[123] vdd gnd cell_6t
Xbit_r124_c64 bl[64] br[64] wl[124] vdd gnd cell_6t
Xbit_r125_c64 bl[64] br[64] wl[125] vdd gnd cell_6t
Xbit_r126_c64 bl[64] br[64] wl[126] vdd gnd cell_6t
Xbit_r127_c64 bl[64] br[64] wl[127] vdd gnd cell_6t
Xbit_r128_c64 bl[64] br[64] wl[128] vdd gnd cell_6t
Xbit_r129_c64 bl[64] br[64] wl[129] vdd gnd cell_6t
Xbit_r130_c64 bl[64] br[64] wl[130] vdd gnd cell_6t
Xbit_r131_c64 bl[64] br[64] wl[131] vdd gnd cell_6t
Xbit_r132_c64 bl[64] br[64] wl[132] vdd gnd cell_6t
Xbit_r133_c64 bl[64] br[64] wl[133] vdd gnd cell_6t
Xbit_r134_c64 bl[64] br[64] wl[134] vdd gnd cell_6t
Xbit_r135_c64 bl[64] br[64] wl[135] vdd gnd cell_6t
Xbit_r136_c64 bl[64] br[64] wl[136] vdd gnd cell_6t
Xbit_r137_c64 bl[64] br[64] wl[137] vdd gnd cell_6t
Xbit_r138_c64 bl[64] br[64] wl[138] vdd gnd cell_6t
Xbit_r139_c64 bl[64] br[64] wl[139] vdd gnd cell_6t
Xbit_r140_c64 bl[64] br[64] wl[140] vdd gnd cell_6t
Xbit_r141_c64 bl[64] br[64] wl[141] vdd gnd cell_6t
Xbit_r142_c64 bl[64] br[64] wl[142] vdd gnd cell_6t
Xbit_r143_c64 bl[64] br[64] wl[143] vdd gnd cell_6t
Xbit_r144_c64 bl[64] br[64] wl[144] vdd gnd cell_6t
Xbit_r145_c64 bl[64] br[64] wl[145] vdd gnd cell_6t
Xbit_r146_c64 bl[64] br[64] wl[146] vdd gnd cell_6t
Xbit_r147_c64 bl[64] br[64] wl[147] vdd gnd cell_6t
Xbit_r148_c64 bl[64] br[64] wl[148] vdd gnd cell_6t
Xbit_r149_c64 bl[64] br[64] wl[149] vdd gnd cell_6t
Xbit_r150_c64 bl[64] br[64] wl[150] vdd gnd cell_6t
Xbit_r151_c64 bl[64] br[64] wl[151] vdd gnd cell_6t
Xbit_r152_c64 bl[64] br[64] wl[152] vdd gnd cell_6t
Xbit_r153_c64 bl[64] br[64] wl[153] vdd gnd cell_6t
Xbit_r154_c64 bl[64] br[64] wl[154] vdd gnd cell_6t
Xbit_r155_c64 bl[64] br[64] wl[155] vdd gnd cell_6t
Xbit_r156_c64 bl[64] br[64] wl[156] vdd gnd cell_6t
Xbit_r157_c64 bl[64] br[64] wl[157] vdd gnd cell_6t
Xbit_r158_c64 bl[64] br[64] wl[158] vdd gnd cell_6t
Xbit_r159_c64 bl[64] br[64] wl[159] vdd gnd cell_6t
Xbit_r160_c64 bl[64] br[64] wl[160] vdd gnd cell_6t
Xbit_r161_c64 bl[64] br[64] wl[161] vdd gnd cell_6t
Xbit_r162_c64 bl[64] br[64] wl[162] vdd gnd cell_6t
Xbit_r163_c64 bl[64] br[64] wl[163] vdd gnd cell_6t
Xbit_r164_c64 bl[64] br[64] wl[164] vdd gnd cell_6t
Xbit_r165_c64 bl[64] br[64] wl[165] vdd gnd cell_6t
Xbit_r166_c64 bl[64] br[64] wl[166] vdd gnd cell_6t
Xbit_r167_c64 bl[64] br[64] wl[167] vdd gnd cell_6t
Xbit_r168_c64 bl[64] br[64] wl[168] vdd gnd cell_6t
Xbit_r169_c64 bl[64] br[64] wl[169] vdd gnd cell_6t
Xbit_r170_c64 bl[64] br[64] wl[170] vdd gnd cell_6t
Xbit_r171_c64 bl[64] br[64] wl[171] vdd gnd cell_6t
Xbit_r172_c64 bl[64] br[64] wl[172] vdd gnd cell_6t
Xbit_r173_c64 bl[64] br[64] wl[173] vdd gnd cell_6t
Xbit_r174_c64 bl[64] br[64] wl[174] vdd gnd cell_6t
Xbit_r175_c64 bl[64] br[64] wl[175] vdd gnd cell_6t
Xbit_r176_c64 bl[64] br[64] wl[176] vdd gnd cell_6t
Xbit_r177_c64 bl[64] br[64] wl[177] vdd gnd cell_6t
Xbit_r178_c64 bl[64] br[64] wl[178] vdd gnd cell_6t
Xbit_r179_c64 bl[64] br[64] wl[179] vdd gnd cell_6t
Xbit_r180_c64 bl[64] br[64] wl[180] vdd gnd cell_6t
Xbit_r181_c64 bl[64] br[64] wl[181] vdd gnd cell_6t
Xbit_r182_c64 bl[64] br[64] wl[182] vdd gnd cell_6t
Xbit_r183_c64 bl[64] br[64] wl[183] vdd gnd cell_6t
Xbit_r184_c64 bl[64] br[64] wl[184] vdd gnd cell_6t
Xbit_r185_c64 bl[64] br[64] wl[185] vdd gnd cell_6t
Xbit_r186_c64 bl[64] br[64] wl[186] vdd gnd cell_6t
Xbit_r187_c64 bl[64] br[64] wl[187] vdd gnd cell_6t
Xbit_r188_c64 bl[64] br[64] wl[188] vdd gnd cell_6t
Xbit_r189_c64 bl[64] br[64] wl[189] vdd gnd cell_6t
Xbit_r190_c64 bl[64] br[64] wl[190] vdd gnd cell_6t
Xbit_r191_c64 bl[64] br[64] wl[191] vdd gnd cell_6t
Xbit_r192_c64 bl[64] br[64] wl[192] vdd gnd cell_6t
Xbit_r193_c64 bl[64] br[64] wl[193] vdd gnd cell_6t
Xbit_r194_c64 bl[64] br[64] wl[194] vdd gnd cell_6t
Xbit_r195_c64 bl[64] br[64] wl[195] vdd gnd cell_6t
Xbit_r196_c64 bl[64] br[64] wl[196] vdd gnd cell_6t
Xbit_r197_c64 bl[64] br[64] wl[197] vdd gnd cell_6t
Xbit_r198_c64 bl[64] br[64] wl[198] vdd gnd cell_6t
Xbit_r199_c64 bl[64] br[64] wl[199] vdd gnd cell_6t
Xbit_r200_c64 bl[64] br[64] wl[200] vdd gnd cell_6t
Xbit_r201_c64 bl[64] br[64] wl[201] vdd gnd cell_6t
Xbit_r202_c64 bl[64] br[64] wl[202] vdd gnd cell_6t
Xbit_r203_c64 bl[64] br[64] wl[203] vdd gnd cell_6t
Xbit_r204_c64 bl[64] br[64] wl[204] vdd gnd cell_6t
Xbit_r205_c64 bl[64] br[64] wl[205] vdd gnd cell_6t
Xbit_r206_c64 bl[64] br[64] wl[206] vdd gnd cell_6t
Xbit_r207_c64 bl[64] br[64] wl[207] vdd gnd cell_6t
Xbit_r208_c64 bl[64] br[64] wl[208] vdd gnd cell_6t
Xbit_r209_c64 bl[64] br[64] wl[209] vdd gnd cell_6t
Xbit_r210_c64 bl[64] br[64] wl[210] vdd gnd cell_6t
Xbit_r211_c64 bl[64] br[64] wl[211] vdd gnd cell_6t
Xbit_r212_c64 bl[64] br[64] wl[212] vdd gnd cell_6t
Xbit_r213_c64 bl[64] br[64] wl[213] vdd gnd cell_6t
Xbit_r214_c64 bl[64] br[64] wl[214] vdd gnd cell_6t
Xbit_r215_c64 bl[64] br[64] wl[215] vdd gnd cell_6t
Xbit_r216_c64 bl[64] br[64] wl[216] vdd gnd cell_6t
Xbit_r217_c64 bl[64] br[64] wl[217] vdd gnd cell_6t
Xbit_r218_c64 bl[64] br[64] wl[218] vdd gnd cell_6t
Xbit_r219_c64 bl[64] br[64] wl[219] vdd gnd cell_6t
Xbit_r220_c64 bl[64] br[64] wl[220] vdd gnd cell_6t
Xbit_r221_c64 bl[64] br[64] wl[221] vdd gnd cell_6t
Xbit_r222_c64 bl[64] br[64] wl[222] vdd gnd cell_6t
Xbit_r223_c64 bl[64] br[64] wl[223] vdd gnd cell_6t
Xbit_r224_c64 bl[64] br[64] wl[224] vdd gnd cell_6t
Xbit_r225_c64 bl[64] br[64] wl[225] vdd gnd cell_6t
Xbit_r226_c64 bl[64] br[64] wl[226] vdd gnd cell_6t
Xbit_r227_c64 bl[64] br[64] wl[227] vdd gnd cell_6t
Xbit_r228_c64 bl[64] br[64] wl[228] vdd gnd cell_6t
Xbit_r229_c64 bl[64] br[64] wl[229] vdd gnd cell_6t
Xbit_r230_c64 bl[64] br[64] wl[230] vdd gnd cell_6t
Xbit_r231_c64 bl[64] br[64] wl[231] vdd gnd cell_6t
Xbit_r232_c64 bl[64] br[64] wl[232] vdd gnd cell_6t
Xbit_r233_c64 bl[64] br[64] wl[233] vdd gnd cell_6t
Xbit_r234_c64 bl[64] br[64] wl[234] vdd gnd cell_6t
Xbit_r235_c64 bl[64] br[64] wl[235] vdd gnd cell_6t
Xbit_r236_c64 bl[64] br[64] wl[236] vdd gnd cell_6t
Xbit_r237_c64 bl[64] br[64] wl[237] vdd gnd cell_6t
Xbit_r238_c64 bl[64] br[64] wl[238] vdd gnd cell_6t
Xbit_r239_c64 bl[64] br[64] wl[239] vdd gnd cell_6t
Xbit_r240_c64 bl[64] br[64] wl[240] vdd gnd cell_6t
Xbit_r241_c64 bl[64] br[64] wl[241] vdd gnd cell_6t
Xbit_r242_c64 bl[64] br[64] wl[242] vdd gnd cell_6t
Xbit_r243_c64 bl[64] br[64] wl[243] vdd gnd cell_6t
Xbit_r244_c64 bl[64] br[64] wl[244] vdd gnd cell_6t
Xbit_r245_c64 bl[64] br[64] wl[245] vdd gnd cell_6t
Xbit_r246_c64 bl[64] br[64] wl[246] vdd gnd cell_6t
Xbit_r247_c64 bl[64] br[64] wl[247] vdd gnd cell_6t
Xbit_r248_c64 bl[64] br[64] wl[248] vdd gnd cell_6t
Xbit_r249_c64 bl[64] br[64] wl[249] vdd gnd cell_6t
Xbit_r250_c64 bl[64] br[64] wl[250] vdd gnd cell_6t
Xbit_r251_c64 bl[64] br[64] wl[251] vdd gnd cell_6t
Xbit_r252_c64 bl[64] br[64] wl[252] vdd gnd cell_6t
Xbit_r253_c64 bl[64] br[64] wl[253] vdd gnd cell_6t
Xbit_r254_c64 bl[64] br[64] wl[254] vdd gnd cell_6t
Xbit_r255_c64 bl[64] br[64] wl[255] vdd gnd cell_6t
Xbit_r0_c65 bl[65] br[65] wl[0] vdd gnd cell_6t
Xbit_r1_c65 bl[65] br[65] wl[1] vdd gnd cell_6t
Xbit_r2_c65 bl[65] br[65] wl[2] vdd gnd cell_6t
Xbit_r3_c65 bl[65] br[65] wl[3] vdd gnd cell_6t
Xbit_r4_c65 bl[65] br[65] wl[4] vdd gnd cell_6t
Xbit_r5_c65 bl[65] br[65] wl[5] vdd gnd cell_6t
Xbit_r6_c65 bl[65] br[65] wl[6] vdd gnd cell_6t
Xbit_r7_c65 bl[65] br[65] wl[7] vdd gnd cell_6t
Xbit_r8_c65 bl[65] br[65] wl[8] vdd gnd cell_6t
Xbit_r9_c65 bl[65] br[65] wl[9] vdd gnd cell_6t
Xbit_r10_c65 bl[65] br[65] wl[10] vdd gnd cell_6t
Xbit_r11_c65 bl[65] br[65] wl[11] vdd gnd cell_6t
Xbit_r12_c65 bl[65] br[65] wl[12] vdd gnd cell_6t
Xbit_r13_c65 bl[65] br[65] wl[13] vdd gnd cell_6t
Xbit_r14_c65 bl[65] br[65] wl[14] vdd gnd cell_6t
Xbit_r15_c65 bl[65] br[65] wl[15] vdd gnd cell_6t
Xbit_r16_c65 bl[65] br[65] wl[16] vdd gnd cell_6t
Xbit_r17_c65 bl[65] br[65] wl[17] vdd gnd cell_6t
Xbit_r18_c65 bl[65] br[65] wl[18] vdd gnd cell_6t
Xbit_r19_c65 bl[65] br[65] wl[19] vdd gnd cell_6t
Xbit_r20_c65 bl[65] br[65] wl[20] vdd gnd cell_6t
Xbit_r21_c65 bl[65] br[65] wl[21] vdd gnd cell_6t
Xbit_r22_c65 bl[65] br[65] wl[22] vdd gnd cell_6t
Xbit_r23_c65 bl[65] br[65] wl[23] vdd gnd cell_6t
Xbit_r24_c65 bl[65] br[65] wl[24] vdd gnd cell_6t
Xbit_r25_c65 bl[65] br[65] wl[25] vdd gnd cell_6t
Xbit_r26_c65 bl[65] br[65] wl[26] vdd gnd cell_6t
Xbit_r27_c65 bl[65] br[65] wl[27] vdd gnd cell_6t
Xbit_r28_c65 bl[65] br[65] wl[28] vdd gnd cell_6t
Xbit_r29_c65 bl[65] br[65] wl[29] vdd gnd cell_6t
Xbit_r30_c65 bl[65] br[65] wl[30] vdd gnd cell_6t
Xbit_r31_c65 bl[65] br[65] wl[31] vdd gnd cell_6t
Xbit_r32_c65 bl[65] br[65] wl[32] vdd gnd cell_6t
Xbit_r33_c65 bl[65] br[65] wl[33] vdd gnd cell_6t
Xbit_r34_c65 bl[65] br[65] wl[34] vdd gnd cell_6t
Xbit_r35_c65 bl[65] br[65] wl[35] vdd gnd cell_6t
Xbit_r36_c65 bl[65] br[65] wl[36] vdd gnd cell_6t
Xbit_r37_c65 bl[65] br[65] wl[37] vdd gnd cell_6t
Xbit_r38_c65 bl[65] br[65] wl[38] vdd gnd cell_6t
Xbit_r39_c65 bl[65] br[65] wl[39] vdd gnd cell_6t
Xbit_r40_c65 bl[65] br[65] wl[40] vdd gnd cell_6t
Xbit_r41_c65 bl[65] br[65] wl[41] vdd gnd cell_6t
Xbit_r42_c65 bl[65] br[65] wl[42] vdd gnd cell_6t
Xbit_r43_c65 bl[65] br[65] wl[43] vdd gnd cell_6t
Xbit_r44_c65 bl[65] br[65] wl[44] vdd gnd cell_6t
Xbit_r45_c65 bl[65] br[65] wl[45] vdd gnd cell_6t
Xbit_r46_c65 bl[65] br[65] wl[46] vdd gnd cell_6t
Xbit_r47_c65 bl[65] br[65] wl[47] vdd gnd cell_6t
Xbit_r48_c65 bl[65] br[65] wl[48] vdd gnd cell_6t
Xbit_r49_c65 bl[65] br[65] wl[49] vdd gnd cell_6t
Xbit_r50_c65 bl[65] br[65] wl[50] vdd gnd cell_6t
Xbit_r51_c65 bl[65] br[65] wl[51] vdd gnd cell_6t
Xbit_r52_c65 bl[65] br[65] wl[52] vdd gnd cell_6t
Xbit_r53_c65 bl[65] br[65] wl[53] vdd gnd cell_6t
Xbit_r54_c65 bl[65] br[65] wl[54] vdd gnd cell_6t
Xbit_r55_c65 bl[65] br[65] wl[55] vdd gnd cell_6t
Xbit_r56_c65 bl[65] br[65] wl[56] vdd gnd cell_6t
Xbit_r57_c65 bl[65] br[65] wl[57] vdd gnd cell_6t
Xbit_r58_c65 bl[65] br[65] wl[58] vdd gnd cell_6t
Xbit_r59_c65 bl[65] br[65] wl[59] vdd gnd cell_6t
Xbit_r60_c65 bl[65] br[65] wl[60] vdd gnd cell_6t
Xbit_r61_c65 bl[65] br[65] wl[61] vdd gnd cell_6t
Xbit_r62_c65 bl[65] br[65] wl[62] vdd gnd cell_6t
Xbit_r63_c65 bl[65] br[65] wl[63] vdd gnd cell_6t
Xbit_r64_c65 bl[65] br[65] wl[64] vdd gnd cell_6t
Xbit_r65_c65 bl[65] br[65] wl[65] vdd gnd cell_6t
Xbit_r66_c65 bl[65] br[65] wl[66] vdd gnd cell_6t
Xbit_r67_c65 bl[65] br[65] wl[67] vdd gnd cell_6t
Xbit_r68_c65 bl[65] br[65] wl[68] vdd gnd cell_6t
Xbit_r69_c65 bl[65] br[65] wl[69] vdd gnd cell_6t
Xbit_r70_c65 bl[65] br[65] wl[70] vdd gnd cell_6t
Xbit_r71_c65 bl[65] br[65] wl[71] vdd gnd cell_6t
Xbit_r72_c65 bl[65] br[65] wl[72] vdd gnd cell_6t
Xbit_r73_c65 bl[65] br[65] wl[73] vdd gnd cell_6t
Xbit_r74_c65 bl[65] br[65] wl[74] vdd gnd cell_6t
Xbit_r75_c65 bl[65] br[65] wl[75] vdd gnd cell_6t
Xbit_r76_c65 bl[65] br[65] wl[76] vdd gnd cell_6t
Xbit_r77_c65 bl[65] br[65] wl[77] vdd gnd cell_6t
Xbit_r78_c65 bl[65] br[65] wl[78] vdd gnd cell_6t
Xbit_r79_c65 bl[65] br[65] wl[79] vdd gnd cell_6t
Xbit_r80_c65 bl[65] br[65] wl[80] vdd gnd cell_6t
Xbit_r81_c65 bl[65] br[65] wl[81] vdd gnd cell_6t
Xbit_r82_c65 bl[65] br[65] wl[82] vdd gnd cell_6t
Xbit_r83_c65 bl[65] br[65] wl[83] vdd gnd cell_6t
Xbit_r84_c65 bl[65] br[65] wl[84] vdd gnd cell_6t
Xbit_r85_c65 bl[65] br[65] wl[85] vdd gnd cell_6t
Xbit_r86_c65 bl[65] br[65] wl[86] vdd gnd cell_6t
Xbit_r87_c65 bl[65] br[65] wl[87] vdd gnd cell_6t
Xbit_r88_c65 bl[65] br[65] wl[88] vdd gnd cell_6t
Xbit_r89_c65 bl[65] br[65] wl[89] vdd gnd cell_6t
Xbit_r90_c65 bl[65] br[65] wl[90] vdd gnd cell_6t
Xbit_r91_c65 bl[65] br[65] wl[91] vdd gnd cell_6t
Xbit_r92_c65 bl[65] br[65] wl[92] vdd gnd cell_6t
Xbit_r93_c65 bl[65] br[65] wl[93] vdd gnd cell_6t
Xbit_r94_c65 bl[65] br[65] wl[94] vdd gnd cell_6t
Xbit_r95_c65 bl[65] br[65] wl[95] vdd gnd cell_6t
Xbit_r96_c65 bl[65] br[65] wl[96] vdd gnd cell_6t
Xbit_r97_c65 bl[65] br[65] wl[97] vdd gnd cell_6t
Xbit_r98_c65 bl[65] br[65] wl[98] vdd gnd cell_6t
Xbit_r99_c65 bl[65] br[65] wl[99] vdd gnd cell_6t
Xbit_r100_c65 bl[65] br[65] wl[100] vdd gnd cell_6t
Xbit_r101_c65 bl[65] br[65] wl[101] vdd gnd cell_6t
Xbit_r102_c65 bl[65] br[65] wl[102] vdd gnd cell_6t
Xbit_r103_c65 bl[65] br[65] wl[103] vdd gnd cell_6t
Xbit_r104_c65 bl[65] br[65] wl[104] vdd gnd cell_6t
Xbit_r105_c65 bl[65] br[65] wl[105] vdd gnd cell_6t
Xbit_r106_c65 bl[65] br[65] wl[106] vdd gnd cell_6t
Xbit_r107_c65 bl[65] br[65] wl[107] vdd gnd cell_6t
Xbit_r108_c65 bl[65] br[65] wl[108] vdd gnd cell_6t
Xbit_r109_c65 bl[65] br[65] wl[109] vdd gnd cell_6t
Xbit_r110_c65 bl[65] br[65] wl[110] vdd gnd cell_6t
Xbit_r111_c65 bl[65] br[65] wl[111] vdd gnd cell_6t
Xbit_r112_c65 bl[65] br[65] wl[112] vdd gnd cell_6t
Xbit_r113_c65 bl[65] br[65] wl[113] vdd gnd cell_6t
Xbit_r114_c65 bl[65] br[65] wl[114] vdd gnd cell_6t
Xbit_r115_c65 bl[65] br[65] wl[115] vdd gnd cell_6t
Xbit_r116_c65 bl[65] br[65] wl[116] vdd gnd cell_6t
Xbit_r117_c65 bl[65] br[65] wl[117] vdd gnd cell_6t
Xbit_r118_c65 bl[65] br[65] wl[118] vdd gnd cell_6t
Xbit_r119_c65 bl[65] br[65] wl[119] vdd gnd cell_6t
Xbit_r120_c65 bl[65] br[65] wl[120] vdd gnd cell_6t
Xbit_r121_c65 bl[65] br[65] wl[121] vdd gnd cell_6t
Xbit_r122_c65 bl[65] br[65] wl[122] vdd gnd cell_6t
Xbit_r123_c65 bl[65] br[65] wl[123] vdd gnd cell_6t
Xbit_r124_c65 bl[65] br[65] wl[124] vdd gnd cell_6t
Xbit_r125_c65 bl[65] br[65] wl[125] vdd gnd cell_6t
Xbit_r126_c65 bl[65] br[65] wl[126] vdd gnd cell_6t
Xbit_r127_c65 bl[65] br[65] wl[127] vdd gnd cell_6t
Xbit_r128_c65 bl[65] br[65] wl[128] vdd gnd cell_6t
Xbit_r129_c65 bl[65] br[65] wl[129] vdd gnd cell_6t
Xbit_r130_c65 bl[65] br[65] wl[130] vdd gnd cell_6t
Xbit_r131_c65 bl[65] br[65] wl[131] vdd gnd cell_6t
Xbit_r132_c65 bl[65] br[65] wl[132] vdd gnd cell_6t
Xbit_r133_c65 bl[65] br[65] wl[133] vdd gnd cell_6t
Xbit_r134_c65 bl[65] br[65] wl[134] vdd gnd cell_6t
Xbit_r135_c65 bl[65] br[65] wl[135] vdd gnd cell_6t
Xbit_r136_c65 bl[65] br[65] wl[136] vdd gnd cell_6t
Xbit_r137_c65 bl[65] br[65] wl[137] vdd gnd cell_6t
Xbit_r138_c65 bl[65] br[65] wl[138] vdd gnd cell_6t
Xbit_r139_c65 bl[65] br[65] wl[139] vdd gnd cell_6t
Xbit_r140_c65 bl[65] br[65] wl[140] vdd gnd cell_6t
Xbit_r141_c65 bl[65] br[65] wl[141] vdd gnd cell_6t
Xbit_r142_c65 bl[65] br[65] wl[142] vdd gnd cell_6t
Xbit_r143_c65 bl[65] br[65] wl[143] vdd gnd cell_6t
Xbit_r144_c65 bl[65] br[65] wl[144] vdd gnd cell_6t
Xbit_r145_c65 bl[65] br[65] wl[145] vdd gnd cell_6t
Xbit_r146_c65 bl[65] br[65] wl[146] vdd gnd cell_6t
Xbit_r147_c65 bl[65] br[65] wl[147] vdd gnd cell_6t
Xbit_r148_c65 bl[65] br[65] wl[148] vdd gnd cell_6t
Xbit_r149_c65 bl[65] br[65] wl[149] vdd gnd cell_6t
Xbit_r150_c65 bl[65] br[65] wl[150] vdd gnd cell_6t
Xbit_r151_c65 bl[65] br[65] wl[151] vdd gnd cell_6t
Xbit_r152_c65 bl[65] br[65] wl[152] vdd gnd cell_6t
Xbit_r153_c65 bl[65] br[65] wl[153] vdd gnd cell_6t
Xbit_r154_c65 bl[65] br[65] wl[154] vdd gnd cell_6t
Xbit_r155_c65 bl[65] br[65] wl[155] vdd gnd cell_6t
Xbit_r156_c65 bl[65] br[65] wl[156] vdd gnd cell_6t
Xbit_r157_c65 bl[65] br[65] wl[157] vdd gnd cell_6t
Xbit_r158_c65 bl[65] br[65] wl[158] vdd gnd cell_6t
Xbit_r159_c65 bl[65] br[65] wl[159] vdd gnd cell_6t
Xbit_r160_c65 bl[65] br[65] wl[160] vdd gnd cell_6t
Xbit_r161_c65 bl[65] br[65] wl[161] vdd gnd cell_6t
Xbit_r162_c65 bl[65] br[65] wl[162] vdd gnd cell_6t
Xbit_r163_c65 bl[65] br[65] wl[163] vdd gnd cell_6t
Xbit_r164_c65 bl[65] br[65] wl[164] vdd gnd cell_6t
Xbit_r165_c65 bl[65] br[65] wl[165] vdd gnd cell_6t
Xbit_r166_c65 bl[65] br[65] wl[166] vdd gnd cell_6t
Xbit_r167_c65 bl[65] br[65] wl[167] vdd gnd cell_6t
Xbit_r168_c65 bl[65] br[65] wl[168] vdd gnd cell_6t
Xbit_r169_c65 bl[65] br[65] wl[169] vdd gnd cell_6t
Xbit_r170_c65 bl[65] br[65] wl[170] vdd gnd cell_6t
Xbit_r171_c65 bl[65] br[65] wl[171] vdd gnd cell_6t
Xbit_r172_c65 bl[65] br[65] wl[172] vdd gnd cell_6t
Xbit_r173_c65 bl[65] br[65] wl[173] vdd gnd cell_6t
Xbit_r174_c65 bl[65] br[65] wl[174] vdd gnd cell_6t
Xbit_r175_c65 bl[65] br[65] wl[175] vdd gnd cell_6t
Xbit_r176_c65 bl[65] br[65] wl[176] vdd gnd cell_6t
Xbit_r177_c65 bl[65] br[65] wl[177] vdd gnd cell_6t
Xbit_r178_c65 bl[65] br[65] wl[178] vdd gnd cell_6t
Xbit_r179_c65 bl[65] br[65] wl[179] vdd gnd cell_6t
Xbit_r180_c65 bl[65] br[65] wl[180] vdd gnd cell_6t
Xbit_r181_c65 bl[65] br[65] wl[181] vdd gnd cell_6t
Xbit_r182_c65 bl[65] br[65] wl[182] vdd gnd cell_6t
Xbit_r183_c65 bl[65] br[65] wl[183] vdd gnd cell_6t
Xbit_r184_c65 bl[65] br[65] wl[184] vdd gnd cell_6t
Xbit_r185_c65 bl[65] br[65] wl[185] vdd gnd cell_6t
Xbit_r186_c65 bl[65] br[65] wl[186] vdd gnd cell_6t
Xbit_r187_c65 bl[65] br[65] wl[187] vdd gnd cell_6t
Xbit_r188_c65 bl[65] br[65] wl[188] vdd gnd cell_6t
Xbit_r189_c65 bl[65] br[65] wl[189] vdd gnd cell_6t
Xbit_r190_c65 bl[65] br[65] wl[190] vdd gnd cell_6t
Xbit_r191_c65 bl[65] br[65] wl[191] vdd gnd cell_6t
Xbit_r192_c65 bl[65] br[65] wl[192] vdd gnd cell_6t
Xbit_r193_c65 bl[65] br[65] wl[193] vdd gnd cell_6t
Xbit_r194_c65 bl[65] br[65] wl[194] vdd gnd cell_6t
Xbit_r195_c65 bl[65] br[65] wl[195] vdd gnd cell_6t
Xbit_r196_c65 bl[65] br[65] wl[196] vdd gnd cell_6t
Xbit_r197_c65 bl[65] br[65] wl[197] vdd gnd cell_6t
Xbit_r198_c65 bl[65] br[65] wl[198] vdd gnd cell_6t
Xbit_r199_c65 bl[65] br[65] wl[199] vdd gnd cell_6t
Xbit_r200_c65 bl[65] br[65] wl[200] vdd gnd cell_6t
Xbit_r201_c65 bl[65] br[65] wl[201] vdd gnd cell_6t
Xbit_r202_c65 bl[65] br[65] wl[202] vdd gnd cell_6t
Xbit_r203_c65 bl[65] br[65] wl[203] vdd gnd cell_6t
Xbit_r204_c65 bl[65] br[65] wl[204] vdd gnd cell_6t
Xbit_r205_c65 bl[65] br[65] wl[205] vdd gnd cell_6t
Xbit_r206_c65 bl[65] br[65] wl[206] vdd gnd cell_6t
Xbit_r207_c65 bl[65] br[65] wl[207] vdd gnd cell_6t
Xbit_r208_c65 bl[65] br[65] wl[208] vdd gnd cell_6t
Xbit_r209_c65 bl[65] br[65] wl[209] vdd gnd cell_6t
Xbit_r210_c65 bl[65] br[65] wl[210] vdd gnd cell_6t
Xbit_r211_c65 bl[65] br[65] wl[211] vdd gnd cell_6t
Xbit_r212_c65 bl[65] br[65] wl[212] vdd gnd cell_6t
Xbit_r213_c65 bl[65] br[65] wl[213] vdd gnd cell_6t
Xbit_r214_c65 bl[65] br[65] wl[214] vdd gnd cell_6t
Xbit_r215_c65 bl[65] br[65] wl[215] vdd gnd cell_6t
Xbit_r216_c65 bl[65] br[65] wl[216] vdd gnd cell_6t
Xbit_r217_c65 bl[65] br[65] wl[217] vdd gnd cell_6t
Xbit_r218_c65 bl[65] br[65] wl[218] vdd gnd cell_6t
Xbit_r219_c65 bl[65] br[65] wl[219] vdd gnd cell_6t
Xbit_r220_c65 bl[65] br[65] wl[220] vdd gnd cell_6t
Xbit_r221_c65 bl[65] br[65] wl[221] vdd gnd cell_6t
Xbit_r222_c65 bl[65] br[65] wl[222] vdd gnd cell_6t
Xbit_r223_c65 bl[65] br[65] wl[223] vdd gnd cell_6t
Xbit_r224_c65 bl[65] br[65] wl[224] vdd gnd cell_6t
Xbit_r225_c65 bl[65] br[65] wl[225] vdd gnd cell_6t
Xbit_r226_c65 bl[65] br[65] wl[226] vdd gnd cell_6t
Xbit_r227_c65 bl[65] br[65] wl[227] vdd gnd cell_6t
Xbit_r228_c65 bl[65] br[65] wl[228] vdd gnd cell_6t
Xbit_r229_c65 bl[65] br[65] wl[229] vdd gnd cell_6t
Xbit_r230_c65 bl[65] br[65] wl[230] vdd gnd cell_6t
Xbit_r231_c65 bl[65] br[65] wl[231] vdd gnd cell_6t
Xbit_r232_c65 bl[65] br[65] wl[232] vdd gnd cell_6t
Xbit_r233_c65 bl[65] br[65] wl[233] vdd gnd cell_6t
Xbit_r234_c65 bl[65] br[65] wl[234] vdd gnd cell_6t
Xbit_r235_c65 bl[65] br[65] wl[235] vdd gnd cell_6t
Xbit_r236_c65 bl[65] br[65] wl[236] vdd gnd cell_6t
Xbit_r237_c65 bl[65] br[65] wl[237] vdd gnd cell_6t
Xbit_r238_c65 bl[65] br[65] wl[238] vdd gnd cell_6t
Xbit_r239_c65 bl[65] br[65] wl[239] vdd gnd cell_6t
Xbit_r240_c65 bl[65] br[65] wl[240] vdd gnd cell_6t
Xbit_r241_c65 bl[65] br[65] wl[241] vdd gnd cell_6t
Xbit_r242_c65 bl[65] br[65] wl[242] vdd gnd cell_6t
Xbit_r243_c65 bl[65] br[65] wl[243] vdd gnd cell_6t
Xbit_r244_c65 bl[65] br[65] wl[244] vdd gnd cell_6t
Xbit_r245_c65 bl[65] br[65] wl[245] vdd gnd cell_6t
Xbit_r246_c65 bl[65] br[65] wl[246] vdd gnd cell_6t
Xbit_r247_c65 bl[65] br[65] wl[247] vdd gnd cell_6t
Xbit_r248_c65 bl[65] br[65] wl[248] vdd gnd cell_6t
Xbit_r249_c65 bl[65] br[65] wl[249] vdd gnd cell_6t
Xbit_r250_c65 bl[65] br[65] wl[250] vdd gnd cell_6t
Xbit_r251_c65 bl[65] br[65] wl[251] vdd gnd cell_6t
Xbit_r252_c65 bl[65] br[65] wl[252] vdd gnd cell_6t
Xbit_r253_c65 bl[65] br[65] wl[253] vdd gnd cell_6t
Xbit_r254_c65 bl[65] br[65] wl[254] vdd gnd cell_6t
Xbit_r255_c65 bl[65] br[65] wl[255] vdd gnd cell_6t
Xbit_r0_c66 bl[66] br[66] wl[0] vdd gnd cell_6t
Xbit_r1_c66 bl[66] br[66] wl[1] vdd gnd cell_6t
Xbit_r2_c66 bl[66] br[66] wl[2] vdd gnd cell_6t
Xbit_r3_c66 bl[66] br[66] wl[3] vdd gnd cell_6t
Xbit_r4_c66 bl[66] br[66] wl[4] vdd gnd cell_6t
Xbit_r5_c66 bl[66] br[66] wl[5] vdd gnd cell_6t
Xbit_r6_c66 bl[66] br[66] wl[6] vdd gnd cell_6t
Xbit_r7_c66 bl[66] br[66] wl[7] vdd gnd cell_6t
Xbit_r8_c66 bl[66] br[66] wl[8] vdd gnd cell_6t
Xbit_r9_c66 bl[66] br[66] wl[9] vdd gnd cell_6t
Xbit_r10_c66 bl[66] br[66] wl[10] vdd gnd cell_6t
Xbit_r11_c66 bl[66] br[66] wl[11] vdd gnd cell_6t
Xbit_r12_c66 bl[66] br[66] wl[12] vdd gnd cell_6t
Xbit_r13_c66 bl[66] br[66] wl[13] vdd gnd cell_6t
Xbit_r14_c66 bl[66] br[66] wl[14] vdd gnd cell_6t
Xbit_r15_c66 bl[66] br[66] wl[15] vdd gnd cell_6t
Xbit_r16_c66 bl[66] br[66] wl[16] vdd gnd cell_6t
Xbit_r17_c66 bl[66] br[66] wl[17] vdd gnd cell_6t
Xbit_r18_c66 bl[66] br[66] wl[18] vdd gnd cell_6t
Xbit_r19_c66 bl[66] br[66] wl[19] vdd gnd cell_6t
Xbit_r20_c66 bl[66] br[66] wl[20] vdd gnd cell_6t
Xbit_r21_c66 bl[66] br[66] wl[21] vdd gnd cell_6t
Xbit_r22_c66 bl[66] br[66] wl[22] vdd gnd cell_6t
Xbit_r23_c66 bl[66] br[66] wl[23] vdd gnd cell_6t
Xbit_r24_c66 bl[66] br[66] wl[24] vdd gnd cell_6t
Xbit_r25_c66 bl[66] br[66] wl[25] vdd gnd cell_6t
Xbit_r26_c66 bl[66] br[66] wl[26] vdd gnd cell_6t
Xbit_r27_c66 bl[66] br[66] wl[27] vdd gnd cell_6t
Xbit_r28_c66 bl[66] br[66] wl[28] vdd gnd cell_6t
Xbit_r29_c66 bl[66] br[66] wl[29] vdd gnd cell_6t
Xbit_r30_c66 bl[66] br[66] wl[30] vdd gnd cell_6t
Xbit_r31_c66 bl[66] br[66] wl[31] vdd gnd cell_6t
Xbit_r32_c66 bl[66] br[66] wl[32] vdd gnd cell_6t
Xbit_r33_c66 bl[66] br[66] wl[33] vdd gnd cell_6t
Xbit_r34_c66 bl[66] br[66] wl[34] vdd gnd cell_6t
Xbit_r35_c66 bl[66] br[66] wl[35] vdd gnd cell_6t
Xbit_r36_c66 bl[66] br[66] wl[36] vdd gnd cell_6t
Xbit_r37_c66 bl[66] br[66] wl[37] vdd gnd cell_6t
Xbit_r38_c66 bl[66] br[66] wl[38] vdd gnd cell_6t
Xbit_r39_c66 bl[66] br[66] wl[39] vdd gnd cell_6t
Xbit_r40_c66 bl[66] br[66] wl[40] vdd gnd cell_6t
Xbit_r41_c66 bl[66] br[66] wl[41] vdd gnd cell_6t
Xbit_r42_c66 bl[66] br[66] wl[42] vdd gnd cell_6t
Xbit_r43_c66 bl[66] br[66] wl[43] vdd gnd cell_6t
Xbit_r44_c66 bl[66] br[66] wl[44] vdd gnd cell_6t
Xbit_r45_c66 bl[66] br[66] wl[45] vdd gnd cell_6t
Xbit_r46_c66 bl[66] br[66] wl[46] vdd gnd cell_6t
Xbit_r47_c66 bl[66] br[66] wl[47] vdd gnd cell_6t
Xbit_r48_c66 bl[66] br[66] wl[48] vdd gnd cell_6t
Xbit_r49_c66 bl[66] br[66] wl[49] vdd gnd cell_6t
Xbit_r50_c66 bl[66] br[66] wl[50] vdd gnd cell_6t
Xbit_r51_c66 bl[66] br[66] wl[51] vdd gnd cell_6t
Xbit_r52_c66 bl[66] br[66] wl[52] vdd gnd cell_6t
Xbit_r53_c66 bl[66] br[66] wl[53] vdd gnd cell_6t
Xbit_r54_c66 bl[66] br[66] wl[54] vdd gnd cell_6t
Xbit_r55_c66 bl[66] br[66] wl[55] vdd gnd cell_6t
Xbit_r56_c66 bl[66] br[66] wl[56] vdd gnd cell_6t
Xbit_r57_c66 bl[66] br[66] wl[57] vdd gnd cell_6t
Xbit_r58_c66 bl[66] br[66] wl[58] vdd gnd cell_6t
Xbit_r59_c66 bl[66] br[66] wl[59] vdd gnd cell_6t
Xbit_r60_c66 bl[66] br[66] wl[60] vdd gnd cell_6t
Xbit_r61_c66 bl[66] br[66] wl[61] vdd gnd cell_6t
Xbit_r62_c66 bl[66] br[66] wl[62] vdd gnd cell_6t
Xbit_r63_c66 bl[66] br[66] wl[63] vdd gnd cell_6t
Xbit_r64_c66 bl[66] br[66] wl[64] vdd gnd cell_6t
Xbit_r65_c66 bl[66] br[66] wl[65] vdd gnd cell_6t
Xbit_r66_c66 bl[66] br[66] wl[66] vdd gnd cell_6t
Xbit_r67_c66 bl[66] br[66] wl[67] vdd gnd cell_6t
Xbit_r68_c66 bl[66] br[66] wl[68] vdd gnd cell_6t
Xbit_r69_c66 bl[66] br[66] wl[69] vdd gnd cell_6t
Xbit_r70_c66 bl[66] br[66] wl[70] vdd gnd cell_6t
Xbit_r71_c66 bl[66] br[66] wl[71] vdd gnd cell_6t
Xbit_r72_c66 bl[66] br[66] wl[72] vdd gnd cell_6t
Xbit_r73_c66 bl[66] br[66] wl[73] vdd gnd cell_6t
Xbit_r74_c66 bl[66] br[66] wl[74] vdd gnd cell_6t
Xbit_r75_c66 bl[66] br[66] wl[75] vdd gnd cell_6t
Xbit_r76_c66 bl[66] br[66] wl[76] vdd gnd cell_6t
Xbit_r77_c66 bl[66] br[66] wl[77] vdd gnd cell_6t
Xbit_r78_c66 bl[66] br[66] wl[78] vdd gnd cell_6t
Xbit_r79_c66 bl[66] br[66] wl[79] vdd gnd cell_6t
Xbit_r80_c66 bl[66] br[66] wl[80] vdd gnd cell_6t
Xbit_r81_c66 bl[66] br[66] wl[81] vdd gnd cell_6t
Xbit_r82_c66 bl[66] br[66] wl[82] vdd gnd cell_6t
Xbit_r83_c66 bl[66] br[66] wl[83] vdd gnd cell_6t
Xbit_r84_c66 bl[66] br[66] wl[84] vdd gnd cell_6t
Xbit_r85_c66 bl[66] br[66] wl[85] vdd gnd cell_6t
Xbit_r86_c66 bl[66] br[66] wl[86] vdd gnd cell_6t
Xbit_r87_c66 bl[66] br[66] wl[87] vdd gnd cell_6t
Xbit_r88_c66 bl[66] br[66] wl[88] vdd gnd cell_6t
Xbit_r89_c66 bl[66] br[66] wl[89] vdd gnd cell_6t
Xbit_r90_c66 bl[66] br[66] wl[90] vdd gnd cell_6t
Xbit_r91_c66 bl[66] br[66] wl[91] vdd gnd cell_6t
Xbit_r92_c66 bl[66] br[66] wl[92] vdd gnd cell_6t
Xbit_r93_c66 bl[66] br[66] wl[93] vdd gnd cell_6t
Xbit_r94_c66 bl[66] br[66] wl[94] vdd gnd cell_6t
Xbit_r95_c66 bl[66] br[66] wl[95] vdd gnd cell_6t
Xbit_r96_c66 bl[66] br[66] wl[96] vdd gnd cell_6t
Xbit_r97_c66 bl[66] br[66] wl[97] vdd gnd cell_6t
Xbit_r98_c66 bl[66] br[66] wl[98] vdd gnd cell_6t
Xbit_r99_c66 bl[66] br[66] wl[99] vdd gnd cell_6t
Xbit_r100_c66 bl[66] br[66] wl[100] vdd gnd cell_6t
Xbit_r101_c66 bl[66] br[66] wl[101] vdd gnd cell_6t
Xbit_r102_c66 bl[66] br[66] wl[102] vdd gnd cell_6t
Xbit_r103_c66 bl[66] br[66] wl[103] vdd gnd cell_6t
Xbit_r104_c66 bl[66] br[66] wl[104] vdd gnd cell_6t
Xbit_r105_c66 bl[66] br[66] wl[105] vdd gnd cell_6t
Xbit_r106_c66 bl[66] br[66] wl[106] vdd gnd cell_6t
Xbit_r107_c66 bl[66] br[66] wl[107] vdd gnd cell_6t
Xbit_r108_c66 bl[66] br[66] wl[108] vdd gnd cell_6t
Xbit_r109_c66 bl[66] br[66] wl[109] vdd gnd cell_6t
Xbit_r110_c66 bl[66] br[66] wl[110] vdd gnd cell_6t
Xbit_r111_c66 bl[66] br[66] wl[111] vdd gnd cell_6t
Xbit_r112_c66 bl[66] br[66] wl[112] vdd gnd cell_6t
Xbit_r113_c66 bl[66] br[66] wl[113] vdd gnd cell_6t
Xbit_r114_c66 bl[66] br[66] wl[114] vdd gnd cell_6t
Xbit_r115_c66 bl[66] br[66] wl[115] vdd gnd cell_6t
Xbit_r116_c66 bl[66] br[66] wl[116] vdd gnd cell_6t
Xbit_r117_c66 bl[66] br[66] wl[117] vdd gnd cell_6t
Xbit_r118_c66 bl[66] br[66] wl[118] vdd gnd cell_6t
Xbit_r119_c66 bl[66] br[66] wl[119] vdd gnd cell_6t
Xbit_r120_c66 bl[66] br[66] wl[120] vdd gnd cell_6t
Xbit_r121_c66 bl[66] br[66] wl[121] vdd gnd cell_6t
Xbit_r122_c66 bl[66] br[66] wl[122] vdd gnd cell_6t
Xbit_r123_c66 bl[66] br[66] wl[123] vdd gnd cell_6t
Xbit_r124_c66 bl[66] br[66] wl[124] vdd gnd cell_6t
Xbit_r125_c66 bl[66] br[66] wl[125] vdd gnd cell_6t
Xbit_r126_c66 bl[66] br[66] wl[126] vdd gnd cell_6t
Xbit_r127_c66 bl[66] br[66] wl[127] vdd gnd cell_6t
Xbit_r128_c66 bl[66] br[66] wl[128] vdd gnd cell_6t
Xbit_r129_c66 bl[66] br[66] wl[129] vdd gnd cell_6t
Xbit_r130_c66 bl[66] br[66] wl[130] vdd gnd cell_6t
Xbit_r131_c66 bl[66] br[66] wl[131] vdd gnd cell_6t
Xbit_r132_c66 bl[66] br[66] wl[132] vdd gnd cell_6t
Xbit_r133_c66 bl[66] br[66] wl[133] vdd gnd cell_6t
Xbit_r134_c66 bl[66] br[66] wl[134] vdd gnd cell_6t
Xbit_r135_c66 bl[66] br[66] wl[135] vdd gnd cell_6t
Xbit_r136_c66 bl[66] br[66] wl[136] vdd gnd cell_6t
Xbit_r137_c66 bl[66] br[66] wl[137] vdd gnd cell_6t
Xbit_r138_c66 bl[66] br[66] wl[138] vdd gnd cell_6t
Xbit_r139_c66 bl[66] br[66] wl[139] vdd gnd cell_6t
Xbit_r140_c66 bl[66] br[66] wl[140] vdd gnd cell_6t
Xbit_r141_c66 bl[66] br[66] wl[141] vdd gnd cell_6t
Xbit_r142_c66 bl[66] br[66] wl[142] vdd gnd cell_6t
Xbit_r143_c66 bl[66] br[66] wl[143] vdd gnd cell_6t
Xbit_r144_c66 bl[66] br[66] wl[144] vdd gnd cell_6t
Xbit_r145_c66 bl[66] br[66] wl[145] vdd gnd cell_6t
Xbit_r146_c66 bl[66] br[66] wl[146] vdd gnd cell_6t
Xbit_r147_c66 bl[66] br[66] wl[147] vdd gnd cell_6t
Xbit_r148_c66 bl[66] br[66] wl[148] vdd gnd cell_6t
Xbit_r149_c66 bl[66] br[66] wl[149] vdd gnd cell_6t
Xbit_r150_c66 bl[66] br[66] wl[150] vdd gnd cell_6t
Xbit_r151_c66 bl[66] br[66] wl[151] vdd gnd cell_6t
Xbit_r152_c66 bl[66] br[66] wl[152] vdd gnd cell_6t
Xbit_r153_c66 bl[66] br[66] wl[153] vdd gnd cell_6t
Xbit_r154_c66 bl[66] br[66] wl[154] vdd gnd cell_6t
Xbit_r155_c66 bl[66] br[66] wl[155] vdd gnd cell_6t
Xbit_r156_c66 bl[66] br[66] wl[156] vdd gnd cell_6t
Xbit_r157_c66 bl[66] br[66] wl[157] vdd gnd cell_6t
Xbit_r158_c66 bl[66] br[66] wl[158] vdd gnd cell_6t
Xbit_r159_c66 bl[66] br[66] wl[159] vdd gnd cell_6t
Xbit_r160_c66 bl[66] br[66] wl[160] vdd gnd cell_6t
Xbit_r161_c66 bl[66] br[66] wl[161] vdd gnd cell_6t
Xbit_r162_c66 bl[66] br[66] wl[162] vdd gnd cell_6t
Xbit_r163_c66 bl[66] br[66] wl[163] vdd gnd cell_6t
Xbit_r164_c66 bl[66] br[66] wl[164] vdd gnd cell_6t
Xbit_r165_c66 bl[66] br[66] wl[165] vdd gnd cell_6t
Xbit_r166_c66 bl[66] br[66] wl[166] vdd gnd cell_6t
Xbit_r167_c66 bl[66] br[66] wl[167] vdd gnd cell_6t
Xbit_r168_c66 bl[66] br[66] wl[168] vdd gnd cell_6t
Xbit_r169_c66 bl[66] br[66] wl[169] vdd gnd cell_6t
Xbit_r170_c66 bl[66] br[66] wl[170] vdd gnd cell_6t
Xbit_r171_c66 bl[66] br[66] wl[171] vdd gnd cell_6t
Xbit_r172_c66 bl[66] br[66] wl[172] vdd gnd cell_6t
Xbit_r173_c66 bl[66] br[66] wl[173] vdd gnd cell_6t
Xbit_r174_c66 bl[66] br[66] wl[174] vdd gnd cell_6t
Xbit_r175_c66 bl[66] br[66] wl[175] vdd gnd cell_6t
Xbit_r176_c66 bl[66] br[66] wl[176] vdd gnd cell_6t
Xbit_r177_c66 bl[66] br[66] wl[177] vdd gnd cell_6t
Xbit_r178_c66 bl[66] br[66] wl[178] vdd gnd cell_6t
Xbit_r179_c66 bl[66] br[66] wl[179] vdd gnd cell_6t
Xbit_r180_c66 bl[66] br[66] wl[180] vdd gnd cell_6t
Xbit_r181_c66 bl[66] br[66] wl[181] vdd gnd cell_6t
Xbit_r182_c66 bl[66] br[66] wl[182] vdd gnd cell_6t
Xbit_r183_c66 bl[66] br[66] wl[183] vdd gnd cell_6t
Xbit_r184_c66 bl[66] br[66] wl[184] vdd gnd cell_6t
Xbit_r185_c66 bl[66] br[66] wl[185] vdd gnd cell_6t
Xbit_r186_c66 bl[66] br[66] wl[186] vdd gnd cell_6t
Xbit_r187_c66 bl[66] br[66] wl[187] vdd gnd cell_6t
Xbit_r188_c66 bl[66] br[66] wl[188] vdd gnd cell_6t
Xbit_r189_c66 bl[66] br[66] wl[189] vdd gnd cell_6t
Xbit_r190_c66 bl[66] br[66] wl[190] vdd gnd cell_6t
Xbit_r191_c66 bl[66] br[66] wl[191] vdd gnd cell_6t
Xbit_r192_c66 bl[66] br[66] wl[192] vdd gnd cell_6t
Xbit_r193_c66 bl[66] br[66] wl[193] vdd gnd cell_6t
Xbit_r194_c66 bl[66] br[66] wl[194] vdd gnd cell_6t
Xbit_r195_c66 bl[66] br[66] wl[195] vdd gnd cell_6t
Xbit_r196_c66 bl[66] br[66] wl[196] vdd gnd cell_6t
Xbit_r197_c66 bl[66] br[66] wl[197] vdd gnd cell_6t
Xbit_r198_c66 bl[66] br[66] wl[198] vdd gnd cell_6t
Xbit_r199_c66 bl[66] br[66] wl[199] vdd gnd cell_6t
Xbit_r200_c66 bl[66] br[66] wl[200] vdd gnd cell_6t
Xbit_r201_c66 bl[66] br[66] wl[201] vdd gnd cell_6t
Xbit_r202_c66 bl[66] br[66] wl[202] vdd gnd cell_6t
Xbit_r203_c66 bl[66] br[66] wl[203] vdd gnd cell_6t
Xbit_r204_c66 bl[66] br[66] wl[204] vdd gnd cell_6t
Xbit_r205_c66 bl[66] br[66] wl[205] vdd gnd cell_6t
Xbit_r206_c66 bl[66] br[66] wl[206] vdd gnd cell_6t
Xbit_r207_c66 bl[66] br[66] wl[207] vdd gnd cell_6t
Xbit_r208_c66 bl[66] br[66] wl[208] vdd gnd cell_6t
Xbit_r209_c66 bl[66] br[66] wl[209] vdd gnd cell_6t
Xbit_r210_c66 bl[66] br[66] wl[210] vdd gnd cell_6t
Xbit_r211_c66 bl[66] br[66] wl[211] vdd gnd cell_6t
Xbit_r212_c66 bl[66] br[66] wl[212] vdd gnd cell_6t
Xbit_r213_c66 bl[66] br[66] wl[213] vdd gnd cell_6t
Xbit_r214_c66 bl[66] br[66] wl[214] vdd gnd cell_6t
Xbit_r215_c66 bl[66] br[66] wl[215] vdd gnd cell_6t
Xbit_r216_c66 bl[66] br[66] wl[216] vdd gnd cell_6t
Xbit_r217_c66 bl[66] br[66] wl[217] vdd gnd cell_6t
Xbit_r218_c66 bl[66] br[66] wl[218] vdd gnd cell_6t
Xbit_r219_c66 bl[66] br[66] wl[219] vdd gnd cell_6t
Xbit_r220_c66 bl[66] br[66] wl[220] vdd gnd cell_6t
Xbit_r221_c66 bl[66] br[66] wl[221] vdd gnd cell_6t
Xbit_r222_c66 bl[66] br[66] wl[222] vdd gnd cell_6t
Xbit_r223_c66 bl[66] br[66] wl[223] vdd gnd cell_6t
Xbit_r224_c66 bl[66] br[66] wl[224] vdd gnd cell_6t
Xbit_r225_c66 bl[66] br[66] wl[225] vdd gnd cell_6t
Xbit_r226_c66 bl[66] br[66] wl[226] vdd gnd cell_6t
Xbit_r227_c66 bl[66] br[66] wl[227] vdd gnd cell_6t
Xbit_r228_c66 bl[66] br[66] wl[228] vdd gnd cell_6t
Xbit_r229_c66 bl[66] br[66] wl[229] vdd gnd cell_6t
Xbit_r230_c66 bl[66] br[66] wl[230] vdd gnd cell_6t
Xbit_r231_c66 bl[66] br[66] wl[231] vdd gnd cell_6t
Xbit_r232_c66 bl[66] br[66] wl[232] vdd gnd cell_6t
Xbit_r233_c66 bl[66] br[66] wl[233] vdd gnd cell_6t
Xbit_r234_c66 bl[66] br[66] wl[234] vdd gnd cell_6t
Xbit_r235_c66 bl[66] br[66] wl[235] vdd gnd cell_6t
Xbit_r236_c66 bl[66] br[66] wl[236] vdd gnd cell_6t
Xbit_r237_c66 bl[66] br[66] wl[237] vdd gnd cell_6t
Xbit_r238_c66 bl[66] br[66] wl[238] vdd gnd cell_6t
Xbit_r239_c66 bl[66] br[66] wl[239] vdd gnd cell_6t
Xbit_r240_c66 bl[66] br[66] wl[240] vdd gnd cell_6t
Xbit_r241_c66 bl[66] br[66] wl[241] vdd gnd cell_6t
Xbit_r242_c66 bl[66] br[66] wl[242] vdd gnd cell_6t
Xbit_r243_c66 bl[66] br[66] wl[243] vdd gnd cell_6t
Xbit_r244_c66 bl[66] br[66] wl[244] vdd gnd cell_6t
Xbit_r245_c66 bl[66] br[66] wl[245] vdd gnd cell_6t
Xbit_r246_c66 bl[66] br[66] wl[246] vdd gnd cell_6t
Xbit_r247_c66 bl[66] br[66] wl[247] vdd gnd cell_6t
Xbit_r248_c66 bl[66] br[66] wl[248] vdd gnd cell_6t
Xbit_r249_c66 bl[66] br[66] wl[249] vdd gnd cell_6t
Xbit_r250_c66 bl[66] br[66] wl[250] vdd gnd cell_6t
Xbit_r251_c66 bl[66] br[66] wl[251] vdd gnd cell_6t
Xbit_r252_c66 bl[66] br[66] wl[252] vdd gnd cell_6t
Xbit_r253_c66 bl[66] br[66] wl[253] vdd gnd cell_6t
Xbit_r254_c66 bl[66] br[66] wl[254] vdd gnd cell_6t
Xbit_r255_c66 bl[66] br[66] wl[255] vdd gnd cell_6t
Xbit_r0_c67 bl[67] br[67] wl[0] vdd gnd cell_6t
Xbit_r1_c67 bl[67] br[67] wl[1] vdd gnd cell_6t
Xbit_r2_c67 bl[67] br[67] wl[2] vdd gnd cell_6t
Xbit_r3_c67 bl[67] br[67] wl[3] vdd gnd cell_6t
Xbit_r4_c67 bl[67] br[67] wl[4] vdd gnd cell_6t
Xbit_r5_c67 bl[67] br[67] wl[5] vdd gnd cell_6t
Xbit_r6_c67 bl[67] br[67] wl[6] vdd gnd cell_6t
Xbit_r7_c67 bl[67] br[67] wl[7] vdd gnd cell_6t
Xbit_r8_c67 bl[67] br[67] wl[8] vdd gnd cell_6t
Xbit_r9_c67 bl[67] br[67] wl[9] vdd gnd cell_6t
Xbit_r10_c67 bl[67] br[67] wl[10] vdd gnd cell_6t
Xbit_r11_c67 bl[67] br[67] wl[11] vdd gnd cell_6t
Xbit_r12_c67 bl[67] br[67] wl[12] vdd gnd cell_6t
Xbit_r13_c67 bl[67] br[67] wl[13] vdd gnd cell_6t
Xbit_r14_c67 bl[67] br[67] wl[14] vdd gnd cell_6t
Xbit_r15_c67 bl[67] br[67] wl[15] vdd gnd cell_6t
Xbit_r16_c67 bl[67] br[67] wl[16] vdd gnd cell_6t
Xbit_r17_c67 bl[67] br[67] wl[17] vdd gnd cell_6t
Xbit_r18_c67 bl[67] br[67] wl[18] vdd gnd cell_6t
Xbit_r19_c67 bl[67] br[67] wl[19] vdd gnd cell_6t
Xbit_r20_c67 bl[67] br[67] wl[20] vdd gnd cell_6t
Xbit_r21_c67 bl[67] br[67] wl[21] vdd gnd cell_6t
Xbit_r22_c67 bl[67] br[67] wl[22] vdd gnd cell_6t
Xbit_r23_c67 bl[67] br[67] wl[23] vdd gnd cell_6t
Xbit_r24_c67 bl[67] br[67] wl[24] vdd gnd cell_6t
Xbit_r25_c67 bl[67] br[67] wl[25] vdd gnd cell_6t
Xbit_r26_c67 bl[67] br[67] wl[26] vdd gnd cell_6t
Xbit_r27_c67 bl[67] br[67] wl[27] vdd gnd cell_6t
Xbit_r28_c67 bl[67] br[67] wl[28] vdd gnd cell_6t
Xbit_r29_c67 bl[67] br[67] wl[29] vdd gnd cell_6t
Xbit_r30_c67 bl[67] br[67] wl[30] vdd gnd cell_6t
Xbit_r31_c67 bl[67] br[67] wl[31] vdd gnd cell_6t
Xbit_r32_c67 bl[67] br[67] wl[32] vdd gnd cell_6t
Xbit_r33_c67 bl[67] br[67] wl[33] vdd gnd cell_6t
Xbit_r34_c67 bl[67] br[67] wl[34] vdd gnd cell_6t
Xbit_r35_c67 bl[67] br[67] wl[35] vdd gnd cell_6t
Xbit_r36_c67 bl[67] br[67] wl[36] vdd gnd cell_6t
Xbit_r37_c67 bl[67] br[67] wl[37] vdd gnd cell_6t
Xbit_r38_c67 bl[67] br[67] wl[38] vdd gnd cell_6t
Xbit_r39_c67 bl[67] br[67] wl[39] vdd gnd cell_6t
Xbit_r40_c67 bl[67] br[67] wl[40] vdd gnd cell_6t
Xbit_r41_c67 bl[67] br[67] wl[41] vdd gnd cell_6t
Xbit_r42_c67 bl[67] br[67] wl[42] vdd gnd cell_6t
Xbit_r43_c67 bl[67] br[67] wl[43] vdd gnd cell_6t
Xbit_r44_c67 bl[67] br[67] wl[44] vdd gnd cell_6t
Xbit_r45_c67 bl[67] br[67] wl[45] vdd gnd cell_6t
Xbit_r46_c67 bl[67] br[67] wl[46] vdd gnd cell_6t
Xbit_r47_c67 bl[67] br[67] wl[47] vdd gnd cell_6t
Xbit_r48_c67 bl[67] br[67] wl[48] vdd gnd cell_6t
Xbit_r49_c67 bl[67] br[67] wl[49] vdd gnd cell_6t
Xbit_r50_c67 bl[67] br[67] wl[50] vdd gnd cell_6t
Xbit_r51_c67 bl[67] br[67] wl[51] vdd gnd cell_6t
Xbit_r52_c67 bl[67] br[67] wl[52] vdd gnd cell_6t
Xbit_r53_c67 bl[67] br[67] wl[53] vdd gnd cell_6t
Xbit_r54_c67 bl[67] br[67] wl[54] vdd gnd cell_6t
Xbit_r55_c67 bl[67] br[67] wl[55] vdd gnd cell_6t
Xbit_r56_c67 bl[67] br[67] wl[56] vdd gnd cell_6t
Xbit_r57_c67 bl[67] br[67] wl[57] vdd gnd cell_6t
Xbit_r58_c67 bl[67] br[67] wl[58] vdd gnd cell_6t
Xbit_r59_c67 bl[67] br[67] wl[59] vdd gnd cell_6t
Xbit_r60_c67 bl[67] br[67] wl[60] vdd gnd cell_6t
Xbit_r61_c67 bl[67] br[67] wl[61] vdd gnd cell_6t
Xbit_r62_c67 bl[67] br[67] wl[62] vdd gnd cell_6t
Xbit_r63_c67 bl[67] br[67] wl[63] vdd gnd cell_6t
Xbit_r64_c67 bl[67] br[67] wl[64] vdd gnd cell_6t
Xbit_r65_c67 bl[67] br[67] wl[65] vdd gnd cell_6t
Xbit_r66_c67 bl[67] br[67] wl[66] vdd gnd cell_6t
Xbit_r67_c67 bl[67] br[67] wl[67] vdd gnd cell_6t
Xbit_r68_c67 bl[67] br[67] wl[68] vdd gnd cell_6t
Xbit_r69_c67 bl[67] br[67] wl[69] vdd gnd cell_6t
Xbit_r70_c67 bl[67] br[67] wl[70] vdd gnd cell_6t
Xbit_r71_c67 bl[67] br[67] wl[71] vdd gnd cell_6t
Xbit_r72_c67 bl[67] br[67] wl[72] vdd gnd cell_6t
Xbit_r73_c67 bl[67] br[67] wl[73] vdd gnd cell_6t
Xbit_r74_c67 bl[67] br[67] wl[74] vdd gnd cell_6t
Xbit_r75_c67 bl[67] br[67] wl[75] vdd gnd cell_6t
Xbit_r76_c67 bl[67] br[67] wl[76] vdd gnd cell_6t
Xbit_r77_c67 bl[67] br[67] wl[77] vdd gnd cell_6t
Xbit_r78_c67 bl[67] br[67] wl[78] vdd gnd cell_6t
Xbit_r79_c67 bl[67] br[67] wl[79] vdd gnd cell_6t
Xbit_r80_c67 bl[67] br[67] wl[80] vdd gnd cell_6t
Xbit_r81_c67 bl[67] br[67] wl[81] vdd gnd cell_6t
Xbit_r82_c67 bl[67] br[67] wl[82] vdd gnd cell_6t
Xbit_r83_c67 bl[67] br[67] wl[83] vdd gnd cell_6t
Xbit_r84_c67 bl[67] br[67] wl[84] vdd gnd cell_6t
Xbit_r85_c67 bl[67] br[67] wl[85] vdd gnd cell_6t
Xbit_r86_c67 bl[67] br[67] wl[86] vdd gnd cell_6t
Xbit_r87_c67 bl[67] br[67] wl[87] vdd gnd cell_6t
Xbit_r88_c67 bl[67] br[67] wl[88] vdd gnd cell_6t
Xbit_r89_c67 bl[67] br[67] wl[89] vdd gnd cell_6t
Xbit_r90_c67 bl[67] br[67] wl[90] vdd gnd cell_6t
Xbit_r91_c67 bl[67] br[67] wl[91] vdd gnd cell_6t
Xbit_r92_c67 bl[67] br[67] wl[92] vdd gnd cell_6t
Xbit_r93_c67 bl[67] br[67] wl[93] vdd gnd cell_6t
Xbit_r94_c67 bl[67] br[67] wl[94] vdd gnd cell_6t
Xbit_r95_c67 bl[67] br[67] wl[95] vdd gnd cell_6t
Xbit_r96_c67 bl[67] br[67] wl[96] vdd gnd cell_6t
Xbit_r97_c67 bl[67] br[67] wl[97] vdd gnd cell_6t
Xbit_r98_c67 bl[67] br[67] wl[98] vdd gnd cell_6t
Xbit_r99_c67 bl[67] br[67] wl[99] vdd gnd cell_6t
Xbit_r100_c67 bl[67] br[67] wl[100] vdd gnd cell_6t
Xbit_r101_c67 bl[67] br[67] wl[101] vdd gnd cell_6t
Xbit_r102_c67 bl[67] br[67] wl[102] vdd gnd cell_6t
Xbit_r103_c67 bl[67] br[67] wl[103] vdd gnd cell_6t
Xbit_r104_c67 bl[67] br[67] wl[104] vdd gnd cell_6t
Xbit_r105_c67 bl[67] br[67] wl[105] vdd gnd cell_6t
Xbit_r106_c67 bl[67] br[67] wl[106] vdd gnd cell_6t
Xbit_r107_c67 bl[67] br[67] wl[107] vdd gnd cell_6t
Xbit_r108_c67 bl[67] br[67] wl[108] vdd gnd cell_6t
Xbit_r109_c67 bl[67] br[67] wl[109] vdd gnd cell_6t
Xbit_r110_c67 bl[67] br[67] wl[110] vdd gnd cell_6t
Xbit_r111_c67 bl[67] br[67] wl[111] vdd gnd cell_6t
Xbit_r112_c67 bl[67] br[67] wl[112] vdd gnd cell_6t
Xbit_r113_c67 bl[67] br[67] wl[113] vdd gnd cell_6t
Xbit_r114_c67 bl[67] br[67] wl[114] vdd gnd cell_6t
Xbit_r115_c67 bl[67] br[67] wl[115] vdd gnd cell_6t
Xbit_r116_c67 bl[67] br[67] wl[116] vdd gnd cell_6t
Xbit_r117_c67 bl[67] br[67] wl[117] vdd gnd cell_6t
Xbit_r118_c67 bl[67] br[67] wl[118] vdd gnd cell_6t
Xbit_r119_c67 bl[67] br[67] wl[119] vdd gnd cell_6t
Xbit_r120_c67 bl[67] br[67] wl[120] vdd gnd cell_6t
Xbit_r121_c67 bl[67] br[67] wl[121] vdd gnd cell_6t
Xbit_r122_c67 bl[67] br[67] wl[122] vdd gnd cell_6t
Xbit_r123_c67 bl[67] br[67] wl[123] vdd gnd cell_6t
Xbit_r124_c67 bl[67] br[67] wl[124] vdd gnd cell_6t
Xbit_r125_c67 bl[67] br[67] wl[125] vdd gnd cell_6t
Xbit_r126_c67 bl[67] br[67] wl[126] vdd gnd cell_6t
Xbit_r127_c67 bl[67] br[67] wl[127] vdd gnd cell_6t
Xbit_r128_c67 bl[67] br[67] wl[128] vdd gnd cell_6t
Xbit_r129_c67 bl[67] br[67] wl[129] vdd gnd cell_6t
Xbit_r130_c67 bl[67] br[67] wl[130] vdd gnd cell_6t
Xbit_r131_c67 bl[67] br[67] wl[131] vdd gnd cell_6t
Xbit_r132_c67 bl[67] br[67] wl[132] vdd gnd cell_6t
Xbit_r133_c67 bl[67] br[67] wl[133] vdd gnd cell_6t
Xbit_r134_c67 bl[67] br[67] wl[134] vdd gnd cell_6t
Xbit_r135_c67 bl[67] br[67] wl[135] vdd gnd cell_6t
Xbit_r136_c67 bl[67] br[67] wl[136] vdd gnd cell_6t
Xbit_r137_c67 bl[67] br[67] wl[137] vdd gnd cell_6t
Xbit_r138_c67 bl[67] br[67] wl[138] vdd gnd cell_6t
Xbit_r139_c67 bl[67] br[67] wl[139] vdd gnd cell_6t
Xbit_r140_c67 bl[67] br[67] wl[140] vdd gnd cell_6t
Xbit_r141_c67 bl[67] br[67] wl[141] vdd gnd cell_6t
Xbit_r142_c67 bl[67] br[67] wl[142] vdd gnd cell_6t
Xbit_r143_c67 bl[67] br[67] wl[143] vdd gnd cell_6t
Xbit_r144_c67 bl[67] br[67] wl[144] vdd gnd cell_6t
Xbit_r145_c67 bl[67] br[67] wl[145] vdd gnd cell_6t
Xbit_r146_c67 bl[67] br[67] wl[146] vdd gnd cell_6t
Xbit_r147_c67 bl[67] br[67] wl[147] vdd gnd cell_6t
Xbit_r148_c67 bl[67] br[67] wl[148] vdd gnd cell_6t
Xbit_r149_c67 bl[67] br[67] wl[149] vdd gnd cell_6t
Xbit_r150_c67 bl[67] br[67] wl[150] vdd gnd cell_6t
Xbit_r151_c67 bl[67] br[67] wl[151] vdd gnd cell_6t
Xbit_r152_c67 bl[67] br[67] wl[152] vdd gnd cell_6t
Xbit_r153_c67 bl[67] br[67] wl[153] vdd gnd cell_6t
Xbit_r154_c67 bl[67] br[67] wl[154] vdd gnd cell_6t
Xbit_r155_c67 bl[67] br[67] wl[155] vdd gnd cell_6t
Xbit_r156_c67 bl[67] br[67] wl[156] vdd gnd cell_6t
Xbit_r157_c67 bl[67] br[67] wl[157] vdd gnd cell_6t
Xbit_r158_c67 bl[67] br[67] wl[158] vdd gnd cell_6t
Xbit_r159_c67 bl[67] br[67] wl[159] vdd gnd cell_6t
Xbit_r160_c67 bl[67] br[67] wl[160] vdd gnd cell_6t
Xbit_r161_c67 bl[67] br[67] wl[161] vdd gnd cell_6t
Xbit_r162_c67 bl[67] br[67] wl[162] vdd gnd cell_6t
Xbit_r163_c67 bl[67] br[67] wl[163] vdd gnd cell_6t
Xbit_r164_c67 bl[67] br[67] wl[164] vdd gnd cell_6t
Xbit_r165_c67 bl[67] br[67] wl[165] vdd gnd cell_6t
Xbit_r166_c67 bl[67] br[67] wl[166] vdd gnd cell_6t
Xbit_r167_c67 bl[67] br[67] wl[167] vdd gnd cell_6t
Xbit_r168_c67 bl[67] br[67] wl[168] vdd gnd cell_6t
Xbit_r169_c67 bl[67] br[67] wl[169] vdd gnd cell_6t
Xbit_r170_c67 bl[67] br[67] wl[170] vdd gnd cell_6t
Xbit_r171_c67 bl[67] br[67] wl[171] vdd gnd cell_6t
Xbit_r172_c67 bl[67] br[67] wl[172] vdd gnd cell_6t
Xbit_r173_c67 bl[67] br[67] wl[173] vdd gnd cell_6t
Xbit_r174_c67 bl[67] br[67] wl[174] vdd gnd cell_6t
Xbit_r175_c67 bl[67] br[67] wl[175] vdd gnd cell_6t
Xbit_r176_c67 bl[67] br[67] wl[176] vdd gnd cell_6t
Xbit_r177_c67 bl[67] br[67] wl[177] vdd gnd cell_6t
Xbit_r178_c67 bl[67] br[67] wl[178] vdd gnd cell_6t
Xbit_r179_c67 bl[67] br[67] wl[179] vdd gnd cell_6t
Xbit_r180_c67 bl[67] br[67] wl[180] vdd gnd cell_6t
Xbit_r181_c67 bl[67] br[67] wl[181] vdd gnd cell_6t
Xbit_r182_c67 bl[67] br[67] wl[182] vdd gnd cell_6t
Xbit_r183_c67 bl[67] br[67] wl[183] vdd gnd cell_6t
Xbit_r184_c67 bl[67] br[67] wl[184] vdd gnd cell_6t
Xbit_r185_c67 bl[67] br[67] wl[185] vdd gnd cell_6t
Xbit_r186_c67 bl[67] br[67] wl[186] vdd gnd cell_6t
Xbit_r187_c67 bl[67] br[67] wl[187] vdd gnd cell_6t
Xbit_r188_c67 bl[67] br[67] wl[188] vdd gnd cell_6t
Xbit_r189_c67 bl[67] br[67] wl[189] vdd gnd cell_6t
Xbit_r190_c67 bl[67] br[67] wl[190] vdd gnd cell_6t
Xbit_r191_c67 bl[67] br[67] wl[191] vdd gnd cell_6t
Xbit_r192_c67 bl[67] br[67] wl[192] vdd gnd cell_6t
Xbit_r193_c67 bl[67] br[67] wl[193] vdd gnd cell_6t
Xbit_r194_c67 bl[67] br[67] wl[194] vdd gnd cell_6t
Xbit_r195_c67 bl[67] br[67] wl[195] vdd gnd cell_6t
Xbit_r196_c67 bl[67] br[67] wl[196] vdd gnd cell_6t
Xbit_r197_c67 bl[67] br[67] wl[197] vdd gnd cell_6t
Xbit_r198_c67 bl[67] br[67] wl[198] vdd gnd cell_6t
Xbit_r199_c67 bl[67] br[67] wl[199] vdd gnd cell_6t
Xbit_r200_c67 bl[67] br[67] wl[200] vdd gnd cell_6t
Xbit_r201_c67 bl[67] br[67] wl[201] vdd gnd cell_6t
Xbit_r202_c67 bl[67] br[67] wl[202] vdd gnd cell_6t
Xbit_r203_c67 bl[67] br[67] wl[203] vdd gnd cell_6t
Xbit_r204_c67 bl[67] br[67] wl[204] vdd gnd cell_6t
Xbit_r205_c67 bl[67] br[67] wl[205] vdd gnd cell_6t
Xbit_r206_c67 bl[67] br[67] wl[206] vdd gnd cell_6t
Xbit_r207_c67 bl[67] br[67] wl[207] vdd gnd cell_6t
Xbit_r208_c67 bl[67] br[67] wl[208] vdd gnd cell_6t
Xbit_r209_c67 bl[67] br[67] wl[209] vdd gnd cell_6t
Xbit_r210_c67 bl[67] br[67] wl[210] vdd gnd cell_6t
Xbit_r211_c67 bl[67] br[67] wl[211] vdd gnd cell_6t
Xbit_r212_c67 bl[67] br[67] wl[212] vdd gnd cell_6t
Xbit_r213_c67 bl[67] br[67] wl[213] vdd gnd cell_6t
Xbit_r214_c67 bl[67] br[67] wl[214] vdd gnd cell_6t
Xbit_r215_c67 bl[67] br[67] wl[215] vdd gnd cell_6t
Xbit_r216_c67 bl[67] br[67] wl[216] vdd gnd cell_6t
Xbit_r217_c67 bl[67] br[67] wl[217] vdd gnd cell_6t
Xbit_r218_c67 bl[67] br[67] wl[218] vdd gnd cell_6t
Xbit_r219_c67 bl[67] br[67] wl[219] vdd gnd cell_6t
Xbit_r220_c67 bl[67] br[67] wl[220] vdd gnd cell_6t
Xbit_r221_c67 bl[67] br[67] wl[221] vdd gnd cell_6t
Xbit_r222_c67 bl[67] br[67] wl[222] vdd gnd cell_6t
Xbit_r223_c67 bl[67] br[67] wl[223] vdd gnd cell_6t
Xbit_r224_c67 bl[67] br[67] wl[224] vdd gnd cell_6t
Xbit_r225_c67 bl[67] br[67] wl[225] vdd gnd cell_6t
Xbit_r226_c67 bl[67] br[67] wl[226] vdd gnd cell_6t
Xbit_r227_c67 bl[67] br[67] wl[227] vdd gnd cell_6t
Xbit_r228_c67 bl[67] br[67] wl[228] vdd gnd cell_6t
Xbit_r229_c67 bl[67] br[67] wl[229] vdd gnd cell_6t
Xbit_r230_c67 bl[67] br[67] wl[230] vdd gnd cell_6t
Xbit_r231_c67 bl[67] br[67] wl[231] vdd gnd cell_6t
Xbit_r232_c67 bl[67] br[67] wl[232] vdd gnd cell_6t
Xbit_r233_c67 bl[67] br[67] wl[233] vdd gnd cell_6t
Xbit_r234_c67 bl[67] br[67] wl[234] vdd gnd cell_6t
Xbit_r235_c67 bl[67] br[67] wl[235] vdd gnd cell_6t
Xbit_r236_c67 bl[67] br[67] wl[236] vdd gnd cell_6t
Xbit_r237_c67 bl[67] br[67] wl[237] vdd gnd cell_6t
Xbit_r238_c67 bl[67] br[67] wl[238] vdd gnd cell_6t
Xbit_r239_c67 bl[67] br[67] wl[239] vdd gnd cell_6t
Xbit_r240_c67 bl[67] br[67] wl[240] vdd gnd cell_6t
Xbit_r241_c67 bl[67] br[67] wl[241] vdd gnd cell_6t
Xbit_r242_c67 bl[67] br[67] wl[242] vdd gnd cell_6t
Xbit_r243_c67 bl[67] br[67] wl[243] vdd gnd cell_6t
Xbit_r244_c67 bl[67] br[67] wl[244] vdd gnd cell_6t
Xbit_r245_c67 bl[67] br[67] wl[245] vdd gnd cell_6t
Xbit_r246_c67 bl[67] br[67] wl[246] vdd gnd cell_6t
Xbit_r247_c67 bl[67] br[67] wl[247] vdd gnd cell_6t
Xbit_r248_c67 bl[67] br[67] wl[248] vdd gnd cell_6t
Xbit_r249_c67 bl[67] br[67] wl[249] vdd gnd cell_6t
Xbit_r250_c67 bl[67] br[67] wl[250] vdd gnd cell_6t
Xbit_r251_c67 bl[67] br[67] wl[251] vdd gnd cell_6t
Xbit_r252_c67 bl[67] br[67] wl[252] vdd gnd cell_6t
Xbit_r253_c67 bl[67] br[67] wl[253] vdd gnd cell_6t
Xbit_r254_c67 bl[67] br[67] wl[254] vdd gnd cell_6t
Xbit_r255_c67 bl[67] br[67] wl[255] vdd gnd cell_6t
Xbit_r0_c68 bl[68] br[68] wl[0] vdd gnd cell_6t
Xbit_r1_c68 bl[68] br[68] wl[1] vdd gnd cell_6t
Xbit_r2_c68 bl[68] br[68] wl[2] vdd gnd cell_6t
Xbit_r3_c68 bl[68] br[68] wl[3] vdd gnd cell_6t
Xbit_r4_c68 bl[68] br[68] wl[4] vdd gnd cell_6t
Xbit_r5_c68 bl[68] br[68] wl[5] vdd gnd cell_6t
Xbit_r6_c68 bl[68] br[68] wl[6] vdd gnd cell_6t
Xbit_r7_c68 bl[68] br[68] wl[7] vdd gnd cell_6t
Xbit_r8_c68 bl[68] br[68] wl[8] vdd gnd cell_6t
Xbit_r9_c68 bl[68] br[68] wl[9] vdd gnd cell_6t
Xbit_r10_c68 bl[68] br[68] wl[10] vdd gnd cell_6t
Xbit_r11_c68 bl[68] br[68] wl[11] vdd gnd cell_6t
Xbit_r12_c68 bl[68] br[68] wl[12] vdd gnd cell_6t
Xbit_r13_c68 bl[68] br[68] wl[13] vdd gnd cell_6t
Xbit_r14_c68 bl[68] br[68] wl[14] vdd gnd cell_6t
Xbit_r15_c68 bl[68] br[68] wl[15] vdd gnd cell_6t
Xbit_r16_c68 bl[68] br[68] wl[16] vdd gnd cell_6t
Xbit_r17_c68 bl[68] br[68] wl[17] vdd gnd cell_6t
Xbit_r18_c68 bl[68] br[68] wl[18] vdd gnd cell_6t
Xbit_r19_c68 bl[68] br[68] wl[19] vdd gnd cell_6t
Xbit_r20_c68 bl[68] br[68] wl[20] vdd gnd cell_6t
Xbit_r21_c68 bl[68] br[68] wl[21] vdd gnd cell_6t
Xbit_r22_c68 bl[68] br[68] wl[22] vdd gnd cell_6t
Xbit_r23_c68 bl[68] br[68] wl[23] vdd gnd cell_6t
Xbit_r24_c68 bl[68] br[68] wl[24] vdd gnd cell_6t
Xbit_r25_c68 bl[68] br[68] wl[25] vdd gnd cell_6t
Xbit_r26_c68 bl[68] br[68] wl[26] vdd gnd cell_6t
Xbit_r27_c68 bl[68] br[68] wl[27] vdd gnd cell_6t
Xbit_r28_c68 bl[68] br[68] wl[28] vdd gnd cell_6t
Xbit_r29_c68 bl[68] br[68] wl[29] vdd gnd cell_6t
Xbit_r30_c68 bl[68] br[68] wl[30] vdd gnd cell_6t
Xbit_r31_c68 bl[68] br[68] wl[31] vdd gnd cell_6t
Xbit_r32_c68 bl[68] br[68] wl[32] vdd gnd cell_6t
Xbit_r33_c68 bl[68] br[68] wl[33] vdd gnd cell_6t
Xbit_r34_c68 bl[68] br[68] wl[34] vdd gnd cell_6t
Xbit_r35_c68 bl[68] br[68] wl[35] vdd gnd cell_6t
Xbit_r36_c68 bl[68] br[68] wl[36] vdd gnd cell_6t
Xbit_r37_c68 bl[68] br[68] wl[37] vdd gnd cell_6t
Xbit_r38_c68 bl[68] br[68] wl[38] vdd gnd cell_6t
Xbit_r39_c68 bl[68] br[68] wl[39] vdd gnd cell_6t
Xbit_r40_c68 bl[68] br[68] wl[40] vdd gnd cell_6t
Xbit_r41_c68 bl[68] br[68] wl[41] vdd gnd cell_6t
Xbit_r42_c68 bl[68] br[68] wl[42] vdd gnd cell_6t
Xbit_r43_c68 bl[68] br[68] wl[43] vdd gnd cell_6t
Xbit_r44_c68 bl[68] br[68] wl[44] vdd gnd cell_6t
Xbit_r45_c68 bl[68] br[68] wl[45] vdd gnd cell_6t
Xbit_r46_c68 bl[68] br[68] wl[46] vdd gnd cell_6t
Xbit_r47_c68 bl[68] br[68] wl[47] vdd gnd cell_6t
Xbit_r48_c68 bl[68] br[68] wl[48] vdd gnd cell_6t
Xbit_r49_c68 bl[68] br[68] wl[49] vdd gnd cell_6t
Xbit_r50_c68 bl[68] br[68] wl[50] vdd gnd cell_6t
Xbit_r51_c68 bl[68] br[68] wl[51] vdd gnd cell_6t
Xbit_r52_c68 bl[68] br[68] wl[52] vdd gnd cell_6t
Xbit_r53_c68 bl[68] br[68] wl[53] vdd gnd cell_6t
Xbit_r54_c68 bl[68] br[68] wl[54] vdd gnd cell_6t
Xbit_r55_c68 bl[68] br[68] wl[55] vdd gnd cell_6t
Xbit_r56_c68 bl[68] br[68] wl[56] vdd gnd cell_6t
Xbit_r57_c68 bl[68] br[68] wl[57] vdd gnd cell_6t
Xbit_r58_c68 bl[68] br[68] wl[58] vdd gnd cell_6t
Xbit_r59_c68 bl[68] br[68] wl[59] vdd gnd cell_6t
Xbit_r60_c68 bl[68] br[68] wl[60] vdd gnd cell_6t
Xbit_r61_c68 bl[68] br[68] wl[61] vdd gnd cell_6t
Xbit_r62_c68 bl[68] br[68] wl[62] vdd gnd cell_6t
Xbit_r63_c68 bl[68] br[68] wl[63] vdd gnd cell_6t
Xbit_r64_c68 bl[68] br[68] wl[64] vdd gnd cell_6t
Xbit_r65_c68 bl[68] br[68] wl[65] vdd gnd cell_6t
Xbit_r66_c68 bl[68] br[68] wl[66] vdd gnd cell_6t
Xbit_r67_c68 bl[68] br[68] wl[67] vdd gnd cell_6t
Xbit_r68_c68 bl[68] br[68] wl[68] vdd gnd cell_6t
Xbit_r69_c68 bl[68] br[68] wl[69] vdd gnd cell_6t
Xbit_r70_c68 bl[68] br[68] wl[70] vdd gnd cell_6t
Xbit_r71_c68 bl[68] br[68] wl[71] vdd gnd cell_6t
Xbit_r72_c68 bl[68] br[68] wl[72] vdd gnd cell_6t
Xbit_r73_c68 bl[68] br[68] wl[73] vdd gnd cell_6t
Xbit_r74_c68 bl[68] br[68] wl[74] vdd gnd cell_6t
Xbit_r75_c68 bl[68] br[68] wl[75] vdd gnd cell_6t
Xbit_r76_c68 bl[68] br[68] wl[76] vdd gnd cell_6t
Xbit_r77_c68 bl[68] br[68] wl[77] vdd gnd cell_6t
Xbit_r78_c68 bl[68] br[68] wl[78] vdd gnd cell_6t
Xbit_r79_c68 bl[68] br[68] wl[79] vdd gnd cell_6t
Xbit_r80_c68 bl[68] br[68] wl[80] vdd gnd cell_6t
Xbit_r81_c68 bl[68] br[68] wl[81] vdd gnd cell_6t
Xbit_r82_c68 bl[68] br[68] wl[82] vdd gnd cell_6t
Xbit_r83_c68 bl[68] br[68] wl[83] vdd gnd cell_6t
Xbit_r84_c68 bl[68] br[68] wl[84] vdd gnd cell_6t
Xbit_r85_c68 bl[68] br[68] wl[85] vdd gnd cell_6t
Xbit_r86_c68 bl[68] br[68] wl[86] vdd gnd cell_6t
Xbit_r87_c68 bl[68] br[68] wl[87] vdd gnd cell_6t
Xbit_r88_c68 bl[68] br[68] wl[88] vdd gnd cell_6t
Xbit_r89_c68 bl[68] br[68] wl[89] vdd gnd cell_6t
Xbit_r90_c68 bl[68] br[68] wl[90] vdd gnd cell_6t
Xbit_r91_c68 bl[68] br[68] wl[91] vdd gnd cell_6t
Xbit_r92_c68 bl[68] br[68] wl[92] vdd gnd cell_6t
Xbit_r93_c68 bl[68] br[68] wl[93] vdd gnd cell_6t
Xbit_r94_c68 bl[68] br[68] wl[94] vdd gnd cell_6t
Xbit_r95_c68 bl[68] br[68] wl[95] vdd gnd cell_6t
Xbit_r96_c68 bl[68] br[68] wl[96] vdd gnd cell_6t
Xbit_r97_c68 bl[68] br[68] wl[97] vdd gnd cell_6t
Xbit_r98_c68 bl[68] br[68] wl[98] vdd gnd cell_6t
Xbit_r99_c68 bl[68] br[68] wl[99] vdd gnd cell_6t
Xbit_r100_c68 bl[68] br[68] wl[100] vdd gnd cell_6t
Xbit_r101_c68 bl[68] br[68] wl[101] vdd gnd cell_6t
Xbit_r102_c68 bl[68] br[68] wl[102] vdd gnd cell_6t
Xbit_r103_c68 bl[68] br[68] wl[103] vdd gnd cell_6t
Xbit_r104_c68 bl[68] br[68] wl[104] vdd gnd cell_6t
Xbit_r105_c68 bl[68] br[68] wl[105] vdd gnd cell_6t
Xbit_r106_c68 bl[68] br[68] wl[106] vdd gnd cell_6t
Xbit_r107_c68 bl[68] br[68] wl[107] vdd gnd cell_6t
Xbit_r108_c68 bl[68] br[68] wl[108] vdd gnd cell_6t
Xbit_r109_c68 bl[68] br[68] wl[109] vdd gnd cell_6t
Xbit_r110_c68 bl[68] br[68] wl[110] vdd gnd cell_6t
Xbit_r111_c68 bl[68] br[68] wl[111] vdd gnd cell_6t
Xbit_r112_c68 bl[68] br[68] wl[112] vdd gnd cell_6t
Xbit_r113_c68 bl[68] br[68] wl[113] vdd gnd cell_6t
Xbit_r114_c68 bl[68] br[68] wl[114] vdd gnd cell_6t
Xbit_r115_c68 bl[68] br[68] wl[115] vdd gnd cell_6t
Xbit_r116_c68 bl[68] br[68] wl[116] vdd gnd cell_6t
Xbit_r117_c68 bl[68] br[68] wl[117] vdd gnd cell_6t
Xbit_r118_c68 bl[68] br[68] wl[118] vdd gnd cell_6t
Xbit_r119_c68 bl[68] br[68] wl[119] vdd gnd cell_6t
Xbit_r120_c68 bl[68] br[68] wl[120] vdd gnd cell_6t
Xbit_r121_c68 bl[68] br[68] wl[121] vdd gnd cell_6t
Xbit_r122_c68 bl[68] br[68] wl[122] vdd gnd cell_6t
Xbit_r123_c68 bl[68] br[68] wl[123] vdd gnd cell_6t
Xbit_r124_c68 bl[68] br[68] wl[124] vdd gnd cell_6t
Xbit_r125_c68 bl[68] br[68] wl[125] vdd gnd cell_6t
Xbit_r126_c68 bl[68] br[68] wl[126] vdd gnd cell_6t
Xbit_r127_c68 bl[68] br[68] wl[127] vdd gnd cell_6t
Xbit_r128_c68 bl[68] br[68] wl[128] vdd gnd cell_6t
Xbit_r129_c68 bl[68] br[68] wl[129] vdd gnd cell_6t
Xbit_r130_c68 bl[68] br[68] wl[130] vdd gnd cell_6t
Xbit_r131_c68 bl[68] br[68] wl[131] vdd gnd cell_6t
Xbit_r132_c68 bl[68] br[68] wl[132] vdd gnd cell_6t
Xbit_r133_c68 bl[68] br[68] wl[133] vdd gnd cell_6t
Xbit_r134_c68 bl[68] br[68] wl[134] vdd gnd cell_6t
Xbit_r135_c68 bl[68] br[68] wl[135] vdd gnd cell_6t
Xbit_r136_c68 bl[68] br[68] wl[136] vdd gnd cell_6t
Xbit_r137_c68 bl[68] br[68] wl[137] vdd gnd cell_6t
Xbit_r138_c68 bl[68] br[68] wl[138] vdd gnd cell_6t
Xbit_r139_c68 bl[68] br[68] wl[139] vdd gnd cell_6t
Xbit_r140_c68 bl[68] br[68] wl[140] vdd gnd cell_6t
Xbit_r141_c68 bl[68] br[68] wl[141] vdd gnd cell_6t
Xbit_r142_c68 bl[68] br[68] wl[142] vdd gnd cell_6t
Xbit_r143_c68 bl[68] br[68] wl[143] vdd gnd cell_6t
Xbit_r144_c68 bl[68] br[68] wl[144] vdd gnd cell_6t
Xbit_r145_c68 bl[68] br[68] wl[145] vdd gnd cell_6t
Xbit_r146_c68 bl[68] br[68] wl[146] vdd gnd cell_6t
Xbit_r147_c68 bl[68] br[68] wl[147] vdd gnd cell_6t
Xbit_r148_c68 bl[68] br[68] wl[148] vdd gnd cell_6t
Xbit_r149_c68 bl[68] br[68] wl[149] vdd gnd cell_6t
Xbit_r150_c68 bl[68] br[68] wl[150] vdd gnd cell_6t
Xbit_r151_c68 bl[68] br[68] wl[151] vdd gnd cell_6t
Xbit_r152_c68 bl[68] br[68] wl[152] vdd gnd cell_6t
Xbit_r153_c68 bl[68] br[68] wl[153] vdd gnd cell_6t
Xbit_r154_c68 bl[68] br[68] wl[154] vdd gnd cell_6t
Xbit_r155_c68 bl[68] br[68] wl[155] vdd gnd cell_6t
Xbit_r156_c68 bl[68] br[68] wl[156] vdd gnd cell_6t
Xbit_r157_c68 bl[68] br[68] wl[157] vdd gnd cell_6t
Xbit_r158_c68 bl[68] br[68] wl[158] vdd gnd cell_6t
Xbit_r159_c68 bl[68] br[68] wl[159] vdd gnd cell_6t
Xbit_r160_c68 bl[68] br[68] wl[160] vdd gnd cell_6t
Xbit_r161_c68 bl[68] br[68] wl[161] vdd gnd cell_6t
Xbit_r162_c68 bl[68] br[68] wl[162] vdd gnd cell_6t
Xbit_r163_c68 bl[68] br[68] wl[163] vdd gnd cell_6t
Xbit_r164_c68 bl[68] br[68] wl[164] vdd gnd cell_6t
Xbit_r165_c68 bl[68] br[68] wl[165] vdd gnd cell_6t
Xbit_r166_c68 bl[68] br[68] wl[166] vdd gnd cell_6t
Xbit_r167_c68 bl[68] br[68] wl[167] vdd gnd cell_6t
Xbit_r168_c68 bl[68] br[68] wl[168] vdd gnd cell_6t
Xbit_r169_c68 bl[68] br[68] wl[169] vdd gnd cell_6t
Xbit_r170_c68 bl[68] br[68] wl[170] vdd gnd cell_6t
Xbit_r171_c68 bl[68] br[68] wl[171] vdd gnd cell_6t
Xbit_r172_c68 bl[68] br[68] wl[172] vdd gnd cell_6t
Xbit_r173_c68 bl[68] br[68] wl[173] vdd gnd cell_6t
Xbit_r174_c68 bl[68] br[68] wl[174] vdd gnd cell_6t
Xbit_r175_c68 bl[68] br[68] wl[175] vdd gnd cell_6t
Xbit_r176_c68 bl[68] br[68] wl[176] vdd gnd cell_6t
Xbit_r177_c68 bl[68] br[68] wl[177] vdd gnd cell_6t
Xbit_r178_c68 bl[68] br[68] wl[178] vdd gnd cell_6t
Xbit_r179_c68 bl[68] br[68] wl[179] vdd gnd cell_6t
Xbit_r180_c68 bl[68] br[68] wl[180] vdd gnd cell_6t
Xbit_r181_c68 bl[68] br[68] wl[181] vdd gnd cell_6t
Xbit_r182_c68 bl[68] br[68] wl[182] vdd gnd cell_6t
Xbit_r183_c68 bl[68] br[68] wl[183] vdd gnd cell_6t
Xbit_r184_c68 bl[68] br[68] wl[184] vdd gnd cell_6t
Xbit_r185_c68 bl[68] br[68] wl[185] vdd gnd cell_6t
Xbit_r186_c68 bl[68] br[68] wl[186] vdd gnd cell_6t
Xbit_r187_c68 bl[68] br[68] wl[187] vdd gnd cell_6t
Xbit_r188_c68 bl[68] br[68] wl[188] vdd gnd cell_6t
Xbit_r189_c68 bl[68] br[68] wl[189] vdd gnd cell_6t
Xbit_r190_c68 bl[68] br[68] wl[190] vdd gnd cell_6t
Xbit_r191_c68 bl[68] br[68] wl[191] vdd gnd cell_6t
Xbit_r192_c68 bl[68] br[68] wl[192] vdd gnd cell_6t
Xbit_r193_c68 bl[68] br[68] wl[193] vdd gnd cell_6t
Xbit_r194_c68 bl[68] br[68] wl[194] vdd gnd cell_6t
Xbit_r195_c68 bl[68] br[68] wl[195] vdd gnd cell_6t
Xbit_r196_c68 bl[68] br[68] wl[196] vdd gnd cell_6t
Xbit_r197_c68 bl[68] br[68] wl[197] vdd gnd cell_6t
Xbit_r198_c68 bl[68] br[68] wl[198] vdd gnd cell_6t
Xbit_r199_c68 bl[68] br[68] wl[199] vdd gnd cell_6t
Xbit_r200_c68 bl[68] br[68] wl[200] vdd gnd cell_6t
Xbit_r201_c68 bl[68] br[68] wl[201] vdd gnd cell_6t
Xbit_r202_c68 bl[68] br[68] wl[202] vdd gnd cell_6t
Xbit_r203_c68 bl[68] br[68] wl[203] vdd gnd cell_6t
Xbit_r204_c68 bl[68] br[68] wl[204] vdd gnd cell_6t
Xbit_r205_c68 bl[68] br[68] wl[205] vdd gnd cell_6t
Xbit_r206_c68 bl[68] br[68] wl[206] vdd gnd cell_6t
Xbit_r207_c68 bl[68] br[68] wl[207] vdd gnd cell_6t
Xbit_r208_c68 bl[68] br[68] wl[208] vdd gnd cell_6t
Xbit_r209_c68 bl[68] br[68] wl[209] vdd gnd cell_6t
Xbit_r210_c68 bl[68] br[68] wl[210] vdd gnd cell_6t
Xbit_r211_c68 bl[68] br[68] wl[211] vdd gnd cell_6t
Xbit_r212_c68 bl[68] br[68] wl[212] vdd gnd cell_6t
Xbit_r213_c68 bl[68] br[68] wl[213] vdd gnd cell_6t
Xbit_r214_c68 bl[68] br[68] wl[214] vdd gnd cell_6t
Xbit_r215_c68 bl[68] br[68] wl[215] vdd gnd cell_6t
Xbit_r216_c68 bl[68] br[68] wl[216] vdd gnd cell_6t
Xbit_r217_c68 bl[68] br[68] wl[217] vdd gnd cell_6t
Xbit_r218_c68 bl[68] br[68] wl[218] vdd gnd cell_6t
Xbit_r219_c68 bl[68] br[68] wl[219] vdd gnd cell_6t
Xbit_r220_c68 bl[68] br[68] wl[220] vdd gnd cell_6t
Xbit_r221_c68 bl[68] br[68] wl[221] vdd gnd cell_6t
Xbit_r222_c68 bl[68] br[68] wl[222] vdd gnd cell_6t
Xbit_r223_c68 bl[68] br[68] wl[223] vdd gnd cell_6t
Xbit_r224_c68 bl[68] br[68] wl[224] vdd gnd cell_6t
Xbit_r225_c68 bl[68] br[68] wl[225] vdd gnd cell_6t
Xbit_r226_c68 bl[68] br[68] wl[226] vdd gnd cell_6t
Xbit_r227_c68 bl[68] br[68] wl[227] vdd gnd cell_6t
Xbit_r228_c68 bl[68] br[68] wl[228] vdd gnd cell_6t
Xbit_r229_c68 bl[68] br[68] wl[229] vdd gnd cell_6t
Xbit_r230_c68 bl[68] br[68] wl[230] vdd gnd cell_6t
Xbit_r231_c68 bl[68] br[68] wl[231] vdd gnd cell_6t
Xbit_r232_c68 bl[68] br[68] wl[232] vdd gnd cell_6t
Xbit_r233_c68 bl[68] br[68] wl[233] vdd gnd cell_6t
Xbit_r234_c68 bl[68] br[68] wl[234] vdd gnd cell_6t
Xbit_r235_c68 bl[68] br[68] wl[235] vdd gnd cell_6t
Xbit_r236_c68 bl[68] br[68] wl[236] vdd gnd cell_6t
Xbit_r237_c68 bl[68] br[68] wl[237] vdd gnd cell_6t
Xbit_r238_c68 bl[68] br[68] wl[238] vdd gnd cell_6t
Xbit_r239_c68 bl[68] br[68] wl[239] vdd gnd cell_6t
Xbit_r240_c68 bl[68] br[68] wl[240] vdd gnd cell_6t
Xbit_r241_c68 bl[68] br[68] wl[241] vdd gnd cell_6t
Xbit_r242_c68 bl[68] br[68] wl[242] vdd gnd cell_6t
Xbit_r243_c68 bl[68] br[68] wl[243] vdd gnd cell_6t
Xbit_r244_c68 bl[68] br[68] wl[244] vdd gnd cell_6t
Xbit_r245_c68 bl[68] br[68] wl[245] vdd gnd cell_6t
Xbit_r246_c68 bl[68] br[68] wl[246] vdd gnd cell_6t
Xbit_r247_c68 bl[68] br[68] wl[247] vdd gnd cell_6t
Xbit_r248_c68 bl[68] br[68] wl[248] vdd gnd cell_6t
Xbit_r249_c68 bl[68] br[68] wl[249] vdd gnd cell_6t
Xbit_r250_c68 bl[68] br[68] wl[250] vdd gnd cell_6t
Xbit_r251_c68 bl[68] br[68] wl[251] vdd gnd cell_6t
Xbit_r252_c68 bl[68] br[68] wl[252] vdd gnd cell_6t
Xbit_r253_c68 bl[68] br[68] wl[253] vdd gnd cell_6t
Xbit_r254_c68 bl[68] br[68] wl[254] vdd gnd cell_6t
Xbit_r255_c68 bl[68] br[68] wl[255] vdd gnd cell_6t
Xbit_r0_c69 bl[69] br[69] wl[0] vdd gnd cell_6t
Xbit_r1_c69 bl[69] br[69] wl[1] vdd gnd cell_6t
Xbit_r2_c69 bl[69] br[69] wl[2] vdd gnd cell_6t
Xbit_r3_c69 bl[69] br[69] wl[3] vdd gnd cell_6t
Xbit_r4_c69 bl[69] br[69] wl[4] vdd gnd cell_6t
Xbit_r5_c69 bl[69] br[69] wl[5] vdd gnd cell_6t
Xbit_r6_c69 bl[69] br[69] wl[6] vdd gnd cell_6t
Xbit_r7_c69 bl[69] br[69] wl[7] vdd gnd cell_6t
Xbit_r8_c69 bl[69] br[69] wl[8] vdd gnd cell_6t
Xbit_r9_c69 bl[69] br[69] wl[9] vdd gnd cell_6t
Xbit_r10_c69 bl[69] br[69] wl[10] vdd gnd cell_6t
Xbit_r11_c69 bl[69] br[69] wl[11] vdd gnd cell_6t
Xbit_r12_c69 bl[69] br[69] wl[12] vdd gnd cell_6t
Xbit_r13_c69 bl[69] br[69] wl[13] vdd gnd cell_6t
Xbit_r14_c69 bl[69] br[69] wl[14] vdd gnd cell_6t
Xbit_r15_c69 bl[69] br[69] wl[15] vdd gnd cell_6t
Xbit_r16_c69 bl[69] br[69] wl[16] vdd gnd cell_6t
Xbit_r17_c69 bl[69] br[69] wl[17] vdd gnd cell_6t
Xbit_r18_c69 bl[69] br[69] wl[18] vdd gnd cell_6t
Xbit_r19_c69 bl[69] br[69] wl[19] vdd gnd cell_6t
Xbit_r20_c69 bl[69] br[69] wl[20] vdd gnd cell_6t
Xbit_r21_c69 bl[69] br[69] wl[21] vdd gnd cell_6t
Xbit_r22_c69 bl[69] br[69] wl[22] vdd gnd cell_6t
Xbit_r23_c69 bl[69] br[69] wl[23] vdd gnd cell_6t
Xbit_r24_c69 bl[69] br[69] wl[24] vdd gnd cell_6t
Xbit_r25_c69 bl[69] br[69] wl[25] vdd gnd cell_6t
Xbit_r26_c69 bl[69] br[69] wl[26] vdd gnd cell_6t
Xbit_r27_c69 bl[69] br[69] wl[27] vdd gnd cell_6t
Xbit_r28_c69 bl[69] br[69] wl[28] vdd gnd cell_6t
Xbit_r29_c69 bl[69] br[69] wl[29] vdd gnd cell_6t
Xbit_r30_c69 bl[69] br[69] wl[30] vdd gnd cell_6t
Xbit_r31_c69 bl[69] br[69] wl[31] vdd gnd cell_6t
Xbit_r32_c69 bl[69] br[69] wl[32] vdd gnd cell_6t
Xbit_r33_c69 bl[69] br[69] wl[33] vdd gnd cell_6t
Xbit_r34_c69 bl[69] br[69] wl[34] vdd gnd cell_6t
Xbit_r35_c69 bl[69] br[69] wl[35] vdd gnd cell_6t
Xbit_r36_c69 bl[69] br[69] wl[36] vdd gnd cell_6t
Xbit_r37_c69 bl[69] br[69] wl[37] vdd gnd cell_6t
Xbit_r38_c69 bl[69] br[69] wl[38] vdd gnd cell_6t
Xbit_r39_c69 bl[69] br[69] wl[39] vdd gnd cell_6t
Xbit_r40_c69 bl[69] br[69] wl[40] vdd gnd cell_6t
Xbit_r41_c69 bl[69] br[69] wl[41] vdd gnd cell_6t
Xbit_r42_c69 bl[69] br[69] wl[42] vdd gnd cell_6t
Xbit_r43_c69 bl[69] br[69] wl[43] vdd gnd cell_6t
Xbit_r44_c69 bl[69] br[69] wl[44] vdd gnd cell_6t
Xbit_r45_c69 bl[69] br[69] wl[45] vdd gnd cell_6t
Xbit_r46_c69 bl[69] br[69] wl[46] vdd gnd cell_6t
Xbit_r47_c69 bl[69] br[69] wl[47] vdd gnd cell_6t
Xbit_r48_c69 bl[69] br[69] wl[48] vdd gnd cell_6t
Xbit_r49_c69 bl[69] br[69] wl[49] vdd gnd cell_6t
Xbit_r50_c69 bl[69] br[69] wl[50] vdd gnd cell_6t
Xbit_r51_c69 bl[69] br[69] wl[51] vdd gnd cell_6t
Xbit_r52_c69 bl[69] br[69] wl[52] vdd gnd cell_6t
Xbit_r53_c69 bl[69] br[69] wl[53] vdd gnd cell_6t
Xbit_r54_c69 bl[69] br[69] wl[54] vdd gnd cell_6t
Xbit_r55_c69 bl[69] br[69] wl[55] vdd gnd cell_6t
Xbit_r56_c69 bl[69] br[69] wl[56] vdd gnd cell_6t
Xbit_r57_c69 bl[69] br[69] wl[57] vdd gnd cell_6t
Xbit_r58_c69 bl[69] br[69] wl[58] vdd gnd cell_6t
Xbit_r59_c69 bl[69] br[69] wl[59] vdd gnd cell_6t
Xbit_r60_c69 bl[69] br[69] wl[60] vdd gnd cell_6t
Xbit_r61_c69 bl[69] br[69] wl[61] vdd gnd cell_6t
Xbit_r62_c69 bl[69] br[69] wl[62] vdd gnd cell_6t
Xbit_r63_c69 bl[69] br[69] wl[63] vdd gnd cell_6t
Xbit_r64_c69 bl[69] br[69] wl[64] vdd gnd cell_6t
Xbit_r65_c69 bl[69] br[69] wl[65] vdd gnd cell_6t
Xbit_r66_c69 bl[69] br[69] wl[66] vdd gnd cell_6t
Xbit_r67_c69 bl[69] br[69] wl[67] vdd gnd cell_6t
Xbit_r68_c69 bl[69] br[69] wl[68] vdd gnd cell_6t
Xbit_r69_c69 bl[69] br[69] wl[69] vdd gnd cell_6t
Xbit_r70_c69 bl[69] br[69] wl[70] vdd gnd cell_6t
Xbit_r71_c69 bl[69] br[69] wl[71] vdd gnd cell_6t
Xbit_r72_c69 bl[69] br[69] wl[72] vdd gnd cell_6t
Xbit_r73_c69 bl[69] br[69] wl[73] vdd gnd cell_6t
Xbit_r74_c69 bl[69] br[69] wl[74] vdd gnd cell_6t
Xbit_r75_c69 bl[69] br[69] wl[75] vdd gnd cell_6t
Xbit_r76_c69 bl[69] br[69] wl[76] vdd gnd cell_6t
Xbit_r77_c69 bl[69] br[69] wl[77] vdd gnd cell_6t
Xbit_r78_c69 bl[69] br[69] wl[78] vdd gnd cell_6t
Xbit_r79_c69 bl[69] br[69] wl[79] vdd gnd cell_6t
Xbit_r80_c69 bl[69] br[69] wl[80] vdd gnd cell_6t
Xbit_r81_c69 bl[69] br[69] wl[81] vdd gnd cell_6t
Xbit_r82_c69 bl[69] br[69] wl[82] vdd gnd cell_6t
Xbit_r83_c69 bl[69] br[69] wl[83] vdd gnd cell_6t
Xbit_r84_c69 bl[69] br[69] wl[84] vdd gnd cell_6t
Xbit_r85_c69 bl[69] br[69] wl[85] vdd gnd cell_6t
Xbit_r86_c69 bl[69] br[69] wl[86] vdd gnd cell_6t
Xbit_r87_c69 bl[69] br[69] wl[87] vdd gnd cell_6t
Xbit_r88_c69 bl[69] br[69] wl[88] vdd gnd cell_6t
Xbit_r89_c69 bl[69] br[69] wl[89] vdd gnd cell_6t
Xbit_r90_c69 bl[69] br[69] wl[90] vdd gnd cell_6t
Xbit_r91_c69 bl[69] br[69] wl[91] vdd gnd cell_6t
Xbit_r92_c69 bl[69] br[69] wl[92] vdd gnd cell_6t
Xbit_r93_c69 bl[69] br[69] wl[93] vdd gnd cell_6t
Xbit_r94_c69 bl[69] br[69] wl[94] vdd gnd cell_6t
Xbit_r95_c69 bl[69] br[69] wl[95] vdd gnd cell_6t
Xbit_r96_c69 bl[69] br[69] wl[96] vdd gnd cell_6t
Xbit_r97_c69 bl[69] br[69] wl[97] vdd gnd cell_6t
Xbit_r98_c69 bl[69] br[69] wl[98] vdd gnd cell_6t
Xbit_r99_c69 bl[69] br[69] wl[99] vdd gnd cell_6t
Xbit_r100_c69 bl[69] br[69] wl[100] vdd gnd cell_6t
Xbit_r101_c69 bl[69] br[69] wl[101] vdd gnd cell_6t
Xbit_r102_c69 bl[69] br[69] wl[102] vdd gnd cell_6t
Xbit_r103_c69 bl[69] br[69] wl[103] vdd gnd cell_6t
Xbit_r104_c69 bl[69] br[69] wl[104] vdd gnd cell_6t
Xbit_r105_c69 bl[69] br[69] wl[105] vdd gnd cell_6t
Xbit_r106_c69 bl[69] br[69] wl[106] vdd gnd cell_6t
Xbit_r107_c69 bl[69] br[69] wl[107] vdd gnd cell_6t
Xbit_r108_c69 bl[69] br[69] wl[108] vdd gnd cell_6t
Xbit_r109_c69 bl[69] br[69] wl[109] vdd gnd cell_6t
Xbit_r110_c69 bl[69] br[69] wl[110] vdd gnd cell_6t
Xbit_r111_c69 bl[69] br[69] wl[111] vdd gnd cell_6t
Xbit_r112_c69 bl[69] br[69] wl[112] vdd gnd cell_6t
Xbit_r113_c69 bl[69] br[69] wl[113] vdd gnd cell_6t
Xbit_r114_c69 bl[69] br[69] wl[114] vdd gnd cell_6t
Xbit_r115_c69 bl[69] br[69] wl[115] vdd gnd cell_6t
Xbit_r116_c69 bl[69] br[69] wl[116] vdd gnd cell_6t
Xbit_r117_c69 bl[69] br[69] wl[117] vdd gnd cell_6t
Xbit_r118_c69 bl[69] br[69] wl[118] vdd gnd cell_6t
Xbit_r119_c69 bl[69] br[69] wl[119] vdd gnd cell_6t
Xbit_r120_c69 bl[69] br[69] wl[120] vdd gnd cell_6t
Xbit_r121_c69 bl[69] br[69] wl[121] vdd gnd cell_6t
Xbit_r122_c69 bl[69] br[69] wl[122] vdd gnd cell_6t
Xbit_r123_c69 bl[69] br[69] wl[123] vdd gnd cell_6t
Xbit_r124_c69 bl[69] br[69] wl[124] vdd gnd cell_6t
Xbit_r125_c69 bl[69] br[69] wl[125] vdd gnd cell_6t
Xbit_r126_c69 bl[69] br[69] wl[126] vdd gnd cell_6t
Xbit_r127_c69 bl[69] br[69] wl[127] vdd gnd cell_6t
Xbit_r128_c69 bl[69] br[69] wl[128] vdd gnd cell_6t
Xbit_r129_c69 bl[69] br[69] wl[129] vdd gnd cell_6t
Xbit_r130_c69 bl[69] br[69] wl[130] vdd gnd cell_6t
Xbit_r131_c69 bl[69] br[69] wl[131] vdd gnd cell_6t
Xbit_r132_c69 bl[69] br[69] wl[132] vdd gnd cell_6t
Xbit_r133_c69 bl[69] br[69] wl[133] vdd gnd cell_6t
Xbit_r134_c69 bl[69] br[69] wl[134] vdd gnd cell_6t
Xbit_r135_c69 bl[69] br[69] wl[135] vdd gnd cell_6t
Xbit_r136_c69 bl[69] br[69] wl[136] vdd gnd cell_6t
Xbit_r137_c69 bl[69] br[69] wl[137] vdd gnd cell_6t
Xbit_r138_c69 bl[69] br[69] wl[138] vdd gnd cell_6t
Xbit_r139_c69 bl[69] br[69] wl[139] vdd gnd cell_6t
Xbit_r140_c69 bl[69] br[69] wl[140] vdd gnd cell_6t
Xbit_r141_c69 bl[69] br[69] wl[141] vdd gnd cell_6t
Xbit_r142_c69 bl[69] br[69] wl[142] vdd gnd cell_6t
Xbit_r143_c69 bl[69] br[69] wl[143] vdd gnd cell_6t
Xbit_r144_c69 bl[69] br[69] wl[144] vdd gnd cell_6t
Xbit_r145_c69 bl[69] br[69] wl[145] vdd gnd cell_6t
Xbit_r146_c69 bl[69] br[69] wl[146] vdd gnd cell_6t
Xbit_r147_c69 bl[69] br[69] wl[147] vdd gnd cell_6t
Xbit_r148_c69 bl[69] br[69] wl[148] vdd gnd cell_6t
Xbit_r149_c69 bl[69] br[69] wl[149] vdd gnd cell_6t
Xbit_r150_c69 bl[69] br[69] wl[150] vdd gnd cell_6t
Xbit_r151_c69 bl[69] br[69] wl[151] vdd gnd cell_6t
Xbit_r152_c69 bl[69] br[69] wl[152] vdd gnd cell_6t
Xbit_r153_c69 bl[69] br[69] wl[153] vdd gnd cell_6t
Xbit_r154_c69 bl[69] br[69] wl[154] vdd gnd cell_6t
Xbit_r155_c69 bl[69] br[69] wl[155] vdd gnd cell_6t
Xbit_r156_c69 bl[69] br[69] wl[156] vdd gnd cell_6t
Xbit_r157_c69 bl[69] br[69] wl[157] vdd gnd cell_6t
Xbit_r158_c69 bl[69] br[69] wl[158] vdd gnd cell_6t
Xbit_r159_c69 bl[69] br[69] wl[159] vdd gnd cell_6t
Xbit_r160_c69 bl[69] br[69] wl[160] vdd gnd cell_6t
Xbit_r161_c69 bl[69] br[69] wl[161] vdd gnd cell_6t
Xbit_r162_c69 bl[69] br[69] wl[162] vdd gnd cell_6t
Xbit_r163_c69 bl[69] br[69] wl[163] vdd gnd cell_6t
Xbit_r164_c69 bl[69] br[69] wl[164] vdd gnd cell_6t
Xbit_r165_c69 bl[69] br[69] wl[165] vdd gnd cell_6t
Xbit_r166_c69 bl[69] br[69] wl[166] vdd gnd cell_6t
Xbit_r167_c69 bl[69] br[69] wl[167] vdd gnd cell_6t
Xbit_r168_c69 bl[69] br[69] wl[168] vdd gnd cell_6t
Xbit_r169_c69 bl[69] br[69] wl[169] vdd gnd cell_6t
Xbit_r170_c69 bl[69] br[69] wl[170] vdd gnd cell_6t
Xbit_r171_c69 bl[69] br[69] wl[171] vdd gnd cell_6t
Xbit_r172_c69 bl[69] br[69] wl[172] vdd gnd cell_6t
Xbit_r173_c69 bl[69] br[69] wl[173] vdd gnd cell_6t
Xbit_r174_c69 bl[69] br[69] wl[174] vdd gnd cell_6t
Xbit_r175_c69 bl[69] br[69] wl[175] vdd gnd cell_6t
Xbit_r176_c69 bl[69] br[69] wl[176] vdd gnd cell_6t
Xbit_r177_c69 bl[69] br[69] wl[177] vdd gnd cell_6t
Xbit_r178_c69 bl[69] br[69] wl[178] vdd gnd cell_6t
Xbit_r179_c69 bl[69] br[69] wl[179] vdd gnd cell_6t
Xbit_r180_c69 bl[69] br[69] wl[180] vdd gnd cell_6t
Xbit_r181_c69 bl[69] br[69] wl[181] vdd gnd cell_6t
Xbit_r182_c69 bl[69] br[69] wl[182] vdd gnd cell_6t
Xbit_r183_c69 bl[69] br[69] wl[183] vdd gnd cell_6t
Xbit_r184_c69 bl[69] br[69] wl[184] vdd gnd cell_6t
Xbit_r185_c69 bl[69] br[69] wl[185] vdd gnd cell_6t
Xbit_r186_c69 bl[69] br[69] wl[186] vdd gnd cell_6t
Xbit_r187_c69 bl[69] br[69] wl[187] vdd gnd cell_6t
Xbit_r188_c69 bl[69] br[69] wl[188] vdd gnd cell_6t
Xbit_r189_c69 bl[69] br[69] wl[189] vdd gnd cell_6t
Xbit_r190_c69 bl[69] br[69] wl[190] vdd gnd cell_6t
Xbit_r191_c69 bl[69] br[69] wl[191] vdd gnd cell_6t
Xbit_r192_c69 bl[69] br[69] wl[192] vdd gnd cell_6t
Xbit_r193_c69 bl[69] br[69] wl[193] vdd gnd cell_6t
Xbit_r194_c69 bl[69] br[69] wl[194] vdd gnd cell_6t
Xbit_r195_c69 bl[69] br[69] wl[195] vdd gnd cell_6t
Xbit_r196_c69 bl[69] br[69] wl[196] vdd gnd cell_6t
Xbit_r197_c69 bl[69] br[69] wl[197] vdd gnd cell_6t
Xbit_r198_c69 bl[69] br[69] wl[198] vdd gnd cell_6t
Xbit_r199_c69 bl[69] br[69] wl[199] vdd gnd cell_6t
Xbit_r200_c69 bl[69] br[69] wl[200] vdd gnd cell_6t
Xbit_r201_c69 bl[69] br[69] wl[201] vdd gnd cell_6t
Xbit_r202_c69 bl[69] br[69] wl[202] vdd gnd cell_6t
Xbit_r203_c69 bl[69] br[69] wl[203] vdd gnd cell_6t
Xbit_r204_c69 bl[69] br[69] wl[204] vdd gnd cell_6t
Xbit_r205_c69 bl[69] br[69] wl[205] vdd gnd cell_6t
Xbit_r206_c69 bl[69] br[69] wl[206] vdd gnd cell_6t
Xbit_r207_c69 bl[69] br[69] wl[207] vdd gnd cell_6t
Xbit_r208_c69 bl[69] br[69] wl[208] vdd gnd cell_6t
Xbit_r209_c69 bl[69] br[69] wl[209] vdd gnd cell_6t
Xbit_r210_c69 bl[69] br[69] wl[210] vdd gnd cell_6t
Xbit_r211_c69 bl[69] br[69] wl[211] vdd gnd cell_6t
Xbit_r212_c69 bl[69] br[69] wl[212] vdd gnd cell_6t
Xbit_r213_c69 bl[69] br[69] wl[213] vdd gnd cell_6t
Xbit_r214_c69 bl[69] br[69] wl[214] vdd gnd cell_6t
Xbit_r215_c69 bl[69] br[69] wl[215] vdd gnd cell_6t
Xbit_r216_c69 bl[69] br[69] wl[216] vdd gnd cell_6t
Xbit_r217_c69 bl[69] br[69] wl[217] vdd gnd cell_6t
Xbit_r218_c69 bl[69] br[69] wl[218] vdd gnd cell_6t
Xbit_r219_c69 bl[69] br[69] wl[219] vdd gnd cell_6t
Xbit_r220_c69 bl[69] br[69] wl[220] vdd gnd cell_6t
Xbit_r221_c69 bl[69] br[69] wl[221] vdd gnd cell_6t
Xbit_r222_c69 bl[69] br[69] wl[222] vdd gnd cell_6t
Xbit_r223_c69 bl[69] br[69] wl[223] vdd gnd cell_6t
Xbit_r224_c69 bl[69] br[69] wl[224] vdd gnd cell_6t
Xbit_r225_c69 bl[69] br[69] wl[225] vdd gnd cell_6t
Xbit_r226_c69 bl[69] br[69] wl[226] vdd gnd cell_6t
Xbit_r227_c69 bl[69] br[69] wl[227] vdd gnd cell_6t
Xbit_r228_c69 bl[69] br[69] wl[228] vdd gnd cell_6t
Xbit_r229_c69 bl[69] br[69] wl[229] vdd gnd cell_6t
Xbit_r230_c69 bl[69] br[69] wl[230] vdd gnd cell_6t
Xbit_r231_c69 bl[69] br[69] wl[231] vdd gnd cell_6t
Xbit_r232_c69 bl[69] br[69] wl[232] vdd gnd cell_6t
Xbit_r233_c69 bl[69] br[69] wl[233] vdd gnd cell_6t
Xbit_r234_c69 bl[69] br[69] wl[234] vdd gnd cell_6t
Xbit_r235_c69 bl[69] br[69] wl[235] vdd gnd cell_6t
Xbit_r236_c69 bl[69] br[69] wl[236] vdd gnd cell_6t
Xbit_r237_c69 bl[69] br[69] wl[237] vdd gnd cell_6t
Xbit_r238_c69 bl[69] br[69] wl[238] vdd gnd cell_6t
Xbit_r239_c69 bl[69] br[69] wl[239] vdd gnd cell_6t
Xbit_r240_c69 bl[69] br[69] wl[240] vdd gnd cell_6t
Xbit_r241_c69 bl[69] br[69] wl[241] vdd gnd cell_6t
Xbit_r242_c69 bl[69] br[69] wl[242] vdd gnd cell_6t
Xbit_r243_c69 bl[69] br[69] wl[243] vdd gnd cell_6t
Xbit_r244_c69 bl[69] br[69] wl[244] vdd gnd cell_6t
Xbit_r245_c69 bl[69] br[69] wl[245] vdd gnd cell_6t
Xbit_r246_c69 bl[69] br[69] wl[246] vdd gnd cell_6t
Xbit_r247_c69 bl[69] br[69] wl[247] vdd gnd cell_6t
Xbit_r248_c69 bl[69] br[69] wl[248] vdd gnd cell_6t
Xbit_r249_c69 bl[69] br[69] wl[249] vdd gnd cell_6t
Xbit_r250_c69 bl[69] br[69] wl[250] vdd gnd cell_6t
Xbit_r251_c69 bl[69] br[69] wl[251] vdd gnd cell_6t
Xbit_r252_c69 bl[69] br[69] wl[252] vdd gnd cell_6t
Xbit_r253_c69 bl[69] br[69] wl[253] vdd gnd cell_6t
Xbit_r254_c69 bl[69] br[69] wl[254] vdd gnd cell_6t
Xbit_r255_c69 bl[69] br[69] wl[255] vdd gnd cell_6t
Xbit_r0_c70 bl[70] br[70] wl[0] vdd gnd cell_6t
Xbit_r1_c70 bl[70] br[70] wl[1] vdd gnd cell_6t
Xbit_r2_c70 bl[70] br[70] wl[2] vdd gnd cell_6t
Xbit_r3_c70 bl[70] br[70] wl[3] vdd gnd cell_6t
Xbit_r4_c70 bl[70] br[70] wl[4] vdd gnd cell_6t
Xbit_r5_c70 bl[70] br[70] wl[5] vdd gnd cell_6t
Xbit_r6_c70 bl[70] br[70] wl[6] vdd gnd cell_6t
Xbit_r7_c70 bl[70] br[70] wl[7] vdd gnd cell_6t
Xbit_r8_c70 bl[70] br[70] wl[8] vdd gnd cell_6t
Xbit_r9_c70 bl[70] br[70] wl[9] vdd gnd cell_6t
Xbit_r10_c70 bl[70] br[70] wl[10] vdd gnd cell_6t
Xbit_r11_c70 bl[70] br[70] wl[11] vdd gnd cell_6t
Xbit_r12_c70 bl[70] br[70] wl[12] vdd gnd cell_6t
Xbit_r13_c70 bl[70] br[70] wl[13] vdd gnd cell_6t
Xbit_r14_c70 bl[70] br[70] wl[14] vdd gnd cell_6t
Xbit_r15_c70 bl[70] br[70] wl[15] vdd gnd cell_6t
Xbit_r16_c70 bl[70] br[70] wl[16] vdd gnd cell_6t
Xbit_r17_c70 bl[70] br[70] wl[17] vdd gnd cell_6t
Xbit_r18_c70 bl[70] br[70] wl[18] vdd gnd cell_6t
Xbit_r19_c70 bl[70] br[70] wl[19] vdd gnd cell_6t
Xbit_r20_c70 bl[70] br[70] wl[20] vdd gnd cell_6t
Xbit_r21_c70 bl[70] br[70] wl[21] vdd gnd cell_6t
Xbit_r22_c70 bl[70] br[70] wl[22] vdd gnd cell_6t
Xbit_r23_c70 bl[70] br[70] wl[23] vdd gnd cell_6t
Xbit_r24_c70 bl[70] br[70] wl[24] vdd gnd cell_6t
Xbit_r25_c70 bl[70] br[70] wl[25] vdd gnd cell_6t
Xbit_r26_c70 bl[70] br[70] wl[26] vdd gnd cell_6t
Xbit_r27_c70 bl[70] br[70] wl[27] vdd gnd cell_6t
Xbit_r28_c70 bl[70] br[70] wl[28] vdd gnd cell_6t
Xbit_r29_c70 bl[70] br[70] wl[29] vdd gnd cell_6t
Xbit_r30_c70 bl[70] br[70] wl[30] vdd gnd cell_6t
Xbit_r31_c70 bl[70] br[70] wl[31] vdd gnd cell_6t
Xbit_r32_c70 bl[70] br[70] wl[32] vdd gnd cell_6t
Xbit_r33_c70 bl[70] br[70] wl[33] vdd gnd cell_6t
Xbit_r34_c70 bl[70] br[70] wl[34] vdd gnd cell_6t
Xbit_r35_c70 bl[70] br[70] wl[35] vdd gnd cell_6t
Xbit_r36_c70 bl[70] br[70] wl[36] vdd gnd cell_6t
Xbit_r37_c70 bl[70] br[70] wl[37] vdd gnd cell_6t
Xbit_r38_c70 bl[70] br[70] wl[38] vdd gnd cell_6t
Xbit_r39_c70 bl[70] br[70] wl[39] vdd gnd cell_6t
Xbit_r40_c70 bl[70] br[70] wl[40] vdd gnd cell_6t
Xbit_r41_c70 bl[70] br[70] wl[41] vdd gnd cell_6t
Xbit_r42_c70 bl[70] br[70] wl[42] vdd gnd cell_6t
Xbit_r43_c70 bl[70] br[70] wl[43] vdd gnd cell_6t
Xbit_r44_c70 bl[70] br[70] wl[44] vdd gnd cell_6t
Xbit_r45_c70 bl[70] br[70] wl[45] vdd gnd cell_6t
Xbit_r46_c70 bl[70] br[70] wl[46] vdd gnd cell_6t
Xbit_r47_c70 bl[70] br[70] wl[47] vdd gnd cell_6t
Xbit_r48_c70 bl[70] br[70] wl[48] vdd gnd cell_6t
Xbit_r49_c70 bl[70] br[70] wl[49] vdd gnd cell_6t
Xbit_r50_c70 bl[70] br[70] wl[50] vdd gnd cell_6t
Xbit_r51_c70 bl[70] br[70] wl[51] vdd gnd cell_6t
Xbit_r52_c70 bl[70] br[70] wl[52] vdd gnd cell_6t
Xbit_r53_c70 bl[70] br[70] wl[53] vdd gnd cell_6t
Xbit_r54_c70 bl[70] br[70] wl[54] vdd gnd cell_6t
Xbit_r55_c70 bl[70] br[70] wl[55] vdd gnd cell_6t
Xbit_r56_c70 bl[70] br[70] wl[56] vdd gnd cell_6t
Xbit_r57_c70 bl[70] br[70] wl[57] vdd gnd cell_6t
Xbit_r58_c70 bl[70] br[70] wl[58] vdd gnd cell_6t
Xbit_r59_c70 bl[70] br[70] wl[59] vdd gnd cell_6t
Xbit_r60_c70 bl[70] br[70] wl[60] vdd gnd cell_6t
Xbit_r61_c70 bl[70] br[70] wl[61] vdd gnd cell_6t
Xbit_r62_c70 bl[70] br[70] wl[62] vdd gnd cell_6t
Xbit_r63_c70 bl[70] br[70] wl[63] vdd gnd cell_6t
Xbit_r64_c70 bl[70] br[70] wl[64] vdd gnd cell_6t
Xbit_r65_c70 bl[70] br[70] wl[65] vdd gnd cell_6t
Xbit_r66_c70 bl[70] br[70] wl[66] vdd gnd cell_6t
Xbit_r67_c70 bl[70] br[70] wl[67] vdd gnd cell_6t
Xbit_r68_c70 bl[70] br[70] wl[68] vdd gnd cell_6t
Xbit_r69_c70 bl[70] br[70] wl[69] vdd gnd cell_6t
Xbit_r70_c70 bl[70] br[70] wl[70] vdd gnd cell_6t
Xbit_r71_c70 bl[70] br[70] wl[71] vdd gnd cell_6t
Xbit_r72_c70 bl[70] br[70] wl[72] vdd gnd cell_6t
Xbit_r73_c70 bl[70] br[70] wl[73] vdd gnd cell_6t
Xbit_r74_c70 bl[70] br[70] wl[74] vdd gnd cell_6t
Xbit_r75_c70 bl[70] br[70] wl[75] vdd gnd cell_6t
Xbit_r76_c70 bl[70] br[70] wl[76] vdd gnd cell_6t
Xbit_r77_c70 bl[70] br[70] wl[77] vdd gnd cell_6t
Xbit_r78_c70 bl[70] br[70] wl[78] vdd gnd cell_6t
Xbit_r79_c70 bl[70] br[70] wl[79] vdd gnd cell_6t
Xbit_r80_c70 bl[70] br[70] wl[80] vdd gnd cell_6t
Xbit_r81_c70 bl[70] br[70] wl[81] vdd gnd cell_6t
Xbit_r82_c70 bl[70] br[70] wl[82] vdd gnd cell_6t
Xbit_r83_c70 bl[70] br[70] wl[83] vdd gnd cell_6t
Xbit_r84_c70 bl[70] br[70] wl[84] vdd gnd cell_6t
Xbit_r85_c70 bl[70] br[70] wl[85] vdd gnd cell_6t
Xbit_r86_c70 bl[70] br[70] wl[86] vdd gnd cell_6t
Xbit_r87_c70 bl[70] br[70] wl[87] vdd gnd cell_6t
Xbit_r88_c70 bl[70] br[70] wl[88] vdd gnd cell_6t
Xbit_r89_c70 bl[70] br[70] wl[89] vdd gnd cell_6t
Xbit_r90_c70 bl[70] br[70] wl[90] vdd gnd cell_6t
Xbit_r91_c70 bl[70] br[70] wl[91] vdd gnd cell_6t
Xbit_r92_c70 bl[70] br[70] wl[92] vdd gnd cell_6t
Xbit_r93_c70 bl[70] br[70] wl[93] vdd gnd cell_6t
Xbit_r94_c70 bl[70] br[70] wl[94] vdd gnd cell_6t
Xbit_r95_c70 bl[70] br[70] wl[95] vdd gnd cell_6t
Xbit_r96_c70 bl[70] br[70] wl[96] vdd gnd cell_6t
Xbit_r97_c70 bl[70] br[70] wl[97] vdd gnd cell_6t
Xbit_r98_c70 bl[70] br[70] wl[98] vdd gnd cell_6t
Xbit_r99_c70 bl[70] br[70] wl[99] vdd gnd cell_6t
Xbit_r100_c70 bl[70] br[70] wl[100] vdd gnd cell_6t
Xbit_r101_c70 bl[70] br[70] wl[101] vdd gnd cell_6t
Xbit_r102_c70 bl[70] br[70] wl[102] vdd gnd cell_6t
Xbit_r103_c70 bl[70] br[70] wl[103] vdd gnd cell_6t
Xbit_r104_c70 bl[70] br[70] wl[104] vdd gnd cell_6t
Xbit_r105_c70 bl[70] br[70] wl[105] vdd gnd cell_6t
Xbit_r106_c70 bl[70] br[70] wl[106] vdd gnd cell_6t
Xbit_r107_c70 bl[70] br[70] wl[107] vdd gnd cell_6t
Xbit_r108_c70 bl[70] br[70] wl[108] vdd gnd cell_6t
Xbit_r109_c70 bl[70] br[70] wl[109] vdd gnd cell_6t
Xbit_r110_c70 bl[70] br[70] wl[110] vdd gnd cell_6t
Xbit_r111_c70 bl[70] br[70] wl[111] vdd gnd cell_6t
Xbit_r112_c70 bl[70] br[70] wl[112] vdd gnd cell_6t
Xbit_r113_c70 bl[70] br[70] wl[113] vdd gnd cell_6t
Xbit_r114_c70 bl[70] br[70] wl[114] vdd gnd cell_6t
Xbit_r115_c70 bl[70] br[70] wl[115] vdd gnd cell_6t
Xbit_r116_c70 bl[70] br[70] wl[116] vdd gnd cell_6t
Xbit_r117_c70 bl[70] br[70] wl[117] vdd gnd cell_6t
Xbit_r118_c70 bl[70] br[70] wl[118] vdd gnd cell_6t
Xbit_r119_c70 bl[70] br[70] wl[119] vdd gnd cell_6t
Xbit_r120_c70 bl[70] br[70] wl[120] vdd gnd cell_6t
Xbit_r121_c70 bl[70] br[70] wl[121] vdd gnd cell_6t
Xbit_r122_c70 bl[70] br[70] wl[122] vdd gnd cell_6t
Xbit_r123_c70 bl[70] br[70] wl[123] vdd gnd cell_6t
Xbit_r124_c70 bl[70] br[70] wl[124] vdd gnd cell_6t
Xbit_r125_c70 bl[70] br[70] wl[125] vdd gnd cell_6t
Xbit_r126_c70 bl[70] br[70] wl[126] vdd gnd cell_6t
Xbit_r127_c70 bl[70] br[70] wl[127] vdd gnd cell_6t
Xbit_r128_c70 bl[70] br[70] wl[128] vdd gnd cell_6t
Xbit_r129_c70 bl[70] br[70] wl[129] vdd gnd cell_6t
Xbit_r130_c70 bl[70] br[70] wl[130] vdd gnd cell_6t
Xbit_r131_c70 bl[70] br[70] wl[131] vdd gnd cell_6t
Xbit_r132_c70 bl[70] br[70] wl[132] vdd gnd cell_6t
Xbit_r133_c70 bl[70] br[70] wl[133] vdd gnd cell_6t
Xbit_r134_c70 bl[70] br[70] wl[134] vdd gnd cell_6t
Xbit_r135_c70 bl[70] br[70] wl[135] vdd gnd cell_6t
Xbit_r136_c70 bl[70] br[70] wl[136] vdd gnd cell_6t
Xbit_r137_c70 bl[70] br[70] wl[137] vdd gnd cell_6t
Xbit_r138_c70 bl[70] br[70] wl[138] vdd gnd cell_6t
Xbit_r139_c70 bl[70] br[70] wl[139] vdd gnd cell_6t
Xbit_r140_c70 bl[70] br[70] wl[140] vdd gnd cell_6t
Xbit_r141_c70 bl[70] br[70] wl[141] vdd gnd cell_6t
Xbit_r142_c70 bl[70] br[70] wl[142] vdd gnd cell_6t
Xbit_r143_c70 bl[70] br[70] wl[143] vdd gnd cell_6t
Xbit_r144_c70 bl[70] br[70] wl[144] vdd gnd cell_6t
Xbit_r145_c70 bl[70] br[70] wl[145] vdd gnd cell_6t
Xbit_r146_c70 bl[70] br[70] wl[146] vdd gnd cell_6t
Xbit_r147_c70 bl[70] br[70] wl[147] vdd gnd cell_6t
Xbit_r148_c70 bl[70] br[70] wl[148] vdd gnd cell_6t
Xbit_r149_c70 bl[70] br[70] wl[149] vdd gnd cell_6t
Xbit_r150_c70 bl[70] br[70] wl[150] vdd gnd cell_6t
Xbit_r151_c70 bl[70] br[70] wl[151] vdd gnd cell_6t
Xbit_r152_c70 bl[70] br[70] wl[152] vdd gnd cell_6t
Xbit_r153_c70 bl[70] br[70] wl[153] vdd gnd cell_6t
Xbit_r154_c70 bl[70] br[70] wl[154] vdd gnd cell_6t
Xbit_r155_c70 bl[70] br[70] wl[155] vdd gnd cell_6t
Xbit_r156_c70 bl[70] br[70] wl[156] vdd gnd cell_6t
Xbit_r157_c70 bl[70] br[70] wl[157] vdd gnd cell_6t
Xbit_r158_c70 bl[70] br[70] wl[158] vdd gnd cell_6t
Xbit_r159_c70 bl[70] br[70] wl[159] vdd gnd cell_6t
Xbit_r160_c70 bl[70] br[70] wl[160] vdd gnd cell_6t
Xbit_r161_c70 bl[70] br[70] wl[161] vdd gnd cell_6t
Xbit_r162_c70 bl[70] br[70] wl[162] vdd gnd cell_6t
Xbit_r163_c70 bl[70] br[70] wl[163] vdd gnd cell_6t
Xbit_r164_c70 bl[70] br[70] wl[164] vdd gnd cell_6t
Xbit_r165_c70 bl[70] br[70] wl[165] vdd gnd cell_6t
Xbit_r166_c70 bl[70] br[70] wl[166] vdd gnd cell_6t
Xbit_r167_c70 bl[70] br[70] wl[167] vdd gnd cell_6t
Xbit_r168_c70 bl[70] br[70] wl[168] vdd gnd cell_6t
Xbit_r169_c70 bl[70] br[70] wl[169] vdd gnd cell_6t
Xbit_r170_c70 bl[70] br[70] wl[170] vdd gnd cell_6t
Xbit_r171_c70 bl[70] br[70] wl[171] vdd gnd cell_6t
Xbit_r172_c70 bl[70] br[70] wl[172] vdd gnd cell_6t
Xbit_r173_c70 bl[70] br[70] wl[173] vdd gnd cell_6t
Xbit_r174_c70 bl[70] br[70] wl[174] vdd gnd cell_6t
Xbit_r175_c70 bl[70] br[70] wl[175] vdd gnd cell_6t
Xbit_r176_c70 bl[70] br[70] wl[176] vdd gnd cell_6t
Xbit_r177_c70 bl[70] br[70] wl[177] vdd gnd cell_6t
Xbit_r178_c70 bl[70] br[70] wl[178] vdd gnd cell_6t
Xbit_r179_c70 bl[70] br[70] wl[179] vdd gnd cell_6t
Xbit_r180_c70 bl[70] br[70] wl[180] vdd gnd cell_6t
Xbit_r181_c70 bl[70] br[70] wl[181] vdd gnd cell_6t
Xbit_r182_c70 bl[70] br[70] wl[182] vdd gnd cell_6t
Xbit_r183_c70 bl[70] br[70] wl[183] vdd gnd cell_6t
Xbit_r184_c70 bl[70] br[70] wl[184] vdd gnd cell_6t
Xbit_r185_c70 bl[70] br[70] wl[185] vdd gnd cell_6t
Xbit_r186_c70 bl[70] br[70] wl[186] vdd gnd cell_6t
Xbit_r187_c70 bl[70] br[70] wl[187] vdd gnd cell_6t
Xbit_r188_c70 bl[70] br[70] wl[188] vdd gnd cell_6t
Xbit_r189_c70 bl[70] br[70] wl[189] vdd gnd cell_6t
Xbit_r190_c70 bl[70] br[70] wl[190] vdd gnd cell_6t
Xbit_r191_c70 bl[70] br[70] wl[191] vdd gnd cell_6t
Xbit_r192_c70 bl[70] br[70] wl[192] vdd gnd cell_6t
Xbit_r193_c70 bl[70] br[70] wl[193] vdd gnd cell_6t
Xbit_r194_c70 bl[70] br[70] wl[194] vdd gnd cell_6t
Xbit_r195_c70 bl[70] br[70] wl[195] vdd gnd cell_6t
Xbit_r196_c70 bl[70] br[70] wl[196] vdd gnd cell_6t
Xbit_r197_c70 bl[70] br[70] wl[197] vdd gnd cell_6t
Xbit_r198_c70 bl[70] br[70] wl[198] vdd gnd cell_6t
Xbit_r199_c70 bl[70] br[70] wl[199] vdd gnd cell_6t
Xbit_r200_c70 bl[70] br[70] wl[200] vdd gnd cell_6t
Xbit_r201_c70 bl[70] br[70] wl[201] vdd gnd cell_6t
Xbit_r202_c70 bl[70] br[70] wl[202] vdd gnd cell_6t
Xbit_r203_c70 bl[70] br[70] wl[203] vdd gnd cell_6t
Xbit_r204_c70 bl[70] br[70] wl[204] vdd gnd cell_6t
Xbit_r205_c70 bl[70] br[70] wl[205] vdd gnd cell_6t
Xbit_r206_c70 bl[70] br[70] wl[206] vdd gnd cell_6t
Xbit_r207_c70 bl[70] br[70] wl[207] vdd gnd cell_6t
Xbit_r208_c70 bl[70] br[70] wl[208] vdd gnd cell_6t
Xbit_r209_c70 bl[70] br[70] wl[209] vdd gnd cell_6t
Xbit_r210_c70 bl[70] br[70] wl[210] vdd gnd cell_6t
Xbit_r211_c70 bl[70] br[70] wl[211] vdd gnd cell_6t
Xbit_r212_c70 bl[70] br[70] wl[212] vdd gnd cell_6t
Xbit_r213_c70 bl[70] br[70] wl[213] vdd gnd cell_6t
Xbit_r214_c70 bl[70] br[70] wl[214] vdd gnd cell_6t
Xbit_r215_c70 bl[70] br[70] wl[215] vdd gnd cell_6t
Xbit_r216_c70 bl[70] br[70] wl[216] vdd gnd cell_6t
Xbit_r217_c70 bl[70] br[70] wl[217] vdd gnd cell_6t
Xbit_r218_c70 bl[70] br[70] wl[218] vdd gnd cell_6t
Xbit_r219_c70 bl[70] br[70] wl[219] vdd gnd cell_6t
Xbit_r220_c70 bl[70] br[70] wl[220] vdd gnd cell_6t
Xbit_r221_c70 bl[70] br[70] wl[221] vdd gnd cell_6t
Xbit_r222_c70 bl[70] br[70] wl[222] vdd gnd cell_6t
Xbit_r223_c70 bl[70] br[70] wl[223] vdd gnd cell_6t
Xbit_r224_c70 bl[70] br[70] wl[224] vdd gnd cell_6t
Xbit_r225_c70 bl[70] br[70] wl[225] vdd gnd cell_6t
Xbit_r226_c70 bl[70] br[70] wl[226] vdd gnd cell_6t
Xbit_r227_c70 bl[70] br[70] wl[227] vdd gnd cell_6t
Xbit_r228_c70 bl[70] br[70] wl[228] vdd gnd cell_6t
Xbit_r229_c70 bl[70] br[70] wl[229] vdd gnd cell_6t
Xbit_r230_c70 bl[70] br[70] wl[230] vdd gnd cell_6t
Xbit_r231_c70 bl[70] br[70] wl[231] vdd gnd cell_6t
Xbit_r232_c70 bl[70] br[70] wl[232] vdd gnd cell_6t
Xbit_r233_c70 bl[70] br[70] wl[233] vdd gnd cell_6t
Xbit_r234_c70 bl[70] br[70] wl[234] vdd gnd cell_6t
Xbit_r235_c70 bl[70] br[70] wl[235] vdd gnd cell_6t
Xbit_r236_c70 bl[70] br[70] wl[236] vdd gnd cell_6t
Xbit_r237_c70 bl[70] br[70] wl[237] vdd gnd cell_6t
Xbit_r238_c70 bl[70] br[70] wl[238] vdd gnd cell_6t
Xbit_r239_c70 bl[70] br[70] wl[239] vdd gnd cell_6t
Xbit_r240_c70 bl[70] br[70] wl[240] vdd gnd cell_6t
Xbit_r241_c70 bl[70] br[70] wl[241] vdd gnd cell_6t
Xbit_r242_c70 bl[70] br[70] wl[242] vdd gnd cell_6t
Xbit_r243_c70 bl[70] br[70] wl[243] vdd gnd cell_6t
Xbit_r244_c70 bl[70] br[70] wl[244] vdd gnd cell_6t
Xbit_r245_c70 bl[70] br[70] wl[245] vdd gnd cell_6t
Xbit_r246_c70 bl[70] br[70] wl[246] vdd gnd cell_6t
Xbit_r247_c70 bl[70] br[70] wl[247] vdd gnd cell_6t
Xbit_r248_c70 bl[70] br[70] wl[248] vdd gnd cell_6t
Xbit_r249_c70 bl[70] br[70] wl[249] vdd gnd cell_6t
Xbit_r250_c70 bl[70] br[70] wl[250] vdd gnd cell_6t
Xbit_r251_c70 bl[70] br[70] wl[251] vdd gnd cell_6t
Xbit_r252_c70 bl[70] br[70] wl[252] vdd gnd cell_6t
Xbit_r253_c70 bl[70] br[70] wl[253] vdd gnd cell_6t
Xbit_r254_c70 bl[70] br[70] wl[254] vdd gnd cell_6t
Xbit_r255_c70 bl[70] br[70] wl[255] vdd gnd cell_6t
Xbit_r0_c71 bl[71] br[71] wl[0] vdd gnd cell_6t
Xbit_r1_c71 bl[71] br[71] wl[1] vdd gnd cell_6t
Xbit_r2_c71 bl[71] br[71] wl[2] vdd gnd cell_6t
Xbit_r3_c71 bl[71] br[71] wl[3] vdd gnd cell_6t
Xbit_r4_c71 bl[71] br[71] wl[4] vdd gnd cell_6t
Xbit_r5_c71 bl[71] br[71] wl[5] vdd gnd cell_6t
Xbit_r6_c71 bl[71] br[71] wl[6] vdd gnd cell_6t
Xbit_r7_c71 bl[71] br[71] wl[7] vdd gnd cell_6t
Xbit_r8_c71 bl[71] br[71] wl[8] vdd gnd cell_6t
Xbit_r9_c71 bl[71] br[71] wl[9] vdd gnd cell_6t
Xbit_r10_c71 bl[71] br[71] wl[10] vdd gnd cell_6t
Xbit_r11_c71 bl[71] br[71] wl[11] vdd gnd cell_6t
Xbit_r12_c71 bl[71] br[71] wl[12] vdd gnd cell_6t
Xbit_r13_c71 bl[71] br[71] wl[13] vdd gnd cell_6t
Xbit_r14_c71 bl[71] br[71] wl[14] vdd gnd cell_6t
Xbit_r15_c71 bl[71] br[71] wl[15] vdd gnd cell_6t
Xbit_r16_c71 bl[71] br[71] wl[16] vdd gnd cell_6t
Xbit_r17_c71 bl[71] br[71] wl[17] vdd gnd cell_6t
Xbit_r18_c71 bl[71] br[71] wl[18] vdd gnd cell_6t
Xbit_r19_c71 bl[71] br[71] wl[19] vdd gnd cell_6t
Xbit_r20_c71 bl[71] br[71] wl[20] vdd gnd cell_6t
Xbit_r21_c71 bl[71] br[71] wl[21] vdd gnd cell_6t
Xbit_r22_c71 bl[71] br[71] wl[22] vdd gnd cell_6t
Xbit_r23_c71 bl[71] br[71] wl[23] vdd gnd cell_6t
Xbit_r24_c71 bl[71] br[71] wl[24] vdd gnd cell_6t
Xbit_r25_c71 bl[71] br[71] wl[25] vdd gnd cell_6t
Xbit_r26_c71 bl[71] br[71] wl[26] vdd gnd cell_6t
Xbit_r27_c71 bl[71] br[71] wl[27] vdd gnd cell_6t
Xbit_r28_c71 bl[71] br[71] wl[28] vdd gnd cell_6t
Xbit_r29_c71 bl[71] br[71] wl[29] vdd gnd cell_6t
Xbit_r30_c71 bl[71] br[71] wl[30] vdd gnd cell_6t
Xbit_r31_c71 bl[71] br[71] wl[31] vdd gnd cell_6t
Xbit_r32_c71 bl[71] br[71] wl[32] vdd gnd cell_6t
Xbit_r33_c71 bl[71] br[71] wl[33] vdd gnd cell_6t
Xbit_r34_c71 bl[71] br[71] wl[34] vdd gnd cell_6t
Xbit_r35_c71 bl[71] br[71] wl[35] vdd gnd cell_6t
Xbit_r36_c71 bl[71] br[71] wl[36] vdd gnd cell_6t
Xbit_r37_c71 bl[71] br[71] wl[37] vdd gnd cell_6t
Xbit_r38_c71 bl[71] br[71] wl[38] vdd gnd cell_6t
Xbit_r39_c71 bl[71] br[71] wl[39] vdd gnd cell_6t
Xbit_r40_c71 bl[71] br[71] wl[40] vdd gnd cell_6t
Xbit_r41_c71 bl[71] br[71] wl[41] vdd gnd cell_6t
Xbit_r42_c71 bl[71] br[71] wl[42] vdd gnd cell_6t
Xbit_r43_c71 bl[71] br[71] wl[43] vdd gnd cell_6t
Xbit_r44_c71 bl[71] br[71] wl[44] vdd gnd cell_6t
Xbit_r45_c71 bl[71] br[71] wl[45] vdd gnd cell_6t
Xbit_r46_c71 bl[71] br[71] wl[46] vdd gnd cell_6t
Xbit_r47_c71 bl[71] br[71] wl[47] vdd gnd cell_6t
Xbit_r48_c71 bl[71] br[71] wl[48] vdd gnd cell_6t
Xbit_r49_c71 bl[71] br[71] wl[49] vdd gnd cell_6t
Xbit_r50_c71 bl[71] br[71] wl[50] vdd gnd cell_6t
Xbit_r51_c71 bl[71] br[71] wl[51] vdd gnd cell_6t
Xbit_r52_c71 bl[71] br[71] wl[52] vdd gnd cell_6t
Xbit_r53_c71 bl[71] br[71] wl[53] vdd gnd cell_6t
Xbit_r54_c71 bl[71] br[71] wl[54] vdd gnd cell_6t
Xbit_r55_c71 bl[71] br[71] wl[55] vdd gnd cell_6t
Xbit_r56_c71 bl[71] br[71] wl[56] vdd gnd cell_6t
Xbit_r57_c71 bl[71] br[71] wl[57] vdd gnd cell_6t
Xbit_r58_c71 bl[71] br[71] wl[58] vdd gnd cell_6t
Xbit_r59_c71 bl[71] br[71] wl[59] vdd gnd cell_6t
Xbit_r60_c71 bl[71] br[71] wl[60] vdd gnd cell_6t
Xbit_r61_c71 bl[71] br[71] wl[61] vdd gnd cell_6t
Xbit_r62_c71 bl[71] br[71] wl[62] vdd gnd cell_6t
Xbit_r63_c71 bl[71] br[71] wl[63] vdd gnd cell_6t
Xbit_r64_c71 bl[71] br[71] wl[64] vdd gnd cell_6t
Xbit_r65_c71 bl[71] br[71] wl[65] vdd gnd cell_6t
Xbit_r66_c71 bl[71] br[71] wl[66] vdd gnd cell_6t
Xbit_r67_c71 bl[71] br[71] wl[67] vdd gnd cell_6t
Xbit_r68_c71 bl[71] br[71] wl[68] vdd gnd cell_6t
Xbit_r69_c71 bl[71] br[71] wl[69] vdd gnd cell_6t
Xbit_r70_c71 bl[71] br[71] wl[70] vdd gnd cell_6t
Xbit_r71_c71 bl[71] br[71] wl[71] vdd gnd cell_6t
Xbit_r72_c71 bl[71] br[71] wl[72] vdd gnd cell_6t
Xbit_r73_c71 bl[71] br[71] wl[73] vdd gnd cell_6t
Xbit_r74_c71 bl[71] br[71] wl[74] vdd gnd cell_6t
Xbit_r75_c71 bl[71] br[71] wl[75] vdd gnd cell_6t
Xbit_r76_c71 bl[71] br[71] wl[76] vdd gnd cell_6t
Xbit_r77_c71 bl[71] br[71] wl[77] vdd gnd cell_6t
Xbit_r78_c71 bl[71] br[71] wl[78] vdd gnd cell_6t
Xbit_r79_c71 bl[71] br[71] wl[79] vdd gnd cell_6t
Xbit_r80_c71 bl[71] br[71] wl[80] vdd gnd cell_6t
Xbit_r81_c71 bl[71] br[71] wl[81] vdd gnd cell_6t
Xbit_r82_c71 bl[71] br[71] wl[82] vdd gnd cell_6t
Xbit_r83_c71 bl[71] br[71] wl[83] vdd gnd cell_6t
Xbit_r84_c71 bl[71] br[71] wl[84] vdd gnd cell_6t
Xbit_r85_c71 bl[71] br[71] wl[85] vdd gnd cell_6t
Xbit_r86_c71 bl[71] br[71] wl[86] vdd gnd cell_6t
Xbit_r87_c71 bl[71] br[71] wl[87] vdd gnd cell_6t
Xbit_r88_c71 bl[71] br[71] wl[88] vdd gnd cell_6t
Xbit_r89_c71 bl[71] br[71] wl[89] vdd gnd cell_6t
Xbit_r90_c71 bl[71] br[71] wl[90] vdd gnd cell_6t
Xbit_r91_c71 bl[71] br[71] wl[91] vdd gnd cell_6t
Xbit_r92_c71 bl[71] br[71] wl[92] vdd gnd cell_6t
Xbit_r93_c71 bl[71] br[71] wl[93] vdd gnd cell_6t
Xbit_r94_c71 bl[71] br[71] wl[94] vdd gnd cell_6t
Xbit_r95_c71 bl[71] br[71] wl[95] vdd gnd cell_6t
Xbit_r96_c71 bl[71] br[71] wl[96] vdd gnd cell_6t
Xbit_r97_c71 bl[71] br[71] wl[97] vdd gnd cell_6t
Xbit_r98_c71 bl[71] br[71] wl[98] vdd gnd cell_6t
Xbit_r99_c71 bl[71] br[71] wl[99] vdd gnd cell_6t
Xbit_r100_c71 bl[71] br[71] wl[100] vdd gnd cell_6t
Xbit_r101_c71 bl[71] br[71] wl[101] vdd gnd cell_6t
Xbit_r102_c71 bl[71] br[71] wl[102] vdd gnd cell_6t
Xbit_r103_c71 bl[71] br[71] wl[103] vdd gnd cell_6t
Xbit_r104_c71 bl[71] br[71] wl[104] vdd gnd cell_6t
Xbit_r105_c71 bl[71] br[71] wl[105] vdd gnd cell_6t
Xbit_r106_c71 bl[71] br[71] wl[106] vdd gnd cell_6t
Xbit_r107_c71 bl[71] br[71] wl[107] vdd gnd cell_6t
Xbit_r108_c71 bl[71] br[71] wl[108] vdd gnd cell_6t
Xbit_r109_c71 bl[71] br[71] wl[109] vdd gnd cell_6t
Xbit_r110_c71 bl[71] br[71] wl[110] vdd gnd cell_6t
Xbit_r111_c71 bl[71] br[71] wl[111] vdd gnd cell_6t
Xbit_r112_c71 bl[71] br[71] wl[112] vdd gnd cell_6t
Xbit_r113_c71 bl[71] br[71] wl[113] vdd gnd cell_6t
Xbit_r114_c71 bl[71] br[71] wl[114] vdd gnd cell_6t
Xbit_r115_c71 bl[71] br[71] wl[115] vdd gnd cell_6t
Xbit_r116_c71 bl[71] br[71] wl[116] vdd gnd cell_6t
Xbit_r117_c71 bl[71] br[71] wl[117] vdd gnd cell_6t
Xbit_r118_c71 bl[71] br[71] wl[118] vdd gnd cell_6t
Xbit_r119_c71 bl[71] br[71] wl[119] vdd gnd cell_6t
Xbit_r120_c71 bl[71] br[71] wl[120] vdd gnd cell_6t
Xbit_r121_c71 bl[71] br[71] wl[121] vdd gnd cell_6t
Xbit_r122_c71 bl[71] br[71] wl[122] vdd gnd cell_6t
Xbit_r123_c71 bl[71] br[71] wl[123] vdd gnd cell_6t
Xbit_r124_c71 bl[71] br[71] wl[124] vdd gnd cell_6t
Xbit_r125_c71 bl[71] br[71] wl[125] vdd gnd cell_6t
Xbit_r126_c71 bl[71] br[71] wl[126] vdd gnd cell_6t
Xbit_r127_c71 bl[71] br[71] wl[127] vdd gnd cell_6t
Xbit_r128_c71 bl[71] br[71] wl[128] vdd gnd cell_6t
Xbit_r129_c71 bl[71] br[71] wl[129] vdd gnd cell_6t
Xbit_r130_c71 bl[71] br[71] wl[130] vdd gnd cell_6t
Xbit_r131_c71 bl[71] br[71] wl[131] vdd gnd cell_6t
Xbit_r132_c71 bl[71] br[71] wl[132] vdd gnd cell_6t
Xbit_r133_c71 bl[71] br[71] wl[133] vdd gnd cell_6t
Xbit_r134_c71 bl[71] br[71] wl[134] vdd gnd cell_6t
Xbit_r135_c71 bl[71] br[71] wl[135] vdd gnd cell_6t
Xbit_r136_c71 bl[71] br[71] wl[136] vdd gnd cell_6t
Xbit_r137_c71 bl[71] br[71] wl[137] vdd gnd cell_6t
Xbit_r138_c71 bl[71] br[71] wl[138] vdd gnd cell_6t
Xbit_r139_c71 bl[71] br[71] wl[139] vdd gnd cell_6t
Xbit_r140_c71 bl[71] br[71] wl[140] vdd gnd cell_6t
Xbit_r141_c71 bl[71] br[71] wl[141] vdd gnd cell_6t
Xbit_r142_c71 bl[71] br[71] wl[142] vdd gnd cell_6t
Xbit_r143_c71 bl[71] br[71] wl[143] vdd gnd cell_6t
Xbit_r144_c71 bl[71] br[71] wl[144] vdd gnd cell_6t
Xbit_r145_c71 bl[71] br[71] wl[145] vdd gnd cell_6t
Xbit_r146_c71 bl[71] br[71] wl[146] vdd gnd cell_6t
Xbit_r147_c71 bl[71] br[71] wl[147] vdd gnd cell_6t
Xbit_r148_c71 bl[71] br[71] wl[148] vdd gnd cell_6t
Xbit_r149_c71 bl[71] br[71] wl[149] vdd gnd cell_6t
Xbit_r150_c71 bl[71] br[71] wl[150] vdd gnd cell_6t
Xbit_r151_c71 bl[71] br[71] wl[151] vdd gnd cell_6t
Xbit_r152_c71 bl[71] br[71] wl[152] vdd gnd cell_6t
Xbit_r153_c71 bl[71] br[71] wl[153] vdd gnd cell_6t
Xbit_r154_c71 bl[71] br[71] wl[154] vdd gnd cell_6t
Xbit_r155_c71 bl[71] br[71] wl[155] vdd gnd cell_6t
Xbit_r156_c71 bl[71] br[71] wl[156] vdd gnd cell_6t
Xbit_r157_c71 bl[71] br[71] wl[157] vdd gnd cell_6t
Xbit_r158_c71 bl[71] br[71] wl[158] vdd gnd cell_6t
Xbit_r159_c71 bl[71] br[71] wl[159] vdd gnd cell_6t
Xbit_r160_c71 bl[71] br[71] wl[160] vdd gnd cell_6t
Xbit_r161_c71 bl[71] br[71] wl[161] vdd gnd cell_6t
Xbit_r162_c71 bl[71] br[71] wl[162] vdd gnd cell_6t
Xbit_r163_c71 bl[71] br[71] wl[163] vdd gnd cell_6t
Xbit_r164_c71 bl[71] br[71] wl[164] vdd gnd cell_6t
Xbit_r165_c71 bl[71] br[71] wl[165] vdd gnd cell_6t
Xbit_r166_c71 bl[71] br[71] wl[166] vdd gnd cell_6t
Xbit_r167_c71 bl[71] br[71] wl[167] vdd gnd cell_6t
Xbit_r168_c71 bl[71] br[71] wl[168] vdd gnd cell_6t
Xbit_r169_c71 bl[71] br[71] wl[169] vdd gnd cell_6t
Xbit_r170_c71 bl[71] br[71] wl[170] vdd gnd cell_6t
Xbit_r171_c71 bl[71] br[71] wl[171] vdd gnd cell_6t
Xbit_r172_c71 bl[71] br[71] wl[172] vdd gnd cell_6t
Xbit_r173_c71 bl[71] br[71] wl[173] vdd gnd cell_6t
Xbit_r174_c71 bl[71] br[71] wl[174] vdd gnd cell_6t
Xbit_r175_c71 bl[71] br[71] wl[175] vdd gnd cell_6t
Xbit_r176_c71 bl[71] br[71] wl[176] vdd gnd cell_6t
Xbit_r177_c71 bl[71] br[71] wl[177] vdd gnd cell_6t
Xbit_r178_c71 bl[71] br[71] wl[178] vdd gnd cell_6t
Xbit_r179_c71 bl[71] br[71] wl[179] vdd gnd cell_6t
Xbit_r180_c71 bl[71] br[71] wl[180] vdd gnd cell_6t
Xbit_r181_c71 bl[71] br[71] wl[181] vdd gnd cell_6t
Xbit_r182_c71 bl[71] br[71] wl[182] vdd gnd cell_6t
Xbit_r183_c71 bl[71] br[71] wl[183] vdd gnd cell_6t
Xbit_r184_c71 bl[71] br[71] wl[184] vdd gnd cell_6t
Xbit_r185_c71 bl[71] br[71] wl[185] vdd gnd cell_6t
Xbit_r186_c71 bl[71] br[71] wl[186] vdd gnd cell_6t
Xbit_r187_c71 bl[71] br[71] wl[187] vdd gnd cell_6t
Xbit_r188_c71 bl[71] br[71] wl[188] vdd gnd cell_6t
Xbit_r189_c71 bl[71] br[71] wl[189] vdd gnd cell_6t
Xbit_r190_c71 bl[71] br[71] wl[190] vdd gnd cell_6t
Xbit_r191_c71 bl[71] br[71] wl[191] vdd gnd cell_6t
Xbit_r192_c71 bl[71] br[71] wl[192] vdd gnd cell_6t
Xbit_r193_c71 bl[71] br[71] wl[193] vdd gnd cell_6t
Xbit_r194_c71 bl[71] br[71] wl[194] vdd gnd cell_6t
Xbit_r195_c71 bl[71] br[71] wl[195] vdd gnd cell_6t
Xbit_r196_c71 bl[71] br[71] wl[196] vdd gnd cell_6t
Xbit_r197_c71 bl[71] br[71] wl[197] vdd gnd cell_6t
Xbit_r198_c71 bl[71] br[71] wl[198] vdd gnd cell_6t
Xbit_r199_c71 bl[71] br[71] wl[199] vdd gnd cell_6t
Xbit_r200_c71 bl[71] br[71] wl[200] vdd gnd cell_6t
Xbit_r201_c71 bl[71] br[71] wl[201] vdd gnd cell_6t
Xbit_r202_c71 bl[71] br[71] wl[202] vdd gnd cell_6t
Xbit_r203_c71 bl[71] br[71] wl[203] vdd gnd cell_6t
Xbit_r204_c71 bl[71] br[71] wl[204] vdd gnd cell_6t
Xbit_r205_c71 bl[71] br[71] wl[205] vdd gnd cell_6t
Xbit_r206_c71 bl[71] br[71] wl[206] vdd gnd cell_6t
Xbit_r207_c71 bl[71] br[71] wl[207] vdd gnd cell_6t
Xbit_r208_c71 bl[71] br[71] wl[208] vdd gnd cell_6t
Xbit_r209_c71 bl[71] br[71] wl[209] vdd gnd cell_6t
Xbit_r210_c71 bl[71] br[71] wl[210] vdd gnd cell_6t
Xbit_r211_c71 bl[71] br[71] wl[211] vdd gnd cell_6t
Xbit_r212_c71 bl[71] br[71] wl[212] vdd gnd cell_6t
Xbit_r213_c71 bl[71] br[71] wl[213] vdd gnd cell_6t
Xbit_r214_c71 bl[71] br[71] wl[214] vdd gnd cell_6t
Xbit_r215_c71 bl[71] br[71] wl[215] vdd gnd cell_6t
Xbit_r216_c71 bl[71] br[71] wl[216] vdd gnd cell_6t
Xbit_r217_c71 bl[71] br[71] wl[217] vdd gnd cell_6t
Xbit_r218_c71 bl[71] br[71] wl[218] vdd gnd cell_6t
Xbit_r219_c71 bl[71] br[71] wl[219] vdd gnd cell_6t
Xbit_r220_c71 bl[71] br[71] wl[220] vdd gnd cell_6t
Xbit_r221_c71 bl[71] br[71] wl[221] vdd gnd cell_6t
Xbit_r222_c71 bl[71] br[71] wl[222] vdd gnd cell_6t
Xbit_r223_c71 bl[71] br[71] wl[223] vdd gnd cell_6t
Xbit_r224_c71 bl[71] br[71] wl[224] vdd gnd cell_6t
Xbit_r225_c71 bl[71] br[71] wl[225] vdd gnd cell_6t
Xbit_r226_c71 bl[71] br[71] wl[226] vdd gnd cell_6t
Xbit_r227_c71 bl[71] br[71] wl[227] vdd gnd cell_6t
Xbit_r228_c71 bl[71] br[71] wl[228] vdd gnd cell_6t
Xbit_r229_c71 bl[71] br[71] wl[229] vdd gnd cell_6t
Xbit_r230_c71 bl[71] br[71] wl[230] vdd gnd cell_6t
Xbit_r231_c71 bl[71] br[71] wl[231] vdd gnd cell_6t
Xbit_r232_c71 bl[71] br[71] wl[232] vdd gnd cell_6t
Xbit_r233_c71 bl[71] br[71] wl[233] vdd gnd cell_6t
Xbit_r234_c71 bl[71] br[71] wl[234] vdd gnd cell_6t
Xbit_r235_c71 bl[71] br[71] wl[235] vdd gnd cell_6t
Xbit_r236_c71 bl[71] br[71] wl[236] vdd gnd cell_6t
Xbit_r237_c71 bl[71] br[71] wl[237] vdd gnd cell_6t
Xbit_r238_c71 bl[71] br[71] wl[238] vdd gnd cell_6t
Xbit_r239_c71 bl[71] br[71] wl[239] vdd gnd cell_6t
Xbit_r240_c71 bl[71] br[71] wl[240] vdd gnd cell_6t
Xbit_r241_c71 bl[71] br[71] wl[241] vdd gnd cell_6t
Xbit_r242_c71 bl[71] br[71] wl[242] vdd gnd cell_6t
Xbit_r243_c71 bl[71] br[71] wl[243] vdd gnd cell_6t
Xbit_r244_c71 bl[71] br[71] wl[244] vdd gnd cell_6t
Xbit_r245_c71 bl[71] br[71] wl[245] vdd gnd cell_6t
Xbit_r246_c71 bl[71] br[71] wl[246] vdd gnd cell_6t
Xbit_r247_c71 bl[71] br[71] wl[247] vdd gnd cell_6t
Xbit_r248_c71 bl[71] br[71] wl[248] vdd gnd cell_6t
Xbit_r249_c71 bl[71] br[71] wl[249] vdd gnd cell_6t
Xbit_r250_c71 bl[71] br[71] wl[250] vdd gnd cell_6t
Xbit_r251_c71 bl[71] br[71] wl[251] vdd gnd cell_6t
Xbit_r252_c71 bl[71] br[71] wl[252] vdd gnd cell_6t
Xbit_r253_c71 bl[71] br[71] wl[253] vdd gnd cell_6t
Xbit_r254_c71 bl[71] br[71] wl[254] vdd gnd cell_6t
Xbit_r255_c71 bl[71] br[71] wl[255] vdd gnd cell_6t
Xbit_r0_c72 bl[72] br[72] wl[0] vdd gnd cell_6t
Xbit_r1_c72 bl[72] br[72] wl[1] vdd gnd cell_6t
Xbit_r2_c72 bl[72] br[72] wl[2] vdd gnd cell_6t
Xbit_r3_c72 bl[72] br[72] wl[3] vdd gnd cell_6t
Xbit_r4_c72 bl[72] br[72] wl[4] vdd gnd cell_6t
Xbit_r5_c72 bl[72] br[72] wl[5] vdd gnd cell_6t
Xbit_r6_c72 bl[72] br[72] wl[6] vdd gnd cell_6t
Xbit_r7_c72 bl[72] br[72] wl[7] vdd gnd cell_6t
Xbit_r8_c72 bl[72] br[72] wl[8] vdd gnd cell_6t
Xbit_r9_c72 bl[72] br[72] wl[9] vdd gnd cell_6t
Xbit_r10_c72 bl[72] br[72] wl[10] vdd gnd cell_6t
Xbit_r11_c72 bl[72] br[72] wl[11] vdd gnd cell_6t
Xbit_r12_c72 bl[72] br[72] wl[12] vdd gnd cell_6t
Xbit_r13_c72 bl[72] br[72] wl[13] vdd gnd cell_6t
Xbit_r14_c72 bl[72] br[72] wl[14] vdd gnd cell_6t
Xbit_r15_c72 bl[72] br[72] wl[15] vdd gnd cell_6t
Xbit_r16_c72 bl[72] br[72] wl[16] vdd gnd cell_6t
Xbit_r17_c72 bl[72] br[72] wl[17] vdd gnd cell_6t
Xbit_r18_c72 bl[72] br[72] wl[18] vdd gnd cell_6t
Xbit_r19_c72 bl[72] br[72] wl[19] vdd gnd cell_6t
Xbit_r20_c72 bl[72] br[72] wl[20] vdd gnd cell_6t
Xbit_r21_c72 bl[72] br[72] wl[21] vdd gnd cell_6t
Xbit_r22_c72 bl[72] br[72] wl[22] vdd gnd cell_6t
Xbit_r23_c72 bl[72] br[72] wl[23] vdd gnd cell_6t
Xbit_r24_c72 bl[72] br[72] wl[24] vdd gnd cell_6t
Xbit_r25_c72 bl[72] br[72] wl[25] vdd gnd cell_6t
Xbit_r26_c72 bl[72] br[72] wl[26] vdd gnd cell_6t
Xbit_r27_c72 bl[72] br[72] wl[27] vdd gnd cell_6t
Xbit_r28_c72 bl[72] br[72] wl[28] vdd gnd cell_6t
Xbit_r29_c72 bl[72] br[72] wl[29] vdd gnd cell_6t
Xbit_r30_c72 bl[72] br[72] wl[30] vdd gnd cell_6t
Xbit_r31_c72 bl[72] br[72] wl[31] vdd gnd cell_6t
Xbit_r32_c72 bl[72] br[72] wl[32] vdd gnd cell_6t
Xbit_r33_c72 bl[72] br[72] wl[33] vdd gnd cell_6t
Xbit_r34_c72 bl[72] br[72] wl[34] vdd gnd cell_6t
Xbit_r35_c72 bl[72] br[72] wl[35] vdd gnd cell_6t
Xbit_r36_c72 bl[72] br[72] wl[36] vdd gnd cell_6t
Xbit_r37_c72 bl[72] br[72] wl[37] vdd gnd cell_6t
Xbit_r38_c72 bl[72] br[72] wl[38] vdd gnd cell_6t
Xbit_r39_c72 bl[72] br[72] wl[39] vdd gnd cell_6t
Xbit_r40_c72 bl[72] br[72] wl[40] vdd gnd cell_6t
Xbit_r41_c72 bl[72] br[72] wl[41] vdd gnd cell_6t
Xbit_r42_c72 bl[72] br[72] wl[42] vdd gnd cell_6t
Xbit_r43_c72 bl[72] br[72] wl[43] vdd gnd cell_6t
Xbit_r44_c72 bl[72] br[72] wl[44] vdd gnd cell_6t
Xbit_r45_c72 bl[72] br[72] wl[45] vdd gnd cell_6t
Xbit_r46_c72 bl[72] br[72] wl[46] vdd gnd cell_6t
Xbit_r47_c72 bl[72] br[72] wl[47] vdd gnd cell_6t
Xbit_r48_c72 bl[72] br[72] wl[48] vdd gnd cell_6t
Xbit_r49_c72 bl[72] br[72] wl[49] vdd gnd cell_6t
Xbit_r50_c72 bl[72] br[72] wl[50] vdd gnd cell_6t
Xbit_r51_c72 bl[72] br[72] wl[51] vdd gnd cell_6t
Xbit_r52_c72 bl[72] br[72] wl[52] vdd gnd cell_6t
Xbit_r53_c72 bl[72] br[72] wl[53] vdd gnd cell_6t
Xbit_r54_c72 bl[72] br[72] wl[54] vdd gnd cell_6t
Xbit_r55_c72 bl[72] br[72] wl[55] vdd gnd cell_6t
Xbit_r56_c72 bl[72] br[72] wl[56] vdd gnd cell_6t
Xbit_r57_c72 bl[72] br[72] wl[57] vdd gnd cell_6t
Xbit_r58_c72 bl[72] br[72] wl[58] vdd gnd cell_6t
Xbit_r59_c72 bl[72] br[72] wl[59] vdd gnd cell_6t
Xbit_r60_c72 bl[72] br[72] wl[60] vdd gnd cell_6t
Xbit_r61_c72 bl[72] br[72] wl[61] vdd gnd cell_6t
Xbit_r62_c72 bl[72] br[72] wl[62] vdd gnd cell_6t
Xbit_r63_c72 bl[72] br[72] wl[63] vdd gnd cell_6t
Xbit_r64_c72 bl[72] br[72] wl[64] vdd gnd cell_6t
Xbit_r65_c72 bl[72] br[72] wl[65] vdd gnd cell_6t
Xbit_r66_c72 bl[72] br[72] wl[66] vdd gnd cell_6t
Xbit_r67_c72 bl[72] br[72] wl[67] vdd gnd cell_6t
Xbit_r68_c72 bl[72] br[72] wl[68] vdd gnd cell_6t
Xbit_r69_c72 bl[72] br[72] wl[69] vdd gnd cell_6t
Xbit_r70_c72 bl[72] br[72] wl[70] vdd gnd cell_6t
Xbit_r71_c72 bl[72] br[72] wl[71] vdd gnd cell_6t
Xbit_r72_c72 bl[72] br[72] wl[72] vdd gnd cell_6t
Xbit_r73_c72 bl[72] br[72] wl[73] vdd gnd cell_6t
Xbit_r74_c72 bl[72] br[72] wl[74] vdd gnd cell_6t
Xbit_r75_c72 bl[72] br[72] wl[75] vdd gnd cell_6t
Xbit_r76_c72 bl[72] br[72] wl[76] vdd gnd cell_6t
Xbit_r77_c72 bl[72] br[72] wl[77] vdd gnd cell_6t
Xbit_r78_c72 bl[72] br[72] wl[78] vdd gnd cell_6t
Xbit_r79_c72 bl[72] br[72] wl[79] vdd gnd cell_6t
Xbit_r80_c72 bl[72] br[72] wl[80] vdd gnd cell_6t
Xbit_r81_c72 bl[72] br[72] wl[81] vdd gnd cell_6t
Xbit_r82_c72 bl[72] br[72] wl[82] vdd gnd cell_6t
Xbit_r83_c72 bl[72] br[72] wl[83] vdd gnd cell_6t
Xbit_r84_c72 bl[72] br[72] wl[84] vdd gnd cell_6t
Xbit_r85_c72 bl[72] br[72] wl[85] vdd gnd cell_6t
Xbit_r86_c72 bl[72] br[72] wl[86] vdd gnd cell_6t
Xbit_r87_c72 bl[72] br[72] wl[87] vdd gnd cell_6t
Xbit_r88_c72 bl[72] br[72] wl[88] vdd gnd cell_6t
Xbit_r89_c72 bl[72] br[72] wl[89] vdd gnd cell_6t
Xbit_r90_c72 bl[72] br[72] wl[90] vdd gnd cell_6t
Xbit_r91_c72 bl[72] br[72] wl[91] vdd gnd cell_6t
Xbit_r92_c72 bl[72] br[72] wl[92] vdd gnd cell_6t
Xbit_r93_c72 bl[72] br[72] wl[93] vdd gnd cell_6t
Xbit_r94_c72 bl[72] br[72] wl[94] vdd gnd cell_6t
Xbit_r95_c72 bl[72] br[72] wl[95] vdd gnd cell_6t
Xbit_r96_c72 bl[72] br[72] wl[96] vdd gnd cell_6t
Xbit_r97_c72 bl[72] br[72] wl[97] vdd gnd cell_6t
Xbit_r98_c72 bl[72] br[72] wl[98] vdd gnd cell_6t
Xbit_r99_c72 bl[72] br[72] wl[99] vdd gnd cell_6t
Xbit_r100_c72 bl[72] br[72] wl[100] vdd gnd cell_6t
Xbit_r101_c72 bl[72] br[72] wl[101] vdd gnd cell_6t
Xbit_r102_c72 bl[72] br[72] wl[102] vdd gnd cell_6t
Xbit_r103_c72 bl[72] br[72] wl[103] vdd gnd cell_6t
Xbit_r104_c72 bl[72] br[72] wl[104] vdd gnd cell_6t
Xbit_r105_c72 bl[72] br[72] wl[105] vdd gnd cell_6t
Xbit_r106_c72 bl[72] br[72] wl[106] vdd gnd cell_6t
Xbit_r107_c72 bl[72] br[72] wl[107] vdd gnd cell_6t
Xbit_r108_c72 bl[72] br[72] wl[108] vdd gnd cell_6t
Xbit_r109_c72 bl[72] br[72] wl[109] vdd gnd cell_6t
Xbit_r110_c72 bl[72] br[72] wl[110] vdd gnd cell_6t
Xbit_r111_c72 bl[72] br[72] wl[111] vdd gnd cell_6t
Xbit_r112_c72 bl[72] br[72] wl[112] vdd gnd cell_6t
Xbit_r113_c72 bl[72] br[72] wl[113] vdd gnd cell_6t
Xbit_r114_c72 bl[72] br[72] wl[114] vdd gnd cell_6t
Xbit_r115_c72 bl[72] br[72] wl[115] vdd gnd cell_6t
Xbit_r116_c72 bl[72] br[72] wl[116] vdd gnd cell_6t
Xbit_r117_c72 bl[72] br[72] wl[117] vdd gnd cell_6t
Xbit_r118_c72 bl[72] br[72] wl[118] vdd gnd cell_6t
Xbit_r119_c72 bl[72] br[72] wl[119] vdd gnd cell_6t
Xbit_r120_c72 bl[72] br[72] wl[120] vdd gnd cell_6t
Xbit_r121_c72 bl[72] br[72] wl[121] vdd gnd cell_6t
Xbit_r122_c72 bl[72] br[72] wl[122] vdd gnd cell_6t
Xbit_r123_c72 bl[72] br[72] wl[123] vdd gnd cell_6t
Xbit_r124_c72 bl[72] br[72] wl[124] vdd gnd cell_6t
Xbit_r125_c72 bl[72] br[72] wl[125] vdd gnd cell_6t
Xbit_r126_c72 bl[72] br[72] wl[126] vdd gnd cell_6t
Xbit_r127_c72 bl[72] br[72] wl[127] vdd gnd cell_6t
Xbit_r128_c72 bl[72] br[72] wl[128] vdd gnd cell_6t
Xbit_r129_c72 bl[72] br[72] wl[129] vdd gnd cell_6t
Xbit_r130_c72 bl[72] br[72] wl[130] vdd gnd cell_6t
Xbit_r131_c72 bl[72] br[72] wl[131] vdd gnd cell_6t
Xbit_r132_c72 bl[72] br[72] wl[132] vdd gnd cell_6t
Xbit_r133_c72 bl[72] br[72] wl[133] vdd gnd cell_6t
Xbit_r134_c72 bl[72] br[72] wl[134] vdd gnd cell_6t
Xbit_r135_c72 bl[72] br[72] wl[135] vdd gnd cell_6t
Xbit_r136_c72 bl[72] br[72] wl[136] vdd gnd cell_6t
Xbit_r137_c72 bl[72] br[72] wl[137] vdd gnd cell_6t
Xbit_r138_c72 bl[72] br[72] wl[138] vdd gnd cell_6t
Xbit_r139_c72 bl[72] br[72] wl[139] vdd gnd cell_6t
Xbit_r140_c72 bl[72] br[72] wl[140] vdd gnd cell_6t
Xbit_r141_c72 bl[72] br[72] wl[141] vdd gnd cell_6t
Xbit_r142_c72 bl[72] br[72] wl[142] vdd gnd cell_6t
Xbit_r143_c72 bl[72] br[72] wl[143] vdd gnd cell_6t
Xbit_r144_c72 bl[72] br[72] wl[144] vdd gnd cell_6t
Xbit_r145_c72 bl[72] br[72] wl[145] vdd gnd cell_6t
Xbit_r146_c72 bl[72] br[72] wl[146] vdd gnd cell_6t
Xbit_r147_c72 bl[72] br[72] wl[147] vdd gnd cell_6t
Xbit_r148_c72 bl[72] br[72] wl[148] vdd gnd cell_6t
Xbit_r149_c72 bl[72] br[72] wl[149] vdd gnd cell_6t
Xbit_r150_c72 bl[72] br[72] wl[150] vdd gnd cell_6t
Xbit_r151_c72 bl[72] br[72] wl[151] vdd gnd cell_6t
Xbit_r152_c72 bl[72] br[72] wl[152] vdd gnd cell_6t
Xbit_r153_c72 bl[72] br[72] wl[153] vdd gnd cell_6t
Xbit_r154_c72 bl[72] br[72] wl[154] vdd gnd cell_6t
Xbit_r155_c72 bl[72] br[72] wl[155] vdd gnd cell_6t
Xbit_r156_c72 bl[72] br[72] wl[156] vdd gnd cell_6t
Xbit_r157_c72 bl[72] br[72] wl[157] vdd gnd cell_6t
Xbit_r158_c72 bl[72] br[72] wl[158] vdd gnd cell_6t
Xbit_r159_c72 bl[72] br[72] wl[159] vdd gnd cell_6t
Xbit_r160_c72 bl[72] br[72] wl[160] vdd gnd cell_6t
Xbit_r161_c72 bl[72] br[72] wl[161] vdd gnd cell_6t
Xbit_r162_c72 bl[72] br[72] wl[162] vdd gnd cell_6t
Xbit_r163_c72 bl[72] br[72] wl[163] vdd gnd cell_6t
Xbit_r164_c72 bl[72] br[72] wl[164] vdd gnd cell_6t
Xbit_r165_c72 bl[72] br[72] wl[165] vdd gnd cell_6t
Xbit_r166_c72 bl[72] br[72] wl[166] vdd gnd cell_6t
Xbit_r167_c72 bl[72] br[72] wl[167] vdd gnd cell_6t
Xbit_r168_c72 bl[72] br[72] wl[168] vdd gnd cell_6t
Xbit_r169_c72 bl[72] br[72] wl[169] vdd gnd cell_6t
Xbit_r170_c72 bl[72] br[72] wl[170] vdd gnd cell_6t
Xbit_r171_c72 bl[72] br[72] wl[171] vdd gnd cell_6t
Xbit_r172_c72 bl[72] br[72] wl[172] vdd gnd cell_6t
Xbit_r173_c72 bl[72] br[72] wl[173] vdd gnd cell_6t
Xbit_r174_c72 bl[72] br[72] wl[174] vdd gnd cell_6t
Xbit_r175_c72 bl[72] br[72] wl[175] vdd gnd cell_6t
Xbit_r176_c72 bl[72] br[72] wl[176] vdd gnd cell_6t
Xbit_r177_c72 bl[72] br[72] wl[177] vdd gnd cell_6t
Xbit_r178_c72 bl[72] br[72] wl[178] vdd gnd cell_6t
Xbit_r179_c72 bl[72] br[72] wl[179] vdd gnd cell_6t
Xbit_r180_c72 bl[72] br[72] wl[180] vdd gnd cell_6t
Xbit_r181_c72 bl[72] br[72] wl[181] vdd gnd cell_6t
Xbit_r182_c72 bl[72] br[72] wl[182] vdd gnd cell_6t
Xbit_r183_c72 bl[72] br[72] wl[183] vdd gnd cell_6t
Xbit_r184_c72 bl[72] br[72] wl[184] vdd gnd cell_6t
Xbit_r185_c72 bl[72] br[72] wl[185] vdd gnd cell_6t
Xbit_r186_c72 bl[72] br[72] wl[186] vdd gnd cell_6t
Xbit_r187_c72 bl[72] br[72] wl[187] vdd gnd cell_6t
Xbit_r188_c72 bl[72] br[72] wl[188] vdd gnd cell_6t
Xbit_r189_c72 bl[72] br[72] wl[189] vdd gnd cell_6t
Xbit_r190_c72 bl[72] br[72] wl[190] vdd gnd cell_6t
Xbit_r191_c72 bl[72] br[72] wl[191] vdd gnd cell_6t
Xbit_r192_c72 bl[72] br[72] wl[192] vdd gnd cell_6t
Xbit_r193_c72 bl[72] br[72] wl[193] vdd gnd cell_6t
Xbit_r194_c72 bl[72] br[72] wl[194] vdd gnd cell_6t
Xbit_r195_c72 bl[72] br[72] wl[195] vdd gnd cell_6t
Xbit_r196_c72 bl[72] br[72] wl[196] vdd gnd cell_6t
Xbit_r197_c72 bl[72] br[72] wl[197] vdd gnd cell_6t
Xbit_r198_c72 bl[72] br[72] wl[198] vdd gnd cell_6t
Xbit_r199_c72 bl[72] br[72] wl[199] vdd gnd cell_6t
Xbit_r200_c72 bl[72] br[72] wl[200] vdd gnd cell_6t
Xbit_r201_c72 bl[72] br[72] wl[201] vdd gnd cell_6t
Xbit_r202_c72 bl[72] br[72] wl[202] vdd gnd cell_6t
Xbit_r203_c72 bl[72] br[72] wl[203] vdd gnd cell_6t
Xbit_r204_c72 bl[72] br[72] wl[204] vdd gnd cell_6t
Xbit_r205_c72 bl[72] br[72] wl[205] vdd gnd cell_6t
Xbit_r206_c72 bl[72] br[72] wl[206] vdd gnd cell_6t
Xbit_r207_c72 bl[72] br[72] wl[207] vdd gnd cell_6t
Xbit_r208_c72 bl[72] br[72] wl[208] vdd gnd cell_6t
Xbit_r209_c72 bl[72] br[72] wl[209] vdd gnd cell_6t
Xbit_r210_c72 bl[72] br[72] wl[210] vdd gnd cell_6t
Xbit_r211_c72 bl[72] br[72] wl[211] vdd gnd cell_6t
Xbit_r212_c72 bl[72] br[72] wl[212] vdd gnd cell_6t
Xbit_r213_c72 bl[72] br[72] wl[213] vdd gnd cell_6t
Xbit_r214_c72 bl[72] br[72] wl[214] vdd gnd cell_6t
Xbit_r215_c72 bl[72] br[72] wl[215] vdd gnd cell_6t
Xbit_r216_c72 bl[72] br[72] wl[216] vdd gnd cell_6t
Xbit_r217_c72 bl[72] br[72] wl[217] vdd gnd cell_6t
Xbit_r218_c72 bl[72] br[72] wl[218] vdd gnd cell_6t
Xbit_r219_c72 bl[72] br[72] wl[219] vdd gnd cell_6t
Xbit_r220_c72 bl[72] br[72] wl[220] vdd gnd cell_6t
Xbit_r221_c72 bl[72] br[72] wl[221] vdd gnd cell_6t
Xbit_r222_c72 bl[72] br[72] wl[222] vdd gnd cell_6t
Xbit_r223_c72 bl[72] br[72] wl[223] vdd gnd cell_6t
Xbit_r224_c72 bl[72] br[72] wl[224] vdd gnd cell_6t
Xbit_r225_c72 bl[72] br[72] wl[225] vdd gnd cell_6t
Xbit_r226_c72 bl[72] br[72] wl[226] vdd gnd cell_6t
Xbit_r227_c72 bl[72] br[72] wl[227] vdd gnd cell_6t
Xbit_r228_c72 bl[72] br[72] wl[228] vdd gnd cell_6t
Xbit_r229_c72 bl[72] br[72] wl[229] vdd gnd cell_6t
Xbit_r230_c72 bl[72] br[72] wl[230] vdd gnd cell_6t
Xbit_r231_c72 bl[72] br[72] wl[231] vdd gnd cell_6t
Xbit_r232_c72 bl[72] br[72] wl[232] vdd gnd cell_6t
Xbit_r233_c72 bl[72] br[72] wl[233] vdd gnd cell_6t
Xbit_r234_c72 bl[72] br[72] wl[234] vdd gnd cell_6t
Xbit_r235_c72 bl[72] br[72] wl[235] vdd gnd cell_6t
Xbit_r236_c72 bl[72] br[72] wl[236] vdd gnd cell_6t
Xbit_r237_c72 bl[72] br[72] wl[237] vdd gnd cell_6t
Xbit_r238_c72 bl[72] br[72] wl[238] vdd gnd cell_6t
Xbit_r239_c72 bl[72] br[72] wl[239] vdd gnd cell_6t
Xbit_r240_c72 bl[72] br[72] wl[240] vdd gnd cell_6t
Xbit_r241_c72 bl[72] br[72] wl[241] vdd gnd cell_6t
Xbit_r242_c72 bl[72] br[72] wl[242] vdd gnd cell_6t
Xbit_r243_c72 bl[72] br[72] wl[243] vdd gnd cell_6t
Xbit_r244_c72 bl[72] br[72] wl[244] vdd gnd cell_6t
Xbit_r245_c72 bl[72] br[72] wl[245] vdd gnd cell_6t
Xbit_r246_c72 bl[72] br[72] wl[246] vdd gnd cell_6t
Xbit_r247_c72 bl[72] br[72] wl[247] vdd gnd cell_6t
Xbit_r248_c72 bl[72] br[72] wl[248] vdd gnd cell_6t
Xbit_r249_c72 bl[72] br[72] wl[249] vdd gnd cell_6t
Xbit_r250_c72 bl[72] br[72] wl[250] vdd gnd cell_6t
Xbit_r251_c72 bl[72] br[72] wl[251] vdd gnd cell_6t
Xbit_r252_c72 bl[72] br[72] wl[252] vdd gnd cell_6t
Xbit_r253_c72 bl[72] br[72] wl[253] vdd gnd cell_6t
Xbit_r254_c72 bl[72] br[72] wl[254] vdd gnd cell_6t
Xbit_r255_c72 bl[72] br[72] wl[255] vdd gnd cell_6t
Xbit_r0_c73 bl[73] br[73] wl[0] vdd gnd cell_6t
Xbit_r1_c73 bl[73] br[73] wl[1] vdd gnd cell_6t
Xbit_r2_c73 bl[73] br[73] wl[2] vdd gnd cell_6t
Xbit_r3_c73 bl[73] br[73] wl[3] vdd gnd cell_6t
Xbit_r4_c73 bl[73] br[73] wl[4] vdd gnd cell_6t
Xbit_r5_c73 bl[73] br[73] wl[5] vdd gnd cell_6t
Xbit_r6_c73 bl[73] br[73] wl[6] vdd gnd cell_6t
Xbit_r7_c73 bl[73] br[73] wl[7] vdd gnd cell_6t
Xbit_r8_c73 bl[73] br[73] wl[8] vdd gnd cell_6t
Xbit_r9_c73 bl[73] br[73] wl[9] vdd gnd cell_6t
Xbit_r10_c73 bl[73] br[73] wl[10] vdd gnd cell_6t
Xbit_r11_c73 bl[73] br[73] wl[11] vdd gnd cell_6t
Xbit_r12_c73 bl[73] br[73] wl[12] vdd gnd cell_6t
Xbit_r13_c73 bl[73] br[73] wl[13] vdd gnd cell_6t
Xbit_r14_c73 bl[73] br[73] wl[14] vdd gnd cell_6t
Xbit_r15_c73 bl[73] br[73] wl[15] vdd gnd cell_6t
Xbit_r16_c73 bl[73] br[73] wl[16] vdd gnd cell_6t
Xbit_r17_c73 bl[73] br[73] wl[17] vdd gnd cell_6t
Xbit_r18_c73 bl[73] br[73] wl[18] vdd gnd cell_6t
Xbit_r19_c73 bl[73] br[73] wl[19] vdd gnd cell_6t
Xbit_r20_c73 bl[73] br[73] wl[20] vdd gnd cell_6t
Xbit_r21_c73 bl[73] br[73] wl[21] vdd gnd cell_6t
Xbit_r22_c73 bl[73] br[73] wl[22] vdd gnd cell_6t
Xbit_r23_c73 bl[73] br[73] wl[23] vdd gnd cell_6t
Xbit_r24_c73 bl[73] br[73] wl[24] vdd gnd cell_6t
Xbit_r25_c73 bl[73] br[73] wl[25] vdd gnd cell_6t
Xbit_r26_c73 bl[73] br[73] wl[26] vdd gnd cell_6t
Xbit_r27_c73 bl[73] br[73] wl[27] vdd gnd cell_6t
Xbit_r28_c73 bl[73] br[73] wl[28] vdd gnd cell_6t
Xbit_r29_c73 bl[73] br[73] wl[29] vdd gnd cell_6t
Xbit_r30_c73 bl[73] br[73] wl[30] vdd gnd cell_6t
Xbit_r31_c73 bl[73] br[73] wl[31] vdd gnd cell_6t
Xbit_r32_c73 bl[73] br[73] wl[32] vdd gnd cell_6t
Xbit_r33_c73 bl[73] br[73] wl[33] vdd gnd cell_6t
Xbit_r34_c73 bl[73] br[73] wl[34] vdd gnd cell_6t
Xbit_r35_c73 bl[73] br[73] wl[35] vdd gnd cell_6t
Xbit_r36_c73 bl[73] br[73] wl[36] vdd gnd cell_6t
Xbit_r37_c73 bl[73] br[73] wl[37] vdd gnd cell_6t
Xbit_r38_c73 bl[73] br[73] wl[38] vdd gnd cell_6t
Xbit_r39_c73 bl[73] br[73] wl[39] vdd gnd cell_6t
Xbit_r40_c73 bl[73] br[73] wl[40] vdd gnd cell_6t
Xbit_r41_c73 bl[73] br[73] wl[41] vdd gnd cell_6t
Xbit_r42_c73 bl[73] br[73] wl[42] vdd gnd cell_6t
Xbit_r43_c73 bl[73] br[73] wl[43] vdd gnd cell_6t
Xbit_r44_c73 bl[73] br[73] wl[44] vdd gnd cell_6t
Xbit_r45_c73 bl[73] br[73] wl[45] vdd gnd cell_6t
Xbit_r46_c73 bl[73] br[73] wl[46] vdd gnd cell_6t
Xbit_r47_c73 bl[73] br[73] wl[47] vdd gnd cell_6t
Xbit_r48_c73 bl[73] br[73] wl[48] vdd gnd cell_6t
Xbit_r49_c73 bl[73] br[73] wl[49] vdd gnd cell_6t
Xbit_r50_c73 bl[73] br[73] wl[50] vdd gnd cell_6t
Xbit_r51_c73 bl[73] br[73] wl[51] vdd gnd cell_6t
Xbit_r52_c73 bl[73] br[73] wl[52] vdd gnd cell_6t
Xbit_r53_c73 bl[73] br[73] wl[53] vdd gnd cell_6t
Xbit_r54_c73 bl[73] br[73] wl[54] vdd gnd cell_6t
Xbit_r55_c73 bl[73] br[73] wl[55] vdd gnd cell_6t
Xbit_r56_c73 bl[73] br[73] wl[56] vdd gnd cell_6t
Xbit_r57_c73 bl[73] br[73] wl[57] vdd gnd cell_6t
Xbit_r58_c73 bl[73] br[73] wl[58] vdd gnd cell_6t
Xbit_r59_c73 bl[73] br[73] wl[59] vdd gnd cell_6t
Xbit_r60_c73 bl[73] br[73] wl[60] vdd gnd cell_6t
Xbit_r61_c73 bl[73] br[73] wl[61] vdd gnd cell_6t
Xbit_r62_c73 bl[73] br[73] wl[62] vdd gnd cell_6t
Xbit_r63_c73 bl[73] br[73] wl[63] vdd gnd cell_6t
Xbit_r64_c73 bl[73] br[73] wl[64] vdd gnd cell_6t
Xbit_r65_c73 bl[73] br[73] wl[65] vdd gnd cell_6t
Xbit_r66_c73 bl[73] br[73] wl[66] vdd gnd cell_6t
Xbit_r67_c73 bl[73] br[73] wl[67] vdd gnd cell_6t
Xbit_r68_c73 bl[73] br[73] wl[68] vdd gnd cell_6t
Xbit_r69_c73 bl[73] br[73] wl[69] vdd gnd cell_6t
Xbit_r70_c73 bl[73] br[73] wl[70] vdd gnd cell_6t
Xbit_r71_c73 bl[73] br[73] wl[71] vdd gnd cell_6t
Xbit_r72_c73 bl[73] br[73] wl[72] vdd gnd cell_6t
Xbit_r73_c73 bl[73] br[73] wl[73] vdd gnd cell_6t
Xbit_r74_c73 bl[73] br[73] wl[74] vdd gnd cell_6t
Xbit_r75_c73 bl[73] br[73] wl[75] vdd gnd cell_6t
Xbit_r76_c73 bl[73] br[73] wl[76] vdd gnd cell_6t
Xbit_r77_c73 bl[73] br[73] wl[77] vdd gnd cell_6t
Xbit_r78_c73 bl[73] br[73] wl[78] vdd gnd cell_6t
Xbit_r79_c73 bl[73] br[73] wl[79] vdd gnd cell_6t
Xbit_r80_c73 bl[73] br[73] wl[80] vdd gnd cell_6t
Xbit_r81_c73 bl[73] br[73] wl[81] vdd gnd cell_6t
Xbit_r82_c73 bl[73] br[73] wl[82] vdd gnd cell_6t
Xbit_r83_c73 bl[73] br[73] wl[83] vdd gnd cell_6t
Xbit_r84_c73 bl[73] br[73] wl[84] vdd gnd cell_6t
Xbit_r85_c73 bl[73] br[73] wl[85] vdd gnd cell_6t
Xbit_r86_c73 bl[73] br[73] wl[86] vdd gnd cell_6t
Xbit_r87_c73 bl[73] br[73] wl[87] vdd gnd cell_6t
Xbit_r88_c73 bl[73] br[73] wl[88] vdd gnd cell_6t
Xbit_r89_c73 bl[73] br[73] wl[89] vdd gnd cell_6t
Xbit_r90_c73 bl[73] br[73] wl[90] vdd gnd cell_6t
Xbit_r91_c73 bl[73] br[73] wl[91] vdd gnd cell_6t
Xbit_r92_c73 bl[73] br[73] wl[92] vdd gnd cell_6t
Xbit_r93_c73 bl[73] br[73] wl[93] vdd gnd cell_6t
Xbit_r94_c73 bl[73] br[73] wl[94] vdd gnd cell_6t
Xbit_r95_c73 bl[73] br[73] wl[95] vdd gnd cell_6t
Xbit_r96_c73 bl[73] br[73] wl[96] vdd gnd cell_6t
Xbit_r97_c73 bl[73] br[73] wl[97] vdd gnd cell_6t
Xbit_r98_c73 bl[73] br[73] wl[98] vdd gnd cell_6t
Xbit_r99_c73 bl[73] br[73] wl[99] vdd gnd cell_6t
Xbit_r100_c73 bl[73] br[73] wl[100] vdd gnd cell_6t
Xbit_r101_c73 bl[73] br[73] wl[101] vdd gnd cell_6t
Xbit_r102_c73 bl[73] br[73] wl[102] vdd gnd cell_6t
Xbit_r103_c73 bl[73] br[73] wl[103] vdd gnd cell_6t
Xbit_r104_c73 bl[73] br[73] wl[104] vdd gnd cell_6t
Xbit_r105_c73 bl[73] br[73] wl[105] vdd gnd cell_6t
Xbit_r106_c73 bl[73] br[73] wl[106] vdd gnd cell_6t
Xbit_r107_c73 bl[73] br[73] wl[107] vdd gnd cell_6t
Xbit_r108_c73 bl[73] br[73] wl[108] vdd gnd cell_6t
Xbit_r109_c73 bl[73] br[73] wl[109] vdd gnd cell_6t
Xbit_r110_c73 bl[73] br[73] wl[110] vdd gnd cell_6t
Xbit_r111_c73 bl[73] br[73] wl[111] vdd gnd cell_6t
Xbit_r112_c73 bl[73] br[73] wl[112] vdd gnd cell_6t
Xbit_r113_c73 bl[73] br[73] wl[113] vdd gnd cell_6t
Xbit_r114_c73 bl[73] br[73] wl[114] vdd gnd cell_6t
Xbit_r115_c73 bl[73] br[73] wl[115] vdd gnd cell_6t
Xbit_r116_c73 bl[73] br[73] wl[116] vdd gnd cell_6t
Xbit_r117_c73 bl[73] br[73] wl[117] vdd gnd cell_6t
Xbit_r118_c73 bl[73] br[73] wl[118] vdd gnd cell_6t
Xbit_r119_c73 bl[73] br[73] wl[119] vdd gnd cell_6t
Xbit_r120_c73 bl[73] br[73] wl[120] vdd gnd cell_6t
Xbit_r121_c73 bl[73] br[73] wl[121] vdd gnd cell_6t
Xbit_r122_c73 bl[73] br[73] wl[122] vdd gnd cell_6t
Xbit_r123_c73 bl[73] br[73] wl[123] vdd gnd cell_6t
Xbit_r124_c73 bl[73] br[73] wl[124] vdd gnd cell_6t
Xbit_r125_c73 bl[73] br[73] wl[125] vdd gnd cell_6t
Xbit_r126_c73 bl[73] br[73] wl[126] vdd gnd cell_6t
Xbit_r127_c73 bl[73] br[73] wl[127] vdd gnd cell_6t
Xbit_r128_c73 bl[73] br[73] wl[128] vdd gnd cell_6t
Xbit_r129_c73 bl[73] br[73] wl[129] vdd gnd cell_6t
Xbit_r130_c73 bl[73] br[73] wl[130] vdd gnd cell_6t
Xbit_r131_c73 bl[73] br[73] wl[131] vdd gnd cell_6t
Xbit_r132_c73 bl[73] br[73] wl[132] vdd gnd cell_6t
Xbit_r133_c73 bl[73] br[73] wl[133] vdd gnd cell_6t
Xbit_r134_c73 bl[73] br[73] wl[134] vdd gnd cell_6t
Xbit_r135_c73 bl[73] br[73] wl[135] vdd gnd cell_6t
Xbit_r136_c73 bl[73] br[73] wl[136] vdd gnd cell_6t
Xbit_r137_c73 bl[73] br[73] wl[137] vdd gnd cell_6t
Xbit_r138_c73 bl[73] br[73] wl[138] vdd gnd cell_6t
Xbit_r139_c73 bl[73] br[73] wl[139] vdd gnd cell_6t
Xbit_r140_c73 bl[73] br[73] wl[140] vdd gnd cell_6t
Xbit_r141_c73 bl[73] br[73] wl[141] vdd gnd cell_6t
Xbit_r142_c73 bl[73] br[73] wl[142] vdd gnd cell_6t
Xbit_r143_c73 bl[73] br[73] wl[143] vdd gnd cell_6t
Xbit_r144_c73 bl[73] br[73] wl[144] vdd gnd cell_6t
Xbit_r145_c73 bl[73] br[73] wl[145] vdd gnd cell_6t
Xbit_r146_c73 bl[73] br[73] wl[146] vdd gnd cell_6t
Xbit_r147_c73 bl[73] br[73] wl[147] vdd gnd cell_6t
Xbit_r148_c73 bl[73] br[73] wl[148] vdd gnd cell_6t
Xbit_r149_c73 bl[73] br[73] wl[149] vdd gnd cell_6t
Xbit_r150_c73 bl[73] br[73] wl[150] vdd gnd cell_6t
Xbit_r151_c73 bl[73] br[73] wl[151] vdd gnd cell_6t
Xbit_r152_c73 bl[73] br[73] wl[152] vdd gnd cell_6t
Xbit_r153_c73 bl[73] br[73] wl[153] vdd gnd cell_6t
Xbit_r154_c73 bl[73] br[73] wl[154] vdd gnd cell_6t
Xbit_r155_c73 bl[73] br[73] wl[155] vdd gnd cell_6t
Xbit_r156_c73 bl[73] br[73] wl[156] vdd gnd cell_6t
Xbit_r157_c73 bl[73] br[73] wl[157] vdd gnd cell_6t
Xbit_r158_c73 bl[73] br[73] wl[158] vdd gnd cell_6t
Xbit_r159_c73 bl[73] br[73] wl[159] vdd gnd cell_6t
Xbit_r160_c73 bl[73] br[73] wl[160] vdd gnd cell_6t
Xbit_r161_c73 bl[73] br[73] wl[161] vdd gnd cell_6t
Xbit_r162_c73 bl[73] br[73] wl[162] vdd gnd cell_6t
Xbit_r163_c73 bl[73] br[73] wl[163] vdd gnd cell_6t
Xbit_r164_c73 bl[73] br[73] wl[164] vdd gnd cell_6t
Xbit_r165_c73 bl[73] br[73] wl[165] vdd gnd cell_6t
Xbit_r166_c73 bl[73] br[73] wl[166] vdd gnd cell_6t
Xbit_r167_c73 bl[73] br[73] wl[167] vdd gnd cell_6t
Xbit_r168_c73 bl[73] br[73] wl[168] vdd gnd cell_6t
Xbit_r169_c73 bl[73] br[73] wl[169] vdd gnd cell_6t
Xbit_r170_c73 bl[73] br[73] wl[170] vdd gnd cell_6t
Xbit_r171_c73 bl[73] br[73] wl[171] vdd gnd cell_6t
Xbit_r172_c73 bl[73] br[73] wl[172] vdd gnd cell_6t
Xbit_r173_c73 bl[73] br[73] wl[173] vdd gnd cell_6t
Xbit_r174_c73 bl[73] br[73] wl[174] vdd gnd cell_6t
Xbit_r175_c73 bl[73] br[73] wl[175] vdd gnd cell_6t
Xbit_r176_c73 bl[73] br[73] wl[176] vdd gnd cell_6t
Xbit_r177_c73 bl[73] br[73] wl[177] vdd gnd cell_6t
Xbit_r178_c73 bl[73] br[73] wl[178] vdd gnd cell_6t
Xbit_r179_c73 bl[73] br[73] wl[179] vdd gnd cell_6t
Xbit_r180_c73 bl[73] br[73] wl[180] vdd gnd cell_6t
Xbit_r181_c73 bl[73] br[73] wl[181] vdd gnd cell_6t
Xbit_r182_c73 bl[73] br[73] wl[182] vdd gnd cell_6t
Xbit_r183_c73 bl[73] br[73] wl[183] vdd gnd cell_6t
Xbit_r184_c73 bl[73] br[73] wl[184] vdd gnd cell_6t
Xbit_r185_c73 bl[73] br[73] wl[185] vdd gnd cell_6t
Xbit_r186_c73 bl[73] br[73] wl[186] vdd gnd cell_6t
Xbit_r187_c73 bl[73] br[73] wl[187] vdd gnd cell_6t
Xbit_r188_c73 bl[73] br[73] wl[188] vdd gnd cell_6t
Xbit_r189_c73 bl[73] br[73] wl[189] vdd gnd cell_6t
Xbit_r190_c73 bl[73] br[73] wl[190] vdd gnd cell_6t
Xbit_r191_c73 bl[73] br[73] wl[191] vdd gnd cell_6t
Xbit_r192_c73 bl[73] br[73] wl[192] vdd gnd cell_6t
Xbit_r193_c73 bl[73] br[73] wl[193] vdd gnd cell_6t
Xbit_r194_c73 bl[73] br[73] wl[194] vdd gnd cell_6t
Xbit_r195_c73 bl[73] br[73] wl[195] vdd gnd cell_6t
Xbit_r196_c73 bl[73] br[73] wl[196] vdd gnd cell_6t
Xbit_r197_c73 bl[73] br[73] wl[197] vdd gnd cell_6t
Xbit_r198_c73 bl[73] br[73] wl[198] vdd gnd cell_6t
Xbit_r199_c73 bl[73] br[73] wl[199] vdd gnd cell_6t
Xbit_r200_c73 bl[73] br[73] wl[200] vdd gnd cell_6t
Xbit_r201_c73 bl[73] br[73] wl[201] vdd gnd cell_6t
Xbit_r202_c73 bl[73] br[73] wl[202] vdd gnd cell_6t
Xbit_r203_c73 bl[73] br[73] wl[203] vdd gnd cell_6t
Xbit_r204_c73 bl[73] br[73] wl[204] vdd gnd cell_6t
Xbit_r205_c73 bl[73] br[73] wl[205] vdd gnd cell_6t
Xbit_r206_c73 bl[73] br[73] wl[206] vdd gnd cell_6t
Xbit_r207_c73 bl[73] br[73] wl[207] vdd gnd cell_6t
Xbit_r208_c73 bl[73] br[73] wl[208] vdd gnd cell_6t
Xbit_r209_c73 bl[73] br[73] wl[209] vdd gnd cell_6t
Xbit_r210_c73 bl[73] br[73] wl[210] vdd gnd cell_6t
Xbit_r211_c73 bl[73] br[73] wl[211] vdd gnd cell_6t
Xbit_r212_c73 bl[73] br[73] wl[212] vdd gnd cell_6t
Xbit_r213_c73 bl[73] br[73] wl[213] vdd gnd cell_6t
Xbit_r214_c73 bl[73] br[73] wl[214] vdd gnd cell_6t
Xbit_r215_c73 bl[73] br[73] wl[215] vdd gnd cell_6t
Xbit_r216_c73 bl[73] br[73] wl[216] vdd gnd cell_6t
Xbit_r217_c73 bl[73] br[73] wl[217] vdd gnd cell_6t
Xbit_r218_c73 bl[73] br[73] wl[218] vdd gnd cell_6t
Xbit_r219_c73 bl[73] br[73] wl[219] vdd gnd cell_6t
Xbit_r220_c73 bl[73] br[73] wl[220] vdd gnd cell_6t
Xbit_r221_c73 bl[73] br[73] wl[221] vdd gnd cell_6t
Xbit_r222_c73 bl[73] br[73] wl[222] vdd gnd cell_6t
Xbit_r223_c73 bl[73] br[73] wl[223] vdd gnd cell_6t
Xbit_r224_c73 bl[73] br[73] wl[224] vdd gnd cell_6t
Xbit_r225_c73 bl[73] br[73] wl[225] vdd gnd cell_6t
Xbit_r226_c73 bl[73] br[73] wl[226] vdd gnd cell_6t
Xbit_r227_c73 bl[73] br[73] wl[227] vdd gnd cell_6t
Xbit_r228_c73 bl[73] br[73] wl[228] vdd gnd cell_6t
Xbit_r229_c73 bl[73] br[73] wl[229] vdd gnd cell_6t
Xbit_r230_c73 bl[73] br[73] wl[230] vdd gnd cell_6t
Xbit_r231_c73 bl[73] br[73] wl[231] vdd gnd cell_6t
Xbit_r232_c73 bl[73] br[73] wl[232] vdd gnd cell_6t
Xbit_r233_c73 bl[73] br[73] wl[233] vdd gnd cell_6t
Xbit_r234_c73 bl[73] br[73] wl[234] vdd gnd cell_6t
Xbit_r235_c73 bl[73] br[73] wl[235] vdd gnd cell_6t
Xbit_r236_c73 bl[73] br[73] wl[236] vdd gnd cell_6t
Xbit_r237_c73 bl[73] br[73] wl[237] vdd gnd cell_6t
Xbit_r238_c73 bl[73] br[73] wl[238] vdd gnd cell_6t
Xbit_r239_c73 bl[73] br[73] wl[239] vdd gnd cell_6t
Xbit_r240_c73 bl[73] br[73] wl[240] vdd gnd cell_6t
Xbit_r241_c73 bl[73] br[73] wl[241] vdd gnd cell_6t
Xbit_r242_c73 bl[73] br[73] wl[242] vdd gnd cell_6t
Xbit_r243_c73 bl[73] br[73] wl[243] vdd gnd cell_6t
Xbit_r244_c73 bl[73] br[73] wl[244] vdd gnd cell_6t
Xbit_r245_c73 bl[73] br[73] wl[245] vdd gnd cell_6t
Xbit_r246_c73 bl[73] br[73] wl[246] vdd gnd cell_6t
Xbit_r247_c73 bl[73] br[73] wl[247] vdd gnd cell_6t
Xbit_r248_c73 bl[73] br[73] wl[248] vdd gnd cell_6t
Xbit_r249_c73 bl[73] br[73] wl[249] vdd gnd cell_6t
Xbit_r250_c73 bl[73] br[73] wl[250] vdd gnd cell_6t
Xbit_r251_c73 bl[73] br[73] wl[251] vdd gnd cell_6t
Xbit_r252_c73 bl[73] br[73] wl[252] vdd gnd cell_6t
Xbit_r253_c73 bl[73] br[73] wl[253] vdd gnd cell_6t
Xbit_r254_c73 bl[73] br[73] wl[254] vdd gnd cell_6t
Xbit_r255_c73 bl[73] br[73] wl[255] vdd gnd cell_6t
Xbit_r0_c74 bl[74] br[74] wl[0] vdd gnd cell_6t
Xbit_r1_c74 bl[74] br[74] wl[1] vdd gnd cell_6t
Xbit_r2_c74 bl[74] br[74] wl[2] vdd gnd cell_6t
Xbit_r3_c74 bl[74] br[74] wl[3] vdd gnd cell_6t
Xbit_r4_c74 bl[74] br[74] wl[4] vdd gnd cell_6t
Xbit_r5_c74 bl[74] br[74] wl[5] vdd gnd cell_6t
Xbit_r6_c74 bl[74] br[74] wl[6] vdd gnd cell_6t
Xbit_r7_c74 bl[74] br[74] wl[7] vdd gnd cell_6t
Xbit_r8_c74 bl[74] br[74] wl[8] vdd gnd cell_6t
Xbit_r9_c74 bl[74] br[74] wl[9] vdd gnd cell_6t
Xbit_r10_c74 bl[74] br[74] wl[10] vdd gnd cell_6t
Xbit_r11_c74 bl[74] br[74] wl[11] vdd gnd cell_6t
Xbit_r12_c74 bl[74] br[74] wl[12] vdd gnd cell_6t
Xbit_r13_c74 bl[74] br[74] wl[13] vdd gnd cell_6t
Xbit_r14_c74 bl[74] br[74] wl[14] vdd gnd cell_6t
Xbit_r15_c74 bl[74] br[74] wl[15] vdd gnd cell_6t
Xbit_r16_c74 bl[74] br[74] wl[16] vdd gnd cell_6t
Xbit_r17_c74 bl[74] br[74] wl[17] vdd gnd cell_6t
Xbit_r18_c74 bl[74] br[74] wl[18] vdd gnd cell_6t
Xbit_r19_c74 bl[74] br[74] wl[19] vdd gnd cell_6t
Xbit_r20_c74 bl[74] br[74] wl[20] vdd gnd cell_6t
Xbit_r21_c74 bl[74] br[74] wl[21] vdd gnd cell_6t
Xbit_r22_c74 bl[74] br[74] wl[22] vdd gnd cell_6t
Xbit_r23_c74 bl[74] br[74] wl[23] vdd gnd cell_6t
Xbit_r24_c74 bl[74] br[74] wl[24] vdd gnd cell_6t
Xbit_r25_c74 bl[74] br[74] wl[25] vdd gnd cell_6t
Xbit_r26_c74 bl[74] br[74] wl[26] vdd gnd cell_6t
Xbit_r27_c74 bl[74] br[74] wl[27] vdd gnd cell_6t
Xbit_r28_c74 bl[74] br[74] wl[28] vdd gnd cell_6t
Xbit_r29_c74 bl[74] br[74] wl[29] vdd gnd cell_6t
Xbit_r30_c74 bl[74] br[74] wl[30] vdd gnd cell_6t
Xbit_r31_c74 bl[74] br[74] wl[31] vdd gnd cell_6t
Xbit_r32_c74 bl[74] br[74] wl[32] vdd gnd cell_6t
Xbit_r33_c74 bl[74] br[74] wl[33] vdd gnd cell_6t
Xbit_r34_c74 bl[74] br[74] wl[34] vdd gnd cell_6t
Xbit_r35_c74 bl[74] br[74] wl[35] vdd gnd cell_6t
Xbit_r36_c74 bl[74] br[74] wl[36] vdd gnd cell_6t
Xbit_r37_c74 bl[74] br[74] wl[37] vdd gnd cell_6t
Xbit_r38_c74 bl[74] br[74] wl[38] vdd gnd cell_6t
Xbit_r39_c74 bl[74] br[74] wl[39] vdd gnd cell_6t
Xbit_r40_c74 bl[74] br[74] wl[40] vdd gnd cell_6t
Xbit_r41_c74 bl[74] br[74] wl[41] vdd gnd cell_6t
Xbit_r42_c74 bl[74] br[74] wl[42] vdd gnd cell_6t
Xbit_r43_c74 bl[74] br[74] wl[43] vdd gnd cell_6t
Xbit_r44_c74 bl[74] br[74] wl[44] vdd gnd cell_6t
Xbit_r45_c74 bl[74] br[74] wl[45] vdd gnd cell_6t
Xbit_r46_c74 bl[74] br[74] wl[46] vdd gnd cell_6t
Xbit_r47_c74 bl[74] br[74] wl[47] vdd gnd cell_6t
Xbit_r48_c74 bl[74] br[74] wl[48] vdd gnd cell_6t
Xbit_r49_c74 bl[74] br[74] wl[49] vdd gnd cell_6t
Xbit_r50_c74 bl[74] br[74] wl[50] vdd gnd cell_6t
Xbit_r51_c74 bl[74] br[74] wl[51] vdd gnd cell_6t
Xbit_r52_c74 bl[74] br[74] wl[52] vdd gnd cell_6t
Xbit_r53_c74 bl[74] br[74] wl[53] vdd gnd cell_6t
Xbit_r54_c74 bl[74] br[74] wl[54] vdd gnd cell_6t
Xbit_r55_c74 bl[74] br[74] wl[55] vdd gnd cell_6t
Xbit_r56_c74 bl[74] br[74] wl[56] vdd gnd cell_6t
Xbit_r57_c74 bl[74] br[74] wl[57] vdd gnd cell_6t
Xbit_r58_c74 bl[74] br[74] wl[58] vdd gnd cell_6t
Xbit_r59_c74 bl[74] br[74] wl[59] vdd gnd cell_6t
Xbit_r60_c74 bl[74] br[74] wl[60] vdd gnd cell_6t
Xbit_r61_c74 bl[74] br[74] wl[61] vdd gnd cell_6t
Xbit_r62_c74 bl[74] br[74] wl[62] vdd gnd cell_6t
Xbit_r63_c74 bl[74] br[74] wl[63] vdd gnd cell_6t
Xbit_r64_c74 bl[74] br[74] wl[64] vdd gnd cell_6t
Xbit_r65_c74 bl[74] br[74] wl[65] vdd gnd cell_6t
Xbit_r66_c74 bl[74] br[74] wl[66] vdd gnd cell_6t
Xbit_r67_c74 bl[74] br[74] wl[67] vdd gnd cell_6t
Xbit_r68_c74 bl[74] br[74] wl[68] vdd gnd cell_6t
Xbit_r69_c74 bl[74] br[74] wl[69] vdd gnd cell_6t
Xbit_r70_c74 bl[74] br[74] wl[70] vdd gnd cell_6t
Xbit_r71_c74 bl[74] br[74] wl[71] vdd gnd cell_6t
Xbit_r72_c74 bl[74] br[74] wl[72] vdd gnd cell_6t
Xbit_r73_c74 bl[74] br[74] wl[73] vdd gnd cell_6t
Xbit_r74_c74 bl[74] br[74] wl[74] vdd gnd cell_6t
Xbit_r75_c74 bl[74] br[74] wl[75] vdd gnd cell_6t
Xbit_r76_c74 bl[74] br[74] wl[76] vdd gnd cell_6t
Xbit_r77_c74 bl[74] br[74] wl[77] vdd gnd cell_6t
Xbit_r78_c74 bl[74] br[74] wl[78] vdd gnd cell_6t
Xbit_r79_c74 bl[74] br[74] wl[79] vdd gnd cell_6t
Xbit_r80_c74 bl[74] br[74] wl[80] vdd gnd cell_6t
Xbit_r81_c74 bl[74] br[74] wl[81] vdd gnd cell_6t
Xbit_r82_c74 bl[74] br[74] wl[82] vdd gnd cell_6t
Xbit_r83_c74 bl[74] br[74] wl[83] vdd gnd cell_6t
Xbit_r84_c74 bl[74] br[74] wl[84] vdd gnd cell_6t
Xbit_r85_c74 bl[74] br[74] wl[85] vdd gnd cell_6t
Xbit_r86_c74 bl[74] br[74] wl[86] vdd gnd cell_6t
Xbit_r87_c74 bl[74] br[74] wl[87] vdd gnd cell_6t
Xbit_r88_c74 bl[74] br[74] wl[88] vdd gnd cell_6t
Xbit_r89_c74 bl[74] br[74] wl[89] vdd gnd cell_6t
Xbit_r90_c74 bl[74] br[74] wl[90] vdd gnd cell_6t
Xbit_r91_c74 bl[74] br[74] wl[91] vdd gnd cell_6t
Xbit_r92_c74 bl[74] br[74] wl[92] vdd gnd cell_6t
Xbit_r93_c74 bl[74] br[74] wl[93] vdd gnd cell_6t
Xbit_r94_c74 bl[74] br[74] wl[94] vdd gnd cell_6t
Xbit_r95_c74 bl[74] br[74] wl[95] vdd gnd cell_6t
Xbit_r96_c74 bl[74] br[74] wl[96] vdd gnd cell_6t
Xbit_r97_c74 bl[74] br[74] wl[97] vdd gnd cell_6t
Xbit_r98_c74 bl[74] br[74] wl[98] vdd gnd cell_6t
Xbit_r99_c74 bl[74] br[74] wl[99] vdd gnd cell_6t
Xbit_r100_c74 bl[74] br[74] wl[100] vdd gnd cell_6t
Xbit_r101_c74 bl[74] br[74] wl[101] vdd gnd cell_6t
Xbit_r102_c74 bl[74] br[74] wl[102] vdd gnd cell_6t
Xbit_r103_c74 bl[74] br[74] wl[103] vdd gnd cell_6t
Xbit_r104_c74 bl[74] br[74] wl[104] vdd gnd cell_6t
Xbit_r105_c74 bl[74] br[74] wl[105] vdd gnd cell_6t
Xbit_r106_c74 bl[74] br[74] wl[106] vdd gnd cell_6t
Xbit_r107_c74 bl[74] br[74] wl[107] vdd gnd cell_6t
Xbit_r108_c74 bl[74] br[74] wl[108] vdd gnd cell_6t
Xbit_r109_c74 bl[74] br[74] wl[109] vdd gnd cell_6t
Xbit_r110_c74 bl[74] br[74] wl[110] vdd gnd cell_6t
Xbit_r111_c74 bl[74] br[74] wl[111] vdd gnd cell_6t
Xbit_r112_c74 bl[74] br[74] wl[112] vdd gnd cell_6t
Xbit_r113_c74 bl[74] br[74] wl[113] vdd gnd cell_6t
Xbit_r114_c74 bl[74] br[74] wl[114] vdd gnd cell_6t
Xbit_r115_c74 bl[74] br[74] wl[115] vdd gnd cell_6t
Xbit_r116_c74 bl[74] br[74] wl[116] vdd gnd cell_6t
Xbit_r117_c74 bl[74] br[74] wl[117] vdd gnd cell_6t
Xbit_r118_c74 bl[74] br[74] wl[118] vdd gnd cell_6t
Xbit_r119_c74 bl[74] br[74] wl[119] vdd gnd cell_6t
Xbit_r120_c74 bl[74] br[74] wl[120] vdd gnd cell_6t
Xbit_r121_c74 bl[74] br[74] wl[121] vdd gnd cell_6t
Xbit_r122_c74 bl[74] br[74] wl[122] vdd gnd cell_6t
Xbit_r123_c74 bl[74] br[74] wl[123] vdd gnd cell_6t
Xbit_r124_c74 bl[74] br[74] wl[124] vdd gnd cell_6t
Xbit_r125_c74 bl[74] br[74] wl[125] vdd gnd cell_6t
Xbit_r126_c74 bl[74] br[74] wl[126] vdd gnd cell_6t
Xbit_r127_c74 bl[74] br[74] wl[127] vdd gnd cell_6t
Xbit_r128_c74 bl[74] br[74] wl[128] vdd gnd cell_6t
Xbit_r129_c74 bl[74] br[74] wl[129] vdd gnd cell_6t
Xbit_r130_c74 bl[74] br[74] wl[130] vdd gnd cell_6t
Xbit_r131_c74 bl[74] br[74] wl[131] vdd gnd cell_6t
Xbit_r132_c74 bl[74] br[74] wl[132] vdd gnd cell_6t
Xbit_r133_c74 bl[74] br[74] wl[133] vdd gnd cell_6t
Xbit_r134_c74 bl[74] br[74] wl[134] vdd gnd cell_6t
Xbit_r135_c74 bl[74] br[74] wl[135] vdd gnd cell_6t
Xbit_r136_c74 bl[74] br[74] wl[136] vdd gnd cell_6t
Xbit_r137_c74 bl[74] br[74] wl[137] vdd gnd cell_6t
Xbit_r138_c74 bl[74] br[74] wl[138] vdd gnd cell_6t
Xbit_r139_c74 bl[74] br[74] wl[139] vdd gnd cell_6t
Xbit_r140_c74 bl[74] br[74] wl[140] vdd gnd cell_6t
Xbit_r141_c74 bl[74] br[74] wl[141] vdd gnd cell_6t
Xbit_r142_c74 bl[74] br[74] wl[142] vdd gnd cell_6t
Xbit_r143_c74 bl[74] br[74] wl[143] vdd gnd cell_6t
Xbit_r144_c74 bl[74] br[74] wl[144] vdd gnd cell_6t
Xbit_r145_c74 bl[74] br[74] wl[145] vdd gnd cell_6t
Xbit_r146_c74 bl[74] br[74] wl[146] vdd gnd cell_6t
Xbit_r147_c74 bl[74] br[74] wl[147] vdd gnd cell_6t
Xbit_r148_c74 bl[74] br[74] wl[148] vdd gnd cell_6t
Xbit_r149_c74 bl[74] br[74] wl[149] vdd gnd cell_6t
Xbit_r150_c74 bl[74] br[74] wl[150] vdd gnd cell_6t
Xbit_r151_c74 bl[74] br[74] wl[151] vdd gnd cell_6t
Xbit_r152_c74 bl[74] br[74] wl[152] vdd gnd cell_6t
Xbit_r153_c74 bl[74] br[74] wl[153] vdd gnd cell_6t
Xbit_r154_c74 bl[74] br[74] wl[154] vdd gnd cell_6t
Xbit_r155_c74 bl[74] br[74] wl[155] vdd gnd cell_6t
Xbit_r156_c74 bl[74] br[74] wl[156] vdd gnd cell_6t
Xbit_r157_c74 bl[74] br[74] wl[157] vdd gnd cell_6t
Xbit_r158_c74 bl[74] br[74] wl[158] vdd gnd cell_6t
Xbit_r159_c74 bl[74] br[74] wl[159] vdd gnd cell_6t
Xbit_r160_c74 bl[74] br[74] wl[160] vdd gnd cell_6t
Xbit_r161_c74 bl[74] br[74] wl[161] vdd gnd cell_6t
Xbit_r162_c74 bl[74] br[74] wl[162] vdd gnd cell_6t
Xbit_r163_c74 bl[74] br[74] wl[163] vdd gnd cell_6t
Xbit_r164_c74 bl[74] br[74] wl[164] vdd gnd cell_6t
Xbit_r165_c74 bl[74] br[74] wl[165] vdd gnd cell_6t
Xbit_r166_c74 bl[74] br[74] wl[166] vdd gnd cell_6t
Xbit_r167_c74 bl[74] br[74] wl[167] vdd gnd cell_6t
Xbit_r168_c74 bl[74] br[74] wl[168] vdd gnd cell_6t
Xbit_r169_c74 bl[74] br[74] wl[169] vdd gnd cell_6t
Xbit_r170_c74 bl[74] br[74] wl[170] vdd gnd cell_6t
Xbit_r171_c74 bl[74] br[74] wl[171] vdd gnd cell_6t
Xbit_r172_c74 bl[74] br[74] wl[172] vdd gnd cell_6t
Xbit_r173_c74 bl[74] br[74] wl[173] vdd gnd cell_6t
Xbit_r174_c74 bl[74] br[74] wl[174] vdd gnd cell_6t
Xbit_r175_c74 bl[74] br[74] wl[175] vdd gnd cell_6t
Xbit_r176_c74 bl[74] br[74] wl[176] vdd gnd cell_6t
Xbit_r177_c74 bl[74] br[74] wl[177] vdd gnd cell_6t
Xbit_r178_c74 bl[74] br[74] wl[178] vdd gnd cell_6t
Xbit_r179_c74 bl[74] br[74] wl[179] vdd gnd cell_6t
Xbit_r180_c74 bl[74] br[74] wl[180] vdd gnd cell_6t
Xbit_r181_c74 bl[74] br[74] wl[181] vdd gnd cell_6t
Xbit_r182_c74 bl[74] br[74] wl[182] vdd gnd cell_6t
Xbit_r183_c74 bl[74] br[74] wl[183] vdd gnd cell_6t
Xbit_r184_c74 bl[74] br[74] wl[184] vdd gnd cell_6t
Xbit_r185_c74 bl[74] br[74] wl[185] vdd gnd cell_6t
Xbit_r186_c74 bl[74] br[74] wl[186] vdd gnd cell_6t
Xbit_r187_c74 bl[74] br[74] wl[187] vdd gnd cell_6t
Xbit_r188_c74 bl[74] br[74] wl[188] vdd gnd cell_6t
Xbit_r189_c74 bl[74] br[74] wl[189] vdd gnd cell_6t
Xbit_r190_c74 bl[74] br[74] wl[190] vdd gnd cell_6t
Xbit_r191_c74 bl[74] br[74] wl[191] vdd gnd cell_6t
Xbit_r192_c74 bl[74] br[74] wl[192] vdd gnd cell_6t
Xbit_r193_c74 bl[74] br[74] wl[193] vdd gnd cell_6t
Xbit_r194_c74 bl[74] br[74] wl[194] vdd gnd cell_6t
Xbit_r195_c74 bl[74] br[74] wl[195] vdd gnd cell_6t
Xbit_r196_c74 bl[74] br[74] wl[196] vdd gnd cell_6t
Xbit_r197_c74 bl[74] br[74] wl[197] vdd gnd cell_6t
Xbit_r198_c74 bl[74] br[74] wl[198] vdd gnd cell_6t
Xbit_r199_c74 bl[74] br[74] wl[199] vdd gnd cell_6t
Xbit_r200_c74 bl[74] br[74] wl[200] vdd gnd cell_6t
Xbit_r201_c74 bl[74] br[74] wl[201] vdd gnd cell_6t
Xbit_r202_c74 bl[74] br[74] wl[202] vdd gnd cell_6t
Xbit_r203_c74 bl[74] br[74] wl[203] vdd gnd cell_6t
Xbit_r204_c74 bl[74] br[74] wl[204] vdd gnd cell_6t
Xbit_r205_c74 bl[74] br[74] wl[205] vdd gnd cell_6t
Xbit_r206_c74 bl[74] br[74] wl[206] vdd gnd cell_6t
Xbit_r207_c74 bl[74] br[74] wl[207] vdd gnd cell_6t
Xbit_r208_c74 bl[74] br[74] wl[208] vdd gnd cell_6t
Xbit_r209_c74 bl[74] br[74] wl[209] vdd gnd cell_6t
Xbit_r210_c74 bl[74] br[74] wl[210] vdd gnd cell_6t
Xbit_r211_c74 bl[74] br[74] wl[211] vdd gnd cell_6t
Xbit_r212_c74 bl[74] br[74] wl[212] vdd gnd cell_6t
Xbit_r213_c74 bl[74] br[74] wl[213] vdd gnd cell_6t
Xbit_r214_c74 bl[74] br[74] wl[214] vdd gnd cell_6t
Xbit_r215_c74 bl[74] br[74] wl[215] vdd gnd cell_6t
Xbit_r216_c74 bl[74] br[74] wl[216] vdd gnd cell_6t
Xbit_r217_c74 bl[74] br[74] wl[217] vdd gnd cell_6t
Xbit_r218_c74 bl[74] br[74] wl[218] vdd gnd cell_6t
Xbit_r219_c74 bl[74] br[74] wl[219] vdd gnd cell_6t
Xbit_r220_c74 bl[74] br[74] wl[220] vdd gnd cell_6t
Xbit_r221_c74 bl[74] br[74] wl[221] vdd gnd cell_6t
Xbit_r222_c74 bl[74] br[74] wl[222] vdd gnd cell_6t
Xbit_r223_c74 bl[74] br[74] wl[223] vdd gnd cell_6t
Xbit_r224_c74 bl[74] br[74] wl[224] vdd gnd cell_6t
Xbit_r225_c74 bl[74] br[74] wl[225] vdd gnd cell_6t
Xbit_r226_c74 bl[74] br[74] wl[226] vdd gnd cell_6t
Xbit_r227_c74 bl[74] br[74] wl[227] vdd gnd cell_6t
Xbit_r228_c74 bl[74] br[74] wl[228] vdd gnd cell_6t
Xbit_r229_c74 bl[74] br[74] wl[229] vdd gnd cell_6t
Xbit_r230_c74 bl[74] br[74] wl[230] vdd gnd cell_6t
Xbit_r231_c74 bl[74] br[74] wl[231] vdd gnd cell_6t
Xbit_r232_c74 bl[74] br[74] wl[232] vdd gnd cell_6t
Xbit_r233_c74 bl[74] br[74] wl[233] vdd gnd cell_6t
Xbit_r234_c74 bl[74] br[74] wl[234] vdd gnd cell_6t
Xbit_r235_c74 bl[74] br[74] wl[235] vdd gnd cell_6t
Xbit_r236_c74 bl[74] br[74] wl[236] vdd gnd cell_6t
Xbit_r237_c74 bl[74] br[74] wl[237] vdd gnd cell_6t
Xbit_r238_c74 bl[74] br[74] wl[238] vdd gnd cell_6t
Xbit_r239_c74 bl[74] br[74] wl[239] vdd gnd cell_6t
Xbit_r240_c74 bl[74] br[74] wl[240] vdd gnd cell_6t
Xbit_r241_c74 bl[74] br[74] wl[241] vdd gnd cell_6t
Xbit_r242_c74 bl[74] br[74] wl[242] vdd gnd cell_6t
Xbit_r243_c74 bl[74] br[74] wl[243] vdd gnd cell_6t
Xbit_r244_c74 bl[74] br[74] wl[244] vdd gnd cell_6t
Xbit_r245_c74 bl[74] br[74] wl[245] vdd gnd cell_6t
Xbit_r246_c74 bl[74] br[74] wl[246] vdd gnd cell_6t
Xbit_r247_c74 bl[74] br[74] wl[247] vdd gnd cell_6t
Xbit_r248_c74 bl[74] br[74] wl[248] vdd gnd cell_6t
Xbit_r249_c74 bl[74] br[74] wl[249] vdd gnd cell_6t
Xbit_r250_c74 bl[74] br[74] wl[250] vdd gnd cell_6t
Xbit_r251_c74 bl[74] br[74] wl[251] vdd gnd cell_6t
Xbit_r252_c74 bl[74] br[74] wl[252] vdd gnd cell_6t
Xbit_r253_c74 bl[74] br[74] wl[253] vdd gnd cell_6t
Xbit_r254_c74 bl[74] br[74] wl[254] vdd gnd cell_6t
Xbit_r255_c74 bl[74] br[74] wl[255] vdd gnd cell_6t
Xbit_r0_c75 bl[75] br[75] wl[0] vdd gnd cell_6t
Xbit_r1_c75 bl[75] br[75] wl[1] vdd gnd cell_6t
Xbit_r2_c75 bl[75] br[75] wl[2] vdd gnd cell_6t
Xbit_r3_c75 bl[75] br[75] wl[3] vdd gnd cell_6t
Xbit_r4_c75 bl[75] br[75] wl[4] vdd gnd cell_6t
Xbit_r5_c75 bl[75] br[75] wl[5] vdd gnd cell_6t
Xbit_r6_c75 bl[75] br[75] wl[6] vdd gnd cell_6t
Xbit_r7_c75 bl[75] br[75] wl[7] vdd gnd cell_6t
Xbit_r8_c75 bl[75] br[75] wl[8] vdd gnd cell_6t
Xbit_r9_c75 bl[75] br[75] wl[9] vdd gnd cell_6t
Xbit_r10_c75 bl[75] br[75] wl[10] vdd gnd cell_6t
Xbit_r11_c75 bl[75] br[75] wl[11] vdd gnd cell_6t
Xbit_r12_c75 bl[75] br[75] wl[12] vdd gnd cell_6t
Xbit_r13_c75 bl[75] br[75] wl[13] vdd gnd cell_6t
Xbit_r14_c75 bl[75] br[75] wl[14] vdd gnd cell_6t
Xbit_r15_c75 bl[75] br[75] wl[15] vdd gnd cell_6t
Xbit_r16_c75 bl[75] br[75] wl[16] vdd gnd cell_6t
Xbit_r17_c75 bl[75] br[75] wl[17] vdd gnd cell_6t
Xbit_r18_c75 bl[75] br[75] wl[18] vdd gnd cell_6t
Xbit_r19_c75 bl[75] br[75] wl[19] vdd gnd cell_6t
Xbit_r20_c75 bl[75] br[75] wl[20] vdd gnd cell_6t
Xbit_r21_c75 bl[75] br[75] wl[21] vdd gnd cell_6t
Xbit_r22_c75 bl[75] br[75] wl[22] vdd gnd cell_6t
Xbit_r23_c75 bl[75] br[75] wl[23] vdd gnd cell_6t
Xbit_r24_c75 bl[75] br[75] wl[24] vdd gnd cell_6t
Xbit_r25_c75 bl[75] br[75] wl[25] vdd gnd cell_6t
Xbit_r26_c75 bl[75] br[75] wl[26] vdd gnd cell_6t
Xbit_r27_c75 bl[75] br[75] wl[27] vdd gnd cell_6t
Xbit_r28_c75 bl[75] br[75] wl[28] vdd gnd cell_6t
Xbit_r29_c75 bl[75] br[75] wl[29] vdd gnd cell_6t
Xbit_r30_c75 bl[75] br[75] wl[30] vdd gnd cell_6t
Xbit_r31_c75 bl[75] br[75] wl[31] vdd gnd cell_6t
Xbit_r32_c75 bl[75] br[75] wl[32] vdd gnd cell_6t
Xbit_r33_c75 bl[75] br[75] wl[33] vdd gnd cell_6t
Xbit_r34_c75 bl[75] br[75] wl[34] vdd gnd cell_6t
Xbit_r35_c75 bl[75] br[75] wl[35] vdd gnd cell_6t
Xbit_r36_c75 bl[75] br[75] wl[36] vdd gnd cell_6t
Xbit_r37_c75 bl[75] br[75] wl[37] vdd gnd cell_6t
Xbit_r38_c75 bl[75] br[75] wl[38] vdd gnd cell_6t
Xbit_r39_c75 bl[75] br[75] wl[39] vdd gnd cell_6t
Xbit_r40_c75 bl[75] br[75] wl[40] vdd gnd cell_6t
Xbit_r41_c75 bl[75] br[75] wl[41] vdd gnd cell_6t
Xbit_r42_c75 bl[75] br[75] wl[42] vdd gnd cell_6t
Xbit_r43_c75 bl[75] br[75] wl[43] vdd gnd cell_6t
Xbit_r44_c75 bl[75] br[75] wl[44] vdd gnd cell_6t
Xbit_r45_c75 bl[75] br[75] wl[45] vdd gnd cell_6t
Xbit_r46_c75 bl[75] br[75] wl[46] vdd gnd cell_6t
Xbit_r47_c75 bl[75] br[75] wl[47] vdd gnd cell_6t
Xbit_r48_c75 bl[75] br[75] wl[48] vdd gnd cell_6t
Xbit_r49_c75 bl[75] br[75] wl[49] vdd gnd cell_6t
Xbit_r50_c75 bl[75] br[75] wl[50] vdd gnd cell_6t
Xbit_r51_c75 bl[75] br[75] wl[51] vdd gnd cell_6t
Xbit_r52_c75 bl[75] br[75] wl[52] vdd gnd cell_6t
Xbit_r53_c75 bl[75] br[75] wl[53] vdd gnd cell_6t
Xbit_r54_c75 bl[75] br[75] wl[54] vdd gnd cell_6t
Xbit_r55_c75 bl[75] br[75] wl[55] vdd gnd cell_6t
Xbit_r56_c75 bl[75] br[75] wl[56] vdd gnd cell_6t
Xbit_r57_c75 bl[75] br[75] wl[57] vdd gnd cell_6t
Xbit_r58_c75 bl[75] br[75] wl[58] vdd gnd cell_6t
Xbit_r59_c75 bl[75] br[75] wl[59] vdd gnd cell_6t
Xbit_r60_c75 bl[75] br[75] wl[60] vdd gnd cell_6t
Xbit_r61_c75 bl[75] br[75] wl[61] vdd gnd cell_6t
Xbit_r62_c75 bl[75] br[75] wl[62] vdd gnd cell_6t
Xbit_r63_c75 bl[75] br[75] wl[63] vdd gnd cell_6t
Xbit_r64_c75 bl[75] br[75] wl[64] vdd gnd cell_6t
Xbit_r65_c75 bl[75] br[75] wl[65] vdd gnd cell_6t
Xbit_r66_c75 bl[75] br[75] wl[66] vdd gnd cell_6t
Xbit_r67_c75 bl[75] br[75] wl[67] vdd gnd cell_6t
Xbit_r68_c75 bl[75] br[75] wl[68] vdd gnd cell_6t
Xbit_r69_c75 bl[75] br[75] wl[69] vdd gnd cell_6t
Xbit_r70_c75 bl[75] br[75] wl[70] vdd gnd cell_6t
Xbit_r71_c75 bl[75] br[75] wl[71] vdd gnd cell_6t
Xbit_r72_c75 bl[75] br[75] wl[72] vdd gnd cell_6t
Xbit_r73_c75 bl[75] br[75] wl[73] vdd gnd cell_6t
Xbit_r74_c75 bl[75] br[75] wl[74] vdd gnd cell_6t
Xbit_r75_c75 bl[75] br[75] wl[75] vdd gnd cell_6t
Xbit_r76_c75 bl[75] br[75] wl[76] vdd gnd cell_6t
Xbit_r77_c75 bl[75] br[75] wl[77] vdd gnd cell_6t
Xbit_r78_c75 bl[75] br[75] wl[78] vdd gnd cell_6t
Xbit_r79_c75 bl[75] br[75] wl[79] vdd gnd cell_6t
Xbit_r80_c75 bl[75] br[75] wl[80] vdd gnd cell_6t
Xbit_r81_c75 bl[75] br[75] wl[81] vdd gnd cell_6t
Xbit_r82_c75 bl[75] br[75] wl[82] vdd gnd cell_6t
Xbit_r83_c75 bl[75] br[75] wl[83] vdd gnd cell_6t
Xbit_r84_c75 bl[75] br[75] wl[84] vdd gnd cell_6t
Xbit_r85_c75 bl[75] br[75] wl[85] vdd gnd cell_6t
Xbit_r86_c75 bl[75] br[75] wl[86] vdd gnd cell_6t
Xbit_r87_c75 bl[75] br[75] wl[87] vdd gnd cell_6t
Xbit_r88_c75 bl[75] br[75] wl[88] vdd gnd cell_6t
Xbit_r89_c75 bl[75] br[75] wl[89] vdd gnd cell_6t
Xbit_r90_c75 bl[75] br[75] wl[90] vdd gnd cell_6t
Xbit_r91_c75 bl[75] br[75] wl[91] vdd gnd cell_6t
Xbit_r92_c75 bl[75] br[75] wl[92] vdd gnd cell_6t
Xbit_r93_c75 bl[75] br[75] wl[93] vdd gnd cell_6t
Xbit_r94_c75 bl[75] br[75] wl[94] vdd gnd cell_6t
Xbit_r95_c75 bl[75] br[75] wl[95] vdd gnd cell_6t
Xbit_r96_c75 bl[75] br[75] wl[96] vdd gnd cell_6t
Xbit_r97_c75 bl[75] br[75] wl[97] vdd gnd cell_6t
Xbit_r98_c75 bl[75] br[75] wl[98] vdd gnd cell_6t
Xbit_r99_c75 bl[75] br[75] wl[99] vdd gnd cell_6t
Xbit_r100_c75 bl[75] br[75] wl[100] vdd gnd cell_6t
Xbit_r101_c75 bl[75] br[75] wl[101] vdd gnd cell_6t
Xbit_r102_c75 bl[75] br[75] wl[102] vdd gnd cell_6t
Xbit_r103_c75 bl[75] br[75] wl[103] vdd gnd cell_6t
Xbit_r104_c75 bl[75] br[75] wl[104] vdd gnd cell_6t
Xbit_r105_c75 bl[75] br[75] wl[105] vdd gnd cell_6t
Xbit_r106_c75 bl[75] br[75] wl[106] vdd gnd cell_6t
Xbit_r107_c75 bl[75] br[75] wl[107] vdd gnd cell_6t
Xbit_r108_c75 bl[75] br[75] wl[108] vdd gnd cell_6t
Xbit_r109_c75 bl[75] br[75] wl[109] vdd gnd cell_6t
Xbit_r110_c75 bl[75] br[75] wl[110] vdd gnd cell_6t
Xbit_r111_c75 bl[75] br[75] wl[111] vdd gnd cell_6t
Xbit_r112_c75 bl[75] br[75] wl[112] vdd gnd cell_6t
Xbit_r113_c75 bl[75] br[75] wl[113] vdd gnd cell_6t
Xbit_r114_c75 bl[75] br[75] wl[114] vdd gnd cell_6t
Xbit_r115_c75 bl[75] br[75] wl[115] vdd gnd cell_6t
Xbit_r116_c75 bl[75] br[75] wl[116] vdd gnd cell_6t
Xbit_r117_c75 bl[75] br[75] wl[117] vdd gnd cell_6t
Xbit_r118_c75 bl[75] br[75] wl[118] vdd gnd cell_6t
Xbit_r119_c75 bl[75] br[75] wl[119] vdd gnd cell_6t
Xbit_r120_c75 bl[75] br[75] wl[120] vdd gnd cell_6t
Xbit_r121_c75 bl[75] br[75] wl[121] vdd gnd cell_6t
Xbit_r122_c75 bl[75] br[75] wl[122] vdd gnd cell_6t
Xbit_r123_c75 bl[75] br[75] wl[123] vdd gnd cell_6t
Xbit_r124_c75 bl[75] br[75] wl[124] vdd gnd cell_6t
Xbit_r125_c75 bl[75] br[75] wl[125] vdd gnd cell_6t
Xbit_r126_c75 bl[75] br[75] wl[126] vdd gnd cell_6t
Xbit_r127_c75 bl[75] br[75] wl[127] vdd gnd cell_6t
Xbit_r128_c75 bl[75] br[75] wl[128] vdd gnd cell_6t
Xbit_r129_c75 bl[75] br[75] wl[129] vdd gnd cell_6t
Xbit_r130_c75 bl[75] br[75] wl[130] vdd gnd cell_6t
Xbit_r131_c75 bl[75] br[75] wl[131] vdd gnd cell_6t
Xbit_r132_c75 bl[75] br[75] wl[132] vdd gnd cell_6t
Xbit_r133_c75 bl[75] br[75] wl[133] vdd gnd cell_6t
Xbit_r134_c75 bl[75] br[75] wl[134] vdd gnd cell_6t
Xbit_r135_c75 bl[75] br[75] wl[135] vdd gnd cell_6t
Xbit_r136_c75 bl[75] br[75] wl[136] vdd gnd cell_6t
Xbit_r137_c75 bl[75] br[75] wl[137] vdd gnd cell_6t
Xbit_r138_c75 bl[75] br[75] wl[138] vdd gnd cell_6t
Xbit_r139_c75 bl[75] br[75] wl[139] vdd gnd cell_6t
Xbit_r140_c75 bl[75] br[75] wl[140] vdd gnd cell_6t
Xbit_r141_c75 bl[75] br[75] wl[141] vdd gnd cell_6t
Xbit_r142_c75 bl[75] br[75] wl[142] vdd gnd cell_6t
Xbit_r143_c75 bl[75] br[75] wl[143] vdd gnd cell_6t
Xbit_r144_c75 bl[75] br[75] wl[144] vdd gnd cell_6t
Xbit_r145_c75 bl[75] br[75] wl[145] vdd gnd cell_6t
Xbit_r146_c75 bl[75] br[75] wl[146] vdd gnd cell_6t
Xbit_r147_c75 bl[75] br[75] wl[147] vdd gnd cell_6t
Xbit_r148_c75 bl[75] br[75] wl[148] vdd gnd cell_6t
Xbit_r149_c75 bl[75] br[75] wl[149] vdd gnd cell_6t
Xbit_r150_c75 bl[75] br[75] wl[150] vdd gnd cell_6t
Xbit_r151_c75 bl[75] br[75] wl[151] vdd gnd cell_6t
Xbit_r152_c75 bl[75] br[75] wl[152] vdd gnd cell_6t
Xbit_r153_c75 bl[75] br[75] wl[153] vdd gnd cell_6t
Xbit_r154_c75 bl[75] br[75] wl[154] vdd gnd cell_6t
Xbit_r155_c75 bl[75] br[75] wl[155] vdd gnd cell_6t
Xbit_r156_c75 bl[75] br[75] wl[156] vdd gnd cell_6t
Xbit_r157_c75 bl[75] br[75] wl[157] vdd gnd cell_6t
Xbit_r158_c75 bl[75] br[75] wl[158] vdd gnd cell_6t
Xbit_r159_c75 bl[75] br[75] wl[159] vdd gnd cell_6t
Xbit_r160_c75 bl[75] br[75] wl[160] vdd gnd cell_6t
Xbit_r161_c75 bl[75] br[75] wl[161] vdd gnd cell_6t
Xbit_r162_c75 bl[75] br[75] wl[162] vdd gnd cell_6t
Xbit_r163_c75 bl[75] br[75] wl[163] vdd gnd cell_6t
Xbit_r164_c75 bl[75] br[75] wl[164] vdd gnd cell_6t
Xbit_r165_c75 bl[75] br[75] wl[165] vdd gnd cell_6t
Xbit_r166_c75 bl[75] br[75] wl[166] vdd gnd cell_6t
Xbit_r167_c75 bl[75] br[75] wl[167] vdd gnd cell_6t
Xbit_r168_c75 bl[75] br[75] wl[168] vdd gnd cell_6t
Xbit_r169_c75 bl[75] br[75] wl[169] vdd gnd cell_6t
Xbit_r170_c75 bl[75] br[75] wl[170] vdd gnd cell_6t
Xbit_r171_c75 bl[75] br[75] wl[171] vdd gnd cell_6t
Xbit_r172_c75 bl[75] br[75] wl[172] vdd gnd cell_6t
Xbit_r173_c75 bl[75] br[75] wl[173] vdd gnd cell_6t
Xbit_r174_c75 bl[75] br[75] wl[174] vdd gnd cell_6t
Xbit_r175_c75 bl[75] br[75] wl[175] vdd gnd cell_6t
Xbit_r176_c75 bl[75] br[75] wl[176] vdd gnd cell_6t
Xbit_r177_c75 bl[75] br[75] wl[177] vdd gnd cell_6t
Xbit_r178_c75 bl[75] br[75] wl[178] vdd gnd cell_6t
Xbit_r179_c75 bl[75] br[75] wl[179] vdd gnd cell_6t
Xbit_r180_c75 bl[75] br[75] wl[180] vdd gnd cell_6t
Xbit_r181_c75 bl[75] br[75] wl[181] vdd gnd cell_6t
Xbit_r182_c75 bl[75] br[75] wl[182] vdd gnd cell_6t
Xbit_r183_c75 bl[75] br[75] wl[183] vdd gnd cell_6t
Xbit_r184_c75 bl[75] br[75] wl[184] vdd gnd cell_6t
Xbit_r185_c75 bl[75] br[75] wl[185] vdd gnd cell_6t
Xbit_r186_c75 bl[75] br[75] wl[186] vdd gnd cell_6t
Xbit_r187_c75 bl[75] br[75] wl[187] vdd gnd cell_6t
Xbit_r188_c75 bl[75] br[75] wl[188] vdd gnd cell_6t
Xbit_r189_c75 bl[75] br[75] wl[189] vdd gnd cell_6t
Xbit_r190_c75 bl[75] br[75] wl[190] vdd gnd cell_6t
Xbit_r191_c75 bl[75] br[75] wl[191] vdd gnd cell_6t
Xbit_r192_c75 bl[75] br[75] wl[192] vdd gnd cell_6t
Xbit_r193_c75 bl[75] br[75] wl[193] vdd gnd cell_6t
Xbit_r194_c75 bl[75] br[75] wl[194] vdd gnd cell_6t
Xbit_r195_c75 bl[75] br[75] wl[195] vdd gnd cell_6t
Xbit_r196_c75 bl[75] br[75] wl[196] vdd gnd cell_6t
Xbit_r197_c75 bl[75] br[75] wl[197] vdd gnd cell_6t
Xbit_r198_c75 bl[75] br[75] wl[198] vdd gnd cell_6t
Xbit_r199_c75 bl[75] br[75] wl[199] vdd gnd cell_6t
Xbit_r200_c75 bl[75] br[75] wl[200] vdd gnd cell_6t
Xbit_r201_c75 bl[75] br[75] wl[201] vdd gnd cell_6t
Xbit_r202_c75 bl[75] br[75] wl[202] vdd gnd cell_6t
Xbit_r203_c75 bl[75] br[75] wl[203] vdd gnd cell_6t
Xbit_r204_c75 bl[75] br[75] wl[204] vdd gnd cell_6t
Xbit_r205_c75 bl[75] br[75] wl[205] vdd gnd cell_6t
Xbit_r206_c75 bl[75] br[75] wl[206] vdd gnd cell_6t
Xbit_r207_c75 bl[75] br[75] wl[207] vdd gnd cell_6t
Xbit_r208_c75 bl[75] br[75] wl[208] vdd gnd cell_6t
Xbit_r209_c75 bl[75] br[75] wl[209] vdd gnd cell_6t
Xbit_r210_c75 bl[75] br[75] wl[210] vdd gnd cell_6t
Xbit_r211_c75 bl[75] br[75] wl[211] vdd gnd cell_6t
Xbit_r212_c75 bl[75] br[75] wl[212] vdd gnd cell_6t
Xbit_r213_c75 bl[75] br[75] wl[213] vdd gnd cell_6t
Xbit_r214_c75 bl[75] br[75] wl[214] vdd gnd cell_6t
Xbit_r215_c75 bl[75] br[75] wl[215] vdd gnd cell_6t
Xbit_r216_c75 bl[75] br[75] wl[216] vdd gnd cell_6t
Xbit_r217_c75 bl[75] br[75] wl[217] vdd gnd cell_6t
Xbit_r218_c75 bl[75] br[75] wl[218] vdd gnd cell_6t
Xbit_r219_c75 bl[75] br[75] wl[219] vdd gnd cell_6t
Xbit_r220_c75 bl[75] br[75] wl[220] vdd gnd cell_6t
Xbit_r221_c75 bl[75] br[75] wl[221] vdd gnd cell_6t
Xbit_r222_c75 bl[75] br[75] wl[222] vdd gnd cell_6t
Xbit_r223_c75 bl[75] br[75] wl[223] vdd gnd cell_6t
Xbit_r224_c75 bl[75] br[75] wl[224] vdd gnd cell_6t
Xbit_r225_c75 bl[75] br[75] wl[225] vdd gnd cell_6t
Xbit_r226_c75 bl[75] br[75] wl[226] vdd gnd cell_6t
Xbit_r227_c75 bl[75] br[75] wl[227] vdd gnd cell_6t
Xbit_r228_c75 bl[75] br[75] wl[228] vdd gnd cell_6t
Xbit_r229_c75 bl[75] br[75] wl[229] vdd gnd cell_6t
Xbit_r230_c75 bl[75] br[75] wl[230] vdd gnd cell_6t
Xbit_r231_c75 bl[75] br[75] wl[231] vdd gnd cell_6t
Xbit_r232_c75 bl[75] br[75] wl[232] vdd gnd cell_6t
Xbit_r233_c75 bl[75] br[75] wl[233] vdd gnd cell_6t
Xbit_r234_c75 bl[75] br[75] wl[234] vdd gnd cell_6t
Xbit_r235_c75 bl[75] br[75] wl[235] vdd gnd cell_6t
Xbit_r236_c75 bl[75] br[75] wl[236] vdd gnd cell_6t
Xbit_r237_c75 bl[75] br[75] wl[237] vdd gnd cell_6t
Xbit_r238_c75 bl[75] br[75] wl[238] vdd gnd cell_6t
Xbit_r239_c75 bl[75] br[75] wl[239] vdd gnd cell_6t
Xbit_r240_c75 bl[75] br[75] wl[240] vdd gnd cell_6t
Xbit_r241_c75 bl[75] br[75] wl[241] vdd gnd cell_6t
Xbit_r242_c75 bl[75] br[75] wl[242] vdd gnd cell_6t
Xbit_r243_c75 bl[75] br[75] wl[243] vdd gnd cell_6t
Xbit_r244_c75 bl[75] br[75] wl[244] vdd gnd cell_6t
Xbit_r245_c75 bl[75] br[75] wl[245] vdd gnd cell_6t
Xbit_r246_c75 bl[75] br[75] wl[246] vdd gnd cell_6t
Xbit_r247_c75 bl[75] br[75] wl[247] vdd gnd cell_6t
Xbit_r248_c75 bl[75] br[75] wl[248] vdd gnd cell_6t
Xbit_r249_c75 bl[75] br[75] wl[249] vdd gnd cell_6t
Xbit_r250_c75 bl[75] br[75] wl[250] vdd gnd cell_6t
Xbit_r251_c75 bl[75] br[75] wl[251] vdd gnd cell_6t
Xbit_r252_c75 bl[75] br[75] wl[252] vdd gnd cell_6t
Xbit_r253_c75 bl[75] br[75] wl[253] vdd gnd cell_6t
Xbit_r254_c75 bl[75] br[75] wl[254] vdd gnd cell_6t
Xbit_r255_c75 bl[75] br[75] wl[255] vdd gnd cell_6t
Xbit_r0_c76 bl[76] br[76] wl[0] vdd gnd cell_6t
Xbit_r1_c76 bl[76] br[76] wl[1] vdd gnd cell_6t
Xbit_r2_c76 bl[76] br[76] wl[2] vdd gnd cell_6t
Xbit_r3_c76 bl[76] br[76] wl[3] vdd gnd cell_6t
Xbit_r4_c76 bl[76] br[76] wl[4] vdd gnd cell_6t
Xbit_r5_c76 bl[76] br[76] wl[5] vdd gnd cell_6t
Xbit_r6_c76 bl[76] br[76] wl[6] vdd gnd cell_6t
Xbit_r7_c76 bl[76] br[76] wl[7] vdd gnd cell_6t
Xbit_r8_c76 bl[76] br[76] wl[8] vdd gnd cell_6t
Xbit_r9_c76 bl[76] br[76] wl[9] vdd gnd cell_6t
Xbit_r10_c76 bl[76] br[76] wl[10] vdd gnd cell_6t
Xbit_r11_c76 bl[76] br[76] wl[11] vdd gnd cell_6t
Xbit_r12_c76 bl[76] br[76] wl[12] vdd gnd cell_6t
Xbit_r13_c76 bl[76] br[76] wl[13] vdd gnd cell_6t
Xbit_r14_c76 bl[76] br[76] wl[14] vdd gnd cell_6t
Xbit_r15_c76 bl[76] br[76] wl[15] vdd gnd cell_6t
Xbit_r16_c76 bl[76] br[76] wl[16] vdd gnd cell_6t
Xbit_r17_c76 bl[76] br[76] wl[17] vdd gnd cell_6t
Xbit_r18_c76 bl[76] br[76] wl[18] vdd gnd cell_6t
Xbit_r19_c76 bl[76] br[76] wl[19] vdd gnd cell_6t
Xbit_r20_c76 bl[76] br[76] wl[20] vdd gnd cell_6t
Xbit_r21_c76 bl[76] br[76] wl[21] vdd gnd cell_6t
Xbit_r22_c76 bl[76] br[76] wl[22] vdd gnd cell_6t
Xbit_r23_c76 bl[76] br[76] wl[23] vdd gnd cell_6t
Xbit_r24_c76 bl[76] br[76] wl[24] vdd gnd cell_6t
Xbit_r25_c76 bl[76] br[76] wl[25] vdd gnd cell_6t
Xbit_r26_c76 bl[76] br[76] wl[26] vdd gnd cell_6t
Xbit_r27_c76 bl[76] br[76] wl[27] vdd gnd cell_6t
Xbit_r28_c76 bl[76] br[76] wl[28] vdd gnd cell_6t
Xbit_r29_c76 bl[76] br[76] wl[29] vdd gnd cell_6t
Xbit_r30_c76 bl[76] br[76] wl[30] vdd gnd cell_6t
Xbit_r31_c76 bl[76] br[76] wl[31] vdd gnd cell_6t
Xbit_r32_c76 bl[76] br[76] wl[32] vdd gnd cell_6t
Xbit_r33_c76 bl[76] br[76] wl[33] vdd gnd cell_6t
Xbit_r34_c76 bl[76] br[76] wl[34] vdd gnd cell_6t
Xbit_r35_c76 bl[76] br[76] wl[35] vdd gnd cell_6t
Xbit_r36_c76 bl[76] br[76] wl[36] vdd gnd cell_6t
Xbit_r37_c76 bl[76] br[76] wl[37] vdd gnd cell_6t
Xbit_r38_c76 bl[76] br[76] wl[38] vdd gnd cell_6t
Xbit_r39_c76 bl[76] br[76] wl[39] vdd gnd cell_6t
Xbit_r40_c76 bl[76] br[76] wl[40] vdd gnd cell_6t
Xbit_r41_c76 bl[76] br[76] wl[41] vdd gnd cell_6t
Xbit_r42_c76 bl[76] br[76] wl[42] vdd gnd cell_6t
Xbit_r43_c76 bl[76] br[76] wl[43] vdd gnd cell_6t
Xbit_r44_c76 bl[76] br[76] wl[44] vdd gnd cell_6t
Xbit_r45_c76 bl[76] br[76] wl[45] vdd gnd cell_6t
Xbit_r46_c76 bl[76] br[76] wl[46] vdd gnd cell_6t
Xbit_r47_c76 bl[76] br[76] wl[47] vdd gnd cell_6t
Xbit_r48_c76 bl[76] br[76] wl[48] vdd gnd cell_6t
Xbit_r49_c76 bl[76] br[76] wl[49] vdd gnd cell_6t
Xbit_r50_c76 bl[76] br[76] wl[50] vdd gnd cell_6t
Xbit_r51_c76 bl[76] br[76] wl[51] vdd gnd cell_6t
Xbit_r52_c76 bl[76] br[76] wl[52] vdd gnd cell_6t
Xbit_r53_c76 bl[76] br[76] wl[53] vdd gnd cell_6t
Xbit_r54_c76 bl[76] br[76] wl[54] vdd gnd cell_6t
Xbit_r55_c76 bl[76] br[76] wl[55] vdd gnd cell_6t
Xbit_r56_c76 bl[76] br[76] wl[56] vdd gnd cell_6t
Xbit_r57_c76 bl[76] br[76] wl[57] vdd gnd cell_6t
Xbit_r58_c76 bl[76] br[76] wl[58] vdd gnd cell_6t
Xbit_r59_c76 bl[76] br[76] wl[59] vdd gnd cell_6t
Xbit_r60_c76 bl[76] br[76] wl[60] vdd gnd cell_6t
Xbit_r61_c76 bl[76] br[76] wl[61] vdd gnd cell_6t
Xbit_r62_c76 bl[76] br[76] wl[62] vdd gnd cell_6t
Xbit_r63_c76 bl[76] br[76] wl[63] vdd gnd cell_6t
Xbit_r64_c76 bl[76] br[76] wl[64] vdd gnd cell_6t
Xbit_r65_c76 bl[76] br[76] wl[65] vdd gnd cell_6t
Xbit_r66_c76 bl[76] br[76] wl[66] vdd gnd cell_6t
Xbit_r67_c76 bl[76] br[76] wl[67] vdd gnd cell_6t
Xbit_r68_c76 bl[76] br[76] wl[68] vdd gnd cell_6t
Xbit_r69_c76 bl[76] br[76] wl[69] vdd gnd cell_6t
Xbit_r70_c76 bl[76] br[76] wl[70] vdd gnd cell_6t
Xbit_r71_c76 bl[76] br[76] wl[71] vdd gnd cell_6t
Xbit_r72_c76 bl[76] br[76] wl[72] vdd gnd cell_6t
Xbit_r73_c76 bl[76] br[76] wl[73] vdd gnd cell_6t
Xbit_r74_c76 bl[76] br[76] wl[74] vdd gnd cell_6t
Xbit_r75_c76 bl[76] br[76] wl[75] vdd gnd cell_6t
Xbit_r76_c76 bl[76] br[76] wl[76] vdd gnd cell_6t
Xbit_r77_c76 bl[76] br[76] wl[77] vdd gnd cell_6t
Xbit_r78_c76 bl[76] br[76] wl[78] vdd gnd cell_6t
Xbit_r79_c76 bl[76] br[76] wl[79] vdd gnd cell_6t
Xbit_r80_c76 bl[76] br[76] wl[80] vdd gnd cell_6t
Xbit_r81_c76 bl[76] br[76] wl[81] vdd gnd cell_6t
Xbit_r82_c76 bl[76] br[76] wl[82] vdd gnd cell_6t
Xbit_r83_c76 bl[76] br[76] wl[83] vdd gnd cell_6t
Xbit_r84_c76 bl[76] br[76] wl[84] vdd gnd cell_6t
Xbit_r85_c76 bl[76] br[76] wl[85] vdd gnd cell_6t
Xbit_r86_c76 bl[76] br[76] wl[86] vdd gnd cell_6t
Xbit_r87_c76 bl[76] br[76] wl[87] vdd gnd cell_6t
Xbit_r88_c76 bl[76] br[76] wl[88] vdd gnd cell_6t
Xbit_r89_c76 bl[76] br[76] wl[89] vdd gnd cell_6t
Xbit_r90_c76 bl[76] br[76] wl[90] vdd gnd cell_6t
Xbit_r91_c76 bl[76] br[76] wl[91] vdd gnd cell_6t
Xbit_r92_c76 bl[76] br[76] wl[92] vdd gnd cell_6t
Xbit_r93_c76 bl[76] br[76] wl[93] vdd gnd cell_6t
Xbit_r94_c76 bl[76] br[76] wl[94] vdd gnd cell_6t
Xbit_r95_c76 bl[76] br[76] wl[95] vdd gnd cell_6t
Xbit_r96_c76 bl[76] br[76] wl[96] vdd gnd cell_6t
Xbit_r97_c76 bl[76] br[76] wl[97] vdd gnd cell_6t
Xbit_r98_c76 bl[76] br[76] wl[98] vdd gnd cell_6t
Xbit_r99_c76 bl[76] br[76] wl[99] vdd gnd cell_6t
Xbit_r100_c76 bl[76] br[76] wl[100] vdd gnd cell_6t
Xbit_r101_c76 bl[76] br[76] wl[101] vdd gnd cell_6t
Xbit_r102_c76 bl[76] br[76] wl[102] vdd gnd cell_6t
Xbit_r103_c76 bl[76] br[76] wl[103] vdd gnd cell_6t
Xbit_r104_c76 bl[76] br[76] wl[104] vdd gnd cell_6t
Xbit_r105_c76 bl[76] br[76] wl[105] vdd gnd cell_6t
Xbit_r106_c76 bl[76] br[76] wl[106] vdd gnd cell_6t
Xbit_r107_c76 bl[76] br[76] wl[107] vdd gnd cell_6t
Xbit_r108_c76 bl[76] br[76] wl[108] vdd gnd cell_6t
Xbit_r109_c76 bl[76] br[76] wl[109] vdd gnd cell_6t
Xbit_r110_c76 bl[76] br[76] wl[110] vdd gnd cell_6t
Xbit_r111_c76 bl[76] br[76] wl[111] vdd gnd cell_6t
Xbit_r112_c76 bl[76] br[76] wl[112] vdd gnd cell_6t
Xbit_r113_c76 bl[76] br[76] wl[113] vdd gnd cell_6t
Xbit_r114_c76 bl[76] br[76] wl[114] vdd gnd cell_6t
Xbit_r115_c76 bl[76] br[76] wl[115] vdd gnd cell_6t
Xbit_r116_c76 bl[76] br[76] wl[116] vdd gnd cell_6t
Xbit_r117_c76 bl[76] br[76] wl[117] vdd gnd cell_6t
Xbit_r118_c76 bl[76] br[76] wl[118] vdd gnd cell_6t
Xbit_r119_c76 bl[76] br[76] wl[119] vdd gnd cell_6t
Xbit_r120_c76 bl[76] br[76] wl[120] vdd gnd cell_6t
Xbit_r121_c76 bl[76] br[76] wl[121] vdd gnd cell_6t
Xbit_r122_c76 bl[76] br[76] wl[122] vdd gnd cell_6t
Xbit_r123_c76 bl[76] br[76] wl[123] vdd gnd cell_6t
Xbit_r124_c76 bl[76] br[76] wl[124] vdd gnd cell_6t
Xbit_r125_c76 bl[76] br[76] wl[125] vdd gnd cell_6t
Xbit_r126_c76 bl[76] br[76] wl[126] vdd gnd cell_6t
Xbit_r127_c76 bl[76] br[76] wl[127] vdd gnd cell_6t
Xbit_r128_c76 bl[76] br[76] wl[128] vdd gnd cell_6t
Xbit_r129_c76 bl[76] br[76] wl[129] vdd gnd cell_6t
Xbit_r130_c76 bl[76] br[76] wl[130] vdd gnd cell_6t
Xbit_r131_c76 bl[76] br[76] wl[131] vdd gnd cell_6t
Xbit_r132_c76 bl[76] br[76] wl[132] vdd gnd cell_6t
Xbit_r133_c76 bl[76] br[76] wl[133] vdd gnd cell_6t
Xbit_r134_c76 bl[76] br[76] wl[134] vdd gnd cell_6t
Xbit_r135_c76 bl[76] br[76] wl[135] vdd gnd cell_6t
Xbit_r136_c76 bl[76] br[76] wl[136] vdd gnd cell_6t
Xbit_r137_c76 bl[76] br[76] wl[137] vdd gnd cell_6t
Xbit_r138_c76 bl[76] br[76] wl[138] vdd gnd cell_6t
Xbit_r139_c76 bl[76] br[76] wl[139] vdd gnd cell_6t
Xbit_r140_c76 bl[76] br[76] wl[140] vdd gnd cell_6t
Xbit_r141_c76 bl[76] br[76] wl[141] vdd gnd cell_6t
Xbit_r142_c76 bl[76] br[76] wl[142] vdd gnd cell_6t
Xbit_r143_c76 bl[76] br[76] wl[143] vdd gnd cell_6t
Xbit_r144_c76 bl[76] br[76] wl[144] vdd gnd cell_6t
Xbit_r145_c76 bl[76] br[76] wl[145] vdd gnd cell_6t
Xbit_r146_c76 bl[76] br[76] wl[146] vdd gnd cell_6t
Xbit_r147_c76 bl[76] br[76] wl[147] vdd gnd cell_6t
Xbit_r148_c76 bl[76] br[76] wl[148] vdd gnd cell_6t
Xbit_r149_c76 bl[76] br[76] wl[149] vdd gnd cell_6t
Xbit_r150_c76 bl[76] br[76] wl[150] vdd gnd cell_6t
Xbit_r151_c76 bl[76] br[76] wl[151] vdd gnd cell_6t
Xbit_r152_c76 bl[76] br[76] wl[152] vdd gnd cell_6t
Xbit_r153_c76 bl[76] br[76] wl[153] vdd gnd cell_6t
Xbit_r154_c76 bl[76] br[76] wl[154] vdd gnd cell_6t
Xbit_r155_c76 bl[76] br[76] wl[155] vdd gnd cell_6t
Xbit_r156_c76 bl[76] br[76] wl[156] vdd gnd cell_6t
Xbit_r157_c76 bl[76] br[76] wl[157] vdd gnd cell_6t
Xbit_r158_c76 bl[76] br[76] wl[158] vdd gnd cell_6t
Xbit_r159_c76 bl[76] br[76] wl[159] vdd gnd cell_6t
Xbit_r160_c76 bl[76] br[76] wl[160] vdd gnd cell_6t
Xbit_r161_c76 bl[76] br[76] wl[161] vdd gnd cell_6t
Xbit_r162_c76 bl[76] br[76] wl[162] vdd gnd cell_6t
Xbit_r163_c76 bl[76] br[76] wl[163] vdd gnd cell_6t
Xbit_r164_c76 bl[76] br[76] wl[164] vdd gnd cell_6t
Xbit_r165_c76 bl[76] br[76] wl[165] vdd gnd cell_6t
Xbit_r166_c76 bl[76] br[76] wl[166] vdd gnd cell_6t
Xbit_r167_c76 bl[76] br[76] wl[167] vdd gnd cell_6t
Xbit_r168_c76 bl[76] br[76] wl[168] vdd gnd cell_6t
Xbit_r169_c76 bl[76] br[76] wl[169] vdd gnd cell_6t
Xbit_r170_c76 bl[76] br[76] wl[170] vdd gnd cell_6t
Xbit_r171_c76 bl[76] br[76] wl[171] vdd gnd cell_6t
Xbit_r172_c76 bl[76] br[76] wl[172] vdd gnd cell_6t
Xbit_r173_c76 bl[76] br[76] wl[173] vdd gnd cell_6t
Xbit_r174_c76 bl[76] br[76] wl[174] vdd gnd cell_6t
Xbit_r175_c76 bl[76] br[76] wl[175] vdd gnd cell_6t
Xbit_r176_c76 bl[76] br[76] wl[176] vdd gnd cell_6t
Xbit_r177_c76 bl[76] br[76] wl[177] vdd gnd cell_6t
Xbit_r178_c76 bl[76] br[76] wl[178] vdd gnd cell_6t
Xbit_r179_c76 bl[76] br[76] wl[179] vdd gnd cell_6t
Xbit_r180_c76 bl[76] br[76] wl[180] vdd gnd cell_6t
Xbit_r181_c76 bl[76] br[76] wl[181] vdd gnd cell_6t
Xbit_r182_c76 bl[76] br[76] wl[182] vdd gnd cell_6t
Xbit_r183_c76 bl[76] br[76] wl[183] vdd gnd cell_6t
Xbit_r184_c76 bl[76] br[76] wl[184] vdd gnd cell_6t
Xbit_r185_c76 bl[76] br[76] wl[185] vdd gnd cell_6t
Xbit_r186_c76 bl[76] br[76] wl[186] vdd gnd cell_6t
Xbit_r187_c76 bl[76] br[76] wl[187] vdd gnd cell_6t
Xbit_r188_c76 bl[76] br[76] wl[188] vdd gnd cell_6t
Xbit_r189_c76 bl[76] br[76] wl[189] vdd gnd cell_6t
Xbit_r190_c76 bl[76] br[76] wl[190] vdd gnd cell_6t
Xbit_r191_c76 bl[76] br[76] wl[191] vdd gnd cell_6t
Xbit_r192_c76 bl[76] br[76] wl[192] vdd gnd cell_6t
Xbit_r193_c76 bl[76] br[76] wl[193] vdd gnd cell_6t
Xbit_r194_c76 bl[76] br[76] wl[194] vdd gnd cell_6t
Xbit_r195_c76 bl[76] br[76] wl[195] vdd gnd cell_6t
Xbit_r196_c76 bl[76] br[76] wl[196] vdd gnd cell_6t
Xbit_r197_c76 bl[76] br[76] wl[197] vdd gnd cell_6t
Xbit_r198_c76 bl[76] br[76] wl[198] vdd gnd cell_6t
Xbit_r199_c76 bl[76] br[76] wl[199] vdd gnd cell_6t
Xbit_r200_c76 bl[76] br[76] wl[200] vdd gnd cell_6t
Xbit_r201_c76 bl[76] br[76] wl[201] vdd gnd cell_6t
Xbit_r202_c76 bl[76] br[76] wl[202] vdd gnd cell_6t
Xbit_r203_c76 bl[76] br[76] wl[203] vdd gnd cell_6t
Xbit_r204_c76 bl[76] br[76] wl[204] vdd gnd cell_6t
Xbit_r205_c76 bl[76] br[76] wl[205] vdd gnd cell_6t
Xbit_r206_c76 bl[76] br[76] wl[206] vdd gnd cell_6t
Xbit_r207_c76 bl[76] br[76] wl[207] vdd gnd cell_6t
Xbit_r208_c76 bl[76] br[76] wl[208] vdd gnd cell_6t
Xbit_r209_c76 bl[76] br[76] wl[209] vdd gnd cell_6t
Xbit_r210_c76 bl[76] br[76] wl[210] vdd gnd cell_6t
Xbit_r211_c76 bl[76] br[76] wl[211] vdd gnd cell_6t
Xbit_r212_c76 bl[76] br[76] wl[212] vdd gnd cell_6t
Xbit_r213_c76 bl[76] br[76] wl[213] vdd gnd cell_6t
Xbit_r214_c76 bl[76] br[76] wl[214] vdd gnd cell_6t
Xbit_r215_c76 bl[76] br[76] wl[215] vdd gnd cell_6t
Xbit_r216_c76 bl[76] br[76] wl[216] vdd gnd cell_6t
Xbit_r217_c76 bl[76] br[76] wl[217] vdd gnd cell_6t
Xbit_r218_c76 bl[76] br[76] wl[218] vdd gnd cell_6t
Xbit_r219_c76 bl[76] br[76] wl[219] vdd gnd cell_6t
Xbit_r220_c76 bl[76] br[76] wl[220] vdd gnd cell_6t
Xbit_r221_c76 bl[76] br[76] wl[221] vdd gnd cell_6t
Xbit_r222_c76 bl[76] br[76] wl[222] vdd gnd cell_6t
Xbit_r223_c76 bl[76] br[76] wl[223] vdd gnd cell_6t
Xbit_r224_c76 bl[76] br[76] wl[224] vdd gnd cell_6t
Xbit_r225_c76 bl[76] br[76] wl[225] vdd gnd cell_6t
Xbit_r226_c76 bl[76] br[76] wl[226] vdd gnd cell_6t
Xbit_r227_c76 bl[76] br[76] wl[227] vdd gnd cell_6t
Xbit_r228_c76 bl[76] br[76] wl[228] vdd gnd cell_6t
Xbit_r229_c76 bl[76] br[76] wl[229] vdd gnd cell_6t
Xbit_r230_c76 bl[76] br[76] wl[230] vdd gnd cell_6t
Xbit_r231_c76 bl[76] br[76] wl[231] vdd gnd cell_6t
Xbit_r232_c76 bl[76] br[76] wl[232] vdd gnd cell_6t
Xbit_r233_c76 bl[76] br[76] wl[233] vdd gnd cell_6t
Xbit_r234_c76 bl[76] br[76] wl[234] vdd gnd cell_6t
Xbit_r235_c76 bl[76] br[76] wl[235] vdd gnd cell_6t
Xbit_r236_c76 bl[76] br[76] wl[236] vdd gnd cell_6t
Xbit_r237_c76 bl[76] br[76] wl[237] vdd gnd cell_6t
Xbit_r238_c76 bl[76] br[76] wl[238] vdd gnd cell_6t
Xbit_r239_c76 bl[76] br[76] wl[239] vdd gnd cell_6t
Xbit_r240_c76 bl[76] br[76] wl[240] vdd gnd cell_6t
Xbit_r241_c76 bl[76] br[76] wl[241] vdd gnd cell_6t
Xbit_r242_c76 bl[76] br[76] wl[242] vdd gnd cell_6t
Xbit_r243_c76 bl[76] br[76] wl[243] vdd gnd cell_6t
Xbit_r244_c76 bl[76] br[76] wl[244] vdd gnd cell_6t
Xbit_r245_c76 bl[76] br[76] wl[245] vdd gnd cell_6t
Xbit_r246_c76 bl[76] br[76] wl[246] vdd gnd cell_6t
Xbit_r247_c76 bl[76] br[76] wl[247] vdd gnd cell_6t
Xbit_r248_c76 bl[76] br[76] wl[248] vdd gnd cell_6t
Xbit_r249_c76 bl[76] br[76] wl[249] vdd gnd cell_6t
Xbit_r250_c76 bl[76] br[76] wl[250] vdd gnd cell_6t
Xbit_r251_c76 bl[76] br[76] wl[251] vdd gnd cell_6t
Xbit_r252_c76 bl[76] br[76] wl[252] vdd gnd cell_6t
Xbit_r253_c76 bl[76] br[76] wl[253] vdd gnd cell_6t
Xbit_r254_c76 bl[76] br[76] wl[254] vdd gnd cell_6t
Xbit_r255_c76 bl[76] br[76] wl[255] vdd gnd cell_6t
Xbit_r0_c77 bl[77] br[77] wl[0] vdd gnd cell_6t
Xbit_r1_c77 bl[77] br[77] wl[1] vdd gnd cell_6t
Xbit_r2_c77 bl[77] br[77] wl[2] vdd gnd cell_6t
Xbit_r3_c77 bl[77] br[77] wl[3] vdd gnd cell_6t
Xbit_r4_c77 bl[77] br[77] wl[4] vdd gnd cell_6t
Xbit_r5_c77 bl[77] br[77] wl[5] vdd gnd cell_6t
Xbit_r6_c77 bl[77] br[77] wl[6] vdd gnd cell_6t
Xbit_r7_c77 bl[77] br[77] wl[7] vdd gnd cell_6t
Xbit_r8_c77 bl[77] br[77] wl[8] vdd gnd cell_6t
Xbit_r9_c77 bl[77] br[77] wl[9] vdd gnd cell_6t
Xbit_r10_c77 bl[77] br[77] wl[10] vdd gnd cell_6t
Xbit_r11_c77 bl[77] br[77] wl[11] vdd gnd cell_6t
Xbit_r12_c77 bl[77] br[77] wl[12] vdd gnd cell_6t
Xbit_r13_c77 bl[77] br[77] wl[13] vdd gnd cell_6t
Xbit_r14_c77 bl[77] br[77] wl[14] vdd gnd cell_6t
Xbit_r15_c77 bl[77] br[77] wl[15] vdd gnd cell_6t
Xbit_r16_c77 bl[77] br[77] wl[16] vdd gnd cell_6t
Xbit_r17_c77 bl[77] br[77] wl[17] vdd gnd cell_6t
Xbit_r18_c77 bl[77] br[77] wl[18] vdd gnd cell_6t
Xbit_r19_c77 bl[77] br[77] wl[19] vdd gnd cell_6t
Xbit_r20_c77 bl[77] br[77] wl[20] vdd gnd cell_6t
Xbit_r21_c77 bl[77] br[77] wl[21] vdd gnd cell_6t
Xbit_r22_c77 bl[77] br[77] wl[22] vdd gnd cell_6t
Xbit_r23_c77 bl[77] br[77] wl[23] vdd gnd cell_6t
Xbit_r24_c77 bl[77] br[77] wl[24] vdd gnd cell_6t
Xbit_r25_c77 bl[77] br[77] wl[25] vdd gnd cell_6t
Xbit_r26_c77 bl[77] br[77] wl[26] vdd gnd cell_6t
Xbit_r27_c77 bl[77] br[77] wl[27] vdd gnd cell_6t
Xbit_r28_c77 bl[77] br[77] wl[28] vdd gnd cell_6t
Xbit_r29_c77 bl[77] br[77] wl[29] vdd gnd cell_6t
Xbit_r30_c77 bl[77] br[77] wl[30] vdd gnd cell_6t
Xbit_r31_c77 bl[77] br[77] wl[31] vdd gnd cell_6t
Xbit_r32_c77 bl[77] br[77] wl[32] vdd gnd cell_6t
Xbit_r33_c77 bl[77] br[77] wl[33] vdd gnd cell_6t
Xbit_r34_c77 bl[77] br[77] wl[34] vdd gnd cell_6t
Xbit_r35_c77 bl[77] br[77] wl[35] vdd gnd cell_6t
Xbit_r36_c77 bl[77] br[77] wl[36] vdd gnd cell_6t
Xbit_r37_c77 bl[77] br[77] wl[37] vdd gnd cell_6t
Xbit_r38_c77 bl[77] br[77] wl[38] vdd gnd cell_6t
Xbit_r39_c77 bl[77] br[77] wl[39] vdd gnd cell_6t
Xbit_r40_c77 bl[77] br[77] wl[40] vdd gnd cell_6t
Xbit_r41_c77 bl[77] br[77] wl[41] vdd gnd cell_6t
Xbit_r42_c77 bl[77] br[77] wl[42] vdd gnd cell_6t
Xbit_r43_c77 bl[77] br[77] wl[43] vdd gnd cell_6t
Xbit_r44_c77 bl[77] br[77] wl[44] vdd gnd cell_6t
Xbit_r45_c77 bl[77] br[77] wl[45] vdd gnd cell_6t
Xbit_r46_c77 bl[77] br[77] wl[46] vdd gnd cell_6t
Xbit_r47_c77 bl[77] br[77] wl[47] vdd gnd cell_6t
Xbit_r48_c77 bl[77] br[77] wl[48] vdd gnd cell_6t
Xbit_r49_c77 bl[77] br[77] wl[49] vdd gnd cell_6t
Xbit_r50_c77 bl[77] br[77] wl[50] vdd gnd cell_6t
Xbit_r51_c77 bl[77] br[77] wl[51] vdd gnd cell_6t
Xbit_r52_c77 bl[77] br[77] wl[52] vdd gnd cell_6t
Xbit_r53_c77 bl[77] br[77] wl[53] vdd gnd cell_6t
Xbit_r54_c77 bl[77] br[77] wl[54] vdd gnd cell_6t
Xbit_r55_c77 bl[77] br[77] wl[55] vdd gnd cell_6t
Xbit_r56_c77 bl[77] br[77] wl[56] vdd gnd cell_6t
Xbit_r57_c77 bl[77] br[77] wl[57] vdd gnd cell_6t
Xbit_r58_c77 bl[77] br[77] wl[58] vdd gnd cell_6t
Xbit_r59_c77 bl[77] br[77] wl[59] vdd gnd cell_6t
Xbit_r60_c77 bl[77] br[77] wl[60] vdd gnd cell_6t
Xbit_r61_c77 bl[77] br[77] wl[61] vdd gnd cell_6t
Xbit_r62_c77 bl[77] br[77] wl[62] vdd gnd cell_6t
Xbit_r63_c77 bl[77] br[77] wl[63] vdd gnd cell_6t
Xbit_r64_c77 bl[77] br[77] wl[64] vdd gnd cell_6t
Xbit_r65_c77 bl[77] br[77] wl[65] vdd gnd cell_6t
Xbit_r66_c77 bl[77] br[77] wl[66] vdd gnd cell_6t
Xbit_r67_c77 bl[77] br[77] wl[67] vdd gnd cell_6t
Xbit_r68_c77 bl[77] br[77] wl[68] vdd gnd cell_6t
Xbit_r69_c77 bl[77] br[77] wl[69] vdd gnd cell_6t
Xbit_r70_c77 bl[77] br[77] wl[70] vdd gnd cell_6t
Xbit_r71_c77 bl[77] br[77] wl[71] vdd gnd cell_6t
Xbit_r72_c77 bl[77] br[77] wl[72] vdd gnd cell_6t
Xbit_r73_c77 bl[77] br[77] wl[73] vdd gnd cell_6t
Xbit_r74_c77 bl[77] br[77] wl[74] vdd gnd cell_6t
Xbit_r75_c77 bl[77] br[77] wl[75] vdd gnd cell_6t
Xbit_r76_c77 bl[77] br[77] wl[76] vdd gnd cell_6t
Xbit_r77_c77 bl[77] br[77] wl[77] vdd gnd cell_6t
Xbit_r78_c77 bl[77] br[77] wl[78] vdd gnd cell_6t
Xbit_r79_c77 bl[77] br[77] wl[79] vdd gnd cell_6t
Xbit_r80_c77 bl[77] br[77] wl[80] vdd gnd cell_6t
Xbit_r81_c77 bl[77] br[77] wl[81] vdd gnd cell_6t
Xbit_r82_c77 bl[77] br[77] wl[82] vdd gnd cell_6t
Xbit_r83_c77 bl[77] br[77] wl[83] vdd gnd cell_6t
Xbit_r84_c77 bl[77] br[77] wl[84] vdd gnd cell_6t
Xbit_r85_c77 bl[77] br[77] wl[85] vdd gnd cell_6t
Xbit_r86_c77 bl[77] br[77] wl[86] vdd gnd cell_6t
Xbit_r87_c77 bl[77] br[77] wl[87] vdd gnd cell_6t
Xbit_r88_c77 bl[77] br[77] wl[88] vdd gnd cell_6t
Xbit_r89_c77 bl[77] br[77] wl[89] vdd gnd cell_6t
Xbit_r90_c77 bl[77] br[77] wl[90] vdd gnd cell_6t
Xbit_r91_c77 bl[77] br[77] wl[91] vdd gnd cell_6t
Xbit_r92_c77 bl[77] br[77] wl[92] vdd gnd cell_6t
Xbit_r93_c77 bl[77] br[77] wl[93] vdd gnd cell_6t
Xbit_r94_c77 bl[77] br[77] wl[94] vdd gnd cell_6t
Xbit_r95_c77 bl[77] br[77] wl[95] vdd gnd cell_6t
Xbit_r96_c77 bl[77] br[77] wl[96] vdd gnd cell_6t
Xbit_r97_c77 bl[77] br[77] wl[97] vdd gnd cell_6t
Xbit_r98_c77 bl[77] br[77] wl[98] vdd gnd cell_6t
Xbit_r99_c77 bl[77] br[77] wl[99] vdd gnd cell_6t
Xbit_r100_c77 bl[77] br[77] wl[100] vdd gnd cell_6t
Xbit_r101_c77 bl[77] br[77] wl[101] vdd gnd cell_6t
Xbit_r102_c77 bl[77] br[77] wl[102] vdd gnd cell_6t
Xbit_r103_c77 bl[77] br[77] wl[103] vdd gnd cell_6t
Xbit_r104_c77 bl[77] br[77] wl[104] vdd gnd cell_6t
Xbit_r105_c77 bl[77] br[77] wl[105] vdd gnd cell_6t
Xbit_r106_c77 bl[77] br[77] wl[106] vdd gnd cell_6t
Xbit_r107_c77 bl[77] br[77] wl[107] vdd gnd cell_6t
Xbit_r108_c77 bl[77] br[77] wl[108] vdd gnd cell_6t
Xbit_r109_c77 bl[77] br[77] wl[109] vdd gnd cell_6t
Xbit_r110_c77 bl[77] br[77] wl[110] vdd gnd cell_6t
Xbit_r111_c77 bl[77] br[77] wl[111] vdd gnd cell_6t
Xbit_r112_c77 bl[77] br[77] wl[112] vdd gnd cell_6t
Xbit_r113_c77 bl[77] br[77] wl[113] vdd gnd cell_6t
Xbit_r114_c77 bl[77] br[77] wl[114] vdd gnd cell_6t
Xbit_r115_c77 bl[77] br[77] wl[115] vdd gnd cell_6t
Xbit_r116_c77 bl[77] br[77] wl[116] vdd gnd cell_6t
Xbit_r117_c77 bl[77] br[77] wl[117] vdd gnd cell_6t
Xbit_r118_c77 bl[77] br[77] wl[118] vdd gnd cell_6t
Xbit_r119_c77 bl[77] br[77] wl[119] vdd gnd cell_6t
Xbit_r120_c77 bl[77] br[77] wl[120] vdd gnd cell_6t
Xbit_r121_c77 bl[77] br[77] wl[121] vdd gnd cell_6t
Xbit_r122_c77 bl[77] br[77] wl[122] vdd gnd cell_6t
Xbit_r123_c77 bl[77] br[77] wl[123] vdd gnd cell_6t
Xbit_r124_c77 bl[77] br[77] wl[124] vdd gnd cell_6t
Xbit_r125_c77 bl[77] br[77] wl[125] vdd gnd cell_6t
Xbit_r126_c77 bl[77] br[77] wl[126] vdd gnd cell_6t
Xbit_r127_c77 bl[77] br[77] wl[127] vdd gnd cell_6t
Xbit_r128_c77 bl[77] br[77] wl[128] vdd gnd cell_6t
Xbit_r129_c77 bl[77] br[77] wl[129] vdd gnd cell_6t
Xbit_r130_c77 bl[77] br[77] wl[130] vdd gnd cell_6t
Xbit_r131_c77 bl[77] br[77] wl[131] vdd gnd cell_6t
Xbit_r132_c77 bl[77] br[77] wl[132] vdd gnd cell_6t
Xbit_r133_c77 bl[77] br[77] wl[133] vdd gnd cell_6t
Xbit_r134_c77 bl[77] br[77] wl[134] vdd gnd cell_6t
Xbit_r135_c77 bl[77] br[77] wl[135] vdd gnd cell_6t
Xbit_r136_c77 bl[77] br[77] wl[136] vdd gnd cell_6t
Xbit_r137_c77 bl[77] br[77] wl[137] vdd gnd cell_6t
Xbit_r138_c77 bl[77] br[77] wl[138] vdd gnd cell_6t
Xbit_r139_c77 bl[77] br[77] wl[139] vdd gnd cell_6t
Xbit_r140_c77 bl[77] br[77] wl[140] vdd gnd cell_6t
Xbit_r141_c77 bl[77] br[77] wl[141] vdd gnd cell_6t
Xbit_r142_c77 bl[77] br[77] wl[142] vdd gnd cell_6t
Xbit_r143_c77 bl[77] br[77] wl[143] vdd gnd cell_6t
Xbit_r144_c77 bl[77] br[77] wl[144] vdd gnd cell_6t
Xbit_r145_c77 bl[77] br[77] wl[145] vdd gnd cell_6t
Xbit_r146_c77 bl[77] br[77] wl[146] vdd gnd cell_6t
Xbit_r147_c77 bl[77] br[77] wl[147] vdd gnd cell_6t
Xbit_r148_c77 bl[77] br[77] wl[148] vdd gnd cell_6t
Xbit_r149_c77 bl[77] br[77] wl[149] vdd gnd cell_6t
Xbit_r150_c77 bl[77] br[77] wl[150] vdd gnd cell_6t
Xbit_r151_c77 bl[77] br[77] wl[151] vdd gnd cell_6t
Xbit_r152_c77 bl[77] br[77] wl[152] vdd gnd cell_6t
Xbit_r153_c77 bl[77] br[77] wl[153] vdd gnd cell_6t
Xbit_r154_c77 bl[77] br[77] wl[154] vdd gnd cell_6t
Xbit_r155_c77 bl[77] br[77] wl[155] vdd gnd cell_6t
Xbit_r156_c77 bl[77] br[77] wl[156] vdd gnd cell_6t
Xbit_r157_c77 bl[77] br[77] wl[157] vdd gnd cell_6t
Xbit_r158_c77 bl[77] br[77] wl[158] vdd gnd cell_6t
Xbit_r159_c77 bl[77] br[77] wl[159] vdd gnd cell_6t
Xbit_r160_c77 bl[77] br[77] wl[160] vdd gnd cell_6t
Xbit_r161_c77 bl[77] br[77] wl[161] vdd gnd cell_6t
Xbit_r162_c77 bl[77] br[77] wl[162] vdd gnd cell_6t
Xbit_r163_c77 bl[77] br[77] wl[163] vdd gnd cell_6t
Xbit_r164_c77 bl[77] br[77] wl[164] vdd gnd cell_6t
Xbit_r165_c77 bl[77] br[77] wl[165] vdd gnd cell_6t
Xbit_r166_c77 bl[77] br[77] wl[166] vdd gnd cell_6t
Xbit_r167_c77 bl[77] br[77] wl[167] vdd gnd cell_6t
Xbit_r168_c77 bl[77] br[77] wl[168] vdd gnd cell_6t
Xbit_r169_c77 bl[77] br[77] wl[169] vdd gnd cell_6t
Xbit_r170_c77 bl[77] br[77] wl[170] vdd gnd cell_6t
Xbit_r171_c77 bl[77] br[77] wl[171] vdd gnd cell_6t
Xbit_r172_c77 bl[77] br[77] wl[172] vdd gnd cell_6t
Xbit_r173_c77 bl[77] br[77] wl[173] vdd gnd cell_6t
Xbit_r174_c77 bl[77] br[77] wl[174] vdd gnd cell_6t
Xbit_r175_c77 bl[77] br[77] wl[175] vdd gnd cell_6t
Xbit_r176_c77 bl[77] br[77] wl[176] vdd gnd cell_6t
Xbit_r177_c77 bl[77] br[77] wl[177] vdd gnd cell_6t
Xbit_r178_c77 bl[77] br[77] wl[178] vdd gnd cell_6t
Xbit_r179_c77 bl[77] br[77] wl[179] vdd gnd cell_6t
Xbit_r180_c77 bl[77] br[77] wl[180] vdd gnd cell_6t
Xbit_r181_c77 bl[77] br[77] wl[181] vdd gnd cell_6t
Xbit_r182_c77 bl[77] br[77] wl[182] vdd gnd cell_6t
Xbit_r183_c77 bl[77] br[77] wl[183] vdd gnd cell_6t
Xbit_r184_c77 bl[77] br[77] wl[184] vdd gnd cell_6t
Xbit_r185_c77 bl[77] br[77] wl[185] vdd gnd cell_6t
Xbit_r186_c77 bl[77] br[77] wl[186] vdd gnd cell_6t
Xbit_r187_c77 bl[77] br[77] wl[187] vdd gnd cell_6t
Xbit_r188_c77 bl[77] br[77] wl[188] vdd gnd cell_6t
Xbit_r189_c77 bl[77] br[77] wl[189] vdd gnd cell_6t
Xbit_r190_c77 bl[77] br[77] wl[190] vdd gnd cell_6t
Xbit_r191_c77 bl[77] br[77] wl[191] vdd gnd cell_6t
Xbit_r192_c77 bl[77] br[77] wl[192] vdd gnd cell_6t
Xbit_r193_c77 bl[77] br[77] wl[193] vdd gnd cell_6t
Xbit_r194_c77 bl[77] br[77] wl[194] vdd gnd cell_6t
Xbit_r195_c77 bl[77] br[77] wl[195] vdd gnd cell_6t
Xbit_r196_c77 bl[77] br[77] wl[196] vdd gnd cell_6t
Xbit_r197_c77 bl[77] br[77] wl[197] vdd gnd cell_6t
Xbit_r198_c77 bl[77] br[77] wl[198] vdd gnd cell_6t
Xbit_r199_c77 bl[77] br[77] wl[199] vdd gnd cell_6t
Xbit_r200_c77 bl[77] br[77] wl[200] vdd gnd cell_6t
Xbit_r201_c77 bl[77] br[77] wl[201] vdd gnd cell_6t
Xbit_r202_c77 bl[77] br[77] wl[202] vdd gnd cell_6t
Xbit_r203_c77 bl[77] br[77] wl[203] vdd gnd cell_6t
Xbit_r204_c77 bl[77] br[77] wl[204] vdd gnd cell_6t
Xbit_r205_c77 bl[77] br[77] wl[205] vdd gnd cell_6t
Xbit_r206_c77 bl[77] br[77] wl[206] vdd gnd cell_6t
Xbit_r207_c77 bl[77] br[77] wl[207] vdd gnd cell_6t
Xbit_r208_c77 bl[77] br[77] wl[208] vdd gnd cell_6t
Xbit_r209_c77 bl[77] br[77] wl[209] vdd gnd cell_6t
Xbit_r210_c77 bl[77] br[77] wl[210] vdd gnd cell_6t
Xbit_r211_c77 bl[77] br[77] wl[211] vdd gnd cell_6t
Xbit_r212_c77 bl[77] br[77] wl[212] vdd gnd cell_6t
Xbit_r213_c77 bl[77] br[77] wl[213] vdd gnd cell_6t
Xbit_r214_c77 bl[77] br[77] wl[214] vdd gnd cell_6t
Xbit_r215_c77 bl[77] br[77] wl[215] vdd gnd cell_6t
Xbit_r216_c77 bl[77] br[77] wl[216] vdd gnd cell_6t
Xbit_r217_c77 bl[77] br[77] wl[217] vdd gnd cell_6t
Xbit_r218_c77 bl[77] br[77] wl[218] vdd gnd cell_6t
Xbit_r219_c77 bl[77] br[77] wl[219] vdd gnd cell_6t
Xbit_r220_c77 bl[77] br[77] wl[220] vdd gnd cell_6t
Xbit_r221_c77 bl[77] br[77] wl[221] vdd gnd cell_6t
Xbit_r222_c77 bl[77] br[77] wl[222] vdd gnd cell_6t
Xbit_r223_c77 bl[77] br[77] wl[223] vdd gnd cell_6t
Xbit_r224_c77 bl[77] br[77] wl[224] vdd gnd cell_6t
Xbit_r225_c77 bl[77] br[77] wl[225] vdd gnd cell_6t
Xbit_r226_c77 bl[77] br[77] wl[226] vdd gnd cell_6t
Xbit_r227_c77 bl[77] br[77] wl[227] vdd gnd cell_6t
Xbit_r228_c77 bl[77] br[77] wl[228] vdd gnd cell_6t
Xbit_r229_c77 bl[77] br[77] wl[229] vdd gnd cell_6t
Xbit_r230_c77 bl[77] br[77] wl[230] vdd gnd cell_6t
Xbit_r231_c77 bl[77] br[77] wl[231] vdd gnd cell_6t
Xbit_r232_c77 bl[77] br[77] wl[232] vdd gnd cell_6t
Xbit_r233_c77 bl[77] br[77] wl[233] vdd gnd cell_6t
Xbit_r234_c77 bl[77] br[77] wl[234] vdd gnd cell_6t
Xbit_r235_c77 bl[77] br[77] wl[235] vdd gnd cell_6t
Xbit_r236_c77 bl[77] br[77] wl[236] vdd gnd cell_6t
Xbit_r237_c77 bl[77] br[77] wl[237] vdd gnd cell_6t
Xbit_r238_c77 bl[77] br[77] wl[238] vdd gnd cell_6t
Xbit_r239_c77 bl[77] br[77] wl[239] vdd gnd cell_6t
Xbit_r240_c77 bl[77] br[77] wl[240] vdd gnd cell_6t
Xbit_r241_c77 bl[77] br[77] wl[241] vdd gnd cell_6t
Xbit_r242_c77 bl[77] br[77] wl[242] vdd gnd cell_6t
Xbit_r243_c77 bl[77] br[77] wl[243] vdd gnd cell_6t
Xbit_r244_c77 bl[77] br[77] wl[244] vdd gnd cell_6t
Xbit_r245_c77 bl[77] br[77] wl[245] vdd gnd cell_6t
Xbit_r246_c77 bl[77] br[77] wl[246] vdd gnd cell_6t
Xbit_r247_c77 bl[77] br[77] wl[247] vdd gnd cell_6t
Xbit_r248_c77 bl[77] br[77] wl[248] vdd gnd cell_6t
Xbit_r249_c77 bl[77] br[77] wl[249] vdd gnd cell_6t
Xbit_r250_c77 bl[77] br[77] wl[250] vdd gnd cell_6t
Xbit_r251_c77 bl[77] br[77] wl[251] vdd gnd cell_6t
Xbit_r252_c77 bl[77] br[77] wl[252] vdd gnd cell_6t
Xbit_r253_c77 bl[77] br[77] wl[253] vdd gnd cell_6t
Xbit_r254_c77 bl[77] br[77] wl[254] vdd gnd cell_6t
Xbit_r255_c77 bl[77] br[77] wl[255] vdd gnd cell_6t
Xbit_r0_c78 bl[78] br[78] wl[0] vdd gnd cell_6t
Xbit_r1_c78 bl[78] br[78] wl[1] vdd gnd cell_6t
Xbit_r2_c78 bl[78] br[78] wl[2] vdd gnd cell_6t
Xbit_r3_c78 bl[78] br[78] wl[3] vdd gnd cell_6t
Xbit_r4_c78 bl[78] br[78] wl[4] vdd gnd cell_6t
Xbit_r5_c78 bl[78] br[78] wl[5] vdd gnd cell_6t
Xbit_r6_c78 bl[78] br[78] wl[6] vdd gnd cell_6t
Xbit_r7_c78 bl[78] br[78] wl[7] vdd gnd cell_6t
Xbit_r8_c78 bl[78] br[78] wl[8] vdd gnd cell_6t
Xbit_r9_c78 bl[78] br[78] wl[9] vdd gnd cell_6t
Xbit_r10_c78 bl[78] br[78] wl[10] vdd gnd cell_6t
Xbit_r11_c78 bl[78] br[78] wl[11] vdd gnd cell_6t
Xbit_r12_c78 bl[78] br[78] wl[12] vdd gnd cell_6t
Xbit_r13_c78 bl[78] br[78] wl[13] vdd gnd cell_6t
Xbit_r14_c78 bl[78] br[78] wl[14] vdd gnd cell_6t
Xbit_r15_c78 bl[78] br[78] wl[15] vdd gnd cell_6t
Xbit_r16_c78 bl[78] br[78] wl[16] vdd gnd cell_6t
Xbit_r17_c78 bl[78] br[78] wl[17] vdd gnd cell_6t
Xbit_r18_c78 bl[78] br[78] wl[18] vdd gnd cell_6t
Xbit_r19_c78 bl[78] br[78] wl[19] vdd gnd cell_6t
Xbit_r20_c78 bl[78] br[78] wl[20] vdd gnd cell_6t
Xbit_r21_c78 bl[78] br[78] wl[21] vdd gnd cell_6t
Xbit_r22_c78 bl[78] br[78] wl[22] vdd gnd cell_6t
Xbit_r23_c78 bl[78] br[78] wl[23] vdd gnd cell_6t
Xbit_r24_c78 bl[78] br[78] wl[24] vdd gnd cell_6t
Xbit_r25_c78 bl[78] br[78] wl[25] vdd gnd cell_6t
Xbit_r26_c78 bl[78] br[78] wl[26] vdd gnd cell_6t
Xbit_r27_c78 bl[78] br[78] wl[27] vdd gnd cell_6t
Xbit_r28_c78 bl[78] br[78] wl[28] vdd gnd cell_6t
Xbit_r29_c78 bl[78] br[78] wl[29] vdd gnd cell_6t
Xbit_r30_c78 bl[78] br[78] wl[30] vdd gnd cell_6t
Xbit_r31_c78 bl[78] br[78] wl[31] vdd gnd cell_6t
Xbit_r32_c78 bl[78] br[78] wl[32] vdd gnd cell_6t
Xbit_r33_c78 bl[78] br[78] wl[33] vdd gnd cell_6t
Xbit_r34_c78 bl[78] br[78] wl[34] vdd gnd cell_6t
Xbit_r35_c78 bl[78] br[78] wl[35] vdd gnd cell_6t
Xbit_r36_c78 bl[78] br[78] wl[36] vdd gnd cell_6t
Xbit_r37_c78 bl[78] br[78] wl[37] vdd gnd cell_6t
Xbit_r38_c78 bl[78] br[78] wl[38] vdd gnd cell_6t
Xbit_r39_c78 bl[78] br[78] wl[39] vdd gnd cell_6t
Xbit_r40_c78 bl[78] br[78] wl[40] vdd gnd cell_6t
Xbit_r41_c78 bl[78] br[78] wl[41] vdd gnd cell_6t
Xbit_r42_c78 bl[78] br[78] wl[42] vdd gnd cell_6t
Xbit_r43_c78 bl[78] br[78] wl[43] vdd gnd cell_6t
Xbit_r44_c78 bl[78] br[78] wl[44] vdd gnd cell_6t
Xbit_r45_c78 bl[78] br[78] wl[45] vdd gnd cell_6t
Xbit_r46_c78 bl[78] br[78] wl[46] vdd gnd cell_6t
Xbit_r47_c78 bl[78] br[78] wl[47] vdd gnd cell_6t
Xbit_r48_c78 bl[78] br[78] wl[48] vdd gnd cell_6t
Xbit_r49_c78 bl[78] br[78] wl[49] vdd gnd cell_6t
Xbit_r50_c78 bl[78] br[78] wl[50] vdd gnd cell_6t
Xbit_r51_c78 bl[78] br[78] wl[51] vdd gnd cell_6t
Xbit_r52_c78 bl[78] br[78] wl[52] vdd gnd cell_6t
Xbit_r53_c78 bl[78] br[78] wl[53] vdd gnd cell_6t
Xbit_r54_c78 bl[78] br[78] wl[54] vdd gnd cell_6t
Xbit_r55_c78 bl[78] br[78] wl[55] vdd gnd cell_6t
Xbit_r56_c78 bl[78] br[78] wl[56] vdd gnd cell_6t
Xbit_r57_c78 bl[78] br[78] wl[57] vdd gnd cell_6t
Xbit_r58_c78 bl[78] br[78] wl[58] vdd gnd cell_6t
Xbit_r59_c78 bl[78] br[78] wl[59] vdd gnd cell_6t
Xbit_r60_c78 bl[78] br[78] wl[60] vdd gnd cell_6t
Xbit_r61_c78 bl[78] br[78] wl[61] vdd gnd cell_6t
Xbit_r62_c78 bl[78] br[78] wl[62] vdd gnd cell_6t
Xbit_r63_c78 bl[78] br[78] wl[63] vdd gnd cell_6t
Xbit_r64_c78 bl[78] br[78] wl[64] vdd gnd cell_6t
Xbit_r65_c78 bl[78] br[78] wl[65] vdd gnd cell_6t
Xbit_r66_c78 bl[78] br[78] wl[66] vdd gnd cell_6t
Xbit_r67_c78 bl[78] br[78] wl[67] vdd gnd cell_6t
Xbit_r68_c78 bl[78] br[78] wl[68] vdd gnd cell_6t
Xbit_r69_c78 bl[78] br[78] wl[69] vdd gnd cell_6t
Xbit_r70_c78 bl[78] br[78] wl[70] vdd gnd cell_6t
Xbit_r71_c78 bl[78] br[78] wl[71] vdd gnd cell_6t
Xbit_r72_c78 bl[78] br[78] wl[72] vdd gnd cell_6t
Xbit_r73_c78 bl[78] br[78] wl[73] vdd gnd cell_6t
Xbit_r74_c78 bl[78] br[78] wl[74] vdd gnd cell_6t
Xbit_r75_c78 bl[78] br[78] wl[75] vdd gnd cell_6t
Xbit_r76_c78 bl[78] br[78] wl[76] vdd gnd cell_6t
Xbit_r77_c78 bl[78] br[78] wl[77] vdd gnd cell_6t
Xbit_r78_c78 bl[78] br[78] wl[78] vdd gnd cell_6t
Xbit_r79_c78 bl[78] br[78] wl[79] vdd gnd cell_6t
Xbit_r80_c78 bl[78] br[78] wl[80] vdd gnd cell_6t
Xbit_r81_c78 bl[78] br[78] wl[81] vdd gnd cell_6t
Xbit_r82_c78 bl[78] br[78] wl[82] vdd gnd cell_6t
Xbit_r83_c78 bl[78] br[78] wl[83] vdd gnd cell_6t
Xbit_r84_c78 bl[78] br[78] wl[84] vdd gnd cell_6t
Xbit_r85_c78 bl[78] br[78] wl[85] vdd gnd cell_6t
Xbit_r86_c78 bl[78] br[78] wl[86] vdd gnd cell_6t
Xbit_r87_c78 bl[78] br[78] wl[87] vdd gnd cell_6t
Xbit_r88_c78 bl[78] br[78] wl[88] vdd gnd cell_6t
Xbit_r89_c78 bl[78] br[78] wl[89] vdd gnd cell_6t
Xbit_r90_c78 bl[78] br[78] wl[90] vdd gnd cell_6t
Xbit_r91_c78 bl[78] br[78] wl[91] vdd gnd cell_6t
Xbit_r92_c78 bl[78] br[78] wl[92] vdd gnd cell_6t
Xbit_r93_c78 bl[78] br[78] wl[93] vdd gnd cell_6t
Xbit_r94_c78 bl[78] br[78] wl[94] vdd gnd cell_6t
Xbit_r95_c78 bl[78] br[78] wl[95] vdd gnd cell_6t
Xbit_r96_c78 bl[78] br[78] wl[96] vdd gnd cell_6t
Xbit_r97_c78 bl[78] br[78] wl[97] vdd gnd cell_6t
Xbit_r98_c78 bl[78] br[78] wl[98] vdd gnd cell_6t
Xbit_r99_c78 bl[78] br[78] wl[99] vdd gnd cell_6t
Xbit_r100_c78 bl[78] br[78] wl[100] vdd gnd cell_6t
Xbit_r101_c78 bl[78] br[78] wl[101] vdd gnd cell_6t
Xbit_r102_c78 bl[78] br[78] wl[102] vdd gnd cell_6t
Xbit_r103_c78 bl[78] br[78] wl[103] vdd gnd cell_6t
Xbit_r104_c78 bl[78] br[78] wl[104] vdd gnd cell_6t
Xbit_r105_c78 bl[78] br[78] wl[105] vdd gnd cell_6t
Xbit_r106_c78 bl[78] br[78] wl[106] vdd gnd cell_6t
Xbit_r107_c78 bl[78] br[78] wl[107] vdd gnd cell_6t
Xbit_r108_c78 bl[78] br[78] wl[108] vdd gnd cell_6t
Xbit_r109_c78 bl[78] br[78] wl[109] vdd gnd cell_6t
Xbit_r110_c78 bl[78] br[78] wl[110] vdd gnd cell_6t
Xbit_r111_c78 bl[78] br[78] wl[111] vdd gnd cell_6t
Xbit_r112_c78 bl[78] br[78] wl[112] vdd gnd cell_6t
Xbit_r113_c78 bl[78] br[78] wl[113] vdd gnd cell_6t
Xbit_r114_c78 bl[78] br[78] wl[114] vdd gnd cell_6t
Xbit_r115_c78 bl[78] br[78] wl[115] vdd gnd cell_6t
Xbit_r116_c78 bl[78] br[78] wl[116] vdd gnd cell_6t
Xbit_r117_c78 bl[78] br[78] wl[117] vdd gnd cell_6t
Xbit_r118_c78 bl[78] br[78] wl[118] vdd gnd cell_6t
Xbit_r119_c78 bl[78] br[78] wl[119] vdd gnd cell_6t
Xbit_r120_c78 bl[78] br[78] wl[120] vdd gnd cell_6t
Xbit_r121_c78 bl[78] br[78] wl[121] vdd gnd cell_6t
Xbit_r122_c78 bl[78] br[78] wl[122] vdd gnd cell_6t
Xbit_r123_c78 bl[78] br[78] wl[123] vdd gnd cell_6t
Xbit_r124_c78 bl[78] br[78] wl[124] vdd gnd cell_6t
Xbit_r125_c78 bl[78] br[78] wl[125] vdd gnd cell_6t
Xbit_r126_c78 bl[78] br[78] wl[126] vdd gnd cell_6t
Xbit_r127_c78 bl[78] br[78] wl[127] vdd gnd cell_6t
Xbit_r128_c78 bl[78] br[78] wl[128] vdd gnd cell_6t
Xbit_r129_c78 bl[78] br[78] wl[129] vdd gnd cell_6t
Xbit_r130_c78 bl[78] br[78] wl[130] vdd gnd cell_6t
Xbit_r131_c78 bl[78] br[78] wl[131] vdd gnd cell_6t
Xbit_r132_c78 bl[78] br[78] wl[132] vdd gnd cell_6t
Xbit_r133_c78 bl[78] br[78] wl[133] vdd gnd cell_6t
Xbit_r134_c78 bl[78] br[78] wl[134] vdd gnd cell_6t
Xbit_r135_c78 bl[78] br[78] wl[135] vdd gnd cell_6t
Xbit_r136_c78 bl[78] br[78] wl[136] vdd gnd cell_6t
Xbit_r137_c78 bl[78] br[78] wl[137] vdd gnd cell_6t
Xbit_r138_c78 bl[78] br[78] wl[138] vdd gnd cell_6t
Xbit_r139_c78 bl[78] br[78] wl[139] vdd gnd cell_6t
Xbit_r140_c78 bl[78] br[78] wl[140] vdd gnd cell_6t
Xbit_r141_c78 bl[78] br[78] wl[141] vdd gnd cell_6t
Xbit_r142_c78 bl[78] br[78] wl[142] vdd gnd cell_6t
Xbit_r143_c78 bl[78] br[78] wl[143] vdd gnd cell_6t
Xbit_r144_c78 bl[78] br[78] wl[144] vdd gnd cell_6t
Xbit_r145_c78 bl[78] br[78] wl[145] vdd gnd cell_6t
Xbit_r146_c78 bl[78] br[78] wl[146] vdd gnd cell_6t
Xbit_r147_c78 bl[78] br[78] wl[147] vdd gnd cell_6t
Xbit_r148_c78 bl[78] br[78] wl[148] vdd gnd cell_6t
Xbit_r149_c78 bl[78] br[78] wl[149] vdd gnd cell_6t
Xbit_r150_c78 bl[78] br[78] wl[150] vdd gnd cell_6t
Xbit_r151_c78 bl[78] br[78] wl[151] vdd gnd cell_6t
Xbit_r152_c78 bl[78] br[78] wl[152] vdd gnd cell_6t
Xbit_r153_c78 bl[78] br[78] wl[153] vdd gnd cell_6t
Xbit_r154_c78 bl[78] br[78] wl[154] vdd gnd cell_6t
Xbit_r155_c78 bl[78] br[78] wl[155] vdd gnd cell_6t
Xbit_r156_c78 bl[78] br[78] wl[156] vdd gnd cell_6t
Xbit_r157_c78 bl[78] br[78] wl[157] vdd gnd cell_6t
Xbit_r158_c78 bl[78] br[78] wl[158] vdd gnd cell_6t
Xbit_r159_c78 bl[78] br[78] wl[159] vdd gnd cell_6t
Xbit_r160_c78 bl[78] br[78] wl[160] vdd gnd cell_6t
Xbit_r161_c78 bl[78] br[78] wl[161] vdd gnd cell_6t
Xbit_r162_c78 bl[78] br[78] wl[162] vdd gnd cell_6t
Xbit_r163_c78 bl[78] br[78] wl[163] vdd gnd cell_6t
Xbit_r164_c78 bl[78] br[78] wl[164] vdd gnd cell_6t
Xbit_r165_c78 bl[78] br[78] wl[165] vdd gnd cell_6t
Xbit_r166_c78 bl[78] br[78] wl[166] vdd gnd cell_6t
Xbit_r167_c78 bl[78] br[78] wl[167] vdd gnd cell_6t
Xbit_r168_c78 bl[78] br[78] wl[168] vdd gnd cell_6t
Xbit_r169_c78 bl[78] br[78] wl[169] vdd gnd cell_6t
Xbit_r170_c78 bl[78] br[78] wl[170] vdd gnd cell_6t
Xbit_r171_c78 bl[78] br[78] wl[171] vdd gnd cell_6t
Xbit_r172_c78 bl[78] br[78] wl[172] vdd gnd cell_6t
Xbit_r173_c78 bl[78] br[78] wl[173] vdd gnd cell_6t
Xbit_r174_c78 bl[78] br[78] wl[174] vdd gnd cell_6t
Xbit_r175_c78 bl[78] br[78] wl[175] vdd gnd cell_6t
Xbit_r176_c78 bl[78] br[78] wl[176] vdd gnd cell_6t
Xbit_r177_c78 bl[78] br[78] wl[177] vdd gnd cell_6t
Xbit_r178_c78 bl[78] br[78] wl[178] vdd gnd cell_6t
Xbit_r179_c78 bl[78] br[78] wl[179] vdd gnd cell_6t
Xbit_r180_c78 bl[78] br[78] wl[180] vdd gnd cell_6t
Xbit_r181_c78 bl[78] br[78] wl[181] vdd gnd cell_6t
Xbit_r182_c78 bl[78] br[78] wl[182] vdd gnd cell_6t
Xbit_r183_c78 bl[78] br[78] wl[183] vdd gnd cell_6t
Xbit_r184_c78 bl[78] br[78] wl[184] vdd gnd cell_6t
Xbit_r185_c78 bl[78] br[78] wl[185] vdd gnd cell_6t
Xbit_r186_c78 bl[78] br[78] wl[186] vdd gnd cell_6t
Xbit_r187_c78 bl[78] br[78] wl[187] vdd gnd cell_6t
Xbit_r188_c78 bl[78] br[78] wl[188] vdd gnd cell_6t
Xbit_r189_c78 bl[78] br[78] wl[189] vdd gnd cell_6t
Xbit_r190_c78 bl[78] br[78] wl[190] vdd gnd cell_6t
Xbit_r191_c78 bl[78] br[78] wl[191] vdd gnd cell_6t
Xbit_r192_c78 bl[78] br[78] wl[192] vdd gnd cell_6t
Xbit_r193_c78 bl[78] br[78] wl[193] vdd gnd cell_6t
Xbit_r194_c78 bl[78] br[78] wl[194] vdd gnd cell_6t
Xbit_r195_c78 bl[78] br[78] wl[195] vdd gnd cell_6t
Xbit_r196_c78 bl[78] br[78] wl[196] vdd gnd cell_6t
Xbit_r197_c78 bl[78] br[78] wl[197] vdd gnd cell_6t
Xbit_r198_c78 bl[78] br[78] wl[198] vdd gnd cell_6t
Xbit_r199_c78 bl[78] br[78] wl[199] vdd gnd cell_6t
Xbit_r200_c78 bl[78] br[78] wl[200] vdd gnd cell_6t
Xbit_r201_c78 bl[78] br[78] wl[201] vdd gnd cell_6t
Xbit_r202_c78 bl[78] br[78] wl[202] vdd gnd cell_6t
Xbit_r203_c78 bl[78] br[78] wl[203] vdd gnd cell_6t
Xbit_r204_c78 bl[78] br[78] wl[204] vdd gnd cell_6t
Xbit_r205_c78 bl[78] br[78] wl[205] vdd gnd cell_6t
Xbit_r206_c78 bl[78] br[78] wl[206] vdd gnd cell_6t
Xbit_r207_c78 bl[78] br[78] wl[207] vdd gnd cell_6t
Xbit_r208_c78 bl[78] br[78] wl[208] vdd gnd cell_6t
Xbit_r209_c78 bl[78] br[78] wl[209] vdd gnd cell_6t
Xbit_r210_c78 bl[78] br[78] wl[210] vdd gnd cell_6t
Xbit_r211_c78 bl[78] br[78] wl[211] vdd gnd cell_6t
Xbit_r212_c78 bl[78] br[78] wl[212] vdd gnd cell_6t
Xbit_r213_c78 bl[78] br[78] wl[213] vdd gnd cell_6t
Xbit_r214_c78 bl[78] br[78] wl[214] vdd gnd cell_6t
Xbit_r215_c78 bl[78] br[78] wl[215] vdd gnd cell_6t
Xbit_r216_c78 bl[78] br[78] wl[216] vdd gnd cell_6t
Xbit_r217_c78 bl[78] br[78] wl[217] vdd gnd cell_6t
Xbit_r218_c78 bl[78] br[78] wl[218] vdd gnd cell_6t
Xbit_r219_c78 bl[78] br[78] wl[219] vdd gnd cell_6t
Xbit_r220_c78 bl[78] br[78] wl[220] vdd gnd cell_6t
Xbit_r221_c78 bl[78] br[78] wl[221] vdd gnd cell_6t
Xbit_r222_c78 bl[78] br[78] wl[222] vdd gnd cell_6t
Xbit_r223_c78 bl[78] br[78] wl[223] vdd gnd cell_6t
Xbit_r224_c78 bl[78] br[78] wl[224] vdd gnd cell_6t
Xbit_r225_c78 bl[78] br[78] wl[225] vdd gnd cell_6t
Xbit_r226_c78 bl[78] br[78] wl[226] vdd gnd cell_6t
Xbit_r227_c78 bl[78] br[78] wl[227] vdd gnd cell_6t
Xbit_r228_c78 bl[78] br[78] wl[228] vdd gnd cell_6t
Xbit_r229_c78 bl[78] br[78] wl[229] vdd gnd cell_6t
Xbit_r230_c78 bl[78] br[78] wl[230] vdd gnd cell_6t
Xbit_r231_c78 bl[78] br[78] wl[231] vdd gnd cell_6t
Xbit_r232_c78 bl[78] br[78] wl[232] vdd gnd cell_6t
Xbit_r233_c78 bl[78] br[78] wl[233] vdd gnd cell_6t
Xbit_r234_c78 bl[78] br[78] wl[234] vdd gnd cell_6t
Xbit_r235_c78 bl[78] br[78] wl[235] vdd gnd cell_6t
Xbit_r236_c78 bl[78] br[78] wl[236] vdd gnd cell_6t
Xbit_r237_c78 bl[78] br[78] wl[237] vdd gnd cell_6t
Xbit_r238_c78 bl[78] br[78] wl[238] vdd gnd cell_6t
Xbit_r239_c78 bl[78] br[78] wl[239] vdd gnd cell_6t
Xbit_r240_c78 bl[78] br[78] wl[240] vdd gnd cell_6t
Xbit_r241_c78 bl[78] br[78] wl[241] vdd gnd cell_6t
Xbit_r242_c78 bl[78] br[78] wl[242] vdd gnd cell_6t
Xbit_r243_c78 bl[78] br[78] wl[243] vdd gnd cell_6t
Xbit_r244_c78 bl[78] br[78] wl[244] vdd gnd cell_6t
Xbit_r245_c78 bl[78] br[78] wl[245] vdd gnd cell_6t
Xbit_r246_c78 bl[78] br[78] wl[246] vdd gnd cell_6t
Xbit_r247_c78 bl[78] br[78] wl[247] vdd gnd cell_6t
Xbit_r248_c78 bl[78] br[78] wl[248] vdd gnd cell_6t
Xbit_r249_c78 bl[78] br[78] wl[249] vdd gnd cell_6t
Xbit_r250_c78 bl[78] br[78] wl[250] vdd gnd cell_6t
Xbit_r251_c78 bl[78] br[78] wl[251] vdd gnd cell_6t
Xbit_r252_c78 bl[78] br[78] wl[252] vdd gnd cell_6t
Xbit_r253_c78 bl[78] br[78] wl[253] vdd gnd cell_6t
Xbit_r254_c78 bl[78] br[78] wl[254] vdd gnd cell_6t
Xbit_r255_c78 bl[78] br[78] wl[255] vdd gnd cell_6t
Xbit_r0_c79 bl[79] br[79] wl[0] vdd gnd cell_6t
Xbit_r1_c79 bl[79] br[79] wl[1] vdd gnd cell_6t
Xbit_r2_c79 bl[79] br[79] wl[2] vdd gnd cell_6t
Xbit_r3_c79 bl[79] br[79] wl[3] vdd gnd cell_6t
Xbit_r4_c79 bl[79] br[79] wl[4] vdd gnd cell_6t
Xbit_r5_c79 bl[79] br[79] wl[5] vdd gnd cell_6t
Xbit_r6_c79 bl[79] br[79] wl[6] vdd gnd cell_6t
Xbit_r7_c79 bl[79] br[79] wl[7] vdd gnd cell_6t
Xbit_r8_c79 bl[79] br[79] wl[8] vdd gnd cell_6t
Xbit_r9_c79 bl[79] br[79] wl[9] vdd gnd cell_6t
Xbit_r10_c79 bl[79] br[79] wl[10] vdd gnd cell_6t
Xbit_r11_c79 bl[79] br[79] wl[11] vdd gnd cell_6t
Xbit_r12_c79 bl[79] br[79] wl[12] vdd gnd cell_6t
Xbit_r13_c79 bl[79] br[79] wl[13] vdd gnd cell_6t
Xbit_r14_c79 bl[79] br[79] wl[14] vdd gnd cell_6t
Xbit_r15_c79 bl[79] br[79] wl[15] vdd gnd cell_6t
Xbit_r16_c79 bl[79] br[79] wl[16] vdd gnd cell_6t
Xbit_r17_c79 bl[79] br[79] wl[17] vdd gnd cell_6t
Xbit_r18_c79 bl[79] br[79] wl[18] vdd gnd cell_6t
Xbit_r19_c79 bl[79] br[79] wl[19] vdd gnd cell_6t
Xbit_r20_c79 bl[79] br[79] wl[20] vdd gnd cell_6t
Xbit_r21_c79 bl[79] br[79] wl[21] vdd gnd cell_6t
Xbit_r22_c79 bl[79] br[79] wl[22] vdd gnd cell_6t
Xbit_r23_c79 bl[79] br[79] wl[23] vdd gnd cell_6t
Xbit_r24_c79 bl[79] br[79] wl[24] vdd gnd cell_6t
Xbit_r25_c79 bl[79] br[79] wl[25] vdd gnd cell_6t
Xbit_r26_c79 bl[79] br[79] wl[26] vdd gnd cell_6t
Xbit_r27_c79 bl[79] br[79] wl[27] vdd gnd cell_6t
Xbit_r28_c79 bl[79] br[79] wl[28] vdd gnd cell_6t
Xbit_r29_c79 bl[79] br[79] wl[29] vdd gnd cell_6t
Xbit_r30_c79 bl[79] br[79] wl[30] vdd gnd cell_6t
Xbit_r31_c79 bl[79] br[79] wl[31] vdd gnd cell_6t
Xbit_r32_c79 bl[79] br[79] wl[32] vdd gnd cell_6t
Xbit_r33_c79 bl[79] br[79] wl[33] vdd gnd cell_6t
Xbit_r34_c79 bl[79] br[79] wl[34] vdd gnd cell_6t
Xbit_r35_c79 bl[79] br[79] wl[35] vdd gnd cell_6t
Xbit_r36_c79 bl[79] br[79] wl[36] vdd gnd cell_6t
Xbit_r37_c79 bl[79] br[79] wl[37] vdd gnd cell_6t
Xbit_r38_c79 bl[79] br[79] wl[38] vdd gnd cell_6t
Xbit_r39_c79 bl[79] br[79] wl[39] vdd gnd cell_6t
Xbit_r40_c79 bl[79] br[79] wl[40] vdd gnd cell_6t
Xbit_r41_c79 bl[79] br[79] wl[41] vdd gnd cell_6t
Xbit_r42_c79 bl[79] br[79] wl[42] vdd gnd cell_6t
Xbit_r43_c79 bl[79] br[79] wl[43] vdd gnd cell_6t
Xbit_r44_c79 bl[79] br[79] wl[44] vdd gnd cell_6t
Xbit_r45_c79 bl[79] br[79] wl[45] vdd gnd cell_6t
Xbit_r46_c79 bl[79] br[79] wl[46] vdd gnd cell_6t
Xbit_r47_c79 bl[79] br[79] wl[47] vdd gnd cell_6t
Xbit_r48_c79 bl[79] br[79] wl[48] vdd gnd cell_6t
Xbit_r49_c79 bl[79] br[79] wl[49] vdd gnd cell_6t
Xbit_r50_c79 bl[79] br[79] wl[50] vdd gnd cell_6t
Xbit_r51_c79 bl[79] br[79] wl[51] vdd gnd cell_6t
Xbit_r52_c79 bl[79] br[79] wl[52] vdd gnd cell_6t
Xbit_r53_c79 bl[79] br[79] wl[53] vdd gnd cell_6t
Xbit_r54_c79 bl[79] br[79] wl[54] vdd gnd cell_6t
Xbit_r55_c79 bl[79] br[79] wl[55] vdd gnd cell_6t
Xbit_r56_c79 bl[79] br[79] wl[56] vdd gnd cell_6t
Xbit_r57_c79 bl[79] br[79] wl[57] vdd gnd cell_6t
Xbit_r58_c79 bl[79] br[79] wl[58] vdd gnd cell_6t
Xbit_r59_c79 bl[79] br[79] wl[59] vdd gnd cell_6t
Xbit_r60_c79 bl[79] br[79] wl[60] vdd gnd cell_6t
Xbit_r61_c79 bl[79] br[79] wl[61] vdd gnd cell_6t
Xbit_r62_c79 bl[79] br[79] wl[62] vdd gnd cell_6t
Xbit_r63_c79 bl[79] br[79] wl[63] vdd gnd cell_6t
Xbit_r64_c79 bl[79] br[79] wl[64] vdd gnd cell_6t
Xbit_r65_c79 bl[79] br[79] wl[65] vdd gnd cell_6t
Xbit_r66_c79 bl[79] br[79] wl[66] vdd gnd cell_6t
Xbit_r67_c79 bl[79] br[79] wl[67] vdd gnd cell_6t
Xbit_r68_c79 bl[79] br[79] wl[68] vdd gnd cell_6t
Xbit_r69_c79 bl[79] br[79] wl[69] vdd gnd cell_6t
Xbit_r70_c79 bl[79] br[79] wl[70] vdd gnd cell_6t
Xbit_r71_c79 bl[79] br[79] wl[71] vdd gnd cell_6t
Xbit_r72_c79 bl[79] br[79] wl[72] vdd gnd cell_6t
Xbit_r73_c79 bl[79] br[79] wl[73] vdd gnd cell_6t
Xbit_r74_c79 bl[79] br[79] wl[74] vdd gnd cell_6t
Xbit_r75_c79 bl[79] br[79] wl[75] vdd gnd cell_6t
Xbit_r76_c79 bl[79] br[79] wl[76] vdd gnd cell_6t
Xbit_r77_c79 bl[79] br[79] wl[77] vdd gnd cell_6t
Xbit_r78_c79 bl[79] br[79] wl[78] vdd gnd cell_6t
Xbit_r79_c79 bl[79] br[79] wl[79] vdd gnd cell_6t
Xbit_r80_c79 bl[79] br[79] wl[80] vdd gnd cell_6t
Xbit_r81_c79 bl[79] br[79] wl[81] vdd gnd cell_6t
Xbit_r82_c79 bl[79] br[79] wl[82] vdd gnd cell_6t
Xbit_r83_c79 bl[79] br[79] wl[83] vdd gnd cell_6t
Xbit_r84_c79 bl[79] br[79] wl[84] vdd gnd cell_6t
Xbit_r85_c79 bl[79] br[79] wl[85] vdd gnd cell_6t
Xbit_r86_c79 bl[79] br[79] wl[86] vdd gnd cell_6t
Xbit_r87_c79 bl[79] br[79] wl[87] vdd gnd cell_6t
Xbit_r88_c79 bl[79] br[79] wl[88] vdd gnd cell_6t
Xbit_r89_c79 bl[79] br[79] wl[89] vdd gnd cell_6t
Xbit_r90_c79 bl[79] br[79] wl[90] vdd gnd cell_6t
Xbit_r91_c79 bl[79] br[79] wl[91] vdd gnd cell_6t
Xbit_r92_c79 bl[79] br[79] wl[92] vdd gnd cell_6t
Xbit_r93_c79 bl[79] br[79] wl[93] vdd gnd cell_6t
Xbit_r94_c79 bl[79] br[79] wl[94] vdd gnd cell_6t
Xbit_r95_c79 bl[79] br[79] wl[95] vdd gnd cell_6t
Xbit_r96_c79 bl[79] br[79] wl[96] vdd gnd cell_6t
Xbit_r97_c79 bl[79] br[79] wl[97] vdd gnd cell_6t
Xbit_r98_c79 bl[79] br[79] wl[98] vdd gnd cell_6t
Xbit_r99_c79 bl[79] br[79] wl[99] vdd gnd cell_6t
Xbit_r100_c79 bl[79] br[79] wl[100] vdd gnd cell_6t
Xbit_r101_c79 bl[79] br[79] wl[101] vdd gnd cell_6t
Xbit_r102_c79 bl[79] br[79] wl[102] vdd gnd cell_6t
Xbit_r103_c79 bl[79] br[79] wl[103] vdd gnd cell_6t
Xbit_r104_c79 bl[79] br[79] wl[104] vdd gnd cell_6t
Xbit_r105_c79 bl[79] br[79] wl[105] vdd gnd cell_6t
Xbit_r106_c79 bl[79] br[79] wl[106] vdd gnd cell_6t
Xbit_r107_c79 bl[79] br[79] wl[107] vdd gnd cell_6t
Xbit_r108_c79 bl[79] br[79] wl[108] vdd gnd cell_6t
Xbit_r109_c79 bl[79] br[79] wl[109] vdd gnd cell_6t
Xbit_r110_c79 bl[79] br[79] wl[110] vdd gnd cell_6t
Xbit_r111_c79 bl[79] br[79] wl[111] vdd gnd cell_6t
Xbit_r112_c79 bl[79] br[79] wl[112] vdd gnd cell_6t
Xbit_r113_c79 bl[79] br[79] wl[113] vdd gnd cell_6t
Xbit_r114_c79 bl[79] br[79] wl[114] vdd gnd cell_6t
Xbit_r115_c79 bl[79] br[79] wl[115] vdd gnd cell_6t
Xbit_r116_c79 bl[79] br[79] wl[116] vdd gnd cell_6t
Xbit_r117_c79 bl[79] br[79] wl[117] vdd gnd cell_6t
Xbit_r118_c79 bl[79] br[79] wl[118] vdd gnd cell_6t
Xbit_r119_c79 bl[79] br[79] wl[119] vdd gnd cell_6t
Xbit_r120_c79 bl[79] br[79] wl[120] vdd gnd cell_6t
Xbit_r121_c79 bl[79] br[79] wl[121] vdd gnd cell_6t
Xbit_r122_c79 bl[79] br[79] wl[122] vdd gnd cell_6t
Xbit_r123_c79 bl[79] br[79] wl[123] vdd gnd cell_6t
Xbit_r124_c79 bl[79] br[79] wl[124] vdd gnd cell_6t
Xbit_r125_c79 bl[79] br[79] wl[125] vdd gnd cell_6t
Xbit_r126_c79 bl[79] br[79] wl[126] vdd gnd cell_6t
Xbit_r127_c79 bl[79] br[79] wl[127] vdd gnd cell_6t
Xbit_r128_c79 bl[79] br[79] wl[128] vdd gnd cell_6t
Xbit_r129_c79 bl[79] br[79] wl[129] vdd gnd cell_6t
Xbit_r130_c79 bl[79] br[79] wl[130] vdd gnd cell_6t
Xbit_r131_c79 bl[79] br[79] wl[131] vdd gnd cell_6t
Xbit_r132_c79 bl[79] br[79] wl[132] vdd gnd cell_6t
Xbit_r133_c79 bl[79] br[79] wl[133] vdd gnd cell_6t
Xbit_r134_c79 bl[79] br[79] wl[134] vdd gnd cell_6t
Xbit_r135_c79 bl[79] br[79] wl[135] vdd gnd cell_6t
Xbit_r136_c79 bl[79] br[79] wl[136] vdd gnd cell_6t
Xbit_r137_c79 bl[79] br[79] wl[137] vdd gnd cell_6t
Xbit_r138_c79 bl[79] br[79] wl[138] vdd gnd cell_6t
Xbit_r139_c79 bl[79] br[79] wl[139] vdd gnd cell_6t
Xbit_r140_c79 bl[79] br[79] wl[140] vdd gnd cell_6t
Xbit_r141_c79 bl[79] br[79] wl[141] vdd gnd cell_6t
Xbit_r142_c79 bl[79] br[79] wl[142] vdd gnd cell_6t
Xbit_r143_c79 bl[79] br[79] wl[143] vdd gnd cell_6t
Xbit_r144_c79 bl[79] br[79] wl[144] vdd gnd cell_6t
Xbit_r145_c79 bl[79] br[79] wl[145] vdd gnd cell_6t
Xbit_r146_c79 bl[79] br[79] wl[146] vdd gnd cell_6t
Xbit_r147_c79 bl[79] br[79] wl[147] vdd gnd cell_6t
Xbit_r148_c79 bl[79] br[79] wl[148] vdd gnd cell_6t
Xbit_r149_c79 bl[79] br[79] wl[149] vdd gnd cell_6t
Xbit_r150_c79 bl[79] br[79] wl[150] vdd gnd cell_6t
Xbit_r151_c79 bl[79] br[79] wl[151] vdd gnd cell_6t
Xbit_r152_c79 bl[79] br[79] wl[152] vdd gnd cell_6t
Xbit_r153_c79 bl[79] br[79] wl[153] vdd gnd cell_6t
Xbit_r154_c79 bl[79] br[79] wl[154] vdd gnd cell_6t
Xbit_r155_c79 bl[79] br[79] wl[155] vdd gnd cell_6t
Xbit_r156_c79 bl[79] br[79] wl[156] vdd gnd cell_6t
Xbit_r157_c79 bl[79] br[79] wl[157] vdd gnd cell_6t
Xbit_r158_c79 bl[79] br[79] wl[158] vdd gnd cell_6t
Xbit_r159_c79 bl[79] br[79] wl[159] vdd gnd cell_6t
Xbit_r160_c79 bl[79] br[79] wl[160] vdd gnd cell_6t
Xbit_r161_c79 bl[79] br[79] wl[161] vdd gnd cell_6t
Xbit_r162_c79 bl[79] br[79] wl[162] vdd gnd cell_6t
Xbit_r163_c79 bl[79] br[79] wl[163] vdd gnd cell_6t
Xbit_r164_c79 bl[79] br[79] wl[164] vdd gnd cell_6t
Xbit_r165_c79 bl[79] br[79] wl[165] vdd gnd cell_6t
Xbit_r166_c79 bl[79] br[79] wl[166] vdd gnd cell_6t
Xbit_r167_c79 bl[79] br[79] wl[167] vdd gnd cell_6t
Xbit_r168_c79 bl[79] br[79] wl[168] vdd gnd cell_6t
Xbit_r169_c79 bl[79] br[79] wl[169] vdd gnd cell_6t
Xbit_r170_c79 bl[79] br[79] wl[170] vdd gnd cell_6t
Xbit_r171_c79 bl[79] br[79] wl[171] vdd gnd cell_6t
Xbit_r172_c79 bl[79] br[79] wl[172] vdd gnd cell_6t
Xbit_r173_c79 bl[79] br[79] wl[173] vdd gnd cell_6t
Xbit_r174_c79 bl[79] br[79] wl[174] vdd gnd cell_6t
Xbit_r175_c79 bl[79] br[79] wl[175] vdd gnd cell_6t
Xbit_r176_c79 bl[79] br[79] wl[176] vdd gnd cell_6t
Xbit_r177_c79 bl[79] br[79] wl[177] vdd gnd cell_6t
Xbit_r178_c79 bl[79] br[79] wl[178] vdd gnd cell_6t
Xbit_r179_c79 bl[79] br[79] wl[179] vdd gnd cell_6t
Xbit_r180_c79 bl[79] br[79] wl[180] vdd gnd cell_6t
Xbit_r181_c79 bl[79] br[79] wl[181] vdd gnd cell_6t
Xbit_r182_c79 bl[79] br[79] wl[182] vdd gnd cell_6t
Xbit_r183_c79 bl[79] br[79] wl[183] vdd gnd cell_6t
Xbit_r184_c79 bl[79] br[79] wl[184] vdd gnd cell_6t
Xbit_r185_c79 bl[79] br[79] wl[185] vdd gnd cell_6t
Xbit_r186_c79 bl[79] br[79] wl[186] vdd gnd cell_6t
Xbit_r187_c79 bl[79] br[79] wl[187] vdd gnd cell_6t
Xbit_r188_c79 bl[79] br[79] wl[188] vdd gnd cell_6t
Xbit_r189_c79 bl[79] br[79] wl[189] vdd gnd cell_6t
Xbit_r190_c79 bl[79] br[79] wl[190] vdd gnd cell_6t
Xbit_r191_c79 bl[79] br[79] wl[191] vdd gnd cell_6t
Xbit_r192_c79 bl[79] br[79] wl[192] vdd gnd cell_6t
Xbit_r193_c79 bl[79] br[79] wl[193] vdd gnd cell_6t
Xbit_r194_c79 bl[79] br[79] wl[194] vdd gnd cell_6t
Xbit_r195_c79 bl[79] br[79] wl[195] vdd gnd cell_6t
Xbit_r196_c79 bl[79] br[79] wl[196] vdd gnd cell_6t
Xbit_r197_c79 bl[79] br[79] wl[197] vdd gnd cell_6t
Xbit_r198_c79 bl[79] br[79] wl[198] vdd gnd cell_6t
Xbit_r199_c79 bl[79] br[79] wl[199] vdd gnd cell_6t
Xbit_r200_c79 bl[79] br[79] wl[200] vdd gnd cell_6t
Xbit_r201_c79 bl[79] br[79] wl[201] vdd gnd cell_6t
Xbit_r202_c79 bl[79] br[79] wl[202] vdd gnd cell_6t
Xbit_r203_c79 bl[79] br[79] wl[203] vdd gnd cell_6t
Xbit_r204_c79 bl[79] br[79] wl[204] vdd gnd cell_6t
Xbit_r205_c79 bl[79] br[79] wl[205] vdd gnd cell_6t
Xbit_r206_c79 bl[79] br[79] wl[206] vdd gnd cell_6t
Xbit_r207_c79 bl[79] br[79] wl[207] vdd gnd cell_6t
Xbit_r208_c79 bl[79] br[79] wl[208] vdd gnd cell_6t
Xbit_r209_c79 bl[79] br[79] wl[209] vdd gnd cell_6t
Xbit_r210_c79 bl[79] br[79] wl[210] vdd gnd cell_6t
Xbit_r211_c79 bl[79] br[79] wl[211] vdd gnd cell_6t
Xbit_r212_c79 bl[79] br[79] wl[212] vdd gnd cell_6t
Xbit_r213_c79 bl[79] br[79] wl[213] vdd gnd cell_6t
Xbit_r214_c79 bl[79] br[79] wl[214] vdd gnd cell_6t
Xbit_r215_c79 bl[79] br[79] wl[215] vdd gnd cell_6t
Xbit_r216_c79 bl[79] br[79] wl[216] vdd gnd cell_6t
Xbit_r217_c79 bl[79] br[79] wl[217] vdd gnd cell_6t
Xbit_r218_c79 bl[79] br[79] wl[218] vdd gnd cell_6t
Xbit_r219_c79 bl[79] br[79] wl[219] vdd gnd cell_6t
Xbit_r220_c79 bl[79] br[79] wl[220] vdd gnd cell_6t
Xbit_r221_c79 bl[79] br[79] wl[221] vdd gnd cell_6t
Xbit_r222_c79 bl[79] br[79] wl[222] vdd gnd cell_6t
Xbit_r223_c79 bl[79] br[79] wl[223] vdd gnd cell_6t
Xbit_r224_c79 bl[79] br[79] wl[224] vdd gnd cell_6t
Xbit_r225_c79 bl[79] br[79] wl[225] vdd gnd cell_6t
Xbit_r226_c79 bl[79] br[79] wl[226] vdd gnd cell_6t
Xbit_r227_c79 bl[79] br[79] wl[227] vdd gnd cell_6t
Xbit_r228_c79 bl[79] br[79] wl[228] vdd gnd cell_6t
Xbit_r229_c79 bl[79] br[79] wl[229] vdd gnd cell_6t
Xbit_r230_c79 bl[79] br[79] wl[230] vdd gnd cell_6t
Xbit_r231_c79 bl[79] br[79] wl[231] vdd gnd cell_6t
Xbit_r232_c79 bl[79] br[79] wl[232] vdd gnd cell_6t
Xbit_r233_c79 bl[79] br[79] wl[233] vdd gnd cell_6t
Xbit_r234_c79 bl[79] br[79] wl[234] vdd gnd cell_6t
Xbit_r235_c79 bl[79] br[79] wl[235] vdd gnd cell_6t
Xbit_r236_c79 bl[79] br[79] wl[236] vdd gnd cell_6t
Xbit_r237_c79 bl[79] br[79] wl[237] vdd gnd cell_6t
Xbit_r238_c79 bl[79] br[79] wl[238] vdd gnd cell_6t
Xbit_r239_c79 bl[79] br[79] wl[239] vdd gnd cell_6t
Xbit_r240_c79 bl[79] br[79] wl[240] vdd gnd cell_6t
Xbit_r241_c79 bl[79] br[79] wl[241] vdd gnd cell_6t
Xbit_r242_c79 bl[79] br[79] wl[242] vdd gnd cell_6t
Xbit_r243_c79 bl[79] br[79] wl[243] vdd gnd cell_6t
Xbit_r244_c79 bl[79] br[79] wl[244] vdd gnd cell_6t
Xbit_r245_c79 bl[79] br[79] wl[245] vdd gnd cell_6t
Xbit_r246_c79 bl[79] br[79] wl[246] vdd gnd cell_6t
Xbit_r247_c79 bl[79] br[79] wl[247] vdd gnd cell_6t
Xbit_r248_c79 bl[79] br[79] wl[248] vdd gnd cell_6t
Xbit_r249_c79 bl[79] br[79] wl[249] vdd gnd cell_6t
Xbit_r250_c79 bl[79] br[79] wl[250] vdd gnd cell_6t
Xbit_r251_c79 bl[79] br[79] wl[251] vdd gnd cell_6t
Xbit_r252_c79 bl[79] br[79] wl[252] vdd gnd cell_6t
Xbit_r253_c79 bl[79] br[79] wl[253] vdd gnd cell_6t
Xbit_r254_c79 bl[79] br[79] wl[254] vdd gnd cell_6t
Xbit_r255_c79 bl[79] br[79] wl[255] vdd gnd cell_6t
Xbit_r0_c80 bl[80] br[80] wl[0] vdd gnd cell_6t
Xbit_r1_c80 bl[80] br[80] wl[1] vdd gnd cell_6t
Xbit_r2_c80 bl[80] br[80] wl[2] vdd gnd cell_6t
Xbit_r3_c80 bl[80] br[80] wl[3] vdd gnd cell_6t
Xbit_r4_c80 bl[80] br[80] wl[4] vdd gnd cell_6t
Xbit_r5_c80 bl[80] br[80] wl[5] vdd gnd cell_6t
Xbit_r6_c80 bl[80] br[80] wl[6] vdd gnd cell_6t
Xbit_r7_c80 bl[80] br[80] wl[7] vdd gnd cell_6t
Xbit_r8_c80 bl[80] br[80] wl[8] vdd gnd cell_6t
Xbit_r9_c80 bl[80] br[80] wl[9] vdd gnd cell_6t
Xbit_r10_c80 bl[80] br[80] wl[10] vdd gnd cell_6t
Xbit_r11_c80 bl[80] br[80] wl[11] vdd gnd cell_6t
Xbit_r12_c80 bl[80] br[80] wl[12] vdd gnd cell_6t
Xbit_r13_c80 bl[80] br[80] wl[13] vdd gnd cell_6t
Xbit_r14_c80 bl[80] br[80] wl[14] vdd gnd cell_6t
Xbit_r15_c80 bl[80] br[80] wl[15] vdd gnd cell_6t
Xbit_r16_c80 bl[80] br[80] wl[16] vdd gnd cell_6t
Xbit_r17_c80 bl[80] br[80] wl[17] vdd gnd cell_6t
Xbit_r18_c80 bl[80] br[80] wl[18] vdd gnd cell_6t
Xbit_r19_c80 bl[80] br[80] wl[19] vdd gnd cell_6t
Xbit_r20_c80 bl[80] br[80] wl[20] vdd gnd cell_6t
Xbit_r21_c80 bl[80] br[80] wl[21] vdd gnd cell_6t
Xbit_r22_c80 bl[80] br[80] wl[22] vdd gnd cell_6t
Xbit_r23_c80 bl[80] br[80] wl[23] vdd gnd cell_6t
Xbit_r24_c80 bl[80] br[80] wl[24] vdd gnd cell_6t
Xbit_r25_c80 bl[80] br[80] wl[25] vdd gnd cell_6t
Xbit_r26_c80 bl[80] br[80] wl[26] vdd gnd cell_6t
Xbit_r27_c80 bl[80] br[80] wl[27] vdd gnd cell_6t
Xbit_r28_c80 bl[80] br[80] wl[28] vdd gnd cell_6t
Xbit_r29_c80 bl[80] br[80] wl[29] vdd gnd cell_6t
Xbit_r30_c80 bl[80] br[80] wl[30] vdd gnd cell_6t
Xbit_r31_c80 bl[80] br[80] wl[31] vdd gnd cell_6t
Xbit_r32_c80 bl[80] br[80] wl[32] vdd gnd cell_6t
Xbit_r33_c80 bl[80] br[80] wl[33] vdd gnd cell_6t
Xbit_r34_c80 bl[80] br[80] wl[34] vdd gnd cell_6t
Xbit_r35_c80 bl[80] br[80] wl[35] vdd gnd cell_6t
Xbit_r36_c80 bl[80] br[80] wl[36] vdd gnd cell_6t
Xbit_r37_c80 bl[80] br[80] wl[37] vdd gnd cell_6t
Xbit_r38_c80 bl[80] br[80] wl[38] vdd gnd cell_6t
Xbit_r39_c80 bl[80] br[80] wl[39] vdd gnd cell_6t
Xbit_r40_c80 bl[80] br[80] wl[40] vdd gnd cell_6t
Xbit_r41_c80 bl[80] br[80] wl[41] vdd gnd cell_6t
Xbit_r42_c80 bl[80] br[80] wl[42] vdd gnd cell_6t
Xbit_r43_c80 bl[80] br[80] wl[43] vdd gnd cell_6t
Xbit_r44_c80 bl[80] br[80] wl[44] vdd gnd cell_6t
Xbit_r45_c80 bl[80] br[80] wl[45] vdd gnd cell_6t
Xbit_r46_c80 bl[80] br[80] wl[46] vdd gnd cell_6t
Xbit_r47_c80 bl[80] br[80] wl[47] vdd gnd cell_6t
Xbit_r48_c80 bl[80] br[80] wl[48] vdd gnd cell_6t
Xbit_r49_c80 bl[80] br[80] wl[49] vdd gnd cell_6t
Xbit_r50_c80 bl[80] br[80] wl[50] vdd gnd cell_6t
Xbit_r51_c80 bl[80] br[80] wl[51] vdd gnd cell_6t
Xbit_r52_c80 bl[80] br[80] wl[52] vdd gnd cell_6t
Xbit_r53_c80 bl[80] br[80] wl[53] vdd gnd cell_6t
Xbit_r54_c80 bl[80] br[80] wl[54] vdd gnd cell_6t
Xbit_r55_c80 bl[80] br[80] wl[55] vdd gnd cell_6t
Xbit_r56_c80 bl[80] br[80] wl[56] vdd gnd cell_6t
Xbit_r57_c80 bl[80] br[80] wl[57] vdd gnd cell_6t
Xbit_r58_c80 bl[80] br[80] wl[58] vdd gnd cell_6t
Xbit_r59_c80 bl[80] br[80] wl[59] vdd gnd cell_6t
Xbit_r60_c80 bl[80] br[80] wl[60] vdd gnd cell_6t
Xbit_r61_c80 bl[80] br[80] wl[61] vdd gnd cell_6t
Xbit_r62_c80 bl[80] br[80] wl[62] vdd gnd cell_6t
Xbit_r63_c80 bl[80] br[80] wl[63] vdd gnd cell_6t
Xbit_r64_c80 bl[80] br[80] wl[64] vdd gnd cell_6t
Xbit_r65_c80 bl[80] br[80] wl[65] vdd gnd cell_6t
Xbit_r66_c80 bl[80] br[80] wl[66] vdd gnd cell_6t
Xbit_r67_c80 bl[80] br[80] wl[67] vdd gnd cell_6t
Xbit_r68_c80 bl[80] br[80] wl[68] vdd gnd cell_6t
Xbit_r69_c80 bl[80] br[80] wl[69] vdd gnd cell_6t
Xbit_r70_c80 bl[80] br[80] wl[70] vdd gnd cell_6t
Xbit_r71_c80 bl[80] br[80] wl[71] vdd gnd cell_6t
Xbit_r72_c80 bl[80] br[80] wl[72] vdd gnd cell_6t
Xbit_r73_c80 bl[80] br[80] wl[73] vdd gnd cell_6t
Xbit_r74_c80 bl[80] br[80] wl[74] vdd gnd cell_6t
Xbit_r75_c80 bl[80] br[80] wl[75] vdd gnd cell_6t
Xbit_r76_c80 bl[80] br[80] wl[76] vdd gnd cell_6t
Xbit_r77_c80 bl[80] br[80] wl[77] vdd gnd cell_6t
Xbit_r78_c80 bl[80] br[80] wl[78] vdd gnd cell_6t
Xbit_r79_c80 bl[80] br[80] wl[79] vdd gnd cell_6t
Xbit_r80_c80 bl[80] br[80] wl[80] vdd gnd cell_6t
Xbit_r81_c80 bl[80] br[80] wl[81] vdd gnd cell_6t
Xbit_r82_c80 bl[80] br[80] wl[82] vdd gnd cell_6t
Xbit_r83_c80 bl[80] br[80] wl[83] vdd gnd cell_6t
Xbit_r84_c80 bl[80] br[80] wl[84] vdd gnd cell_6t
Xbit_r85_c80 bl[80] br[80] wl[85] vdd gnd cell_6t
Xbit_r86_c80 bl[80] br[80] wl[86] vdd gnd cell_6t
Xbit_r87_c80 bl[80] br[80] wl[87] vdd gnd cell_6t
Xbit_r88_c80 bl[80] br[80] wl[88] vdd gnd cell_6t
Xbit_r89_c80 bl[80] br[80] wl[89] vdd gnd cell_6t
Xbit_r90_c80 bl[80] br[80] wl[90] vdd gnd cell_6t
Xbit_r91_c80 bl[80] br[80] wl[91] vdd gnd cell_6t
Xbit_r92_c80 bl[80] br[80] wl[92] vdd gnd cell_6t
Xbit_r93_c80 bl[80] br[80] wl[93] vdd gnd cell_6t
Xbit_r94_c80 bl[80] br[80] wl[94] vdd gnd cell_6t
Xbit_r95_c80 bl[80] br[80] wl[95] vdd gnd cell_6t
Xbit_r96_c80 bl[80] br[80] wl[96] vdd gnd cell_6t
Xbit_r97_c80 bl[80] br[80] wl[97] vdd gnd cell_6t
Xbit_r98_c80 bl[80] br[80] wl[98] vdd gnd cell_6t
Xbit_r99_c80 bl[80] br[80] wl[99] vdd gnd cell_6t
Xbit_r100_c80 bl[80] br[80] wl[100] vdd gnd cell_6t
Xbit_r101_c80 bl[80] br[80] wl[101] vdd gnd cell_6t
Xbit_r102_c80 bl[80] br[80] wl[102] vdd gnd cell_6t
Xbit_r103_c80 bl[80] br[80] wl[103] vdd gnd cell_6t
Xbit_r104_c80 bl[80] br[80] wl[104] vdd gnd cell_6t
Xbit_r105_c80 bl[80] br[80] wl[105] vdd gnd cell_6t
Xbit_r106_c80 bl[80] br[80] wl[106] vdd gnd cell_6t
Xbit_r107_c80 bl[80] br[80] wl[107] vdd gnd cell_6t
Xbit_r108_c80 bl[80] br[80] wl[108] vdd gnd cell_6t
Xbit_r109_c80 bl[80] br[80] wl[109] vdd gnd cell_6t
Xbit_r110_c80 bl[80] br[80] wl[110] vdd gnd cell_6t
Xbit_r111_c80 bl[80] br[80] wl[111] vdd gnd cell_6t
Xbit_r112_c80 bl[80] br[80] wl[112] vdd gnd cell_6t
Xbit_r113_c80 bl[80] br[80] wl[113] vdd gnd cell_6t
Xbit_r114_c80 bl[80] br[80] wl[114] vdd gnd cell_6t
Xbit_r115_c80 bl[80] br[80] wl[115] vdd gnd cell_6t
Xbit_r116_c80 bl[80] br[80] wl[116] vdd gnd cell_6t
Xbit_r117_c80 bl[80] br[80] wl[117] vdd gnd cell_6t
Xbit_r118_c80 bl[80] br[80] wl[118] vdd gnd cell_6t
Xbit_r119_c80 bl[80] br[80] wl[119] vdd gnd cell_6t
Xbit_r120_c80 bl[80] br[80] wl[120] vdd gnd cell_6t
Xbit_r121_c80 bl[80] br[80] wl[121] vdd gnd cell_6t
Xbit_r122_c80 bl[80] br[80] wl[122] vdd gnd cell_6t
Xbit_r123_c80 bl[80] br[80] wl[123] vdd gnd cell_6t
Xbit_r124_c80 bl[80] br[80] wl[124] vdd gnd cell_6t
Xbit_r125_c80 bl[80] br[80] wl[125] vdd gnd cell_6t
Xbit_r126_c80 bl[80] br[80] wl[126] vdd gnd cell_6t
Xbit_r127_c80 bl[80] br[80] wl[127] vdd gnd cell_6t
Xbit_r128_c80 bl[80] br[80] wl[128] vdd gnd cell_6t
Xbit_r129_c80 bl[80] br[80] wl[129] vdd gnd cell_6t
Xbit_r130_c80 bl[80] br[80] wl[130] vdd gnd cell_6t
Xbit_r131_c80 bl[80] br[80] wl[131] vdd gnd cell_6t
Xbit_r132_c80 bl[80] br[80] wl[132] vdd gnd cell_6t
Xbit_r133_c80 bl[80] br[80] wl[133] vdd gnd cell_6t
Xbit_r134_c80 bl[80] br[80] wl[134] vdd gnd cell_6t
Xbit_r135_c80 bl[80] br[80] wl[135] vdd gnd cell_6t
Xbit_r136_c80 bl[80] br[80] wl[136] vdd gnd cell_6t
Xbit_r137_c80 bl[80] br[80] wl[137] vdd gnd cell_6t
Xbit_r138_c80 bl[80] br[80] wl[138] vdd gnd cell_6t
Xbit_r139_c80 bl[80] br[80] wl[139] vdd gnd cell_6t
Xbit_r140_c80 bl[80] br[80] wl[140] vdd gnd cell_6t
Xbit_r141_c80 bl[80] br[80] wl[141] vdd gnd cell_6t
Xbit_r142_c80 bl[80] br[80] wl[142] vdd gnd cell_6t
Xbit_r143_c80 bl[80] br[80] wl[143] vdd gnd cell_6t
Xbit_r144_c80 bl[80] br[80] wl[144] vdd gnd cell_6t
Xbit_r145_c80 bl[80] br[80] wl[145] vdd gnd cell_6t
Xbit_r146_c80 bl[80] br[80] wl[146] vdd gnd cell_6t
Xbit_r147_c80 bl[80] br[80] wl[147] vdd gnd cell_6t
Xbit_r148_c80 bl[80] br[80] wl[148] vdd gnd cell_6t
Xbit_r149_c80 bl[80] br[80] wl[149] vdd gnd cell_6t
Xbit_r150_c80 bl[80] br[80] wl[150] vdd gnd cell_6t
Xbit_r151_c80 bl[80] br[80] wl[151] vdd gnd cell_6t
Xbit_r152_c80 bl[80] br[80] wl[152] vdd gnd cell_6t
Xbit_r153_c80 bl[80] br[80] wl[153] vdd gnd cell_6t
Xbit_r154_c80 bl[80] br[80] wl[154] vdd gnd cell_6t
Xbit_r155_c80 bl[80] br[80] wl[155] vdd gnd cell_6t
Xbit_r156_c80 bl[80] br[80] wl[156] vdd gnd cell_6t
Xbit_r157_c80 bl[80] br[80] wl[157] vdd gnd cell_6t
Xbit_r158_c80 bl[80] br[80] wl[158] vdd gnd cell_6t
Xbit_r159_c80 bl[80] br[80] wl[159] vdd gnd cell_6t
Xbit_r160_c80 bl[80] br[80] wl[160] vdd gnd cell_6t
Xbit_r161_c80 bl[80] br[80] wl[161] vdd gnd cell_6t
Xbit_r162_c80 bl[80] br[80] wl[162] vdd gnd cell_6t
Xbit_r163_c80 bl[80] br[80] wl[163] vdd gnd cell_6t
Xbit_r164_c80 bl[80] br[80] wl[164] vdd gnd cell_6t
Xbit_r165_c80 bl[80] br[80] wl[165] vdd gnd cell_6t
Xbit_r166_c80 bl[80] br[80] wl[166] vdd gnd cell_6t
Xbit_r167_c80 bl[80] br[80] wl[167] vdd gnd cell_6t
Xbit_r168_c80 bl[80] br[80] wl[168] vdd gnd cell_6t
Xbit_r169_c80 bl[80] br[80] wl[169] vdd gnd cell_6t
Xbit_r170_c80 bl[80] br[80] wl[170] vdd gnd cell_6t
Xbit_r171_c80 bl[80] br[80] wl[171] vdd gnd cell_6t
Xbit_r172_c80 bl[80] br[80] wl[172] vdd gnd cell_6t
Xbit_r173_c80 bl[80] br[80] wl[173] vdd gnd cell_6t
Xbit_r174_c80 bl[80] br[80] wl[174] vdd gnd cell_6t
Xbit_r175_c80 bl[80] br[80] wl[175] vdd gnd cell_6t
Xbit_r176_c80 bl[80] br[80] wl[176] vdd gnd cell_6t
Xbit_r177_c80 bl[80] br[80] wl[177] vdd gnd cell_6t
Xbit_r178_c80 bl[80] br[80] wl[178] vdd gnd cell_6t
Xbit_r179_c80 bl[80] br[80] wl[179] vdd gnd cell_6t
Xbit_r180_c80 bl[80] br[80] wl[180] vdd gnd cell_6t
Xbit_r181_c80 bl[80] br[80] wl[181] vdd gnd cell_6t
Xbit_r182_c80 bl[80] br[80] wl[182] vdd gnd cell_6t
Xbit_r183_c80 bl[80] br[80] wl[183] vdd gnd cell_6t
Xbit_r184_c80 bl[80] br[80] wl[184] vdd gnd cell_6t
Xbit_r185_c80 bl[80] br[80] wl[185] vdd gnd cell_6t
Xbit_r186_c80 bl[80] br[80] wl[186] vdd gnd cell_6t
Xbit_r187_c80 bl[80] br[80] wl[187] vdd gnd cell_6t
Xbit_r188_c80 bl[80] br[80] wl[188] vdd gnd cell_6t
Xbit_r189_c80 bl[80] br[80] wl[189] vdd gnd cell_6t
Xbit_r190_c80 bl[80] br[80] wl[190] vdd gnd cell_6t
Xbit_r191_c80 bl[80] br[80] wl[191] vdd gnd cell_6t
Xbit_r192_c80 bl[80] br[80] wl[192] vdd gnd cell_6t
Xbit_r193_c80 bl[80] br[80] wl[193] vdd gnd cell_6t
Xbit_r194_c80 bl[80] br[80] wl[194] vdd gnd cell_6t
Xbit_r195_c80 bl[80] br[80] wl[195] vdd gnd cell_6t
Xbit_r196_c80 bl[80] br[80] wl[196] vdd gnd cell_6t
Xbit_r197_c80 bl[80] br[80] wl[197] vdd gnd cell_6t
Xbit_r198_c80 bl[80] br[80] wl[198] vdd gnd cell_6t
Xbit_r199_c80 bl[80] br[80] wl[199] vdd gnd cell_6t
Xbit_r200_c80 bl[80] br[80] wl[200] vdd gnd cell_6t
Xbit_r201_c80 bl[80] br[80] wl[201] vdd gnd cell_6t
Xbit_r202_c80 bl[80] br[80] wl[202] vdd gnd cell_6t
Xbit_r203_c80 bl[80] br[80] wl[203] vdd gnd cell_6t
Xbit_r204_c80 bl[80] br[80] wl[204] vdd gnd cell_6t
Xbit_r205_c80 bl[80] br[80] wl[205] vdd gnd cell_6t
Xbit_r206_c80 bl[80] br[80] wl[206] vdd gnd cell_6t
Xbit_r207_c80 bl[80] br[80] wl[207] vdd gnd cell_6t
Xbit_r208_c80 bl[80] br[80] wl[208] vdd gnd cell_6t
Xbit_r209_c80 bl[80] br[80] wl[209] vdd gnd cell_6t
Xbit_r210_c80 bl[80] br[80] wl[210] vdd gnd cell_6t
Xbit_r211_c80 bl[80] br[80] wl[211] vdd gnd cell_6t
Xbit_r212_c80 bl[80] br[80] wl[212] vdd gnd cell_6t
Xbit_r213_c80 bl[80] br[80] wl[213] vdd gnd cell_6t
Xbit_r214_c80 bl[80] br[80] wl[214] vdd gnd cell_6t
Xbit_r215_c80 bl[80] br[80] wl[215] vdd gnd cell_6t
Xbit_r216_c80 bl[80] br[80] wl[216] vdd gnd cell_6t
Xbit_r217_c80 bl[80] br[80] wl[217] vdd gnd cell_6t
Xbit_r218_c80 bl[80] br[80] wl[218] vdd gnd cell_6t
Xbit_r219_c80 bl[80] br[80] wl[219] vdd gnd cell_6t
Xbit_r220_c80 bl[80] br[80] wl[220] vdd gnd cell_6t
Xbit_r221_c80 bl[80] br[80] wl[221] vdd gnd cell_6t
Xbit_r222_c80 bl[80] br[80] wl[222] vdd gnd cell_6t
Xbit_r223_c80 bl[80] br[80] wl[223] vdd gnd cell_6t
Xbit_r224_c80 bl[80] br[80] wl[224] vdd gnd cell_6t
Xbit_r225_c80 bl[80] br[80] wl[225] vdd gnd cell_6t
Xbit_r226_c80 bl[80] br[80] wl[226] vdd gnd cell_6t
Xbit_r227_c80 bl[80] br[80] wl[227] vdd gnd cell_6t
Xbit_r228_c80 bl[80] br[80] wl[228] vdd gnd cell_6t
Xbit_r229_c80 bl[80] br[80] wl[229] vdd gnd cell_6t
Xbit_r230_c80 bl[80] br[80] wl[230] vdd gnd cell_6t
Xbit_r231_c80 bl[80] br[80] wl[231] vdd gnd cell_6t
Xbit_r232_c80 bl[80] br[80] wl[232] vdd gnd cell_6t
Xbit_r233_c80 bl[80] br[80] wl[233] vdd gnd cell_6t
Xbit_r234_c80 bl[80] br[80] wl[234] vdd gnd cell_6t
Xbit_r235_c80 bl[80] br[80] wl[235] vdd gnd cell_6t
Xbit_r236_c80 bl[80] br[80] wl[236] vdd gnd cell_6t
Xbit_r237_c80 bl[80] br[80] wl[237] vdd gnd cell_6t
Xbit_r238_c80 bl[80] br[80] wl[238] vdd gnd cell_6t
Xbit_r239_c80 bl[80] br[80] wl[239] vdd gnd cell_6t
Xbit_r240_c80 bl[80] br[80] wl[240] vdd gnd cell_6t
Xbit_r241_c80 bl[80] br[80] wl[241] vdd gnd cell_6t
Xbit_r242_c80 bl[80] br[80] wl[242] vdd gnd cell_6t
Xbit_r243_c80 bl[80] br[80] wl[243] vdd gnd cell_6t
Xbit_r244_c80 bl[80] br[80] wl[244] vdd gnd cell_6t
Xbit_r245_c80 bl[80] br[80] wl[245] vdd gnd cell_6t
Xbit_r246_c80 bl[80] br[80] wl[246] vdd gnd cell_6t
Xbit_r247_c80 bl[80] br[80] wl[247] vdd gnd cell_6t
Xbit_r248_c80 bl[80] br[80] wl[248] vdd gnd cell_6t
Xbit_r249_c80 bl[80] br[80] wl[249] vdd gnd cell_6t
Xbit_r250_c80 bl[80] br[80] wl[250] vdd gnd cell_6t
Xbit_r251_c80 bl[80] br[80] wl[251] vdd gnd cell_6t
Xbit_r252_c80 bl[80] br[80] wl[252] vdd gnd cell_6t
Xbit_r253_c80 bl[80] br[80] wl[253] vdd gnd cell_6t
Xbit_r254_c80 bl[80] br[80] wl[254] vdd gnd cell_6t
Xbit_r255_c80 bl[80] br[80] wl[255] vdd gnd cell_6t
Xbit_r0_c81 bl[81] br[81] wl[0] vdd gnd cell_6t
Xbit_r1_c81 bl[81] br[81] wl[1] vdd gnd cell_6t
Xbit_r2_c81 bl[81] br[81] wl[2] vdd gnd cell_6t
Xbit_r3_c81 bl[81] br[81] wl[3] vdd gnd cell_6t
Xbit_r4_c81 bl[81] br[81] wl[4] vdd gnd cell_6t
Xbit_r5_c81 bl[81] br[81] wl[5] vdd gnd cell_6t
Xbit_r6_c81 bl[81] br[81] wl[6] vdd gnd cell_6t
Xbit_r7_c81 bl[81] br[81] wl[7] vdd gnd cell_6t
Xbit_r8_c81 bl[81] br[81] wl[8] vdd gnd cell_6t
Xbit_r9_c81 bl[81] br[81] wl[9] vdd gnd cell_6t
Xbit_r10_c81 bl[81] br[81] wl[10] vdd gnd cell_6t
Xbit_r11_c81 bl[81] br[81] wl[11] vdd gnd cell_6t
Xbit_r12_c81 bl[81] br[81] wl[12] vdd gnd cell_6t
Xbit_r13_c81 bl[81] br[81] wl[13] vdd gnd cell_6t
Xbit_r14_c81 bl[81] br[81] wl[14] vdd gnd cell_6t
Xbit_r15_c81 bl[81] br[81] wl[15] vdd gnd cell_6t
Xbit_r16_c81 bl[81] br[81] wl[16] vdd gnd cell_6t
Xbit_r17_c81 bl[81] br[81] wl[17] vdd gnd cell_6t
Xbit_r18_c81 bl[81] br[81] wl[18] vdd gnd cell_6t
Xbit_r19_c81 bl[81] br[81] wl[19] vdd gnd cell_6t
Xbit_r20_c81 bl[81] br[81] wl[20] vdd gnd cell_6t
Xbit_r21_c81 bl[81] br[81] wl[21] vdd gnd cell_6t
Xbit_r22_c81 bl[81] br[81] wl[22] vdd gnd cell_6t
Xbit_r23_c81 bl[81] br[81] wl[23] vdd gnd cell_6t
Xbit_r24_c81 bl[81] br[81] wl[24] vdd gnd cell_6t
Xbit_r25_c81 bl[81] br[81] wl[25] vdd gnd cell_6t
Xbit_r26_c81 bl[81] br[81] wl[26] vdd gnd cell_6t
Xbit_r27_c81 bl[81] br[81] wl[27] vdd gnd cell_6t
Xbit_r28_c81 bl[81] br[81] wl[28] vdd gnd cell_6t
Xbit_r29_c81 bl[81] br[81] wl[29] vdd gnd cell_6t
Xbit_r30_c81 bl[81] br[81] wl[30] vdd gnd cell_6t
Xbit_r31_c81 bl[81] br[81] wl[31] vdd gnd cell_6t
Xbit_r32_c81 bl[81] br[81] wl[32] vdd gnd cell_6t
Xbit_r33_c81 bl[81] br[81] wl[33] vdd gnd cell_6t
Xbit_r34_c81 bl[81] br[81] wl[34] vdd gnd cell_6t
Xbit_r35_c81 bl[81] br[81] wl[35] vdd gnd cell_6t
Xbit_r36_c81 bl[81] br[81] wl[36] vdd gnd cell_6t
Xbit_r37_c81 bl[81] br[81] wl[37] vdd gnd cell_6t
Xbit_r38_c81 bl[81] br[81] wl[38] vdd gnd cell_6t
Xbit_r39_c81 bl[81] br[81] wl[39] vdd gnd cell_6t
Xbit_r40_c81 bl[81] br[81] wl[40] vdd gnd cell_6t
Xbit_r41_c81 bl[81] br[81] wl[41] vdd gnd cell_6t
Xbit_r42_c81 bl[81] br[81] wl[42] vdd gnd cell_6t
Xbit_r43_c81 bl[81] br[81] wl[43] vdd gnd cell_6t
Xbit_r44_c81 bl[81] br[81] wl[44] vdd gnd cell_6t
Xbit_r45_c81 bl[81] br[81] wl[45] vdd gnd cell_6t
Xbit_r46_c81 bl[81] br[81] wl[46] vdd gnd cell_6t
Xbit_r47_c81 bl[81] br[81] wl[47] vdd gnd cell_6t
Xbit_r48_c81 bl[81] br[81] wl[48] vdd gnd cell_6t
Xbit_r49_c81 bl[81] br[81] wl[49] vdd gnd cell_6t
Xbit_r50_c81 bl[81] br[81] wl[50] vdd gnd cell_6t
Xbit_r51_c81 bl[81] br[81] wl[51] vdd gnd cell_6t
Xbit_r52_c81 bl[81] br[81] wl[52] vdd gnd cell_6t
Xbit_r53_c81 bl[81] br[81] wl[53] vdd gnd cell_6t
Xbit_r54_c81 bl[81] br[81] wl[54] vdd gnd cell_6t
Xbit_r55_c81 bl[81] br[81] wl[55] vdd gnd cell_6t
Xbit_r56_c81 bl[81] br[81] wl[56] vdd gnd cell_6t
Xbit_r57_c81 bl[81] br[81] wl[57] vdd gnd cell_6t
Xbit_r58_c81 bl[81] br[81] wl[58] vdd gnd cell_6t
Xbit_r59_c81 bl[81] br[81] wl[59] vdd gnd cell_6t
Xbit_r60_c81 bl[81] br[81] wl[60] vdd gnd cell_6t
Xbit_r61_c81 bl[81] br[81] wl[61] vdd gnd cell_6t
Xbit_r62_c81 bl[81] br[81] wl[62] vdd gnd cell_6t
Xbit_r63_c81 bl[81] br[81] wl[63] vdd gnd cell_6t
Xbit_r64_c81 bl[81] br[81] wl[64] vdd gnd cell_6t
Xbit_r65_c81 bl[81] br[81] wl[65] vdd gnd cell_6t
Xbit_r66_c81 bl[81] br[81] wl[66] vdd gnd cell_6t
Xbit_r67_c81 bl[81] br[81] wl[67] vdd gnd cell_6t
Xbit_r68_c81 bl[81] br[81] wl[68] vdd gnd cell_6t
Xbit_r69_c81 bl[81] br[81] wl[69] vdd gnd cell_6t
Xbit_r70_c81 bl[81] br[81] wl[70] vdd gnd cell_6t
Xbit_r71_c81 bl[81] br[81] wl[71] vdd gnd cell_6t
Xbit_r72_c81 bl[81] br[81] wl[72] vdd gnd cell_6t
Xbit_r73_c81 bl[81] br[81] wl[73] vdd gnd cell_6t
Xbit_r74_c81 bl[81] br[81] wl[74] vdd gnd cell_6t
Xbit_r75_c81 bl[81] br[81] wl[75] vdd gnd cell_6t
Xbit_r76_c81 bl[81] br[81] wl[76] vdd gnd cell_6t
Xbit_r77_c81 bl[81] br[81] wl[77] vdd gnd cell_6t
Xbit_r78_c81 bl[81] br[81] wl[78] vdd gnd cell_6t
Xbit_r79_c81 bl[81] br[81] wl[79] vdd gnd cell_6t
Xbit_r80_c81 bl[81] br[81] wl[80] vdd gnd cell_6t
Xbit_r81_c81 bl[81] br[81] wl[81] vdd gnd cell_6t
Xbit_r82_c81 bl[81] br[81] wl[82] vdd gnd cell_6t
Xbit_r83_c81 bl[81] br[81] wl[83] vdd gnd cell_6t
Xbit_r84_c81 bl[81] br[81] wl[84] vdd gnd cell_6t
Xbit_r85_c81 bl[81] br[81] wl[85] vdd gnd cell_6t
Xbit_r86_c81 bl[81] br[81] wl[86] vdd gnd cell_6t
Xbit_r87_c81 bl[81] br[81] wl[87] vdd gnd cell_6t
Xbit_r88_c81 bl[81] br[81] wl[88] vdd gnd cell_6t
Xbit_r89_c81 bl[81] br[81] wl[89] vdd gnd cell_6t
Xbit_r90_c81 bl[81] br[81] wl[90] vdd gnd cell_6t
Xbit_r91_c81 bl[81] br[81] wl[91] vdd gnd cell_6t
Xbit_r92_c81 bl[81] br[81] wl[92] vdd gnd cell_6t
Xbit_r93_c81 bl[81] br[81] wl[93] vdd gnd cell_6t
Xbit_r94_c81 bl[81] br[81] wl[94] vdd gnd cell_6t
Xbit_r95_c81 bl[81] br[81] wl[95] vdd gnd cell_6t
Xbit_r96_c81 bl[81] br[81] wl[96] vdd gnd cell_6t
Xbit_r97_c81 bl[81] br[81] wl[97] vdd gnd cell_6t
Xbit_r98_c81 bl[81] br[81] wl[98] vdd gnd cell_6t
Xbit_r99_c81 bl[81] br[81] wl[99] vdd gnd cell_6t
Xbit_r100_c81 bl[81] br[81] wl[100] vdd gnd cell_6t
Xbit_r101_c81 bl[81] br[81] wl[101] vdd gnd cell_6t
Xbit_r102_c81 bl[81] br[81] wl[102] vdd gnd cell_6t
Xbit_r103_c81 bl[81] br[81] wl[103] vdd gnd cell_6t
Xbit_r104_c81 bl[81] br[81] wl[104] vdd gnd cell_6t
Xbit_r105_c81 bl[81] br[81] wl[105] vdd gnd cell_6t
Xbit_r106_c81 bl[81] br[81] wl[106] vdd gnd cell_6t
Xbit_r107_c81 bl[81] br[81] wl[107] vdd gnd cell_6t
Xbit_r108_c81 bl[81] br[81] wl[108] vdd gnd cell_6t
Xbit_r109_c81 bl[81] br[81] wl[109] vdd gnd cell_6t
Xbit_r110_c81 bl[81] br[81] wl[110] vdd gnd cell_6t
Xbit_r111_c81 bl[81] br[81] wl[111] vdd gnd cell_6t
Xbit_r112_c81 bl[81] br[81] wl[112] vdd gnd cell_6t
Xbit_r113_c81 bl[81] br[81] wl[113] vdd gnd cell_6t
Xbit_r114_c81 bl[81] br[81] wl[114] vdd gnd cell_6t
Xbit_r115_c81 bl[81] br[81] wl[115] vdd gnd cell_6t
Xbit_r116_c81 bl[81] br[81] wl[116] vdd gnd cell_6t
Xbit_r117_c81 bl[81] br[81] wl[117] vdd gnd cell_6t
Xbit_r118_c81 bl[81] br[81] wl[118] vdd gnd cell_6t
Xbit_r119_c81 bl[81] br[81] wl[119] vdd gnd cell_6t
Xbit_r120_c81 bl[81] br[81] wl[120] vdd gnd cell_6t
Xbit_r121_c81 bl[81] br[81] wl[121] vdd gnd cell_6t
Xbit_r122_c81 bl[81] br[81] wl[122] vdd gnd cell_6t
Xbit_r123_c81 bl[81] br[81] wl[123] vdd gnd cell_6t
Xbit_r124_c81 bl[81] br[81] wl[124] vdd gnd cell_6t
Xbit_r125_c81 bl[81] br[81] wl[125] vdd gnd cell_6t
Xbit_r126_c81 bl[81] br[81] wl[126] vdd gnd cell_6t
Xbit_r127_c81 bl[81] br[81] wl[127] vdd gnd cell_6t
Xbit_r128_c81 bl[81] br[81] wl[128] vdd gnd cell_6t
Xbit_r129_c81 bl[81] br[81] wl[129] vdd gnd cell_6t
Xbit_r130_c81 bl[81] br[81] wl[130] vdd gnd cell_6t
Xbit_r131_c81 bl[81] br[81] wl[131] vdd gnd cell_6t
Xbit_r132_c81 bl[81] br[81] wl[132] vdd gnd cell_6t
Xbit_r133_c81 bl[81] br[81] wl[133] vdd gnd cell_6t
Xbit_r134_c81 bl[81] br[81] wl[134] vdd gnd cell_6t
Xbit_r135_c81 bl[81] br[81] wl[135] vdd gnd cell_6t
Xbit_r136_c81 bl[81] br[81] wl[136] vdd gnd cell_6t
Xbit_r137_c81 bl[81] br[81] wl[137] vdd gnd cell_6t
Xbit_r138_c81 bl[81] br[81] wl[138] vdd gnd cell_6t
Xbit_r139_c81 bl[81] br[81] wl[139] vdd gnd cell_6t
Xbit_r140_c81 bl[81] br[81] wl[140] vdd gnd cell_6t
Xbit_r141_c81 bl[81] br[81] wl[141] vdd gnd cell_6t
Xbit_r142_c81 bl[81] br[81] wl[142] vdd gnd cell_6t
Xbit_r143_c81 bl[81] br[81] wl[143] vdd gnd cell_6t
Xbit_r144_c81 bl[81] br[81] wl[144] vdd gnd cell_6t
Xbit_r145_c81 bl[81] br[81] wl[145] vdd gnd cell_6t
Xbit_r146_c81 bl[81] br[81] wl[146] vdd gnd cell_6t
Xbit_r147_c81 bl[81] br[81] wl[147] vdd gnd cell_6t
Xbit_r148_c81 bl[81] br[81] wl[148] vdd gnd cell_6t
Xbit_r149_c81 bl[81] br[81] wl[149] vdd gnd cell_6t
Xbit_r150_c81 bl[81] br[81] wl[150] vdd gnd cell_6t
Xbit_r151_c81 bl[81] br[81] wl[151] vdd gnd cell_6t
Xbit_r152_c81 bl[81] br[81] wl[152] vdd gnd cell_6t
Xbit_r153_c81 bl[81] br[81] wl[153] vdd gnd cell_6t
Xbit_r154_c81 bl[81] br[81] wl[154] vdd gnd cell_6t
Xbit_r155_c81 bl[81] br[81] wl[155] vdd gnd cell_6t
Xbit_r156_c81 bl[81] br[81] wl[156] vdd gnd cell_6t
Xbit_r157_c81 bl[81] br[81] wl[157] vdd gnd cell_6t
Xbit_r158_c81 bl[81] br[81] wl[158] vdd gnd cell_6t
Xbit_r159_c81 bl[81] br[81] wl[159] vdd gnd cell_6t
Xbit_r160_c81 bl[81] br[81] wl[160] vdd gnd cell_6t
Xbit_r161_c81 bl[81] br[81] wl[161] vdd gnd cell_6t
Xbit_r162_c81 bl[81] br[81] wl[162] vdd gnd cell_6t
Xbit_r163_c81 bl[81] br[81] wl[163] vdd gnd cell_6t
Xbit_r164_c81 bl[81] br[81] wl[164] vdd gnd cell_6t
Xbit_r165_c81 bl[81] br[81] wl[165] vdd gnd cell_6t
Xbit_r166_c81 bl[81] br[81] wl[166] vdd gnd cell_6t
Xbit_r167_c81 bl[81] br[81] wl[167] vdd gnd cell_6t
Xbit_r168_c81 bl[81] br[81] wl[168] vdd gnd cell_6t
Xbit_r169_c81 bl[81] br[81] wl[169] vdd gnd cell_6t
Xbit_r170_c81 bl[81] br[81] wl[170] vdd gnd cell_6t
Xbit_r171_c81 bl[81] br[81] wl[171] vdd gnd cell_6t
Xbit_r172_c81 bl[81] br[81] wl[172] vdd gnd cell_6t
Xbit_r173_c81 bl[81] br[81] wl[173] vdd gnd cell_6t
Xbit_r174_c81 bl[81] br[81] wl[174] vdd gnd cell_6t
Xbit_r175_c81 bl[81] br[81] wl[175] vdd gnd cell_6t
Xbit_r176_c81 bl[81] br[81] wl[176] vdd gnd cell_6t
Xbit_r177_c81 bl[81] br[81] wl[177] vdd gnd cell_6t
Xbit_r178_c81 bl[81] br[81] wl[178] vdd gnd cell_6t
Xbit_r179_c81 bl[81] br[81] wl[179] vdd gnd cell_6t
Xbit_r180_c81 bl[81] br[81] wl[180] vdd gnd cell_6t
Xbit_r181_c81 bl[81] br[81] wl[181] vdd gnd cell_6t
Xbit_r182_c81 bl[81] br[81] wl[182] vdd gnd cell_6t
Xbit_r183_c81 bl[81] br[81] wl[183] vdd gnd cell_6t
Xbit_r184_c81 bl[81] br[81] wl[184] vdd gnd cell_6t
Xbit_r185_c81 bl[81] br[81] wl[185] vdd gnd cell_6t
Xbit_r186_c81 bl[81] br[81] wl[186] vdd gnd cell_6t
Xbit_r187_c81 bl[81] br[81] wl[187] vdd gnd cell_6t
Xbit_r188_c81 bl[81] br[81] wl[188] vdd gnd cell_6t
Xbit_r189_c81 bl[81] br[81] wl[189] vdd gnd cell_6t
Xbit_r190_c81 bl[81] br[81] wl[190] vdd gnd cell_6t
Xbit_r191_c81 bl[81] br[81] wl[191] vdd gnd cell_6t
Xbit_r192_c81 bl[81] br[81] wl[192] vdd gnd cell_6t
Xbit_r193_c81 bl[81] br[81] wl[193] vdd gnd cell_6t
Xbit_r194_c81 bl[81] br[81] wl[194] vdd gnd cell_6t
Xbit_r195_c81 bl[81] br[81] wl[195] vdd gnd cell_6t
Xbit_r196_c81 bl[81] br[81] wl[196] vdd gnd cell_6t
Xbit_r197_c81 bl[81] br[81] wl[197] vdd gnd cell_6t
Xbit_r198_c81 bl[81] br[81] wl[198] vdd gnd cell_6t
Xbit_r199_c81 bl[81] br[81] wl[199] vdd gnd cell_6t
Xbit_r200_c81 bl[81] br[81] wl[200] vdd gnd cell_6t
Xbit_r201_c81 bl[81] br[81] wl[201] vdd gnd cell_6t
Xbit_r202_c81 bl[81] br[81] wl[202] vdd gnd cell_6t
Xbit_r203_c81 bl[81] br[81] wl[203] vdd gnd cell_6t
Xbit_r204_c81 bl[81] br[81] wl[204] vdd gnd cell_6t
Xbit_r205_c81 bl[81] br[81] wl[205] vdd gnd cell_6t
Xbit_r206_c81 bl[81] br[81] wl[206] vdd gnd cell_6t
Xbit_r207_c81 bl[81] br[81] wl[207] vdd gnd cell_6t
Xbit_r208_c81 bl[81] br[81] wl[208] vdd gnd cell_6t
Xbit_r209_c81 bl[81] br[81] wl[209] vdd gnd cell_6t
Xbit_r210_c81 bl[81] br[81] wl[210] vdd gnd cell_6t
Xbit_r211_c81 bl[81] br[81] wl[211] vdd gnd cell_6t
Xbit_r212_c81 bl[81] br[81] wl[212] vdd gnd cell_6t
Xbit_r213_c81 bl[81] br[81] wl[213] vdd gnd cell_6t
Xbit_r214_c81 bl[81] br[81] wl[214] vdd gnd cell_6t
Xbit_r215_c81 bl[81] br[81] wl[215] vdd gnd cell_6t
Xbit_r216_c81 bl[81] br[81] wl[216] vdd gnd cell_6t
Xbit_r217_c81 bl[81] br[81] wl[217] vdd gnd cell_6t
Xbit_r218_c81 bl[81] br[81] wl[218] vdd gnd cell_6t
Xbit_r219_c81 bl[81] br[81] wl[219] vdd gnd cell_6t
Xbit_r220_c81 bl[81] br[81] wl[220] vdd gnd cell_6t
Xbit_r221_c81 bl[81] br[81] wl[221] vdd gnd cell_6t
Xbit_r222_c81 bl[81] br[81] wl[222] vdd gnd cell_6t
Xbit_r223_c81 bl[81] br[81] wl[223] vdd gnd cell_6t
Xbit_r224_c81 bl[81] br[81] wl[224] vdd gnd cell_6t
Xbit_r225_c81 bl[81] br[81] wl[225] vdd gnd cell_6t
Xbit_r226_c81 bl[81] br[81] wl[226] vdd gnd cell_6t
Xbit_r227_c81 bl[81] br[81] wl[227] vdd gnd cell_6t
Xbit_r228_c81 bl[81] br[81] wl[228] vdd gnd cell_6t
Xbit_r229_c81 bl[81] br[81] wl[229] vdd gnd cell_6t
Xbit_r230_c81 bl[81] br[81] wl[230] vdd gnd cell_6t
Xbit_r231_c81 bl[81] br[81] wl[231] vdd gnd cell_6t
Xbit_r232_c81 bl[81] br[81] wl[232] vdd gnd cell_6t
Xbit_r233_c81 bl[81] br[81] wl[233] vdd gnd cell_6t
Xbit_r234_c81 bl[81] br[81] wl[234] vdd gnd cell_6t
Xbit_r235_c81 bl[81] br[81] wl[235] vdd gnd cell_6t
Xbit_r236_c81 bl[81] br[81] wl[236] vdd gnd cell_6t
Xbit_r237_c81 bl[81] br[81] wl[237] vdd gnd cell_6t
Xbit_r238_c81 bl[81] br[81] wl[238] vdd gnd cell_6t
Xbit_r239_c81 bl[81] br[81] wl[239] vdd gnd cell_6t
Xbit_r240_c81 bl[81] br[81] wl[240] vdd gnd cell_6t
Xbit_r241_c81 bl[81] br[81] wl[241] vdd gnd cell_6t
Xbit_r242_c81 bl[81] br[81] wl[242] vdd gnd cell_6t
Xbit_r243_c81 bl[81] br[81] wl[243] vdd gnd cell_6t
Xbit_r244_c81 bl[81] br[81] wl[244] vdd gnd cell_6t
Xbit_r245_c81 bl[81] br[81] wl[245] vdd gnd cell_6t
Xbit_r246_c81 bl[81] br[81] wl[246] vdd gnd cell_6t
Xbit_r247_c81 bl[81] br[81] wl[247] vdd gnd cell_6t
Xbit_r248_c81 bl[81] br[81] wl[248] vdd gnd cell_6t
Xbit_r249_c81 bl[81] br[81] wl[249] vdd gnd cell_6t
Xbit_r250_c81 bl[81] br[81] wl[250] vdd gnd cell_6t
Xbit_r251_c81 bl[81] br[81] wl[251] vdd gnd cell_6t
Xbit_r252_c81 bl[81] br[81] wl[252] vdd gnd cell_6t
Xbit_r253_c81 bl[81] br[81] wl[253] vdd gnd cell_6t
Xbit_r254_c81 bl[81] br[81] wl[254] vdd gnd cell_6t
Xbit_r255_c81 bl[81] br[81] wl[255] vdd gnd cell_6t
Xbit_r0_c82 bl[82] br[82] wl[0] vdd gnd cell_6t
Xbit_r1_c82 bl[82] br[82] wl[1] vdd gnd cell_6t
Xbit_r2_c82 bl[82] br[82] wl[2] vdd gnd cell_6t
Xbit_r3_c82 bl[82] br[82] wl[3] vdd gnd cell_6t
Xbit_r4_c82 bl[82] br[82] wl[4] vdd gnd cell_6t
Xbit_r5_c82 bl[82] br[82] wl[5] vdd gnd cell_6t
Xbit_r6_c82 bl[82] br[82] wl[6] vdd gnd cell_6t
Xbit_r7_c82 bl[82] br[82] wl[7] vdd gnd cell_6t
Xbit_r8_c82 bl[82] br[82] wl[8] vdd gnd cell_6t
Xbit_r9_c82 bl[82] br[82] wl[9] vdd gnd cell_6t
Xbit_r10_c82 bl[82] br[82] wl[10] vdd gnd cell_6t
Xbit_r11_c82 bl[82] br[82] wl[11] vdd gnd cell_6t
Xbit_r12_c82 bl[82] br[82] wl[12] vdd gnd cell_6t
Xbit_r13_c82 bl[82] br[82] wl[13] vdd gnd cell_6t
Xbit_r14_c82 bl[82] br[82] wl[14] vdd gnd cell_6t
Xbit_r15_c82 bl[82] br[82] wl[15] vdd gnd cell_6t
Xbit_r16_c82 bl[82] br[82] wl[16] vdd gnd cell_6t
Xbit_r17_c82 bl[82] br[82] wl[17] vdd gnd cell_6t
Xbit_r18_c82 bl[82] br[82] wl[18] vdd gnd cell_6t
Xbit_r19_c82 bl[82] br[82] wl[19] vdd gnd cell_6t
Xbit_r20_c82 bl[82] br[82] wl[20] vdd gnd cell_6t
Xbit_r21_c82 bl[82] br[82] wl[21] vdd gnd cell_6t
Xbit_r22_c82 bl[82] br[82] wl[22] vdd gnd cell_6t
Xbit_r23_c82 bl[82] br[82] wl[23] vdd gnd cell_6t
Xbit_r24_c82 bl[82] br[82] wl[24] vdd gnd cell_6t
Xbit_r25_c82 bl[82] br[82] wl[25] vdd gnd cell_6t
Xbit_r26_c82 bl[82] br[82] wl[26] vdd gnd cell_6t
Xbit_r27_c82 bl[82] br[82] wl[27] vdd gnd cell_6t
Xbit_r28_c82 bl[82] br[82] wl[28] vdd gnd cell_6t
Xbit_r29_c82 bl[82] br[82] wl[29] vdd gnd cell_6t
Xbit_r30_c82 bl[82] br[82] wl[30] vdd gnd cell_6t
Xbit_r31_c82 bl[82] br[82] wl[31] vdd gnd cell_6t
Xbit_r32_c82 bl[82] br[82] wl[32] vdd gnd cell_6t
Xbit_r33_c82 bl[82] br[82] wl[33] vdd gnd cell_6t
Xbit_r34_c82 bl[82] br[82] wl[34] vdd gnd cell_6t
Xbit_r35_c82 bl[82] br[82] wl[35] vdd gnd cell_6t
Xbit_r36_c82 bl[82] br[82] wl[36] vdd gnd cell_6t
Xbit_r37_c82 bl[82] br[82] wl[37] vdd gnd cell_6t
Xbit_r38_c82 bl[82] br[82] wl[38] vdd gnd cell_6t
Xbit_r39_c82 bl[82] br[82] wl[39] vdd gnd cell_6t
Xbit_r40_c82 bl[82] br[82] wl[40] vdd gnd cell_6t
Xbit_r41_c82 bl[82] br[82] wl[41] vdd gnd cell_6t
Xbit_r42_c82 bl[82] br[82] wl[42] vdd gnd cell_6t
Xbit_r43_c82 bl[82] br[82] wl[43] vdd gnd cell_6t
Xbit_r44_c82 bl[82] br[82] wl[44] vdd gnd cell_6t
Xbit_r45_c82 bl[82] br[82] wl[45] vdd gnd cell_6t
Xbit_r46_c82 bl[82] br[82] wl[46] vdd gnd cell_6t
Xbit_r47_c82 bl[82] br[82] wl[47] vdd gnd cell_6t
Xbit_r48_c82 bl[82] br[82] wl[48] vdd gnd cell_6t
Xbit_r49_c82 bl[82] br[82] wl[49] vdd gnd cell_6t
Xbit_r50_c82 bl[82] br[82] wl[50] vdd gnd cell_6t
Xbit_r51_c82 bl[82] br[82] wl[51] vdd gnd cell_6t
Xbit_r52_c82 bl[82] br[82] wl[52] vdd gnd cell_6t
Xbit_r53_c82 bl[82] br[82] wl[53] vdd gnd cell_6t
Xbit_r54_c82 bl[82] br[82] wl[54] vdd gnd cell_6t
Xbit_r55_c82 bl[82] br[82] wl[55] vdd gnd cell_6t
Xbit_r56_c82 bl[82] br[82] wl[56] vdd gnd cell_6t
Xbit_r57_c82 bl[82] br[82] wl[57] vdd gnd cell_6t
Xbit_r58_c82 bl[82] br[82] wl[58] vdd gnd cell_6t
Xbit_r59_c82 bl[82] br[82] wl[59] vdd gnd cell_6t
Xbit_r60_c82 bl[82] br[82] wl[60] vdd gnd cell_6t
Xbit_r61_c82 bl[82] br[82] wl[61] vdd gnd cell_6t
Xbit_r62_c82 bl[82] br[82] wl[62] vdd gnd cell_6t
Xbit_r63_c82 bl[82] br[82] wl[63] vdd gnd cell_6t
Xbit_r64_c82 bl[82] br[82] wl[64] vdd gnd cell_6t
Xbit_r65_c82 bl[82] br[82] wl[65] vdd gnd cell_6t
Xbit_r66_c82 bl[82] br[82] wl[66] vdd gnd cell_6t
Xbit_r67_c82 bl[82] br[82] wl[67] vdd gnd cell_6t
Xbit_r68_c82 bl[82] br[82] wl[68] vdd gnd cell_6t
Xbit_r69_c82 bl[82] br[82] wl[69] vdd gnd cell_6t
Xbit_r70_c82 bl[82] br[82] wl[70] vdd gnd cell_6t
Xbit_r71_c82 bl[82] br[82] wl[71] vdd gnd cell_6t
Xbit_r72_c82 bl[82] br[82] wl[72] vdd gnd cell_6t
Xbit_r73_c82 bl[82] br[82] wl[73] vdd gnd cell_6t
Xbit_r74_c82 bl[82] br[82] wl[74] vdd gnd cell_6t
Xbit_r75_c82 bl[82] br[82] wl[75] vdd gnd cell_6t
Xbit_r76_c82 bl[82] br[82] wl[76] vdd gnd cell_6t
Xbit_r77_c82 bl[82] br[82] wl[77] vdd gnd cell_6t
Xbit_r78_c82 bl[82] br[82] wl[78] vdd gnd cell_6t
Xbit_r79_c82 bl[82] br[82] wl[79] vdd gnd cell_6t
Xbit_r80_c82 bl[82] br[82] wl[80] vdd gnd cell_6t
Xbit_r81_c82 bl[82] br[82] wl[81] vdd gnd cell_6t
Xbit_r82_c82 bl[82] br[82] wl[82] vdd gnd cell_6t
Xbit_r83_c82 bl[82] br[82] wl[83] vdd gnd cell_6t
Xbit_r84_c82 bl[82] br[82] wl[84] vdd gnd cell_6t
Xbit_r85_c82 bl[82] br[82] wl[85] vdd gnd cell_6t
Xbit_r86_c82 bl[82] br[82] wl[86] vdd gnd cell_6t
Xbit_r87_c82 bl[82] br[82] wl[87] vdd gnd cell_6t
Xbit_r88_c82 bl[82] br[82] wl[88] vdd gnd cell_6t
Xbit_r89_c82 bl[82] br[82] wl[89] vdd gnd cell_6t
Xbit_r90_c82 bl[82] br[82] wl[90] vdd gnd cell_6t
Xbit_r91_c82 bl[82] br[82] wl[91] vdd gnd cell_6t
Xbit_r92_c82 bl[82] br[82] wl[92] vdd gnd cell_6t
Xbit_r93_c82 bl[82] br[82] wl[93] vdd gnd cell_6t
Xbit_r94_c82 bl[82] br[82] wl[94] vdd gnd cell_6t
Xbit_r95_c82 bl[82] br[82] wl[95] vdd gnd cell_6t
Xbit_r96_c82 bl[82] br[82] wl[96] vdd gnd cell_6t
Xbit_r97_c82 bl[82] br[82] wl[97] vdd gnd cell_6t
Xbit_r98_c82 bl[82] br[82] wl[98] vdd gnd cell_6t
Xbit_r99_c82 bl[82] br[82] wl[99] vdd gnd cell_6t
Xbit_r100_c82 bl[82] br[82] wl[100] vdd gnd cell_6t
Xbit_r101_c82 bl[82] br[82] wl[101] vdd gnd cell_6t
Xbit_r102_c82 bl[82] br[82] wl[102] vdd gnd cell_6t
Xbit_r103_c82 bl[82] br[82] wl[103] vdd gnd cell_6t
Xbit_r104_c82 bl[82] br[82] wl[104] vdd gnd cell_6t
Xbit_r105_c82 bl[82] br[82] wl[105] vdd gnd cell_6t
Xbit_r106_c82 bl[82] br[82] wl[106] vdd gnd cell_6t
Xbit_r107_c82 bl[82] br[82] wl[107] vdd gnd cell_6t
Xbit_r108_c82 bl[82] br[82] wl[108] vdd gnd cell_6t
Xbit_r109_c82 bl[82] br[82] wl[109] vdd gnd cell_6t
Xbit_r110_c82 bl[82] br[82] wl[110] vdd gnd cell_6t
Xbit_r111_c82 bl[82] br[82] wl[111] vdd gnd cell_6t
Xbit_r112_c82 bl[82] br[82] wl[112] vdd gnd cell_6t
Xbit_r113_c82 bl[82] br[82] wl[113] vdd gnd cell_6t
Xbit_r114_c82 bl[82] br[82] wl[114] vdd gnd cell_6t
Xbit_r115_c82 bl[82] br[82] wl[115] vdd gnd cell_6t
Xbit_r116_c82 bl[82] br[82] wl[116] vdd gnd cell_6t
Xbit_r117_c82 bl[82] br[82] wl[117] vdd gnd cell_6t
Xbit_r118_c82 bl[82] br[82] wl[118] vdd gnd cell_6t
Xbit_r119_c82 bl[82] br[82] wl[119] vdd gnd cell_6t
Xbit_r120_c82 bl[82] br[82] wl[120] vdd gnd cell_6t
Xbit_r121_c82 bl[82] br[82] wl[121] vdd gnd cell_6t
Xbit_r122_c82 bl[82] br[82] wl[122] vdd gnd cell_6t
Xbit_r123_c82 bl[82] br[82] wl[123] vdd gnd cell_6t
Xbit_r124_c82 bl[82] br[82] wl[124] vdd gnd cell_6t
Xbit_r125_c82 bl[82] br[82] wl[125] vdd gnd cell_6t
Xbit_r126_c82 bl[82] br[82] wl[126] vdd gnd cell_6t
Xbit_r127_c82 bl[82] br[82] wl[127] vdd gnd cell_6t
Xbit_r128_c82 bl[82] br[82] wl[128] vdd gnd cell_6t
Xbit_r129_c82 bl[82] br[82] wl[129] vdd gnd cell_6t
Xbit_r130_c82 bl[82] br[82] wl[130] vdd gnd cell_6t
Xbit_r131_c82 bl[82] br[82] wl[131] vdd gnd cell_6t
Xbit_r132_c82 bl[82] br[82] wl[132] vdd gnd cell_6t
Xbit_r133_c82 bl[82] br[82] wl[133] vdd gnd cell_6t
Xbit_r134_c82 bl[82] br[82] wl[134] vdd gnd cell_6t
Xbit_r135_c82 bl[82] br[82] wl[135] vdd gnd cell_6t
Xbit_r136_c82 bl[82] br[82] wl[136] vdd gnd cell_6t
Xbit_r137_c82 bl[82] br[82] wl[137] vdd gnd cell_6t
Xbit_r138_c82 bl[82] br[82] wl[138] vdd gnd cell_6t
Xbit_r139_c82 bl[82] br[82] wl[139] vdd gnd cell_6t
Xbit_r140_c82 bl[82] br[82] wl[140] vdd gnd cell_6t
Xbit_r141_c82 bl[82] br[82] wl[141] vdd gnd cell_6t
Xbit_r142_c82 bl[82] br[82] wl[142] vdd gnd cell_6t
Xbit_r143_c82 bl[82] br[82] wl[143] vdd gnd cell_6t
Xbit_r144_c82 bl[82] br[82] wl[144] vdd gnd cell_6t
Xbit_r145_c82 bl[82] br[82] wl[145] vdd gnd cell_6t
Xbit_r146_c82 bl[82] br[82] wl[146] vdd gnd cell_6t
Xbit_r147_c82 bl[82] br[82] wl[147] vdd gnd cell_6t
Xbit_r148_c82 bl[82] br[82] wl[148] vdd gnd cell_6t
Xbit_r149_c82 bl[82] br[82] wl[149] vdd gnd cell_6t
Xbit_r150_c82 bl[82] br[82] wl[150] vdd gnd cell_6t
Xbit_r151_c82 bl[82] br[82] wl[151] vdd gnd cell_6t
Xbit_r152_c82 bl[82] br[82] wl[152] vdd gnd cell_6t
Xbit_r153_c82 bl[82] br[82] wl[153] vdd gnd cell_6t
Xbit_r154_c82 bl[82] br[82] wl[154] vdd gnd cell_6t
Xbit_r155_c82 bl[82] br[82] wl[155] vdd gnd cell_6t
Xbit_r156_c82 bl[82] br[82] wl[156] vdd gnd cell_6t
Xbit_r157_c82 bl[82] br[82] wl[157] vdd gnd cell_6t
Xbit_r158_c82 bl[82] br[82] wl[158] vdd gnd cell_6t
Xbit_r159_c82 bl[82] br[82] wl[159] vdd gnd cell_6t
Xbit_r160_c82 bl[82] br[82] wl[160] vdd gnd cell_6t
Xbit_r161_c82 bl[82] br[82] wl[161] vdd gnd cell_6t
Xbit_r162_c82 bl[82] br[82] wl[162] vdd gnd cell_6t
Xbit_r163_c82 bl[82] br[82] wl[163] vdd gnd cell_6t
Xbit_r164_c82 bl[82] br[82] wl[164] vdd gnd cell_6t
Xbit_r165_c82 bl[82] br[82] wl[165] vdd gnd cell_6t
Xbit_r166_c82 bl[82] br[82] wl[166] vdd gnd cell_6t
Xbit_r167_c82 bl[82] br[82] wl[167] vdd gnd cell_6t
Xbit_r168_c82 bl[82] br[82] wl[168] vdd gnd cell_6t
Xbit_r169_c82 bl[82] br[82] wl[169] vdd gnd cell_6t
Xbit_r170_c82 bl[82] br[82] wl[170] vdd gnd cell_6t
Xbit_r171_c82 bl[82] br[82] wl[171] vdd gnd cell_6t
Xbit_r172_c82 bl[82] br[82] wl[172] vdd gnd cell_6t
Xbit_r173_c82 bl[82] br[82] wl[173] vdd gnd cell_6t
Xbit_r174_c82 bl[82] br[82] wl[174] vdd gnd cell_6t
Xbit_r175_c82 bl[82] br[82] wl[175] vdd gnd cell_6t
Xbit_r176_c82 bl[82] br[82] wl[176] vdd gnd cell_6t
Xbit_r177_c82 bl[82] br[82] wl[177] vdd gnd cell_6t
Xbit_r178_c82 bl[82] br[82] wl[178] vdd gnd cell_6t
Xbit_r179_c82 bl[82] br[82] wl[179] vdd gnd cell_6t
Xbit_r180_c82 bl[82] br[82] wl[180] vdd gnd cell_6t
Xbit_r181_c82 bl[82] br[82] wl[181] vdd gnd cell_6t
Xbit_r182_c82 bl[82] br[82] wl[182] vdd gnd cell_6t
Xbit_r183_c82 bl[82] br[82] wl[183] vdd gnd cell_6t
Xbit_r184_c82 bl[82] br[82] wl[184] vdd gnd cell_6t
Xbit_r185_c82 bl[82] br[82] wl[185] vdd gnd cell_6t
Xbit_r186_c82 bl[82] br[82] wl[186] vdd gnd cell_6t
Xbit_r187_c82 bl[82] br[82] wl[187] vdd gnd cell_6t
Xbit_r188_c82 bl[82] br[82] wl[188] vdd gnd cell_6t
Xbit_r189_c82 bl[82] br[82] wl[189] vdd gnd cell_6t
Xbit_r190_c82 bl[82] br[82] wl[190] vdd gnd cell_6t
Xbit_r191_c82 bl[82] br[82] wl[191] vdd gnd cell_6t
Xbit_r192_c82 bl[82] br[82] wl[192] vdd gnd cell_6t
Xbit_r193_c82 bl[82] br[82] wl[193] vdd gnd cell_6t
Xbit_r194_c82 bl[82] br[82] wl[194] vdd gnd cell_6t
Xbit_r195_c82 bl[82] br[82] wl[195] vdd gnd cell_6t
Xbit_r196_c82 bl[82] br[82] wl[196] vdd gnd cell_6t
Xbit_r197_c82 bl[82] br[82] wl[197] vdd gnd cell_6t
Xbit_r198_c82 bl[82] br[82] wl[198] vdd gnd cell_6t
Xbit_r199_c82 bl[82] br[82] wl[199] vdd gnd cell_6t
Xbit_r200_c82 bl[82] br[82] wl[200] vdd gnd cell_6t
Xbit_r201_c82 bl[82] br[82] wl[201] vdd gnd cell_6t
Xbit_r202_c82 bl[82] br[82] wl[202] vdd gnd cell_6t
Xbit_r203_c82 bl[82] br[82] wl[203] vdd gnd cell_6t
Xbit_r204_c82 bl[82] br[82] wl[204] vdd gnd cell_6t
Xbit_r205_c82 bl[82] br[82] wl[205] vdd gnd cell_6t
Xbit_r206_c82 bl[82] br[82] wl[206] vdd gnd cell_6t
Xbit_r207_c82 bl[82] br[82] wl[207] vdd gnd cell_6t
Xbit_r208_c82 bl[82] br[82] wl[208] vdd gnd cell_6t
Xbit_r209_c82 bl[82] br[82] wl[209] vdd gnd cell_6t
Xbit_r210_c82 bl[82] br[82] wl[210] vdd gnd cell_6t
Xbit_r211_c82 bl[82] br[82] wl[211] vdd gnd cell_6t
Xbit_r212_c82 bl[82] br[82] wl[212] vdd gnd cell_6t
Xbit_r213_c82 bl[82] br[82] wl[213] vdd gnd cell_6t
Xbit_r214_c82 bl[82] br[82] wl[214] vdd gnd cell_6t
Xbit_r215_c82 bl[82] br[82] wl[215] vdd gnd cell_6t
Xbit_r216_c82 bl[82] br[82] wl[216] vdd gnd cell_6t
Xbit_r217_c82 bl[82] br[82] wl[217] vdd gnd cell_6t
Xbit_r218_c82 bl[82] br[82] wl[218] vdd gnd cell_6t
Xbit_r219_c82 bl[82] br[82] wl[219] vdd gnd cell_6t
Xbit_r220_c82 bl[82] br[82] wl[220] vdd gnd cell_6t
Xbit_r221_c82 bl[82] br[82] wl[221] vdd gnd cell_6t
Xbit_r222_c82 bl[82] br[82] wl[222] vdd gnd cell_6t
Xbit_r223_c82 bl[82] br[82] wl[223] vdd gnd cell_6t
Xbit_r224_c82 bl[82] br[82] wl[224] vdd gnd cell_6t
Xbit_r225_c82 bl[82] br[82] wl[225] vdd gnd cell_6t
Xbit_r226_c82 bl[82] br[82] wl[226] vdd gnd cell_6t
Xbit_r227_c82 bl[82] br[82] wl[227] vdd gnd cell_6t
Xbit_r228_c82 bl[82] br[82] wl[228] vdd gnd cell_6t
Xbit_r229_c82 bl[82] br[82] wl[229] vdd gnd cell_6t
Xbit_r230_c82 bl[82] br[82] wl[230] vdd gnd cell_6t
Xbit_r231_c82 bl[82] br[82] wl[231] vdd gnd cell_6t
Xbit_r232_c82 bl[82] br[82] wl[232] vdd gnd cell_6t
Xbit_r233_c82 bl[82] br[82] wl[233] vdd gnd cell_6t
Xbit_r234_c82 bl[82] br[82] wl[234] vdd gnd cell_6t
Xbit_r235_c82 bl[82] br[82] wl[235] vdd gnd cell_6t
Xbit_r236_c82 bl[82] br[82] wl[236] vdd gnd cell_6t
Xbit_r237_c82 bl[82] br[82] wl[237] vdd gnd cell_6t
Xbit_r238_c82 bl[82] br[82] wl[238] vdd gnd cell_6t
Xbit_r239_c82 bl[82] br[82] wl[239] vdd gnd cell_6t
Xbit_r240_c82 bl[82] br[82] wl[240] vdd gnd cell_6t
Xbit_r241_c82 bl[82] br[82] wl[241] vdd gnd cell_6t
Xbit_r242_c82 bl[82] br[82] wl[242] vdd gnd cell_6t
Xbit_r243_c82 bl[82] br[82] wl[243] vdd gnd cell_6t
Xbit_r244_c82 bl[82] br[82] wl[244] vdd gnd cell_6t
Xbit_r245_c82 bl[82] br[82] wl[245] vdd gnd cell_6t
Xbit_r246_c82 bl[82] br[82] wl[246] vdd gnd cell_6t
Xbit_r247_c82 bl[82] br[82] wl[247] vdd gnd cell_6t
Xbit_r248_c82 bl[82] br[82] wl[248] vdd gnd cell_6t
Xbit_r249_c82 bl[82] br[82] wl[249] vdd gnd cell_6t
Xbit_r250_c82 bl[82] br[82] wl[250] vdd gnd cell_6t
Xbit_r251_c82 bl[82] br[82] wl[251] vdd gnd cell_6t
Xbit_r252_c82 bl[82] br[82] wl[252] vdd gnd cell_6t
Xbit_r253_c82 bl[82] br[82] wl[253] vdd gnd cell_6t
Xbit_r254_c82 bl[82] br[82] wl[254] vdd gnd cell_6t
Xbit_r255_c82 bl[82] br[82] wl[255] vdd gnd cell_6t
Xbit_r0_c83 bl[83] br[83] wl[0] vdd gnd cell_6t
Xbit_r1_c83 bl[83] br[83] wl[1] vdd gnd cell_6t
Xbit_r2_c83 bl[83] br[83] wl[2] vdd gnd cell_6t
Xbit_r3_c83 bl[83] br[83] wl[3] vdd gnd cell_6t
Xbit_r4_c83 bl[83] br[83] wl[4] vdd gnd cell_6t
Xbit_r5_c83 bl[83] br[83] wl[5] vdd gnd cell_6t
Xbit_r6_c83 bl[83] br[83] wl[6] vdd gnd cell_6t
Xbit_r7_c83 bl[83] br[83] wl[7] vdd gnd cell_6t
Xbit_r8_c83 bl[83] br[83] wl[8] vdd gnd cell_6t
Xbit_r9_c83 bl[83] br[83] wl[9] vdd gnd cell_6t
Xbit_r10_c83 bl[83] br[83] wl[10] vdd gnd cell_6t
Xbit_r11_c83 bl[83] br[83] wl[11] vdd gnd cell_6t
Xbit_r12_c83 bl[83] br[83] wl[12] vdd gnd cell_6t
Xbit_r13_c83 bl[83] br[83] wl[13] vdd gnd cell_6t
Xbit_r14_c83 bl[83] br[83] wl[14] vdd gnd cell_6t
Xbit_r15_c83 bl[83] br[83] wl[15] vdd gnd cell_6t
Xbit_r16_c83 bl[83] br[83] wl[16] vdd gnd cell_6t
Xbit_r17_c83 bl[83] br[83] wl[17] vdd gnd cell_6t
Xbit_r18_c83 bl[83] br[83] wl[18] vdd gnd cell_6t
Xbit_r19_c83 bl[83] br[83] wl[19] vdd gnd cell_6t
Xbit_r20_c83 bl[83] br[83] wl[20] vdd gnd cell_6t
Xbit_r21_c83 bl[83] br[83] wl[21] vdd gnd cell_6t
Xbit_r22_c83 bl[83] br[83] wl[22] vdd gnd cell_6t
Xbit_r23_c83 bl[83] br[83] wl[23] vdd gnd cell_6t
Xbit_r24_c83 bl[83] br[83] wl[24] vdd gnd cell_6t
Xbit_r25_c83 bl[83] br[83] wl[25] vdd gnd cell_6t
Xbit_r26_c83 bl[83] br[83] wl[26] vdd gnd cell_6t
Xbit_r27_c83 bl[83] br[83] wl[27] vdd gnd cell_6t
Xbit_r28_c83 bl[83] br[83] wl[28] vdd gnd cell_6t
Xbit_r29_c83 bl[83] br[83] wl[29] vdd gnd cell_6t
Xbit_r30_c83 bl[83] br[83] wl[30] vdd gnd cell_6t
Xbit_r31_c83 bl[83] br[83] wl[31] vdd gnd cell_6t
Xbit_r32_c83 bl[83] br[83] wl[32] vdd gnd cell_6t
Xbit_r33_c83 bl[83] br[83] wl[33] vdd gnd cell_6t
Xbit_r34_c83 bl[83] br[83] wl[34] vdd gnd cell_6t
Xbit_r35_c83 bl[83] br[83] wl[35] vdd gnd cell_6t
Xbit_r36_c83 bl[83] br[83] wl[36] vdd gnd cell_6t
Xbit_r37_c83 bl[83] br[83] wl[37] vdd gnd cell_6t
Xbit_r38_c83 bl[83] br[83] wl[38] vdd gnd cell_6t
Xbit_r39_c83 bl[83] br[83] wl[39] vdd gnd cell_6t
Xbit_r40_c83 bl[83] br[83] wl[40] vdd gnd cell_6t
Xbit_r41_c83 bl[83] br[83] wl[41] vdd gnd cell_6t
Xbit_r42_c83 bl[83] br[83] wl[42] vdd gnd cell_6t
Xbit_r43_c83 bl[83] br[83] wl[43] vdd gnd cell_6t
Xbit_r44_c83 bl[83] br[83] wl[44] vdd gnd cell_6t
Xbit_r45_c83 bl[83] br[83] wl[45] vdd gnd cell_6t
Xbit_r46_c83 bl[83] br[83] wl[46] vdd gnd cell_6t
Xbit_r47_c83 bl[83] br[83] wl[47] vdd gnd cell_6t
Xbit_r48_c83 bl[83] br[83] wl[48] vdd gnd cell_6t
Xbit_r49_c83 bl[83] br[83] wl[49] vdd gnd cell_6t
Xbit_r50_c83 bl[83] br[83] wl[50] vdd gnd cell_6t
Xbit_r51_c83 bl[83] br[83] wl[51] vdd gnd cell_6t
Xbit_r52_c83 bl[83] br[83] wl[52] vdd gnd cell_6t
Xbit_r53_c83 bl[83] br[83] wl[53] vdd gnd cell_6t
Xbit_r54_c83 bl[83] br[83] wl[54] vdd gnd cell_6t
Xbit_r55_c83 bl[83] br[83] wl[55] vdd gnd cell_6t
Xbit_r56_c83 bl[83] br[83] wl[56] vdd gnd cell_6t
Xbit_r57_c83 bl[83] br[83] wl[57] vdd gnd cell_6t
Xbit_r58_c83 bl[83] br[83] wl[58] vdd gnd cell_6t
Xbit_r59_c83 bl[83] br[83] wl[59] vdd gnd cell_6t
Xbit_r60_c83 bl[83] br[83] wl[60] vdd gnd cell_6t
Xbit_r61_c83 bl[83] br[83] wl[61] vdd gnd cell_6t
Xbit_r62_c83 bl[83] br[83] wl[62] vdd gnd cell_6t
Xbit_r63_c83 bl[83] br[83] wl[63] vdd gnd cell_6t
Xbit_r64_c83 bl[83] br[83] wl[64] vdd gnd cell_6t
Xbit_r65_c83 bl[83] br[83] wl[65] vdd gnd cell_6t
Xbit_r66_c83 bl[83] br[83] wl[66] vdd gnd cell_6t
Xbit_r67_c83 bl[83] br[83] wl[67] vdd gnd cell_6t
Xbit_r68_c83 bl[83] br[83] wl[68] vdd gnd cell_6t
Xbit_r69_c83 bl[83] br[83] wl[69] vdd gnd cell_6t
Xbit_r70_c83 bl[83] br[83] wl[70] vdd gnd cell_6t
Xbit_r71_c83 bl[83] br[83] wl[71] vdd gnd cell_6t
Xbit_r72_c83 bl[83] br[83] wl[72] vdd gnd cell_6t
Xbit_r73_c83 bl[83] br[83] wl[73] vdd gnd cell_6t
Xbit_r74_c83 bl[83] br[83] wl[74] vdd gnd cell_6t
Xbit_r75_c83 bl[83] br[83] wl[75] vdd gnd cell_6t
Xbit_r76_c83 bl[83] br[83] wl[76] vdd gnd cell_6t
Xbit_r77_c83 bl[83] br[83] wl[77] vdd gnd cell_6t
Xbit_r78_c83 bl[83] br[83] wl[78] vdd gnd cell_6t
Xbit_r79_c83 bl[83] br[83] wl[79] vdd gnd cell_6t
Xbit_r80_c83 bl[83] br[83] wl[80] vdd gnd cell_6t
Xbit_r81_c83 bl[83] br[83] wl[81] vdd gnd cell_6t
Xbit_r82_c83 bl[83] br[83] wl[82] vdd gnd cell_6t
Xbit_r83_c83 bl[83] br[83] wl[83] vdd gnd cell_6t
Xbit_r84_c83 bl[83] br[83] wl[84] vdd gnd cell_6t
Xbit_r85_c83 bl[83] br[83] wl[85] vdd gnd cell_6t
Xbit_r86_c83 bl[83] br[83] wl[86] vdd gnd cell_6t
Xbit_r87_c83 bl[83] br[83] wl[87] vdd gnd cell_6t
Xbit_r88_c83 bl[83] br[83] wl[88] vdd gnd cell_6t
Xbit_r89_c83 bl[83] br[83] wl[89] vdd gnd cell_6t
Xbit_r90_c83 bl[83] br[83] wl[90] vdd gnd cell_6t
Xbit_r91_c83 bl[83] br[83] wl[91] vdd gnd cell_6t
Xbit_r92_c83 bl[83] br[83] wl[92] vdd gnd cell_6t
Xbit_r93_c83 bl[83] br[83] wl[93] vdd gnd cell_6t
Xbit_r94_c83 bl[83] br[83] wl[94] vdd gnd cell_6t
Xbit_r95_c83 bl[83] br[83] wl[95] vdd gnd cell_6t
Xbit_r96_c83 bl[83] br[83] wl[96] vdd gnd cell_6t
Xbit_r97_c83 bl[83] br[83] wl[97] vdd gnd cell_6t
Xbit_r98_c83 bl[83] br[83] wl[98] vdd gnd cell_6t
Xbit_r99_c83 bl[83] br[83] wl[99] vdd gnd cell_6t
Xbit_r100_c83 bl[83] br[83] wl[100] vdd gnd cell_6t
Xbit_r101_c83 bl[83] br[83] wl[101] vdd gnd cell_6t
Xbit_r102_c83 bl[83] br[83] wl[102] vdd gnd cell_6t
Xbit_r103_c83 bl[83] br[83] wl[103] vdd gnd cell_6t
Xbit_r104_c83 bl[83] br[83] wl[104] vdd gnd cell_6t
Xbit_r105_c83 bl[83] br[83] wl[105] vdd gnd cell_6t
Xbit_r106_c83 bl[83] br[83] wl[106] vdd gnd cell_6t
Xbit_r107_c83 bl[83] br[83] wl[107] vdd gnd cell_6t
Xbit_r108_c83 bl[83] br[83] wl[108] vdd gnd cell_6t
Xbit_r109_c83 bl[83] br[83] wl[109] vdd gnd cell_6t
Xbit_r110_c83 bl[83] br[83] wl[110] vdd gnd cell_6t
Xbit_r111_c83 bl[83] br[83] wl[111] vdd gnd cell_6t
Xbit_r112_c83 bl[83] br[83] wl[112] vdd gnd cell_6t
Xbit_r113_c83 bl[83] br[83] wl[113] vdd gnd cell_6t
Xbit_r114_c83 bl[83] br[83] wl[114] vdd gnd cell_6t
Xbit_r115_c83 bl[83] br[83] wl[115] vdd gnd cell_6t
Xbit_r116_c83 bl[83] br[83] wl[116] vdd gnd cell_6t
Xbit_r117_c83 bl[83] br[83] wl[117] vdd gnd cell_6t
Xbit_r118_c83 bl[83] br[83] wl[118] vdd gnd cell_6t
Xbit_r119_c83 bl[83] br[83] wl[119] vdd gnd cell_6t
Xbit_r120_c83 bl[83] br[83] wl[120] vdd gnd cell_6t
Xbit_r121_c83 bl[83] br[83] wl[121] vdd gnd cell_6t
Xbit_r122_c83 bl[83] br[83] wl[122] vdd gnd cell_6t
Xbit_r123_c83 bl[83] br[83] wl[123] vdd gnd cell_6t
Xbit_r124_c83 bl[83] br[83] wl[124] vdd gnd cell_6t
Xbit_r125_c83 bl[83] br[83] wl[125] vdd gnd cell_6t
Xbit_r126_c83 bl[83] br[83] wl[126] vdd gnd cell_6t
Xbit_r127_c83 bl[83] br[83] wl[127] vdd gnd cell_6t
Xbit_r128_c83 bl[83] br[83] wl[128] vdd gnd cell_6t
Xbit_r129_c83 bl[83] br[83] wl[129] vdd gnd cell_6t
Xbit_r130_c83 bl[83] br[83] wl[130] vdd gnd cell_6t
Xbit_r131_c83 bl[83] br[83] wl[131] vdd gnd cell_6t
Xbit_r132_c83 bl[83] br[83] wl[132] vdd gnd cell_6t
Xbit_r133_c83 bl[83] br[83] wl[133] vdd gnd cell_6t
Xbit_r134_c83 bl[83] br[83] wl[134] vdd gnd cell_6t
Xbit_r135_c83 bl[83] br[83] wl[135] vdd gnd cell_6t
Xbit_r136_c83 bl[83] br[83] wl[136] vdd gnd cell_6t
Xbit_r137_c83 bl[83] br[83] wl[137] vdd gnd cell_6t
Xbit_r138_c83 bl[83] br[83] wl[138] vdd gnd cell_6t
Xbit_r139_c83 bl[83] br[83] wl[139] vdd gnd cell_6t
Xbit_r140_c83 bl[83] br[83] wl[140] vdd gnd cell_6t
Xbit_r141_c83 bl[83] br[83] wl[141] vdd gnd cell_6t
Xbit_r142_c83 bl[83] br[83] wl[142] vdd gnd cell_6t
Xbit_r143_c83 bl[83] br[83] wl[143] vdd gnd cell_6t
Xbit_r144_c83 bl[83] br[83] wl[144] vdd gnd cell_6t
Xbit_r145_c83 bl[83] br[83] wl[145] vdd gnd cell_6t
Xbit_r146_c83 bl[83] br[83] wl[146] vdd gnd cell_6t
Xbit_r147_c83 bl[83] br[83] wl[147] vdd gnd cell_6t
Xbit_r148_c83 bl[83] br[83] wl[148] vdd gnd cell_6t
Xbit_r149_c83 bl[83] br[83] wl[149] vdd gnd cell_6t
Xbit_r150_c83 bl[83] br[83] wl[150] vdd gnd cell_6t
Xbit_r151_c83 bl[83] br[83] wl[151] vdd gnd cell_6t
Xbit_r152_c83 bl[83] br[83] wl[152] vdd gnd cell_6t
Xbit_r153_c83 bl[83] br[83] wl[153] vdd gnd cell_6t
Xbit_r154_c83 bl[83] br[83] wl[154] vdd gnd cell_6t
Xbit_r155_c83 bl[83] br[83] wl[155] vdd gnd cell_6t
Xbit_r156_c83 bl[83] br[83] wl[156] vdd gnd cell_6t
Xbit_r157_c83 bl[83] br[83] wl[157] vdd gnd cell_6t
Xbit_r158_c83 bl[83] br[83] wl[158] vdd gnd cell_6t
Xbit_r159_c83 bl[83] br[83] wl[159] vdd gnd cell_6t
Xbit_r160_c83 bl[83] br[83] wl[160] vdd gnd cell_6t
Xbit_r161_c83 bl[83] br[83] wl[161] vdd gnd cell_6t
Xbit_r162_c83 bl[83] br[83] wl[162] vdd gnd cell_6t
Xbit_r163_c83 bl[83] br[83] wl[163] vdd gnd cell_6t
Xbit_r164_c83 bl[83] br[83] wl[164] vdd gnd cell_6t
Xbit_r165_c83 bl[83] br[83] wl[165] vdd gnd cell_6t
Xbit_r166_c83 bl[83] br[83] wl[166] vdd gnd cell_6t
Xbit_r167_c83 bl[83] br[83] wl[167] vdd gnd cell_6t
Xbit_r168_c83 bl[83] br[83] wl[168] vdd gnd cell_6t
Xbit_r169_c83 bl[83] br[83] wl[169] vdd gnd cell_6t
Xbit_r170_c83 bl[83] br[83] wl[170] vdd gnd cell_6t
Xbit_r171_c83 bl[83] br[83] wl[171] vdd gnd cell_6t
Xbit_r172_c83 bl[83] br[83] wl[172] vdd gnd cell_6t
Xbit_r173_c83 bl[83] br[83] wl[173] vdd gnd cell_6t
Xbit_r174_c83 bl[83] br[83] wl[174] vdd gnd cell_6t
Xbit_r175_c83 bl[83] br[83] wl[175] vdd gnd cell_6t
Xbit_r176_c83 bl[83] br[83] wl[176] vdd gnd cell_6t
Xbit_r177_c83 bl[83] br[83] wl[177] vdd gnd cell_6t
Xbit_r178_c83 bl[83] br[83] wl[178] vdd gnd cell_6t
Xbit_r179_c83 bl[83] br[83] wl[179] vdd gnd cell_6t
Xbit_r180_c83 bl[83] br[83] wl[180] vdd gnd cell_6t
Xbit_r181_c83 bl[83] br[83] wl[181] vdd gnd cell_6t
Xbit_r182_c83 bl[83] br[83] wl[182] vdd gnd cell_6t
Xbit_r183_c83 bl[83] br[83] wl[183] vdd gnd cell_6t
Xbit_r184_c83 bl[83] br[83] wl[184] vdd gnd cell_6t
Xbit_r185_c83 bl[83] br[83] wl[185] vdd gnd cell_6t
Xbit_r186_c83 bl[83] br[83] wl[186] vdd gnd cell_6t
Xbit_r187_c83 bl[83] br[83] wl[187] vdd gnd cell_6t
Xbit_r188_c83 bl[83] br[83] wl[188] vdd gnd cell_6t
Xbit_r189_c83 bl[83] br[83] wl[189] vdd gnd cell_6t
Xbit_r190_c83 bl[83] br[83] wl[190] vdd gnd cell_6t
Xbit_r191_c83 bl[83] br[83] wl[191] vdd gnd cell_6t
Xbit_r192_c83 bl[83] br[83] wl[192] vdd gnd cell_6t
Xbit_r193_c83 bl[83] br[83] wl[193] vdd gnd cell_6t
Xbit_r194_c83 bl[83] br[83] wl[194] vdd gnd cell_6t
Xbit_r195_c83 bl[83] br[83] wl[195] vdd gnd cell_6t
Xbit_r196_c83 bl[83] br[83] wl[196] vdd gnd cell_6t
Xbit_r197_c83 bl[83] br[83] wl[197] vdd gnd cell_6t
Xbit_r198_c83 bl[83] br[83] wl[198] vdd gnd cell_6t
Xbit_r199_c83 bl[83] br[83] wl[199] vdd gnd cell_6t
Xbit_r200_c83 bl[83] br[83] wl[200] vdd gnd cell_6t
Xbit_r201_c83 bl[83] br[83] wl[201] vdd gnd cell_6t
Xbit_r202_c83 bl[83] br[83] wl[202] vdd gnd cell_6t
Xbit_r203_c83 bl[83] br[83] wl[203] vdd gnd cell_6t
Xbit_r204_c83 bl[83] br[83] wl[204] vdd gnd cell_6t
Xbit_r205_c83 bl[83] br[83] wl[205] vdd gnd cell_6t
Xbit_r206_c83 bl[83] br[83] wl[206] vdd gnd cell_6t
Xbit_r207_c83 bl[83] br[83] wl[207] vdd gnd cell_6t
Xbit_r208_c83 bl[83] br[83] wl[208] vdd gnd cell_6t
Xbit_r209_c83 bl[83] br[83] wl[209] vdd gnd cell_6t
Xbit_r210_c83 bl[83] br[83] wl[210] vdd gnd cell_6t
Xbit_r211_c83 bl[83] br[83] wl[211] vdd gnd cell_6t
Xbit_r212_c83 bl[83] br[83] wl[212] vdd gnd cell_6t
Xbit_r213_c83 bl[83] br[83] wl[213] vdd gnd cell_6t
Xbit_r214_c83 bl[83] br[83] wl[214] vdd gnd cell_6t
Xbit_r215_c83 bl[83] br[83] wl[215] vdd gnd cell_6t
Xbit_r216_c83 bl[83] br[83] wl[216] vdd gnd cell_6t
Xbit_r217_c83 bl[83] br[83] wl[217] vdd gnd cell_6t
Xbit_r218_c83 bl[83] br[83] wl[218] vdd gnd cell_6t
Xbit_r219_c83 bl[83] br[83] wl[219] vdd gnd cell_6t
Xbit_r220_c83 bl[83] br[83] wl[220] vdd gnd cell_6t
Xbit_r221_c83 bl[83] br[83] wl[221] vdd gnd cell_6t
Xbit_r222_c83 bl[83] br[83] wl[222] vdd gnd cell_6t
Xbit_r223_c83 bl[83] br[83] wl[223] vdd gnd cell_6t
Xbit_r224_c83 bl[83] br[83] wl[224] vdd gnd cell_6t
Xbit_r225_c83 bl[83] br[83] wl[225] vdd gnd cell_6t
Xbit_r226_c83 bl[83] br[83] wl[226] vdd gnd cell_6t
Xbit_r227_c83 bl[83] br[83] wl[227] vdd gnd cell_6t
Xbit_r228_c83 bl[83] br[83] wl[228] vdd gnd cell_6t
Xbit_r229_c83 bl[83] br[83] wl[229] vdd gnd cell_6t
Xbit_r230_c83 bl[83] br[83] wl[230] vdd gnd cell_6t
Xbit_r231_c83 bl[83] br[83] wl[231] vdd gnd cell_6t
Xbit_r232_c83 bl[83] br[83] wl[232] vdd gnd cell_6t
Xbit_r233_c83 bl[83] br[83] wl[233] vdd gnd cell_6t
Xbit_r234_c83 bl[83] br[83] wl[234] vdd gnd cell_6t
Xbit_r235_c83 bl[83] br[83] wl[235] vdd gnd cell_6t
Xbit_r236_c83 bl[83] br[83] wl[236] vdd gnd cell_6t
Xbit_r237_c83 bl[83] br[83] wl[237] vdd gnd cell_6t
Xbit_r238_c83 bl[83] br[83] wl[238] vdd gnd cell_6t
Xbit_r239_c83 bl[83] br[83] wl[239] vdd gnd cell_6t
Xbit_r240_c83 bl[83] br[83] wl[240] vdd gnd cell_6t
Xbit_r241_c83 bl[83] br[83] wl[241] vdd gnd cell_6t
Xbit_r242_c83 bl[83] br[83] wl[242] vdd gnd cell_6t
Xbit_r243_c83 bl[83] br[83] wl[243] vdd gnd cell_6t
Xbit_r244_c83 bl[83] br[83] wl[244] vdd gnd cell_6t
Xbit_r245_c83 bl[83] br[83] wl[245] vdd gnd cell_6t
Xbit_r246_c83 bl[83] br[83] wl[246] vdd gnd cell_6t
Xbit_r247_c83 bl[83] br[83] wl[247] vdd gnd cell_6t
Xbit_r248_c83 bl[83] br[83] wl[248] vdd gnd cell_6t
Xbit_r249_c83 bl[83] br[83] wl[249] vdd gnd cell_6t
Xbit_r250_c83 bl[83] br[83] wl[250] vdd gnd cell_6t
Xbit_r251_c83 bl[83] br[83] wl[251] vdd gnd cell_6t
Xbit_r252_c83 bl[83] br[83] wl[252] vdd gnd cell_6t
Xbit_r253_c83 bl[83] br[83] wl[253] vdd gnd cell_6t
Xbit_r254_c83 bl[83] br[83] wl[254] vdd gnd cell_6t
Xbit_r255_c83 bl[83] br[83] wl[255] vdd gnd cell_6t
Xbit_r0_c84 bl[84] br[84] wl[0] vdd gnd cell_6t
Xbit_r1_c84 bl[84] br[84] wl[1] vdd gnd cell_6t
Xbit_r2_c84 bl[84] br[84] wl[2] vdd gnd cell_6t
Xbit_r3_c84 bl[84] br[84] wl[3] vdd gnd cell_6t
Xbit_r4_c84 bl[84] br[84] wl[4] vdd gnd cell_6t
Xbit_r5_c84 bl[84] br[84] wl[5] vdd gnd cell_6t
Xbit_r6_c84 bl[84] br[84] wl[6] vdd gnd cell_6t
Xbit_r7_c84 bl[84] br[84] wl[7] vdd gnd cell_6t
Xbit_r8_c84 bl[84] br[84] wl[8] vdd gnd cell_6t
Xbit_r9_c84 bl[84] br[84] wl[9] vdd gnd cell_6t
Xbit_r10_c84 bl[84] br[84] wl[10] vdd gnd cell_6t
Xbit_r11_c84 bl[84] br[84] wl[11] vdd gnd cell_6t
Xbit_r12_c84 bl[84] br[84] wl[12] vdd gnd cell_6t
Xbit_r13_c84 bl[84] br[84] wl[13] vdd gnd cell_6t
Xbit_r14_c84 bl[84] br[84] wl[14] vdd gnd cell_6t
Xbit_r15_c84 bl[84] br[84] wl[15] vdd gnd cell_6t
Xbit_r16_c84 bl[84] br[84] wl[16] vdd gnd cell_6t
Xbit_r17_c84 bl[84] br[84] wl[17] vdd gnd cell_6t
Xbit_r18_c84 bl[84] br[84] wl[18] vdd gnd cell_6t
Xbit_r19_c84 bl[84] br[84] wl[19] vdd gnd cell_6t
Xbit_r20_c84 bl[84] br[84] wl[20] vdd gnd cell_6t
Xbit_r21_c84 bl[84] br[84] wl[21] vdd gnd cell_6t
Xbit_r22_c84 bl[84] br[84] wl[22] vdd gnd cell_6t
Xbit_r23_c84 bl[84] br[84] wl[23] vdd gnd cell_6t
Xbit_r24_c84 bl[84] br[84] wl[24] vdd gnd cell_6t
Xbit_r25_c84 bl[84] br[84] wl[25] vdd gnd cell_6t
Xbit_r26_c84 bl[84] br[84] wl[26] vdd gnd cell_6t
Xbit_r27_c84 bl[84] br[84] wl[27] vdd gnd cell_6t
Xbit_r28_c84 bl[84] br[84] wl[28] vdd gnd cell_6t
Xbit_r29_c84 bl[84] br[84] wl[29] vdd gnd cell_6t
Xbit_r30_c84 bl[84] br[84] wl[30] vdd gnd cell_6t
Xbit_r31_c84 bl[84] br[84] wl[31] vdd gnd cell_6t
Xbit_r32_c84 bl[84] br[84] wl[32] vdd gnd cell_6t
Xbit_r33_c84 bl[84] br[84] wl[33] vdd gnd cell_6t
Xbit_r34_c84 bl[84] br[84] wl[34] vdd gnd cell_6t
Xbit_r35_c84 bl[84] br[84] wl[35] vdd gnd cell_6t
Xbit_r36_c84 bl[84] br[84] wl[36] vdd gnd cell_6t
Xbit_r37_c84 bl[84] br[84] wl[37] vdd gnd cell_6t
Xbit_r38_c84 bl[84] br[84] wl[38] vdd gnd cell_6t
Xbit_r39_c84 bl[84] br[84] wl[39] vdd gnd cell_6t
Xbit_r40_c84 bl[84] br[84] wl[40] vdd gnd cell_6t
Xbit_r41_c84 bl[84] br[84] wl[41] vdd gnd cell_6t
Xbit_r42_c84 bl[84] br[84] wl[42] vdd gnd cell_6t
Xbit_r43_c84 bl[84] br[84] wl[43] vdd gnd cell_6t
Xbit_r44_c84 bl[84] br[84] wl[44] vdd gnd cell_6t
Xbit_r45_c84 bl[84] br[84] wl[45] vdd gnd cell_6t
Xbit_r46_c84 bl[84] br[84] wl[46] vdd gnd cell_6t
Xbit_r47_c84 bl[84] br[84] wl[47] vdd gnd cell_6t
Xbit_r48_c84 bl[84] br[84] wl[48] vdd gnd cell_6t
Xbit_r49_c84 bl[84] br[84] wl[49] vdd gnd cell_6t
Xbit_r50_c84 bl[84] br[84] wl[50] vdd gnd cell_6t
Xbit_r51_c84 bl[84] br[84] wl[51] vdd gnd cell_6t
Xbit_r52_c84 bl[84] br[84] wl[52] vdd gnd cell_6t
Xbit_r53_c84 bl[84] br[84] wl[53] vdd gnd cell_6t
Xbit_r54_c84 bl[84] br[84] wl[54] vdd gnd cell_6t
Xbit_r55_c84 bl[84] br[84] wl[55] vdd gnd cell_6t
Xbit_r56_c84 bl[84] br[84] wl[56] vdd gnd cell_6t
Xbit_r57_c84 bl[84] br[84] wl[57] vdd gnd cell_6t
Xbit_r58_c84 bl[84] br[84] wl[58] vdd gnd cell_6t
Xbit_r59_c84 bl[84] br[84] wl[59] vdd gnd cell_6t
Xbit_r60_c84 bl[84] br[84] wl[60] vdd gnd cell_6t
Xbit_r61_c84 bl[84] br[84] wl[61] vdd gnd cell_6t
Xbit_r62_c84 bl[84] br[84] wl[62] vdd gnd cell_6t
Xbit_r63_c84 bl[84] br[84] wl[63] vdd gnd cell_6t
Xbit_r64_c84 bl[84] br[84] wl[64] vdd gnd cell_6t
Xbit_r65_c84 bl[84] br[84] wl[65] vdd gnd cell_6t
Xbit_r66_c84 bl[84] br[84] wl[66] vdd gnd cell_6t
Xbit_r67_c84 bl[84] br[84] wl[67] vdd gnd cell_6t
Xbit_r68_c84 bl[84] br[84] wl[68] vdd gnd cell_6t
Xbit_r69_c84 bl[84] br[84] wl[69] vdd gnd cell_6t
Xbit_r70_c84 bl[84] br[84] wl[70] vdd gnd cell_6t
Xbit_r71_c84 bl[84] br[84] wl[71] vdd gnd cell_6t
Xbit_r72_c84 bl[84] br[84] wl[72] vdd gnd cell_6t
Xbit_r73_c84 bl[84] br[84] wl[73] vdd gnd cell_6t
Xbit_r74_c84 bl[84] br[84] wl[74] vdd gnd cell_6t
Xbit_r75_c84 bl[84] br[84] wl[75] vdd gnd cell_6t
Xbit_r76_c84 bl[84] br[84] wl[76] vdd gnd cell_6t
Xbit_r77_c84 bl[84] br[84] wl[77] vdd gnd cell_6t
Xbit_r78_c84 bl[84] br[84] wl[78] vdd gnd cell_6t
Xbit_r79_c84 bl[84] br[84] wl[79] vdd gnd cell_6t
Xbit_r80_c84 bl[84] br[84] wl[80] vdd gnd cell_6t
Xbit_r81_c84 bl[84] br[84] wl[81] vdd gnd cell_6t
Xbit_r82_c84 bl[84] br[84] wl[82] vdd gnd cell_6t
Xbit_r83_c84 bl[84] br[84] wl[83] vdd gnd cell_6t
Xbit_r84_c84 bl[84] br[84] wl[84] vdd gnd cell_6t
Xbit_r85_c84 bl[84] br[84] wl[85] vdd gnd cell_6t
Xbit_r86_c84 bl[84] br[84] wl[86] vdd gnd cell_6t
Xbit_r87_c84 bl[84] br[84] wl[87] vdd gnd cell_6t
Xbit_r88_c84 bl[84] br[84] wl[88] vdd gnd cell_6t
Xbit_r89_c84 bl[84] br[84] wl[89] vdd gnd cell_6t
Xbit_r90_c84 bl[84] br[84] wl[90] vdd gnd cell_6t
Xbit_r91_c84 bl[84] br[84] wl[91] vdd gnd cell_6t
Xbit_r92_c84 bl[84] br[84] wl[92] vdd gnd cell_6t
Xbit_r93_c84 bl[84] br[84] wl[93] vdd gnd cell_6t
Xbit_r94_c84 bl[84] br[84] wl[94] vdd gnd cell_6t
Xbit_r95_c84 bl[84] br[84] wl[95] vdd gnd cell_6t
Xbit_r96_c84 bl[84] br[84] wl[96] vdd gnd cell_6t
Xbit_r97_c84 bl[84] br[84] wl[97] vdd gnd cell_6t
Xbit_r98_c84 bl[84] br[84] wl[98] vdd gnd cell_6t
Xbit_r99_c84 bl[84] br[84] wl[99] vdd gnd cell_6t
Xbit_r100_c84 bl[84] br[84] wl[100] vdd gnd cell_6t
Xbit_r101_c84 bl[84] br[84] wl[101] vdd gnd cell_6t
Xbit_r102_c84 bl[84] br[84] wl[102] vdd gnd cell_6t
Xbit_r103_c84 bl[84] br[84] wl[103] vdd gnd cell_6t
Xbit_r104_c84 bl[84] br[84] wl[104] vdd gnd cell_6t
Xbit_r105_c84 bl[84] br[84] wl[105] vdd gnd cell_6t
Xbit_r106_c84 bl[84] br[84] wl[106] vdd gnd cell_6t
Xbit_r107_c84 bl[84] br[84] wl[107] vdd gnd cell_6t
Xbit_r108_c84 bl[84] br[84] wl[108] vdd gnd cell_6t
Xbit_r109_c84 bl[84] br[84] wl[109] vdd gnd cell_6t
Xbit_r110_c84 bl[84] br[84] wl[110] vdd gnd cell_6t
Xbit_r111_c84 bl[84] br[84] wl[111] vdd gnd cell_6t
Xbit_r112_c84 bl[84] br[84] wl[112] vdd gnd cell_6t
Xbit_r113_c84 bl[84] br[84] wl[113] vdd gnd cell_6t
Xbit_r114_c84 bl[84] br[84] wl[114] vdd gnd cell_6t
Xbit_r115_c84 bl[84] br[84] wl[115] vdd gnd cell_6t
Xbit_r116_c84 bl[84] br[84] wl[116] vdd gnd cell_6t
Xbit_r117_c84 bl[84] br[84] wl[117] vdd gnd cell_6t
Xbit_r118_c84 bl[84] br[84] wl[118] vdd gnd cell_6t
Xbit_r119_c84 bl[84] br[84] wl[119] vdd gnd cell_6t
Xbit_r120_c84 bl[84] br[84] wl[120] vdd gnd cell_6t
Xbit_r121_c84 bl[84] br[84] wl[121] vdd gnd cell_6t
Xbit_r122_c84 bl[84] br[84] wl[122] vdd gnd cell_6t
Xbit_r123_c84 bl[84] br[84] wl[123] vdd gnd cell_6t
Xbit_r124_c84 bl[84] br[84] wl[124] vdd gnd cell_6t
Xbit_r125_c84 bl[84] br[84] wl[125] vdd gnd cell_6t
Xbit_r126_c84 bl[84] br[84] wl[126] vdd gnd cell_6t
Xbit_r127_c84 bl[84] br[84] wl[127] vdd gnd cell_6t
Xbit_r128_c84 bl[84] br[84] wl[128] vdd gnd cell_6t
Xbit_r129_c84 bl[84] br[84] wl[129] vdd gnd cell_6t
Xbit_r130_c84 bl[84] br[84] wl[130] vdd gnd cell_6t
Xbit_r131_c84 bl[84] br[84] wl[131] vdd gnd cell_6t
Xbit_r132_c84 bl[84] br[84] wl[132] vdd gnd cell_6t
Xbit_r133_c84 bl[84] br[84] wl[133] vdd gnd cell_6t
Xbit_r134_c84 bl[84] br[84] wl[134] vdd gnd cell_6t
Xbit_r135_c84 bl[84] br[84] wl[135] vdd gnd cell_6t
Xbit_r136_c84 bl[84] br[84] wl[136] vdd gnd cell_6t
Xbit_r137_c84 bl[84] br[84] wl[137] vdd gnd cell_6t
Xbit_r138_c84 bl[84] br[84] wl[138] vdd gnd cell_6t
Xbit_r139_c84 bl[84] br[84] wl[139] vdd gnd cell_6t
Xbit_r140_c84 bl[84] br[84] wl[140] vdd gnd cell_6t
Xbit_r141_c84 bl[84] br[84] wl[141] vdd gnd cell_6t
Xbit_r142_c84 bl[84] br[84] wl[142] vdd gnd cell_6t
Xbit_r143_c84 bl[84] br[84] wl[143] vdd gnd cell_6t
Xbit_r144_c84 bl[84] br[84] wl[144] vdd gnd cell_6t
Xbit_r145_c84 bl[84] br[84] wl[145] vdd gnd cell_6t
Xbit_r146_c84 bl[84] br[84] wl[146] vdd gnd cell_6t
Xbit_r147_c84 bl[84] br[84] wl[147] vdd gnd cell_6t
Xbit_r148_c84 bl[84] br[84] wl[148] vdd gnd cell_6t
Xbit_r149_c84 bl[84] br[84] wl[149] vdd gnd cell_6t
Xbit_r150_c84 bl[84] br[84] wl[150] vdd gnd cell_6t
Xbit_r151_c84 bl[84] br[84] wl[151] vdd gnd cell_6t
Xbit_r152_c84 bl[84] br[84] wl[152] vdd gnd cell_6t
Xbit_r153_c84 bl[84] br[84] wl[153] vdd gnd cell_6t
Xbit_r154_c84 bl[84] br[84] wl[154] vdd gnd cell_6t
Xbit_r155_c84 bl[84] br[84] wl[155] vdd gnd cell_6t
Xbit_r156_c84 bl[84] br[84] wl[156] vdd gnd cell_6t
Xbit_r157_c84 bl[84] br[84] wl[157] vdd gnd cell_6t
Xbit_r158_c84 bl[84] br[84] wl[158] vdd gnd cell_6t
Xbit_r159_c84 bl[84] br[84] wl[159] vdd gnd cell_6t
Xbit_r160_c84 bl[84] br[84] wl[160] vdd gnd cell_6t
Xbit_r161_c84 bl[84] br[84] wl[161] vdd gnd cell_6t
Xbit_r162_c84 bl[84] br[84] wl[162] vdd gnd cell_6t
Xbit_r163_c84 bl[84] br[84] wl[163] vdd gnd cell_6t
Xbit_r164_c84 bl[84] br[84] wl[164] vdd gnd cell_6t
Xbit_r165_c84 bl[84] br[84] wl[165] vdd gnd cell_6t
Xbit_r166_c84 bl[84] br[84] wl[166] vdd gnd cell_6t
Xbit_r167_c84 bl[84] br[84] wl[167] vdd gnd cell_6t
Xbit_r168_c84 bl[84] br[84] wl[168] vdd gnd cell_6t
Xbit_r169_c84 bl[84] br[84] wl[169] vdd gnd cell_6t
Xbit_r170_c84 bl[84] br[84] wl[170] vdd gnd cell_6t
Xbit_r171_c84 bl[84] br[84] wl[171] vdd gnd cell_6t
Xbit_r172_c84 bl[84] br[84] wl[172] vdd gnd cell_6t
Xbit_r173_c84 bl[84] br[84] wl[173] vdd gnd cell_6t
Xbit_r174_c84 bl[84] br[84] wl[174] vdd gnd cell_6t
Xbit_r175_c84 bl[84] br[84] wl[175] vdd gnd cell_6t
Xbit_r176_c84 bl[84] br[84] wl[176] vdd gnd cell_6t
Xbit_r177_c84 bl[84] br[84] wl[177] vdd gnd cell_6t
Xbit_r178_c84 bl[84] br[84] wl[178] vdd gnd cell_6t
Xbit_r179_c84 bl[84] br[84] wl[179] vdd gnd cell_6t
Xbit_r180_c84 bl[84] br[84] wl[180] vdd gnd cell_6t
Xbit_r181_c84 bl[84] br[84] wl[181] vdd gnd cell_6t
Xbit_r182_c84 bl[84] br[84] wl[182] vdd gnd cell_6t
Xbit_r183_c84 bl[84] br[84] wl[183] vdd gnd cell_6t
Xbit_r184_c84 bl[84] br[84] wl[184] vdd gnd cell_6t
Xbit_r185_c84 bl[84] br[84] wl[185] vdd gnd cell_6t
Xbit_r186_c84 bl[84] br[84] wl[186] vdd gnd cell_6t
Xbit_r187_c84 bl[84] br[84] wl[187] vdd gnd cell_6t
Xbit_r188_c84 bl[84] br[84] wl[188] vdd gnd cell_6t
Xbit_r189_c84 bl[84] br[84] wl[189] vdd gnd cell_6t
Xbit_r190_c84 bl[84] br[84] wl[190] vdd gnd cell_6t
Xbit_r191_c84 bl[84] br[84] wl[191] vdd gnd cell_6t
Xbit_r192_c84 bl[84] br[84] wl[192] vdd gnd cell_6t
Xbit_r193_c84 bl[84] br[84] wl[193] vdd gnd cell_6t
Xbit_r194_c84 bl[84] br[84] wl[194] vdd gnd cell_6t
Xbit_r195_c84 bl[84] br[84] wl[195] vdd gnd cell_6t
Xbit_r196_c84 bl[84] br[84] wl[196] vdd gnd cell_6t
Xbit_r197_c84 bl[84] br[84] wl[197] vdd gnd cell_6t
Xbit_r198_c84 bl[84] br[84] wl[198] vdd gnd cell_6t
Xbit_r199_c84 bl[84] br[84] wl[199] vdd gnd cell_6t
Xbit_r200_c84 bl[84] br[84] wl[200] vdd gnd cell_6t
Xbit_r201_c84 bl[84] br[84] wl[201] vdd gnd cell_6t
Xbit_r202_c84 bl[84] br[84] wl[202] vdd gnd cell_6t
Xbit_r203_c84 bl[84] br[84] wl[203] vdd gnd cell_6t
Xbit_r204_c84 bl[84] br[84] wl[204] vdd gnd cell_6t
Xbit_r205_c84 bl[84] br[84] wl[205] vdd gnd cell_6t
Xbit_r206_c84 bl[84] br[84] wl[206] vdd gnd cell_6t
Xbit_r207_c84 bl[84] br[84] wl[207] vdd gnd cell_6t
Xbit_r208_c84 bl[84] br[84] wl[208] vdd gnd cell_6t
Xbit_r209_c84 bl[84] br[84] wl[209] vdd gnd cell_6t
Xbit_r210_c84 bl[84] br[84] wl[210] vdd gnd cell_6t
Xbit_r211_c84 bl[84] br[84] wl[211] vdd gnd cell_6t
Xbit_r212_c84 bl[84] br[84] wl[212] vdd gnd cell_6t
Xbit_r213_c84 bl[84] br[84] wl[213] vdd gnd cell_6t
Xbit_r214_c84 bl[84] br[84] wl[214] vdd gnd cell_6t
Xbit_r215_c84 bl[84] br[84] wl[215] vdd gnd cell_6t
Xbit_r216_c84 bl[84] br[84] wl[216] vdd gnd cell_6t
Xbit_r217_c84 bl[84] br[84] wl[217] vdd gnd cell_6t
Xbit_r218_c84 bl[84] br[84] wl[218] vdd gnd cell_6t
Xbit_r219_c84 bl[84] br[84] wl[219] vdd gnd cell_6t
Xbit_r220_c84 bl[84] br[84] wl[220] vdd gnd cell_6t
Xbit_r221_c84 bl[84] br[84] wl[221] vdd gnd cell_6t
Xbit_r222_c84 bl[84] br[84] wl[222] vdd gnd cell_6t
Xbit_r223_c84 bl[84] br[84] wl[223] vdd gnd cell_6t
Xbit_r224_c84 bl[84] br[84] wl[224] vdd gnd cell_6t
Xbit_r225_c84 bl[84] br[84] wl[225] vdd gnd cell_6t
Xbit_r226_c84 bl[84] br[84] wl[226] vdd gnd cell_6t
Xbit_r227_c84 bl[84] br[84] wl[227] vdd gnd cell_6t
Xbit_r228_c84 bl[84] br[84] wl[228] vdd gnd cell_6t
Xbit_r229_c84 bl[84] br[84] wl[229] vdd gnd cell_6t
Xbit_r230_c84 bl[84] br[84] wl[230] vdd gnd cell_6t
Xbit_r231_c84 bl[84] br[84] wl[231] vdd gnd cell_6t
Xbit_r232_c84 bl[84] br[84] wl[232] vdd gnd cell_6t
Xbit_r233_c84 bl[84] br[84] wl[233] vdd gnd cell_6t
Xbit_r234_c84 bl[84] br[84] wl[234] vdd gnd cell_6t
Xbit_r235_c84 bl[84] br[84] wl[235] vdd gnd cell_6t
Xbit_r236_c84 bl[84] br[84] wl[236] vdd gnd cell_6t
Xbit_r237_c84 bl[84] br[84] wl[237] vdd gnd cell_6t
Xbit_r238_c84 bl[84] br[84] wl[238] vdd gnd cell_6t
Xbit_r239_c84 bl[84] br[84] wl[239] vdd gnd cell_6t
Xbit_r240_c84 bl[84] br[84] wl[240] vdd gnd cell_6t
Xbit_r241_c84 bl[84] br[84] wl[241] vdd gnd cell_6t
Xbit_r242_c84 bl[84] br[84] wl[242] vdd gnd cell_6t
Xbit_r243_c84 bl[84] br[84] wl[243] vdd gnd cell_6t
Xbit_r244_c84 bl[84] br[84] wl[244] vdd gnd cell_6t
Xbit_r245_c84 bl[84] br[84] wl[245] vdd gnd cell_6t
Xbit_r246_c84 bl[84] br[84] wl[246] vdd gnd cell_6t
Xbit_r247_c84 bl[84] br[84] wl[247] vdd gnd cell_6t
Xbit_r248_c84 bl[84] br[84] wl[248] vdd gnd cell_6t
Xbit_r249_c84 bl[84] br[84] wl[249] vdd gnd cell_6t
Xbit_r250_c84 bl[84] br[84] wl[250] vdd gnd cell_6t
Xbit_r251_c84 bl[84] br[84] wl[251] vdd gnd cell_6t
Xbit_r252_c84 bl[84] br[84] wl[252] vdd gnd cell_6t
Xbit_r253_c84 bl[84] br[84] wl[253] vdd gnd cell_6t
Xbit_r254_c84 bl[84] br[84] wl[254] vdd gnd cell_6t
Xbit_r255_c84 bl[84] br[84] wl[255] vdd gnd cell_6t
Xbit_r0_c85 bl[85] br[85] wl[0] vdd gnd cell_6t
Xbit_r1_c85 bl[85] br[85] wl[1] vdd gnd cell_6t
Xbit_r2_c85 bl[85] br[85] wl[2] vdd gnd cell_6t
Xbit_r3_c85 bl[85] br[85] wl[3] vdd gnd cell_6t
Xbit_r4_c85 bl[85] br[85] wl[4] vdd gnd cell_6t
Xbit_r5_c85 bl[85] br[85] wl[5] vdd gnd cell_6t
Xbit_r6_c85 bl[85] br[85] wl[6] vdd gnd cell_6t
Xbit_r7_c85 bl[85] br[85] wl[7] vdd gnd cell_6t
Xbit_r8_c85 bl[85] br[85] wl[8] vdd gnd cell_6t
Xbit_r9_c85 bl[85] br[85] wl[9] vdd gnd cell_6t
Xbit_r10_c85 bl[85] br[85] wl[10] vdd gnd cell_6t
Xbit_r11_c85 bl[85] br[85] wl[11] vdd gnd cell_6t
Xbit_r12_c85 bl[85] br[85] wl[12] vdd gnd cell_6t
Xbit_r13_c85 bl[85] br[85] wl[13] vdd gnd cell_6t
Xbit_r14_c85 bl[85] br[85] wl[14] vdd gnd cell_6t
Xbit_r15_c85 bl[85] br[85] wl[15] vdd gnd cell_6t
Xbit_r16_c85 bl[85] br[85] wl[16] vdd gnd cell_6t
Xbit_r17_c85 bl[85] br[85] wl[17] vdd gnd cell_6t
Xbit_r18_c85 bl[85] br[85] wl[18] vdd gnd cell_6t
Xbit_r19_c85 bl[85] br[85] wl[19] vdd gnd cell_6t
Xbit_r20_c85 bl[85] br[85] wl[20] vdd gnd cell_6t
Xbit_r21_c85 bl[85] br[85] wl[21] vdd gnd cell_6t
Xbit_r22_c85 bl[85] br[85] wl[22] vdd gnd cell_6t
Xbit_r23_c85 bl[85] br[85] wl[23] vdd gnd cell_6t
Xbit_r24_c85 bl[85] br[85] wl[24] vdd gnd cell_6t
Xbit_r25_c85 bl[85] br[85] wl[25] vdd gnd cell_6t
Xbit_r26_c85 bl[85] br[85] wl[26] vdd gnd cell_6t
Xbit_r27_c85 bl[85] br[85] wl[27] vdd gnd cell_6t
Xbit_r28_c85 bl[85] br[85] wl[28] vdd gnd cell_6t
Xbit_r29_c85 bl[85] br[85] wl[29] vdd gnd cell_6t
Xbit_r30_c85 bl[85] br[85] wl[30] vdd gnd cell_6t
Xbit_r31_c85 bl[85] br[85] wl[31] vdd gnd cell_6t
Xbit_r32_c85 bl[85] br[85] wl[32] vdd gnd cell_6t
Xbit_r33_c85 bl[85] br[85] wl[33] vdd gnd cell_6t
Xbit_r34_c85 bl[85] br[85] wl[34] vdd gnd cell_6t
Xbit_r35_c85 bl[85] br[85] wl[35] vdd gnd cell_6t
Xbit_r36_c85 bl[85] br[85] wl[36] vdd gnd cell_6t
Xbit_r37_c85 bl[85] br[85] wl[37] vdd gnd cell_6t
Xbit_r38_c85 bl[85] br[85] wl[38] vdd gnd cell_6t
Xbit_r39_c85 bl[85] br[85] wl[39] vdd gnd cell_6t
Xbit_r40_c85 bl[85] br[85] wl[40] vdd gnd cell_6t
Xbit_r41_c85 bl[85] br[85] wl[41] vdd gnd cell_6t
Xbit_r42_c85 bl[85] br[85] wl[42] vdd gnd cell_6t
Xbit_r43_c85 bl[85] br[85] wl[43] vdd gnd cell_6t
Xbit_r44_c85 bl[85] br[85] wl[44] vdd gnd cell_6t
Xbit_r45_c85 bl[85] br[85] wl[45] vdd gnd cell_6t
Xbit_r46_c85 bl[85] br[85] wl[46] vdd gnd cell_6t
Xbit_r47_c85 bl[85] br[85] wl[47] vdd gnd cell_6t
Xbit_r48_c85 bl[85] br[85] wl[48] vdd gnd cell_6t
Xbit_r49_c85 bl[85] br[85] wl[49] vdd gnd cell_6t
Xbit_r50_c85 bl[85] br[85] wl[50] vdd gnd cell_6t
Xbit_r51_c85 bl[85] br[85] wl[51] vdd gnd cell_6t
Xbit_r52_c85 bl[85] br[85] wl[52] vdd gnd cell_6t
Xbit_r53_c85 bl[85] br[85] wl[53] vdd gnd cell_6t
Xbit_r54_c85 bl[85] br[85] wl[54] vdd gnd cell_6t
Xbit_r55_c85 bl[85] br[85] wl[55] vdd gnd cell_6t
Xbit_r56_c85 bl[85] br[85] wl[56] vdd gnd cell_6t
Xbit_r57_c85 bl[85] br[85] wl[57] vdd gnd cell_6t
Xbit_r58_c85 bl[85] br[85] wl[58] vdd gnd cell_6t
Xbit_r59_c85 bl[85] br[85] wl[59] vdd gnd cell_6t
Xbit_r60_c85 bl[85] br[85] wl[60] vdd gnd cell_6t
Xbit_r61_c85 bl[85] br[85] wl[61] vdd gnd cell_6t
Xbit_r62_c85 bl[85] br[85] wl[62] vdd gnd cell_6t
Xbit_r63_c85 bl[85] br[85] wl[63] vdd gnd cell_6t
Xbit_r64_c85 bl[85] br[85] wl[64] vdd gnd cell_6t
Xbit_r65_c85 bl[85] br[85] wl[65] vdd gnd cell_6t
Xbit_r66_c85 bl[85] br[85] wl[66] vdd gnd cell_6t
Xbit_r67_c85 bl[85] br[85] wl[67] vdd gnd cell_6t
Xbit_r68_c85 bl[85] br[85] wl[68] vdd gnd cell_6t
Xbit_r69_c85 bl[85] br[85] wl[69] vdd gnd cell_6t
Xbit_r70_c85 bl[85] br[85] wl[70] vdd gnd cell_6t
Xbit_r71_c85 bl[85] br[85] wl[71] vdd gnd cell_6t
Xbit_r72_c85 bl[85] br[85] wl[72] vdd gnd cell_6t
Xbit_r73_c85 bl[85] br[85] wl[73] vdd gnd cell_6t
Xbit_r74_c85 bl[85] br[85] wl[74] vdd gnd cell_6t
Xbit_r75_c85 bl[85] br[85] wl[75] vdd gnd cell_6t
Xbit_r76_c85 bl[85] br[85] wl[76] vdd gnd cell_6t
Xbit_r77_c85 bl[85] br[85] wl[77] vdd gnd cell_6t
Xbit_r78_c85 bl[85] br[85] wl[78] vdd gnd cell_6t
Xbit_r79_c85 bl[85] br[85] wl[79] vdd gnd cell_6t
Xbit_r80_c85 bl[85] br[85] wl[80] vdd gnd cell_6t
Xbit_r81_c85 bl[85] br[85] wl[81] vdd gnd cell_6t
Xbit_r82_c85 bl[85] br[85] wl[82] vdd gnd cell_6t
Xbit_r83_c85 bl[85] br[85] wl[83] vdd gnd cell_6t
Xbit_r84_c85 bl[85] br[85] wl[84] vdd gnd cell_6t
Xbit_r85_c85 bl[85] br[85] wl[85] vdd gnd cell_6t
Xbit_r86_c85 bl[85] br[85] wl[86] vdd gnd cell_6t
Xbit_r87_c85 bl[85] br[85] wl[87] vdd gnd cell_6t
Xbit_r88_c85 bl[85] br[85] wl[88] vdd gnd cell_6t
Xbit_r89_c85 bl[85] br[85] wl[89] vdd gnd cell_6t
Xbit_r90_c85 bl[85] br[85] wl[90] vdd gnd cell_6t
Xbit_r91_c85 bl[85] br[85] wl[91] vdd gnd cell_6t
Xbit_r92_c85 bl[85] br[85] wl[92] vdd gnd cell_6t
Xbit_r93_c85 bl[85] br[85] wl[93] vdd gnd cell_6t
Xbit_r94_c85 bl[85] br[85] wl[94] vdd gnd cell_6t
Xbit_r95_c85 bl[85] br[85] wl[95] vdd gnd cell_6t
Xbit_r96_c85 bl[85] br[85] wl[96] vdd gnd cell_6t
Xbit_r97_c85 bl[85] br[85] wl[97] vdd gnd cell_6t
Xbit_r98_c85 bl[85] br[85] wl[98] vdd gnd cell_6t
Xbit_r99_c85 bl[85] br[85] wl[99] vdd gnd cell_6t
Xbit_r100_c85 bl[85] br[85] wl[100] vdd gnd cell_6t
Xbit_r101_c85 bl[85] br[85] wl[101] vdd gnd cell_6t
Xbit_r102_c85 bl[85] br[85] wl[102] vdd gnd cell_6t
Xbit_r103_c85 bl[85] br[85] wl[103] vdd gnd cell_6t
Xbit_r104_c85 bl[85] br[85] wl[104] vdd gnd cell_6t
Xbit_r105_c85 bl[85] br[85] wl[105] vdd gnd cell_6t
Xbit_r106_c85 bl[85] br[85] wl[106] vdd gnd cell_6t
Xbit_r107_c85 bl[85] br[85] wl[107] vdd gnd cell_6t
Xbit_r108_c85 bl[85] br[85] wl[108] vdd gnd cell_6t
Xbit_r109_c85 bl[85] br[85] wl[109] vdd gnd cell_6t
Xbit_r110_c85 bl[85] br[85] wl[110] vdd gnd cell_6t
Xbit_r111_c85 bl[85] br[85] wl[111] vdd gnd cell_6t
Xbit_r112_c85 bl[85] br[85] wl[112] vdd gnd cell_6t
Xbit_r113_c85 bl[85] br[85] wl[113] vdd gnd cell_6t
Xbit_r114_c85 bl[85] br[85] wl[114] vdd gnd cell_6t
Xbit_r115_c85 bl[85] br[85] wl[115] vdd gnd cell_6t
Xbit_r116_c85 bl[85] br[85] wl[116] vdd gnd cell_6t
Xbit_r117_c85 bl[85] br[85] wl[117] vdd gnd cell_6t
Xbit_r118_c85 bl[85] br[85] wl[118] vdd gnd cell_6t
Xbit_r119_c85 bl[85] br[85] wl[119] vdd gnd cell_6t
Xbit_r120_c85 bl[85] br[85] wl[120] vdd gnd cell_6t
Xbit_r121_c85 bl[85] br[85] wl[121] vdd gnd cell_6t
Xbit_r122_c85 bl[85] br[85] wl[122] vdd gnd cell_6t
Xbit_r123_c85 bl[85] br[85] wl[123] vdd gnd cell_6t
Xbit_r124_c85 bl[85] br[85] wl[124] vdd gnd cell_6t
Xbit_r125_c85 bl[85] br[85] wl[125] vdd gnd cell_6t
Xbit_r126_c85 bl[85] br[85] wl[126] vdd gnd cell_6t
Xbit_r127_c85 bl[85] br[85] wl[127] vdd gnd cell_6t
Xbit_r128_c85 bl[85] br[85] wl[128] vdd gnd cell_6t
Xbit_r129_c85 bl[85] br[85] wl[129] vdd gnd cell_6t
Xbit_r130_c85 bl[85] br[85] wl[130] vdd gnd cell_6t
Xbit_r131_c85 bl[85] br[85] wl[131] vdd gnd cell_6t
Xbit_r132_c85 bl[85] br[85] wl[132] vdd gnd cell_6t
Xbit_r133_c85 bl[85] br[85] wl[133] vdd gnd cell_6t
Xbit_r134_c85 bl[85] br[85] wl[134] vdd gnd cell_6t
Xbit_r135_c85 bl[85] br[85] wl[135] vdd gnd cell_6t
Xbit_r136_c85 bl[85] br[85] wl[136] vdd gnd cell_6t
Xbit_r137_c85 bl[85] br[85] wl[137] vdd gnd cell_6t
Xbit_r138_c85 bl[85] br[85] wl[138] vdd gnd cell_6t
Xbit_r139_c85 bl[85] br[85] wl[139] vdd gnd cell_6t
Xbit_r140_c85 bl[85] br[85] wl[140] vdd gnd cell_6t
Xbit_r141_c85 bl[85] br[85] wl[141] vdd gnd cell_6t
Xbit_r142_c85 bl[85] br[85] wl[142] vdd gnd cell_6t
Xbit_r143_c85 bl[85] br[85] wl[143] vdd gnd cell_6t
Xbit_r144_c85 bl[85] br[85] wl[144] vdd gnd cell_6t
Xbit_r145_c85 bl[85] br[85] wl[145] vdd gnd cell_6t
Xbit_r146_c85 bl[85] br[85] wl[146] vdd gnd cell_6t
Xbit_r147_c85 bl[85] br[85] wl[147] vdd gnd cell_6t
Xbit_r148_c85 bl[85] br[85] wl[148] vdd gnd cell_6t
Xbit_r149_c85 bl[85] br[85] wl[149] vdd gnd cell_6t
Xbit_r150_c85 bl[85] br[85] wl[150] vdd gnd cell_6t
Xbit_r151_c85 bl[85] br[85] wl[151] vdd gnd cell_6t
Xbit_r152_c85 bl[85] br[85] wl[152] vdd gnd cell_6t
Xbit_r153_c85 bl[85] br[85] wl[153] vdd gnd cell_6t
Xbit_r154_c85 bl[85] br[85] wl[154] vdd gnd cell_6t
Xbit_r155_c85 bl[85] br[85] wl[155] vdd gnd cell_6t
Xbit_r156_c85 bl[85] br[85] wl[156] vdd gnd cell_6t
Xbit_r157_c85 bl[85] br[85] wl[157] vdd gnd cell_6t
Xbit_r158_c85 bl[85] br[85] wl[158] vdd gnd cell_6t
Xbit_r159_c85 bl[85] br[85] wl[159] vdd gnd cell_6t
Xbit_r160_c85 bl[85] br[85] wl[160] vdd gnd cell_6t
Xbit_r161_c85 bl[85] br[85] wl[161] vdd gnd cell_6t
Xbit_r162_c85 bl[85] br[85] wl[162] vdd gnd cell_6t
Xbit_r163_c85 bl[85] br[85] wl[163] vdd gnd cell_6t
Xbit_r164_c85 bl[85] br[85] wl[164] vdd gnd cell_6t
Xbit_r165_c85 bl[85] br[85] wl[165] vdd gnd cell_6t
Xbit_r166_c85 bl[85] br[85] wl[166] vdd gnd cell_6t
Xbit_r167_c85 bl[85] br[85] wl[167] vdd gnd cell_6t
Xbit_r168_c85 bl[85] br[85] wl[168] vdd gnd cell_6t
Xbit_r169_c85 bl[85] br[85] wl[169] vdd gnd cell_6t
Xbit_r170_c85 bl[85] br[85] wl[170] vdd gnd cell_6t
Xbit_r171_c85 bl[85] br[85] wl[171] vdd gnd cell_6t
Xbit_r172_c85 bl[85] br[85] wl[172] vdd gnd cell_6t
Xbit_r173_c85 bl[85] br[85] wl[173] vdd gnd cell_6t
Xbit_r174_c85 bl[85] br[85] wl[174] vdd gnd cell_6t
Xbit_r175_c85 bl[85] br[85] wl[175] vdd gnd cell_6t
Xbit_r176_c85 bl[85] br[85] wl[176] vdd gnd cell_6t
Xbit_r177_c85 bl[85] br[85] wl[177] vdd gnd cell_6t
Xbit_r178_c85 bl[85] br[85] wl[178] vdd gnd cell_6t
Xbit_r179_c85 bl[85] br[85] wl[179] vdd gnd cell_6t
Xbit_r180_c85 bl[85] br[85] wl[180] vdd gnd cell_6t
Xbit_r181_c85 bl[85] br[85] wl[181] vdd gnd cell_6t
Xbit_r182_c85 bl[85] br[85] wl[182] vdd gnd cell_6t
Xbit_r183_c85 bl[85] br[85] wl[183] vdd gnd cell_6t
Xbit_r184_c85 bl[85] br[85] wl[184] vdd gnd cell_6t
Xbit_r185_c85 bl[85] br[85] wl[185] vdd gnd cell_6t
Xbit_r186_c85 bl[85] br[85] wl[186] vdd gnd cell_6t
Xbit_r187_c85 bl[85] br[85] wl[187] vdd gnd cell_6t
Xbit_r188_c85 bl[85] br[85] wl[188] vdd gnd cell_6t
Xbit_r189_c85 bl[85] br[85] wl[189] vdd gnd cell_6t
Xbit_r190_c85 bl[85] br[85] wl[190] vdd gnd cell_6t
Xbit_r191_c85 bl[85] br[85] wl[191] vdd gnd cell_6t
Xbit_r192_c85 bl[85] br[85] wl[192] vdd gnd cell_6t
Xbit_r193_c85 bl[85] br[85] wl[193] vdd gnd cell_6t
Xbit_r194_c85 bl[85] br[85] wl[194] vdd gnd cell_6t
Xbit_r195_c85 bl[85] br[85] wl[195] vdd gnd cell_6t
Xbit_r196_c85 bl[85] br[85] wl[196] vdd gnd cell_6t
Xbit_r197_c85 bl[85] br[85] wl[197] vdd gnd cell_6t
Xbit_r198_c85 bl[85] br[85] wl[198] vdd gnd cell_6t
Xbit_r199_c85 bl[85] br[85] wl[199] vdd gnd cell_6t
Xbit_r200_c85 bl[85] br[85] wl[200] vdd gnd cell_6t
Xbit_r201_c85 bl[85] br[85] wl[201] vdd gnd cell_6t
Xbit_r202_c85 bl[85] br[85] wl[202] vdd gnd cell_6t
Xbit_r203_c85 bl[85] br[85] wl[203] vdd gnd cell_6t
Xbit_r204_c85 bl[85] br[85] wl[204] vdd gnd cell_6t
Xbit_r205_c85 bl[85] br[85] wl[205] vdd gnd cell_6t
Xbit_r206_c85 bl[85] br[85] wl[206] vdd gnd cell_6t
Xbit_r207_c85 bl[85] br[85] wl[207] vdd gnd cell_6t
Xbit_r208_c85 bl[85] br[85] wl[208] vdd gnd cell_6t
Xbit_r209_c85 bl[85] br[85] wl[209] vdd gnd cell_6t
Xbit_r210_c85 bl[85] br[85] wl[210] vdd gnd cell_6t
Xbit_r211_c85 bl[85] br[85] wl[211] vdd gnd cell_6t
Xbit_r212_c85 bl[85] br[85] wl[212] vdd gnd cell_6t
Xbit_r213_c85 bl[85] br[85] wl[213] vdd gnd cell_6t
Xbit_r214_c85 bl[85] br[85] wl[214] vdd gnd cell_6t
Xbit_r215_c85 bl[85] br[85] wl[215] vdd gnd cell_6t
Xbit_r216_c85 bl[85] br[85] wl[216] vdd gnd cell_6t
Xbit_r217_c85 bl[85] br[85] wl[217] vdd gnd cell_6t
Xbit_r218_c85 bl[85] br[85] wl[218] vdd gnd cell_6t
Xbit_r219_c85 bl[85] br[85] wl[219] vdd gnd cell_6t
Xbit_r220_c85 bl[85] br[85] wl[220] vdd gnd cell_6t
Xbit_r221_c85 bl[85] br[85] wl[221] vdd gnd cell_6t
Xbit_r222_c85 bl[85] br[85] wl[222] vdd gnd cell_6t
Xbit_r223_c85 bl[85] br[85] wl[223] vdd gnd cell_6t
Xbit_r224_c85 bl[85] br[85] wl[224] vdd gnd cell_6t
Xbit_r225_c85 bl[85] br[85] wl[225] vdd gnd cell_6t
Xbit_r226_c85 bl[85] br[85] wl[226] vdd gnd cell_6t
Xbit_r227_c85 bl[85] br[85] wl[227] vdd gnd cell_6t
Xbit_r228_c85 bl[85] br[85] wl[228] vdd gnd cell_6t
Xbit_r229_c85 bl[85] br[85] wl[229] vdd gnd cell_6t
Xbit_r230_c85 bl[85] br[85] wl[230] vdd gnd cell_6t
Xbit_r231_c85 bl[85] br[85] wl[231] vdd gnd cell_6t
Xbit_r232_c85 bl[85] br[85] wl[232] vdd gnd cell_6t
Xbit_r233_c85 bl[85] br[85] wl[233] vdd gnd cell_6t
Xbit_r234_c85 bl[85] br[85] wl[234] vdd gnd cell_6t
Xbit_r235_c85 bl[85] br[85] wl[235] vdd gnd cell_6t
Xbit_r236_c85 bl[85] br[85] wl[236] vdd gnd cell_6t
Xbit_r237_c85 bl[85] br[85] wl[237] vdd gnd cell_6t
Xbit_r238_c85 bl[85] br[85] wl[238] vdd gnd cell_6t
Xbit_r239_c85 bl[85] br[85] wl[239] vdd gnd cell_6t
Xbit_r240_c85 bl[85] br[85] wl[240] vdd gnd cell_6t
Xbit_r241_c85 bl[85] br[85] wl[241] vdd gnd cell_6t
Xbit_r242_c85 bl[85] br[85] wl[242] vdd gnd cell_6t
Xbit_r243_c85 bl[85] br[85] wl[243] vdd gnd cell_6t
Xbit_r244_c85 bl[85] br[85] wl[244] vdd gnd cell_6t
Xbit_r245_c85 bl[85] br[85] wl[245] vdd gnd cell_6t
Xbit_r246_c85 bl[85] br[85] wl[246] vdd gnd cell_6t
Xbit_r247_c85 bl[85] br[85] wl[247] vdd gnd cell_6t
Xbit_r248_c85 bl[85] br[85] wl[248] vdd gnd cell_6t
Xbit_r249_c85 bl[85] br[85] wl[249] vdd gnd cell_6t
Xbit_r250_c85 bl[85] br[85] wl[250] vdd gnd cell_6t
Xbit_r251_c85 bl[85] br[85] wl[251] vdd gnd cell_6t
Xbit_r252_c85 bl[85] br[85] wl[252] vdd gnd cell_6t
Xbit_r253_c85 bl[85] br[85] wl[253] vdd gnd cell_6t
Xbit_r254_c85 bl[85] br[85] wl[254] vdd gnd cell_6t
Xbit_r255_c85 bl[85] br[85] wl[255] vdd gnd cell_6t
Xbit_r0_c86 bl[86] br[86] wl[0] vdd gnd cell_6t
Xbit_r1_c86 bl[86] br[86] wl[1] vdd gnd cell_6t
Xbit_r2_c86 bl[86] br[86] wl[2] vdd gnd cell_6t
Xbit_r3_c86 bl[86] br[86] wl[3] vdd gnd cell_6t
Xbit_r4_c86 bl[86] br[86] wl[4] vdd gnd cell_6t
Xbit_r5_c86 bl[86] br[86] wl[5] vdd gnd cell_6t
Xbit_r6_c86 bl[86] br[86] wl[6] vdd gnd cell_6t
Xbit_r7_c86 bl[86] br[86] wl[7] vdd gnd cell_6t
Xbit_r8_c86 bl[86] br[86] wl[8] vdd gnd cell_6t
Xbit_r9_c86 bl[86] br[86] wl[9] vdd gnd cell_6t
Xbit_r10_c86 bl[86] br[86] wl[10] vdd gnd cell_6t
Xbit_r11_c86 bl[86] br[86] wl[11] vdd gnd cell_6t
Xbit_r12_c86 bl[86] br[86] wl[12] vdd gnd cell_6t
Xbit_r13_c86 bl[86] br[86] wl[13] vdd gnd cell_6t
Xbit_r14_c86 bl[86] br[86] wl[14] vdd gnd cell_6t
Xbit_r15_c86 bl[86] br[86] wl[15] vdd gnd cell_6t
Xbit_r16_c86 bl[86] br[86] wl[16] vdd gnd cell_6t
Xbit_r17_c86 bl[86] br[86] wl[17] vdd gnd cell_6t
Xbit_r18_c86 bl[86] br[86] wl[18] vdd gnd cell_6t
Xbit_r19_c86 bl[86] br[86] wl[19] vdd gnd cell_6t
Xbit_r20_c86 bl[86] br[86] wl[20] vdd gnd cell_6t
Xbit_r21_c86 bl[86] br[86] wl[21] vdd gnd cell_6t
Xbit_r22_c86 bl[86] br[86] wl[22] vdd gnd cell_6t
Xbit_r23_c86 bl[86] br[86] wl[23] vdd gnd cell_6t
Xbit_r24_c86 bl[86] br[86] wl[24] vdd gnd cell_6t
Xbit_r25_c86 bl[86] br[86] wl[25] vdd gnd cell_6t
Xbit_r26_c86 bl[86] br[86] wl[26] vdd gnd cell_6t
Xbit_r27_c86 bl[86] br[86] wl[27] vdd gnd cell_6t
Xbit_r28_c86 bl[86] br[86] wl[28] vdd gnd cell_6t
Xbit_r29_c86 bl[86] br[86] wl[29] vdd gnd cell_6t
Xbit_r30_c86 bl[86] br[86] wl[30] vdd gnd cell_6t
Xbit_r31_c86 bl[86] br[86] wl[31] vdd gnd cell_6t
Xbit_r32_c86 bl[86] br[86] wl[32] vdd gnd cell_6t
Xbit_r33_c86 bl[86] br[86] wl[33] vdd gnd cell_6t
Xbit_r34_c86 bl[86] br[86] wl[34] vdd gnd cell_6t
Xbit_r35_c86 bl[86] br[86] wl[35] vdd gnd cell_6t
Xbit_r36_c86 bl[86] br[86] wl[36] vdd gnd cell_6t
Xbit_r37_c86 bl[86] br[86] wl[37] vdd gnd cell_6t
Xbit_r38_c86 bl[86] br[86] wl[38] vdd gnd cell_6t
Xbit_r39_c86 bl[86] br[86] wl[39] vdd gnd cell_6t
Xbit_r40_c86 bl[86] br[86] wl[40] vdd gnd cell_6t
Xbit_r41_c86 bl[86] br[86] wl[41] vdd gnd cell_6t
Xbit_r42_c86 bl[86] br[86] wl[42] vdd gnd cell_6t
Xbit_r43_c86 bl[86] br[86] wl[43] vdd gnd cell_6t
Xbit_r44_c86 bl[86] br[86] wl[44] vdd gnd cell_6t
Xbit_r45_c86 bl[86] br[86] wl[45] vdd gnd cell_6t
Xbit_r46_c86 bl[86] br[86] wl[46] vdd gnd cell_6t
Xbit_r47_c86 bl[86] br[86] wl[47] vdd gnd cell_6t
Xbit_r48_c86 bl[86] br[86] wl[48] vdd gnd cell_6t
Xbit_r49_c86 bl[86] br[86] wl[49] vdd gnd cell_6t
Xbit_r50_c86 bl[86] br[86] wl[50] vdd gnd cell_6t
Xbit_r51_c86 bl[86] br[86] wl[51] vdd gnd cell_6t
Xbit_r52_c86 bl[86] br[86] wl[52] vdd gnd cell_6t
Xbit_r53_c86 bl[86] br[86] wl[53] vdd gnd cell_6t
Xbit_r54_c86 bl[86] br[86] wl[54] vdd gnd cell_6t
Xbit_r55_c86 bl[86] br[86] wl[55] vdd gnd cell_6t
Xbit_r56_c86 bl[86] br[86] wl[56] vdd gnd cell_6t
Xbit_r57_c86 bl[86] br[86] wl[57] vdd gnd cell_6t
Xbit_r58_c86 bl[86] br[86] wl[58] vdd gnd cell_6t
Xbit_r59_c86 bl[86] br[86] wl[59] vdd gnd cell_6t
Xbit_r60_c86 bl[86] br[86] wl[60] vdd gnd cell_6t
Xbit_r61_c86 bl[86] br[86] wl[61] vdd gnd cell_6t
Xbit_r62_c86 bl[86] br[86] wl[62] vdd gnd cell_6t
Xbit_r63_c86 bl[86] br[86] wl[63] vdd gnd cell_6t
Xbit_r64_c86 bl[86] br[86] wl[64] vdd gnd cell_6t
Xbit_r65_c86 bl[86] br[86] wl[65] vdd gnd cell_6t
Xbit_r66_c86 bl[86] br[86] wl[66] vdd gnd cell_6t
Xbit_r67_c86 bl[86] br[86] wl[67] vdd gnd cell_6t
Xbit_r68_c86 bl[86] br[86] wl[68] vdd gnd cell_6t
Xbit_r69_c86 bl[86] br[86] wl[69] vdd gnd cell_6t
Xbit_r70_c86 bl[86] br[86] wl[70] vdd gnd cell_6t
Xbit_r71_c86 bl[86] br[86] wl[71] vdd gnd cell_6t
Xbit_r72_c86 bl[86] br[86] wl[72] vdd gnd cell_6t
Xbit_r73_c86 bl[86] br[86] wl[73] vdd gnd cell_6t
Xbit_r74_c86 bl[86] br[86] wl[74] vdd gnd cell_6t
Xbit_r75_c86 bl[86] br[86] wl[75] vdd gnd cell_6t
Xbit_r76_c86 bl[86] br[86] wl[76] vdd gnd cell_6t
Xbit_r77_c86 bl[86] br[86] wl[77] vdd gnd cell_6t
Xbit_r78_c86 bl[86] br[86] wl[78] vdd gnd cell_6t
Xbit_r79_c86 bl[86] br[86] wl[79] vdd gnd cell_6t
Xbit_r80_c86 bl[86] br[86] wl[80] vdd gnd cell_6t
Xbit_r81_c86 bl[86] br[86] wl[81] vdd gnd cell_6t
Xbit_r82_c86 bl[86] br[86] wl[82] vdd gnd cell_6t
Xbit_r83_c86 bl[86] br[86] wl[83] vdd gnd cell_6t
Xbit_r84_c86 bl[86] br[86] wl[84] vdd gnd cell_6t
Xbit_r85_c86 bl[86] br[86] wl[85] vdd gnd cell_6t
Xbit_r86_c86 bl[86] br[86] wl[86] vdd gnd cell_6t
Xbit_r87_c86 bl[86] br[86] wl[87] vdd gnd cell_6t
Xbit_r88_c86 bl[86] br[86] wl[88] vdd gnd cell_6t
Xbit_r89_c86 bl[86] br[86] wl[89] vdd gnd cell_6t
Xbit_r90_c86 bl[86] br[86] wl[90] vdd gnd cell_6t
Xbit_r91_c86 bl[86] br[86] wl[91] vdd gnd cell_6t
Xbit_r92_c86 bl[86] br[86] wl[92] vdd gnd cell_6t
Xbit_r93_c86 bl[86] br[86] wl[93] vdd gnd cell_6t
Xbit_r94_c86 bl[86] br[86] wl[94] vdd gnd cell_6t
Xbit_r95_c86 bl[86] br[86] wl[95] vdd gnd cell_6t
Xbit_r96_c86 bl[86] br[86] wl[96] vdd gnd cell_6t
Xbit_r97_c86 bl[86] br[86] wl[97] vdd gnd cell_6t
Xbit_r98_c86 bl[86] br[86] wl[98] vdd gnd cell_6t
Xbit_r99_c86 bl[86] br[86] wl[99] vdd gnd cell_6t
Xbit_r100_c86 bl[86] br[86] wl[100] vdd gnd cell_6t
Xbit_r101_c86 bl[86] br[86] wl[101] vdd gnd cell_6t
Xbit_r102_c86 bl[86] br[86] wl[102] vdd gnd cell_6t
Xbit_r103_c86 bl[86] br[86] wl[103] vdd gnd cell_6t
Xbit_r104_c86 bl[86] br[86] wl[104] vdd gnd cell_6t
Xbit_r105_c86 bl[86] br[86] wl[105] vdd gnd cell_6t
Xbit_r106_c86 bl[86] br[86] wl[106] vdd gnd cell_6t
Xbit_r107_c86 bl[86] br[86] wl[107] vdd gnd cell_6t
Xbit_r108_c86 bl[86] br[86] wl[108] vdd gnd cell_6t
Xbit_r109_c86 bl[86] br[86] wl[109] vdd gnd cell_6t
Xbit_r110_c86 bl[86] br[86] wl[110] vdd gnd cell_6t
Xbit_r111_c86 bl[86] br[86] wl[111] vdd gnd cell_6t
Xbit_r112_c86 bl[86] br[86] wl[112] vdd gnd cell_6t
Xbit_r113_c86 bl[86] br[86] wl[113] vdd gnd cell_6t
Xbit_r114_c86 bl[86] br[86] wl[114] vdd gnd cell_6t
Xbit_r115_c86 bl[86] br[86] wl[115] vdd gnd cell_6t
Xbit_r116_c86 bl[86] br[86] wl[116] vdd gnd cell_6t
Xbit_r117_c86 bl[86] br[86] wl[117] vdd gnd cell_6t
Xbit_r118_c86 bl[86] br[86] wl[118] vdd gnd cell_6t
Xbit_r119_c86 bl[86] br[86] wl[119] vdd gnd cell_6t
Xbit_r120_c86 bl[86] br[86] wl[120] vdd gnd cell_6t
Xbit_r121_c86 bl[86] br[86] wl[121] vdd gnd cell_6t
Xbit_r122_c86 bl[86] br[86] wl[122] vdd gnd cell_6t
Xbit_r123_c86 bl[86] br[86] wl[123] vdd gnd cell_6t
Xbit_r124_c86 bl[86] br[86] wl[124] vdd gnd cell_6t
Xbit_r125_c86 bl[86] br[86] wl[125] vdd gnd cell_6t
Xbit_r126_c86 bl[86] br[86] wl[126] vdd gnd cell_6t
Xbit_r127_c86 bl[86] br[86] wl[127] vdd gnd cell_6t
Xbit_r128_c86 bl[86] br[86] wl[128] vdd gnd cell_6t
Xbit_r129_c86 bl[86] br[86] wl[129] vdd gnd cell_6t
Xbit_r130_c86 bl[86] br[86] wl[130] vdd gnd cell_6t
Xbit_r131_c86 bl[86] br[86] wl[131] vdd gnd cell_6t
Xbit_r132_c86 bl[86] br[86] wl[132] vdd gnd cell_6t
Xbit_r133_c86 bl[86] br[86] wl[133] vdd gnd cell_6t
Xbit_r134_c86 bl[86] br[86] wl[134] vdd gnd cell_6t
Xbit_r135_c86 bl[86] br[86] wl[135] vdd gnd cell_6t
Xbit_r136_c86 bl[86] br[86] wl[136] vdd gnd cell_6t
Xbit_r137_c86 bl[86] br[86] wl[137] vdd gnd cell_6t
Xbit_r138_c86 bl[86] br[86] wl[138] vdd gnd cell_6t
Xbit_r139_c86 bl[86] br[86] wl[139] vdd gnd cell_6t
Xbit_r140_c86 bl[86] br[86] wl[140] vdd gnd cell_6t
Xbit_r141_c86 bl[86] br[86] wl[141] vdd gnd cell_6t
Xbit_r142_c86 bl[86] br[86] wl[142] vdd gnd cell_6t
Xbit_r143_c86 bl[86] br[86] wl[143] vdd gnd cell_6t
Xbit_r144_c86 bl[86] br[86] wl[144] vdd gnd cell_6t
Xbit_r145_c86 bl[86] br[86] wl[145] vdd gnd cell_6t
Xbit_r146_c86 bl[86] br[86] wl[146] vdd gnd cell_6t
Xbit_r147_c86 bl[86] br[86] wl[147] vdd gnd cell_6t
Xbit_r148_c86 bl[86] br[86] wl[148] vdd gnd cell_6t
Xbit_r149_c86 bl[86] br[86] wl[149] vdd gnd cell_6t
Xbit_r150_c86 bl[86] br[86] wl[150] vdd gnd cell_6t
Xbit_r151_c86 bl[86] br[86] wl[151] vdd gnd cell_6t
Xbit_r152_c86 bl[86] br[86] wl[152] vdd gnd cell_6t
Xbit_r153_c86 bl[86] br[86] wl[153] vdd gnd cell_6t
Xbit_r154_c86 bl[86] br[86] wl[154] vdd gnd cell_6t
Xbit_r155_c86 bl[86] br[86] wl[155] vdd gnd cell_6t
Xbit_r156_c86 bl[86] br[86] wl[156] vdd gnd cell_6t
Xbit_r157_c86 bl[86] br[86] wl[157] vdd gnd cell_6t
Xbit_r158_c86 bl[86] br[86] wl[158] vdd gnd cell_6t
Xbit_r159_c86 bl[86] br[86] wl[159] vdd gnd cell_6t
Xbit_r160_c86 bl[86] br[86] wl[160] vdd gnd cell_6t
Xbit_r161_c86 bl[86] br[86] wl[161] vdd gnd cell_6t
Xbit_r162_c86 bl[86] br[86] wl[162] vdd gnd cell_6t
Xbit_r163_c86 bl[86] br[86] wl[163] vdd gnd cell_6t
Xbit_r164_c86 bl[86] br[86] wl[164] vdd gnd cell_6t
Xbit_r165_c86 bl[86] br[86] wl[165] vdd gnd cell_6t
Xbit_r166_c86 bl[86] br[86] wl[166] vdd gnd cell_6t
Xbit_r167_c86 bl[86] br[86] wl[167] vdd gnd cell_6t
Xbit_r168_c86 bl[86] br[86] wl[168] vdd gnd cell_6t
Xbit_r169_c86 bl[86] br[86] wl[169] vdd gnd cell_6t
Xbit_r170_c86 bl[86] br[86] wl[170] vdd gnd cell_6t
Xbit_r171_c86 bl[86] br[86] wl[171] vdd gnd cell_6t
Xbit_r172_c86 bl[86] br[86] wl[172] vdd gnd cell_6t
Xbit_r173_c86 bl[86] br[86] wl[173] vdd gnd cell_6t
Xbit_r174_c86 bl[86] br[86] wl[174] vdd gnd cell_6t
Xbit_r175_c86 bl[86] br[86] wl[175] vdd gnd cell_6t
Xbit_r176_c86 bl[86] br[86] wl[176] vdd gnd cell_6t
Xbit_r177_c86 bl[86] br[86] wl[177] vdd gnd cell_6t
Xbit_r178_c86 bl[86] br[86] wl[178] vdd gnd cell_6t
Xbit_r179_c86 bl[86] br[86] wl[179] vdd gnd cell_6t
Xbit_r180_c86 bl[86] br[86] wl[180] vdd gnd cell_6t
Xbit_r181_c86 bl[86] br[86] wl[181] vdd gnd cell_6t
Xbit_r182_c86 bl[86] br[86] wl[182] vdd gnd cell_6t
Xbit_r183_c86 bl[86] br[86] wl[183] vdd gnd cell_6t
Xbit_r184_c86 bl[86] br[86] wl[184] vdd gnd cell_6t
Xbit_r185_c86 bl[86] br[86] wl[185] vdd gnd cell_6t
Xbit_r186_c86 bl[86] br[86] wl[186] vdd gnd cell_6t
Xbit_r187_c86 bl[86] br[86] wl[187] vdd gnd cell_6t
Xbit_r188_c86 bl[86] br[86] wl[188] vdd gnd cell_6t
Xbit_r189_c86 bl[86] br[86] wl[189] vdd gnd cell_6t
Xbit_r190_c86 bl[86] br[86] wl[190] vdd gnd cell_6t
Xbit_r191_c86 bl[86] br[86] wl[191] vdd gnd cell_6t
Xbit_r192_c86 bl[86] br[86] wl[192] vdd gnd cell_6t
Xbit_r193_c86 bl[86] br[86] wl[193] vdd gnd cell_6t
Xbit_r194_c86 bl[86] br[86] wl[194] vdd gnd cell_6t
Xbit_r195_c86 bl[86] br[86] wl[195] vdd gnd cell_6t
Xbit_r196_c86 bl[86] br[86] wl[196] vdd gnd cell_6t
Xbit_r197_c86 bl[86] br[86] wl[197] vdd gnd cell_6t
Xbit_r198_c86 bl[86] br[86] wl[198] vdd gnd cell_6t
Xbit_r199_c86 bl[86] br[86] wl[199] vdd gnd cell_6t
Xbit_r200_c86 bl[86] br[86] wl[200] vdd gnd cell_6t
Xbit_r201_c86 bl[86] br[86] wl[201] vdd gnd cell_6t
Xbit_r202_c86 bl[86] br[86] wl[202] vdd gnd cell_6t
Xbit_r203_c86 bl[86] br[86] wl[203] vdd gnd cell_6t
Xbit_r204_c86 bl[86] br[86] wl[204] vdd gnd cell_6t
Xbit_r205_c86 bl[86] br[86] wl[205] vdd gnd cell_6t
Xbit_r206_c86 bl[86] br[86] wl[206] vdd gnd cell_6t
Xbit_r207_c86 bl[86] br[86] wl[207] vdd gnd cell_6t
Xbit_r208_c86 bl[86] br[86] wl[208] vdd gnd cell_6t
Xbit_r209_c86 bl[86] br[86] wl[209] vdd gnd cell_6t
Xbit_r210_c86 bl[86] br[86] wl[210] vdd gnd cell_6t
Xbit_r211_c86 bl[86] br[86] wl[211] vdd gnd cell_6t
Xbit_r212_c86 bl[86] br[86] wl[212] vdd gnd cell_6t
Xbit_r213_c86 bl[86] br[86] wl[213] vdd gnd cell_6t
Xbit_r214_c86 bl[86] br[86] wl[214] vdd gnd cell_6t
Xbit_r215_c86 bl[86] br[86] wl[215] vdd gnd cell_6t
Xbit_r216_c86 bl[86] br[86] wl[216] vdd gnd cell_6t
Xbit_r217_c86 bl[86] br[86] wl[217] vdd gnd cell_6t
Xbit_r218_c86 bl[86] br[86] wl[218] vdd gnd cell_6t
Xbit_r219_c86 bl[86] br[86] wl[219] vdd gnd cell_6t
Xbit_r220_c86 bl[86] br[86] wl[220] vdd gnd cell_6t
Xbit_r221_c86 bl[86] br[86] wl[221] vdd gnd cell_6t
Xbit_r222_c86 bl[86] br[86] wl[222] vdd gnd cell_6t
Xbit_r223_c86 bl[86] br[86] wl[223] vdd gnd cell_6t
Xbit_r224_c86 bl[86] br[86] wl[224] vdd gnd cell_6t
Xbit_r225_c86 bl[86] br[86] wl[225] vdd gnd cell_6t
Xbit_r226_c86 bl[86] br[86] wl[226] vdd gnd cell_6t
Xbit_r227_c86 bl[86] br[86] wl[227] vdd gnd cell_6t
Xbit_r228_c86 bl[86] br[86] wl[228] vdd gnd cell_6t
Xbit_r229_c86 bl[86] br[86] wl[229] vdd gnd cell_6t
Xbit_r230_c86 bl[86] br[86] wl[230] vdd gnd cell_6t
Xbit_r231_c86 bl[86] br[86] wl[231] vdd gnd cell_6t
Xbit_r232_c86 bl[86] br[86] wl[232] vdd gnd cell_6t
Xbit_r233_c86 bl[86] br[86] wl[233] vdd gnd cell_6t
Xbit_r234_c86 bl[86] br[86] wl[234] vdd gnd cell_6t
Xbit_r235_c86 bl[86] br[86] wl[235] vdd gnd cell_6t
Xbit_r236_c86 bl[86] br[86] wl[236] vdd gnd cell_6t
Xbit_r237_c86 bl[86] br[86] wl[237] vdd gnd cell_6t
Xbit_r238_c86 bl[86] br[86] wl[238] vdd gnd cell_6t
Xbit_r239_c86 bl[86] br[86] wl[239] vdd gnd cell_6t
Xbit_r240_c86 bl[86] br[86] wl[240] vdd gnd cell_6t
Xbit_r241_c86 bl[86] br[86] wl[241] vdd gnd cell_6t
Xbit_r242_c86 bl[86] br[86] wl[242] vdd gnd cell_6t
Xbit_r243_c86 bl[86] br[86] wl[243] vdd gnd cell_6t
Xbit_r244_c86 bl[86] br[86] wl[244] vdd gnd cell_6t
Xbit_r245_c86 bl[86] br[86] wl[245] vdd gnd cell_6t
Xbit_r246_c86 bl[86] br[86] wl[246] vdd gnd cell_6t
Xbit_r247_c86 bl[86] br[86] wl[247] vdd gnd cell_6t
Xbit_r248_c86 bl[86] br[86] wl[248] vdd gnd cell_6t
Xbit_r249_c86 bl[86] br[86] wl[249] vdd gnd cell_6t
Xbit_r250_c86 bl[86] br[86] wl[250] vdd gnd cell_6t
Xbit_r251_c86 bl[86] br[86] wl[251] vdd gnd cell_6t
Xbit_r252_c86 bl[86] br[86] wl[252] vdd gnd cell_6t
Xbit_r253_c86 bl[86] br[86] wl[253] vdd gnd cell_6t
Xbit_r254_c86 bl[86] br[86] wl[254] vdd gnd cell_6t
Xbit_r255_c86 bl[86] br[86] wl[255] vdd gnd cell_6t
Xbit_r0_c87 bl[87] br[87] wl[0] vdd gnd cell_6t
Xbit_r1_c87 bl[87] br[87] wl[1] vdd gnd cell_6t
Xbit_r2_c87 bl[87] br[87] wl[2] vdd gnd cell_6t
Xbit_r3_c87 bl[87] br[87] wl[3] vdd gnd cell_6t
Xbit_r4_c87 bl[87] br[87] wl[4] vdd gnd cell_6t
Xbit_r5_c87 bl[87] br[87] wl[5] vdd gnd cell_6t
Xbit_r6_c87 bl[87] br[87] wl[6] vdd gnd cell_6t
Xbit_r7_c87 bl[87] br[87] wl[7] vdd gnd cell_6t
Xbit_r8_c87 bl[87] br[87] wl[8] vdd gnd cell_6t
Xbit_r9_c87 bl[87] br[87] wl[9] vdd gnd cell_6t
Xbit_r10_c87 bl[87] br[87] wl[10] vdd gnd cell_6t
Xbit_r11_c87 bl[87] br[87] wl[11] vdd gnd cell_6t
Xbit_r12_c87 bl[87] br[87] wl[12] vdd gnd cell_6t
Xbit_r13_c87 bl[87] br[87] wl[13] vdd gnd cell_6t
Xbit_r14_c87 bl[87] br[87] wl[14] vdd gnd cell_6t
Xbit_r15_c87 bl[87] br[87] wl[15] vdd gnd cell_6t
Xbit_r16_c87 bl[87] br[87] wl[16] vdd gnd cell_6t
Xbit_r17_c87 bl[87] br[87] wl[17] vdd gnd cell_6t
Xbit_r18_c87 bl[87] br[87] wl[18] vdd gnd cell_6t
Xbit_r19_c87 bl[87] br[87] wl[19] vdd gnd cell_6t
Xbit_r20_c87 bl[87] br[87] wl[20] vdd gnd cell_6t
Xbit_r21_c87 bl[87] br[87] wl[21] vdd gnd cell_6t
Xbit_r22_c87 bl[87] br[87] wl[22] vdd gnd cell_6t
Xbit_r23_c87 bl[87] br[87] wl[23] vdd gnd cell_6t
Xbit_r24_c87 bl[87] br[87] wl[24] vdd gnd cell_6t
Xbit_r25_c87 bl[87] br[87] wl[25] vdd gnd cell_6t
Xbit_r26_c87 bl[87] br[87] wl[26] vdd gnd cell_6t
Xbit_r27_c87 bl[87] br[87] wl[27] vdd gnd cell_6t
Xbit_r28_c87 bl[87] br[87] wl[28] vdd gnd cell_6t
Xbit_r29_c87 bl[87] br[87] wl[29] vdd gnd cell_6t
Xbit_r30_c87 bl[87] br[87] wl[30] vdd gnd cell_6t
Xbit_r31_c87 bl[87] br[87] wl[31] vdd gnd cell_6t
Xbit_r32_c87 bl[87] br[87] wl[32] vdd gnd cell_6t
Xbit_r33_c87 bl[87] br[87] wl[33] vdd gnd cell_6t
Xbit_r34_c87 bl[87] br[87] wl[34] vdd gnd cell_6t
Xbit_r35_c87 bl[87] br[87] wl[35] vdd gnd cell_6t
Xbit_r36_c87 bl[87] br[87] wl[36] vdd gnd cell_6t
Xbit_r37_c87 bl[87] br[87] wl[37] vdd gnd cell_6t
Xbit_r38_c87 bl[87] br[87] wl[38] vdd gnd cell_6t
Xbit_r39_c87 bl[87] br[87] wl[39] vdd gnd cell_6t
Xbit_r40_c87 bl[87] br[87] wl[40] vdd gnd cell_6t
Xbit_r41_c87 bl[87] br[87] wl[41] vdd gnd cell_6t
Xbit_r42_c87 bl[87] br[87] wl[42] vdd gnd cell_6t
Xbit_r43_c87 bl[87] br[87] wl[43] vdd gnd cell_6t
Xbit_r44_c87 bl[87] br[87] wl[44] vdd gnd cell_6t
Xbit_r45_c87 bl[87] br[87] wl[45] vdd gnd cell_6t
Xbit_r46_c87 bl[87] br[87] wl[46] vdd gnd cell_6t
Xbit_r47_c87 bl[87] br[87] wl[47] vdd gnd cell_6t
Xbit_r48_c87 bl[87] br[87] wl[48] vdd gnd cell_6t
Xbit_r49_c87 bl[87] br[87] wl[49] vdd gnd cell_6t
Xbit_r50_c87 bl[87] br[87] wl[50] vdd gnd cell_6t
Xbit_r51_c87 bl[87] br[87] wl[51] vdd gnd cell_6t
Xbit_r52_c87 bl[87] br[87] wl[52] vdd gnd cell_6t
Xbit_r53_c87 bl[87] br[87] wl[53] vdd gnd cell_6t
Xbit_r54_c87 bl[87] br[87] wl[54] vdd gnd cell_6t
Xbit_r55_c87 bl[87] br[87] wl[55] vdd gnd cell_6t
Xbit_r56_c87 bl[87] br[87] wl[56] vdd gnd cell_6t
Xbit_r57_c87 bl[87] br[87] wl[57] vdd gnd cell_6t
Xbit_r58_c87 bl[87] br[87] wl[58] vdd gnd cell_6t
Xbit_r59_c87 bl[87] br[87] wl[59] vdd gnd cell_6t
Xbit_r60_c87 bl[87] br[87] wl[60] vdd gnd cell_6t
Xbit_r61_c87 bl[87] br[87] wl[61] vdd gnd cell_6t
Xbit_r62_c87 bl[87] br[87] wl[62] vdd gnd cell_6t
Xbit_r63_c87 bl[87] br[87] wl[63] vdd gnd cell_6t
Xbit_r64_c87 bl[87] br[87] wl[64] vdd gnd cell_6t
Xbit_r65_c87 bl[87] br[87] wl[65] vdd gnd cell_6t
Xbit_r66_c87 bl[87] br[87] wl[66] vdd gnd cell_6t
Xbit_r67_c87 bl[87] br[87] wl[67] vdd gnd cell_6t
Xbit_r68_c87 bl[87] br[87] wl[68] vdd gnd cell_6t
Xbit_r69_c87 bl[87] br[87] wl[69] vdd gnd cell_6t
Xbit_r70_c87 bl[87] br[87] wl[70] vdd gnd cell_6t
Xbit_r71_c87 bl[87] br[87] wl[71] vdd gnd cell_6t
Xbit_r72_c87 bl[87] br[87] wl[72] vdd gnd cell_6t
Xbit_r73_c87 bl[87] br[87] wl[73] vdd gnd cell_6t
Xbit_r74_c87 bl[87] br[87] wl[74] vdd gnd cell_6t
Xbit_r75_c87 bl[87] br[87] wl[75] vdd gnd cell_6t
Xbit_r76_c87 bl[87] br[87] wl[76] vdd gnd cell_6t
Xbit_r77_c87 bl[87] br[87] wl[77] vdd gnd cell_6t
Xbit_r78_c87 bl[87] br[87] wl[78] vdd gnd cell_6t
Xbit_r79_c87 bl[87] br[87] wl[79] vdd gnd cell_6t
Xbit_r80_c87 bl[87] br[87] wl[80] vdd gnd cell_6t
Xbit_r81_c87 bl[87] br[87] wl[81] vdd gnd cell_6t
Xbit_r82_c87 bl[87] br[87] wl[82] vdd gnd cell_6t
Xbit_r83_c87 bl[87] br[87] wl[83] vdd gnd cell_6t
Xbit_r84_c87 bl[87] br[87] wl[84] vdd gnd cell_6t
Xbit_r85_c87 bl[87] br[87] wl[85] vdd gnd cell_6t
Xbit_r86_c87 bl[87] br[87] wl[86] vdd gnd cell_6t
Xbit_r87_c87 bl[87] br[87] wl[87] vdd gnd cell_6t
Xbit_r88_c87 bl[87] br[87] wl[88] vdd gnd cell_6t
Xbit_r89_c87 bl[87] br[87] wl[89] vdd gnd cell_6t
Xbit_r90_c87 bl[87] br[87] wl[90] vdd gnd cell_6t
Xbit_r91_c87 bl[87] br[87] wl[91] vdd gnd cell_6t
Xbit_r92_c87 bl[87] br[87] wl[92] vdd gnd cell_6t
Xbit_r93_c87 bl[87] br[87] wl[93] vdd gnd cell_6t
Xbit_r94_c87 bl[87] br[87] wl[94] vdd gnd cell_6t
Xbit_r95_c87 bl[87] br[87] wl[95] vdd gnd cell_6t
Xbit_r96_c87 bl[87] br[87] wl[96] vdd gnd cell_6t
Xbit_r97_c87 bl[87] br[87] wl[97] vdd gnd cell_6t
Xbit_r98_c87 bl[87] br[87] wl[98] vdd gnd cell_6t
Xbit_r99_c87 bl[87] br[87] wl[99] vdd gnd cell_6t
Xbit_r100_c87 bl[87] br[87] wl[100] vdd gnd cell_6t
Xbit_r101_c87 bl[87] br[87] wl[101] vdd gnd cell_6t
Xbit_r102_c87 bl[87] br[87] wl[102] vdd gnd cell_6t
Xbit_r103_c87 bl[87] br[87] wl[103] vdd gnd cell_6t
Xbit_r104_c87 bl[87] br[87] wl[104] vdd gnd cell_6t
Xbit_r105_c87 bl[87] br[87] wl[105] vdd gnd cell_6t
Xbit_r106_c87 bl[87] br[87] wl[106] vdd gnd cell_6t
Xbit_r107_c87 bl[87] br[87] wl[107] vdd gnd cell_6t
Xbit_r108_c87 bl[87] br[87] wl[108] vdd gnd cell_6t
Xbit_r109_c87 bl[87] br[87] wl[109] vdd gnd cell_6t
Xbit_r110_c87 bl[87] br[87] wl[110] vdd gnd cell_6t
Xbit_r111_c87 bl[87] br[87] wl[111] vdd gnd cell_6t
Xbit_r112_c87 bl[87] br[87] wl[112] vdd gnd cell_6t
Xbit_r113_c87 bl[87] br[87] wl[113] vdd gnd cell_6t
Xbit_r114_c87 bl[87] br[87] wl[114] vdd gnd cell_6t
Xbit_r115_c87 bl[87] br[87] wl[115] vdd gnd cell_6t
Xbit_r116_c87 bl[87] br[87] wl[116] vdd gnd cell_6t
Xbit_r117_c87 bl[87] br[87] wl[117] vdd gnd cell_6t
Xbit_r118_c87 bl[87] br[87] wl[118] vdd gnd cell_6t
Xbit_r119_c87 bl[87] br[87] wl[119] vdd gnd cell_6t
Xbit_r120_c87 bl[87] br[87] wl[120] vdd gnd cell_6t
Xbit_r121_c87 bl[87] br[87] wl[121] vdd gnd cell_6t
Xbit_r122_c87 bl[87] br[87] wl[122] vdd gnd cell_6t
Xbit_r123_c87 bl[87] br[87] wl[123] vdd gnd cell_6t
Xbit_r124_c87 bl[87] br[87] wl[124] vdd gnd cell_6t
Xbit_r125_c87 bl[87] br[87] wl[125] vdd gnd cell_6t
Xbit_r126_c87 bl[87] br[87] wl[126] vdd gnd cell_6t
Xbit_r127_c87 bl[87] br[87] wl[127] vdd gnd cell_6t
Xbit_r128_c87 bl[87] br[87] wl[128] vdd gnd cell_6t
Xbit_r129_c87 bl[87] br[87] wl[129] vdd gnd cell_6t
Xbit_r130_c87 bl[87] br[87] wl[130] vdd gnd cell_6t
Xbit_r131_c87 bl[87] br[87] wl[131] vdd gnd cell_6t
Xbit_r132_c87 bl[87] br[87] wl[132] vdd gnd cell_6t
Xbit_r133_c87 bl[87] br[87] wl[133] vdd gnd cell_6t
Xbit_r134_c87 bl[87] br[87] wl[134] vdd gnd cell_6t
Xbit_r135_c87 bl[87] br[87] wl[135] vdd gnd cell_6t
Xbit_r136_c87 bl[87] br[87] wl[136] vdd gnd cell_6t
Xbit_r137_c87 bl[87] br[87] wl[137] vdd gnd cell_6t
Xbit_r138_c87 bl[87] br[87] wl[138] vdd gnd cell_6t
Xbit_r139_c87 bl[87] br[87] wl[139] vdd gnd cell_6t
Xbit_r140_c87 bl[87] br[87] wl[140] vdd gnd cell_6t
Xbit_r141_c87 bl[87] br[87] wl[141] vdd gnd cell_6t
Xbit_r142_c87 bl[87] br[87] wl[142] vdd gnd cell_6t
Xbit_r143_c87 bl[87] br[87] wl[143] vdd gnd cell_6t
Xbit_r144_c87 bl[87] br[87] wl[144] vdd gnd cell_6t
Xbit_r145_c87 bl[87] br[87] wl[145] vdd gnd cell_6t
Xbit_r146_c87 bl[87] br[87] wl[146] vdd gnd cell_6t
Xbit_r147_c87 bl[87] br[87] wl[147] vdd gnd cell_6t
Xbit_r148_c87 bl[87] br[87] wl[148] vdd gnd cell_6t
Xbit_r149_c87 bl[87] br[87] wl[149] vdd gnd cell_6t
Xbit_r150_c87 bl[87] br[87] wl[150] vdd gnd cell_6t
Xbit_r151_c87 bl[87] br[87] wl[151] vdd gnd cell_6t
Xbit_r152_c87 bl[87] br[87] wl[152] vdd gnd cell_6t
Xbit_r153_c87 bl[87] br[87] wl[153] vdd gnd cell_6t
Xbit_r154_c87 bl[87] br[87] wl[154] vdd gnd cell_6t
Xbit_r155_c87 bl[87] br[87] wl[155] vdd gnd cell_6t
Xbit_r156_c87 bl[87] br[87] wl[156] vdd gnd cell_6t
Xbit_r157_c87 bl[87] br[87] wl[157] vdd gnd cell_6t
Xbit_r158_c87 bl[87] br[87] wl[158] vdd gnd cell_6t
Xbit_r159_c87 bl[87] br[87] wl[159] vdd gnd cell_6t
Xbit_r160_c87 bl[87] br[87] wl[160] vdd gnd cell_6t
Xbit_r161_c87 bl[87] br[87] wl[161] vdd gnd cell_6t
Xbit_r162_c87 bl[87] br[87] wl[162] vdd gnd cell_6t
Xbit_r163_c87 bl[87] br[87] wl[163] vdd gnd cell_6t
Xbit_r164_c87 bl[87] br[87] wl[164] vdd gnd cell_6t
Xbit_r165_c87 bl[87] br[87] wl[165] vdd gnd cell_6t
Xbit_r166_c87 bl[87] br[87] wl[166] vdd gnd cell_6t
Xbit_r167_c87 bl[87] br[87] wl[167] vdd gnd cell_6t
Xbit_r168_c87 bl[87] br[87] wl[168] vdd gnd cell_6t
Xbit_r169_c87 bl[87] br[87] wl[169] vdd gnd cell_6t
Xbit_r170_c87 bl[87] br[87] wl[170] vdd gnd cell_6t
Xbit_r171_c87 bl[87] br[87] wl[171] vdd gnd cell_6t
Xbit_r172_c87 bl[87] br[87] wl[172] vdd gnd cell_6t
Xbit_r173_c87 bl[87] br[87] wl[173] vdd gnd cell_6t
Xbit_r174_c87 bl[87] br[87] wl[174] vdd gnd cell_6t
Xbit_r175_c87 bl[87] br[87] wl[175] vdd gnd cell_6t
Xbit_r176_c87 bl[87] br[87] wl[176] vdd gnd cell_6t
Xbit_r177_c87 bl[87] br[87] wl[177] vdd gnd cell_6t
Xbit_r178_c87 bl[87] br[87] wl[178] vdd gnd cell_6t
Xbit_r179_c87 bl[87] br[87] wl[179] vdd gnd cell_6t
Xbit_r180_c87 bl[87] br[87] wl[180] vdd gnd cell_6t
Xbit_r181_c87 bl[87] br[87] wl[181] vdd gnd cell_6t
Xbit_r182_c87 bl[87] br[87] wl[182] vdd gnd cell_6t
Xbit_r183_c87 bl[87] br[87] wl[183] vdd gnd cell_6t
Xbit_r184_c87 bl[87] br[87] wl[184] vdd gnd cell_6t
Xbit_r185_c87 bl[87] br[87] wl[185] vdd gnd cell_6t
Xbit_r186_c87 bl[87] br[87] wl[186] vdd gnd cell_6t
Xbit_r187_c87 bl[87] br[87] wl[187] vdd gnd cell_6t
Xbit_r188_c87 bl[87] br[87] wl[188] vdd gnd cell_6t
Xbit_r189_c87 bl[87] br[87] wl[189] vdd gnd cell_6t
Xbit_r190_c87 bl[87] br[87] wl[190] vdd gnd cell_6t
Xbit_r191_c87 bl[87] br[87] wl[191] vdd gnd cell_6t
Xbit_r192_c87 bl[87] br[87] wl[192] vdd gnd cell_6t
Xbit_r193_c87 bl[87] br[87] wl[193] vdd gnd cell_6t
Xbit_r194_c87 bl[87] br[87] wl[194] vdd gnd cell_6t
Xbit_r195_c87 bl[87] br[87] wl[195] vdd gnd cell_6t
Xbit_r196_c87 bl[87] br[87] wl[196] vdd gnd cell_6t
Xbit_r197_c87 bl[87] br[87] wl[197] vdd gnd cell_6t
Xbit_r198_c87 bl[87] br[87] wl[198] vdd gnd cell_6t
Xbit_r199_c87 bl[87] br[87] wl[199] vdd gnd cell_6t
Xbit_r200_c87 bl[87] br[87] wl[200] vdd gnd cell_6t
Xbit_r201_c87 bl[87] br[87] wl[201] vdd gnd cell_6t
Xbit_r202_c87 bl[87] br[87] wl[202] vdd gnd cell_6t
Xbit_r203_c87 bl[87] br[87] wl[203] vdd gnd cell_6t
Xbit_r204_c87 bl[87] br[87] wl[204] vdd gnd cell_6t
Xbit_r205_c87 bl[87] br[87] wl[205] vdd gnd cell_6t
Xbit_r206_c87 bl[87] br[87] wl[206] vdd gnd cell_6t
Xbit_r207_c87 bl[87] br[87] wl[207] vdd gnd cell_6t
Xbit_r208_c87 bl[87] br[87] wl[208] vdd gnd cell_6t
Xbit_r209_c87 bl[87] br[87] wl[209] vdd gnd cell_6t
Xbit_r210_c87 bl[87] br[87] wl[210] vdd gnd cell_6t
Xbit_r211_c87 bl[87] br[87] wl[211] vdd gnd cell_6t
Xbit_r212_c87 bl[87] br[87] wl[212] vdd gnd cell_6t
Xbit_r213_c87 bl[87] br[87] wl[213] vdd gnd cell_6t
Xbit_r214_c87 bl[87] br[87] wl[214] vdd gnd cell_6t
Xbit_r215_c87 bl[87] br[87] wl[215] vdd gnd cell_6t
Xbit_r216_c87 bl[87] br[87] wl[216] vdd gnd cell_6t
Xbit_r217_c87 bl[87] br[87] wl[217] vdd gnd cell_6t
Xbit_r218_c87 bl[87] br[87] wl[218] vdd gnd cell_6t
Xbit_r219_c87 bl[87] br[87] wl[219] vdd gnd cell_6t
Xbit_r220_c87 bl[87] br[87] wl[220] vdd gnd cell_6t
Xbit_r221_c87 bl[87] br[87] wl[221] vdd gnd cell_6t
Xbit_r222_c87 bl[87] br[87] wl[222] vdd gnd cell_6t
Xbit_r223_c87 bl[87] br[87] wl[223] vdd gnd cell_6t
Xbit_r224_c87 bl[87] br[87] wl[224] vdd gnd cell_6t
Xbit_r225_c87 bl[87] br[87] wl[225] vdd gnd cell_6t
Xbit_r226_c87 bl[87] br[87] wl[226] vdd gnd cell_6t
Xbit_r227_c87 bl[87] br[87] wl[227] vdd gnd cell_6t
Xbit_r228_c87 bl[87] br[87] wl[228] vdd gnd cell_6t
Xbit_r229_c87 bl[87] br[87] wl[229] vdd gnd cell_6t
Xbit_r230_c87 bl[87] br[87] wl[230] vdd gnd cell_6t
Xbit_r231_c87 bl[87] br[87] wl[231] vdd gnd cell_6t
Xbit_r232_c87 bl[87] br[87] wl[232] vdd gnd cell_6t
Xbit_r233_c87 bl[87] br[87] wl[233] vdd gnd cell_6t
Xbit_r234_c87 bl[87] br[87] wl[234] vdd gnd cell_6t
Xbit_r235_c87 bl[87] br[87] wl[235] vdd gnd cell_6t
Xbit_r236_c87 bl[87] br[87] wl[236] vdd gnd cell_6t
Xbit_r237_c87 bl[87] br[87] wl[237] vdd gnd cell_6t
Xbit_r238_c87 bl[87] br[87] wl[238] vdd gnd cell_6t
Xbit_r239_c87 bl[87] br[87] wl[239] vdd gnd cell_6t
Xbit_r240_c87 bl[87] br[87] wl[240] vdd gnd cell_6t
Xbit_r241_c87 bl[87] br[87] wl[241] vdd gnd cell_6t
Xbit_r242_c87 bl[87] br[87] wl[242] vdd gnd cell_6t
Xbit_r243_c87 bl[87] br[87] wl[243] vdd gnd cell_6t
Xbit_r244_c87 bl[87] br[87] wl[244] vdd gnd cell_6t
Xbit_r245_c87 bl[87] br[87] wl[245] vdd gnd cell_6t
Xbit_r246_c87 bl[87] br[87] wl[246] vdd gnd cell_6t
Xbit_r247_c87 bl[87] br[87] wl[247] vdd gnd cell_6t
Xbit_r248_c87 bl[87] br[87] wl[248] vdd gnd cell_6t
Xbit_r249_c87 bl[87] br[87] wl[249] vdd gnd cell_6t
Xbit_r250_c87 bl[87] br[87] wl[250] vdd gnd cell_6t
Xbit_r251_c87 bl[87] br[87] wl[251] vdd gnd cell_6t
Xbit_r252_c87 bl[87] br[87] wl[252] vdd gnd cell_6t
Xbit_r253_c87 bl[87] br[87] wl[253] vdd gnd cell_6t
Xbit_r254_c87 bl[87] br[87] wl[254] vdd gnd cell_6t
Xbit_r255_c87 bl[87] br[87] wl[255] vdd gnd cell_6t
Xbit_r0_c88 bl[88] br[88] wl[0] vdd gnd cell_6t
Xbit_r1_c88 bl[88] br[88] wl[1] vdd gnd cell_6t
Xbit_r2_c88 bl[88] br[88] wl[2] vdd gnd cell_6t
Xbit_r3_c88 bl[88] br[88] wl[3] vdd gnd cell_6t
Xbit_r4_c88 bl[88] br[88] wl[4] vdd gnd cell_6t
Xbit_r5_c88 bl[88] br[88] wl[5] vdd gnd cell_6t
Xbit_r6_c88 bl[88] br[88] wl[6] vdd gnd cell_6t
Xbit_r7_c88 bl[88] br[88] wl[7] vdd gnd cell_6t
Xbit_r8_c88 bl[88] br[88] wl[8] vdd gnd cell_6t
Xbit_r9_c88 bl[88] br[88] wl[9] vdd gnd cell_6t
Xbit_r10_c88 bl[88] br[88] wl[10] vdd gnd cell_6t
Xbit_r11_c88 bl[88] br[88] wl[11] vdd gnd cell_6t
Xbit_r12_c88 bl[88] br[88] wl[12] vdd gnd cell_6t
Xbit_r13_c88 bl[88] br[88] wl[13] vdd gnd cell_6t
Xbit_r14_c88 bl[88] br[88] wl[14] vdd gnd cell_6t
Xbit_r15_c88 bl[88] br[88] wl[15] vdd gnd cell_6t
Xbit_r16_c88 bl[88] br[88] wl[16] vdd gnd cell_6t
Xbit_r17_c88 bl[88] br[88] wl[17] vdd gnd cell_6t
Xbit_r18_c88 bl[88] br[88] wl[18] vdd gnd cell_6t
Xbit_r19_c88 bl[88] br[88] wl[19] vdd gnd cell_6t
Xbit_r20_c88 bl[88] br[88] wl[20] vdd gnd cell_6t
Xbit_r21_c88 bl[88] br[88] wl[21] vdd gnd cell_6t
Xbit_r22_c88 bl[88] br[88] wl[22] vdd gnd cell_6t
Xbit_r23_c88 bl[88] br[88] wl[23] vdd gnd cell_6t
Xbit_r24_c88 bl[88] br[88] wl[24] vdd gnd cell_6t
Xbit_r25_c88 bl[88] br[88] wl[25] vdd gnd cell_6t
Xbit_r26_c88 bl[88] br[88] wl[26] vdd gnd cell_6t
Xbit_r27_c88 bl[88] br[88] wl[27] vdd gnd cell_6t
Xbit_r28_c88 bl[88] br[88] wl[28] vdd gnd cell_6t
Xbit_r29_c88 bl[88] br[88] wl[29] vdd gnd cell_6t
Xbit_r30_c88 bl[88] br[88] wl[30] vdd gnd cell_6t
Xbit_r31_c88 bl[88] br[88] wl[31] vdd gnd cell_6t
Xbit_r32_c88 bl[88] br[88] wl[32] vdd gnd cell_6t
Xbit_r33_c88 bl[88] br[88] wl[33] vdd gnd cell_6t
Xbit_r34_c88 bl[88] br[88] wl[34] vdd gnd cell_6t
Xbit_r35_c88 bl[88] br[88] wl[35] vdd gnd cell_6t
Xbit_r36_c88 bl[88] br[88] wl[36] vdd gnd cell_6t
Xbit_r37_c88 bl[88] br[88] wl[37] vdd gnd cell_6t
Xbit_r38_c88 bl[88] br[88] wl[38] vdd gnd cell_6t
Xbit_r39_c88 bl[88] br[88] wl[39] vdd gnd cell_6t
Xbit_r40_c88 bl[88] br[88] wl[40] vdd gnd cell_6t
Xbit_r41_c88 bl[88] br[88] wl[41] vdd gnd cell_6t
Xbit_r42_c88 bl[88] br[88] wl[42] vdd gnd cell_6t
Xbit_r43_c88 bl[88] br[88] wl[43] vdd gnd cell_6t
Xbit_r44_c88 bl[88] br[88] wl[44] vdd gnd cell_6t
Xbit_r45_c88 bl[88] br[88] wl[45] vdd gnd cell_6t
Xbit_r46_c88 bl[88] br[88] wl[46] vdd gnd cell_6t
Xbit_r47_c88 bl[88] br[88] wl[47] vdd gnd cell_6t
Xbit_r48_c88 bl[88] br[88] wl[48] vdd gnd cell_6t
Xbit_r49_c88 bl[88] br[88] wl[49] vdd gnd cell_6t
Xbit_r50_c88 bl[88] br[88] wl[50] vdd gnd cell_6t
Xbit_r51_c88 bl[88] br[88] wl[51] vdd gnd cell_6t
Xbit_r52_c88 bl[88] br[88] wl[52] vdd gnd cell_6t
Xbit_r53_c88 bl[88] br[88] wl[53] vdd gnd cell_6t
Xbit_r54_c88 bl[88] br[88] wl[54] vdd gnd cell_6t
Xbit_r55_c88 bl[88] br[88] wl[55] vdd gnd cell_6t
Xbit_r56_c88 bl[88] br[88] wl[56] vdd gnd cell_6t
Xbit_r57_c88 bl[88] br[88] wl[57] vdd gnd cell_6t
Xbit_r58_c88 bl[88] br[88] wl[58] vdd gnd cell_6t
Xbit_r59_c88 bl[88] br[88] wl[59] vdd gnd cell_6t
Xbit_r60_c88 bl[88] br[88] wl[60] vdd gnd cell_6t
Xbit_r61_c88 bl[88] br[88] wl[61] vdd gnd cell_6t
Xbit_r62_c88 bl[88] br[88] wl[62] vdd gnd cell_6t
Xbit_r63_c88 bl[88] br[88] wl[63] vdd gnd cell_6t
Xbit_r64_c88 bl[88] br[88] wl[64] vdd gnd cell_6t
Xbit_r65_c88 bl[88] br[88] wl[65] vdd gnd cell_6t
Xbit_r66_c88 bl[88] br[88] wl[66] vdd gnd cell_6t
Xbit_r67_c88 bl[88] br[88] wl[67] vdd gnd cell_6t
Xbit_r68_c88 bl[88] br[88] wl[68] vdd gnd cell_6t
Xbit_r69_c88 bl[88] br[88] wl[69] vdd gnd cell_6t
Xbit_r70_c88 bl[88] br[88] wl[70] vdd gnd cell_6t
Xbit_r71_c88 bl[88] br[88] wl[71] vdd gnd cell_6t
Xbit_r72_c88 bl[88] br[88] wl[72] vdd gnd cell_6t
Xbit_r73_c88 bl[88] br[88] wl[73] vdd gnd cell_6t
Xbit_r74_c88 bl[88] br[88] wl[74] vdd gnd cell_6t
Xbit_r75_c88 bl[88] br[88] wl[75] vdd gnd cell_6t
Xbit_r76_c88 bl[88] br[88] wl[76] vdd gnd cell_6t
Xbit_r77_c88 bl[88] br[88] wl[77] vdd gnd cell_6t
Xbit_r78_c88 bl[88] br[88] wl[78] vdd gnd cell_6t
Xbit_r79_c88 bl[88] br[88] wl[79] vdd gnd cell_6t
Xbit_r80_c88 bl[88] br[88] wl[80] vdd gnd cell_6t
Xbit_r81_c88 bl[88] br[88] wl[81] vdd gnd cell_6t
Xbit_r82_c88 bl[88] br[88] wl[82] vdd gnd cell_6t
Xbit_r83_c88 bl[88] br[88] wl[83] vdd gnd cell_6t
Xbit_r84_c88 bl[88] br[88] wl[84] vdd gnd cell_6t
Xbit_r85_c88 bl[88] br[88] wl[85] vdd gnd cell_6t
Xbit_r86_c88 bl[88] br[88] wl[86] vdd gnd cell_6t
Xbit_r87_c88 bl[88] br[88] wl[87] vdd gnd cell_6t
Xbit_r88_c88 bl[88] br[88] wl[88] vdd gnd cell_6t
Xbit_r89_c88 bl[88] br[88] wl[89] vdd gnd cell_6t
Xbit_r90_c88 bl[88] br[88] wl[90] vdd gnd cell_6t
Xbit_r91_c88 bl[88] br[88] wl[91] vdd gnd cell_6t
Xbit_r92_c88 bl[88] br[88] wl[92] vdd gnd cell_6t
Xbit_r93_c88 bl[88] br[88] wl[93] vdd gnd cell_6t
Xbit_r94_c88 bl[88] br[88] wl[94] vdd gnd cell_6t
Xbit_r95_c88 bl[88] br[88] wl[95] vdd gnd cell_6t
Xbit_r96_c88 bl[88] br[88] wl[96] vdd gnd cell_6t
Xbit_r97_c88 bl[88] br[88] wl[97] vdd gnd cell_6t
Xbit_r98_c88 bl[88] br[88] wl[98] vdd gnd cell_6t
Xbit_r99_c88 bl[88] br[88] wl[99] vdd gnd cell_6t
Xbit_r100_c88 bl[88] br[88] wl[100] vdd gnd cell_6t
Xbit_r101_c88 bl[88] br[88] wl[101] vdd gnd cell_6t
Xbit_r102_c88 bl[88] br[88] wl[102] vdd gnd cell_6t
Xbit_r103_c88 bl[88] br[88] wl[103] vdd gnd cell_6t
Xbit_r104_c88 bl[88] br[88] wl[104] vdd gnd cell_6t
Xbit_r105_c88 bl[88] br[88] wl[105] vdd gnd cell_6t
Xbit_r106_c88 bl[88] br[88] wl[106] vdd gnd cell_6t
Xbit_r107_c88 bl[88] br[88] wl[107] vdd gnd cell_6t
Xbit_r108_c88 bl[88] br[88] wl[108] vdd gnd cell_6t
Xbit_r109_c88 bl[88] br[88] wl[109] vdd gnd cell_6t
Xbit_r110_c88 bl[88] br[88] wl[110] vdd gnd cell_6t
Xbit_r111_c88 bl[88] br[88] wl[111] vdd gnd cell_6t
Xbit_r112_c88 bl[88] br[88] wl[112] vdd gnd cell_6t
Xbit_r113_c88 bl[88] br[88] wl[113] vdd gnd cell_6t
Xbit_r114_c88 bl[88] br[88] wl[114] vdd gnd cell_6t
Xbit_r115_c88 bl[88] br[88] wl[115] vdd gnd cell_6t
Xbit_r116_c88 bl[88] br[88] wl[116] vdd gnd cell_6t
Xbit_r117_c88 bl[88] br[88] wl[117] vdd gnd cell_6t
Xbit_r118_c88 bl[88] br[88] wl[118] vdd gnd cell_6t
Xbit_r119_c88 bl[88] br[88] wl[119] vdd gnd cell_6t
Xbit_r120_c88 bl[88] br[88] wl[120] vdd gnd cell_6t
Xbit_r121_c88 bl[88] br[88] wl[121] vdd gnd cell_6t
Xbit_r122_c88 bl[88] br[88] wl[122] vdd gnd cell_6t
Xbit_r123_c88 bl[88] br[88] wl[123] vdd gnd cell_6t
Xbit_r124_c88 bl[88] br[88] wl[124] vdd gnd cell_6t
Xbit_r125_c88 bl[88] br[88] wl[125] vdd gnd cell_6t
Xbit_r126_c88 bl[88] br[88] wl[126] vdd gnd cell_6t
Xbit_r127_c88 bl[88] br[88] wl[127] vdd gnd cell_6t
Xbit_r128_c88 bl[88] br[88] wl[128] vdd gnd cell_6t
Xbit_r129_c88 bl[88] br[88] wl[129] vdd gnd cell_6t
Xbit_r130_c88 bl[88] br[88] wl[130] vdd gnd cell_6t
Xbit_r131_c88 bl[88] br[88] wl[131] vdd gnd cell_6t
Xbit_r132_c88 bl[88] br[88] wl[132] vdd gnd cell_6t
Xbit_r133_c88 bl[88] br[88] wl[133] vdd gnd cell_6t
Xbit_r134_c88 bl[88] br[88] wl[134] vdd gnd cell_6t
Xbit_r135_c88 bl[88] br[88] wl[135] vdd gnd cell_6t
Xbit_r136_c88 bl[88] br[88] wl[136] vdd gnd cell_6t
Xbit_r137_c88 bl[88] br[88] wl[137] vdd gnd cell_6t
Xbit_r138_c88 bl[88] br[88] wl[138] vdd gnd cell_6t
Xbit_r139_c88 bl[88] br[88] wl[139] vdd gnd cell_6t
Xbit_r140_c88 bl[88] br[88] wl[140] vdd gnd cell_6t
Xbit_r141_c88 bl[88] br[88] wl[141] vdd gnd cell_6t
Xbit_r142_c88 bl[88] br[88] wl[142] vdd gnd cell_6t
Xbit_r143_c88 bl[88] br[88] wl[143] vdd gnd cell_6t
Xbit_r144_c88 bl[88] br[88] wl[144] vdd gnd cell_6t
Xbit_r145_c88 bl[88] br[88] wl[145] vdd gnd cell_6t
Xbit_r146_c88 bl[88] br[88] wl[146] vdd gnd cell_6t
Xbit_r147_c88 bl[88] br[88] wl[147] vdd gnd cell_6t
Xbit_r148_c88 bl[88] br[88] wl[148] vdd gnd cell_6t
Xbit_r149_c88 bl[88] br[88] wl[149] vdd gnd cell_6t
Xbit_r150_c88 bl[88] br[88] wl[150] vdd gnd cell_6t
Xbit_r151_c88 bl[88] br[88] wl[151] vdd gnd cell_6t
Xbit_r152_c88 bl[88] br[88] wl[152] vdd gnd cell_6t
Xbit_r153_c88 bl[88] br[88] wl[153] vdd gnd cell_6t
Xbit_r154_c88 bl[88] br[88] wl[154] vdd gnd cell_6t
Xbit_r155_c88 bl[88] br[88] wl[155] vdd gnd cell_6t
Xbit_r156_c88 bl[88] br[88] wl[156] vdd gnd cell_6t
Xbit_r157_c88 bl[88] br[88] wl[157] vdd gnd cell_6t
Xbit_r158_c88 bl[88] br[88] wl[158] vdd gnd cell_6t
Xbit_r159_c88 bl[88] br[88] wl[159] vdd gnd cell_6t
Xbit_r160_c88 bl[88] br[88] wl[160] vdd gnd cell_6t
Xbit_r161_c88 bl[88] br[88] wl[161] vdd gnd cell_6t
Xbit_r162_c88 bl[88] br[88] wl[162] vdd gnd cell_6t
Xbit_r163_c88 bl[88] br[88] wl[163] vdd gnd cell_6t
Xbit_r164_c88 bl[88] br[88] wl[164] vdd gnd cell_6t
Xbit_r165_c88 bl[88] br[88] wl[165] vdd gnd cell_6t
Xbit_r166_c88 bl[88] br[88] wl[166] vdd gnd cell_6t
Xbit_r167_c88 bl[88] br[88] wl[167] vdd gnd cell_6t
Xbit_r168_c88 bl[88] br[88] wl[168] vdd gnd cell_6t
Xbit_r169_c88 bl[88] br[88] wl[169] vdd gnd cell_6t
Xbit_r170_c88 bl[88] br[88] wl[170] vdd gnd cell_6t
Xbit_r171_c88 bl[88] br[88] wl[171] vdd gnd cell_6t
Xbit_r172_c88 bl[88] br[88] wl[172] vdd gnd cell_6t
Xbit_r173_c88 bl[88] br[88] wl[173] vdd gnd cell_6t
Xbit_r174_c88 bl[88] br[88] wl[174] vdd gnd cell_6t
Xbit_r175_c88 bl[88] br[88] wl[175] vdd gnd cell_6t
Xbit_r176_c88 bl[88] br[88] wl[176] vdd gnd cell_6t
Xbit_r177_c88 bl[88] br[88] wl[177] vdd gnd cell_6t
Xbit_r178_c88 bl[88] br[88] wl[178] vdd gnd cell_6t
Xbit_r179_c88 bl[88] br[88] wl[179] vdd gnd cell_6t
Xbit_r180_c88 bl[88] br[88] wl[180] vdd gnd cell_6t
Xbit_r181_c88 bl[88] br[88] wl[181] vdd gnd cell_6t
Xbit_r182_c88 bl[88] br[88] wl[182] vdd gnd cell_6t
Xbit_r183_c88 bl[88] br[88] wl[183] vdd gnd cell_6t
Xbit_r184_c88 bl[88] br[88] wl[184] vdd gnd cell_6t
Xbit_r185_c88 bl[88] br[88] wl[185] vdd gnd cell_6t
Xbit_r186_c88 bl[88] br[88] wl[186] vdd gnd cell_6t
Xbit_r187_c88 bl[88] br[88] wl[187] vdd gnd cell_6t
Xbit_r188_c88 bl[88] br[88] wl[188] vdd gnd cell_6t
Xbit_r189_c88 bl[88] br[88] wl[189] vdd gnd cell_6t
Xbit_r190_c88 bl[88] br[88] wl[190] vdd gnd cell_6t
Xbit_r191_c88 bl[88] br[88] wl[191] vdd gnd cell_6t
Xbit_r192_c88 bl[88] br[88] wl[192] vdd gnd cell_6t
Xbit_r193_c88 bl[88] br[88] wl[193] vdd gnd cell_6t
Xbit_r194_c88 bl[88] br[88] wl[194] vdd gnd cell_6t
Xbit_r195_c88 bl[88] br[88] wl[195] vdd gnd cell_6t
Xbit_r196_c88 bl[88] br[88] wl[196] vdd gnd cell_6t
Xbit_r197_c88 bl[88] br[88] wl[197] vdd gnd cell_6t
Xbit_r198_c88 bl[88] br[88] wl[198] vdd gnd cell_6t
Xbit_r199_c88 bl[88] br[88] wl[199] vdd gnd cell_6t
Xbit_r200_c88 bl[88] br[88] wl[200] vdd gnd cell_6t
Xbit_r201_c88 bl[88] br[88] wl[201] vdd gnd cell_6t
Xbit_r202_c88 bl[88] br[88] wl[202] vdd gnd cell_6t
Xbit_r203_c88 bl[88] br[88] wl[203] vdd gnd cell_6t
Xbit_r204_c88 bl[88] br[88] wl[204] vdd gnd cell_6t
Xbit_r205_c88 bl[88] br[88] wl[205] vdd gnd cell_6t
Xbit_r206_c88 bl[88] br[88] wl[206] vdd gnd cell_6t
Xbit_r207_c88 bl[88] br[88] wl[207] vdd gnd cell_6t
Xbit_r208_c88 bl[88] br[88] wl[208] vdd gnd cell_6t
Xbit_r209_c88 bl[88] br[88] wl[209] vdd gnd cell_6t
Xbit_r210_c88 bl[88] br[88] wl[210] vdd gnd cell_6t
Xbit_r211_c88 bl[88] br[88] wl[211] vdd gnd cell_6t
Xbit_r212_c88 bl[88] br[88] wl[212] vdd gnd cell_6t
Xbit_r213_c88 bl[88] br[88] wl[213] vdd gnd cell_6t
Xbit_r214_c88 bl[88] br[88] wl[214] vdd gnd cell_6t
Xbit_r215_c88 bl[88] br[88] wl[215] vdd gnd cell_6t
Xbit_r216_c88 bl[88] br[88] wl[216] vdd gnd cell_6t
Xbit_r217_c88 bl[88] br[88] wl[217] vdd gnd cell_6t
Xbit_r218_c88 bl[88] br[88] wl[218] vdd gnd cell_6t
Xbit_r219_c88 bl[88] br[88] wl[219] vdd gnd cell_6t
Xbit_r220_c88 bl[88] br[88] wl[220] vdd gnd cell_6t
Xbit_r221_c88 bl[88] br[88] wl[221] vdd gnd cell_6t
Xbit_r222_c88 bl[88] br[88] wl[222] vdd gnd cell_6t
Xbit_r223_c88 bl[88] br[88] wl[223] vdd gnd cell_6t
Xbit_r224_c88 bl[88] br[88] wl[224] vdd gnd cell_6t
Xbit_r225_c88 bl[88] br[88] wl[225] vdd gnd cell_6t
Xbit_r226_c88 bl[88] br[88] wl[226] vdd gnd cell_6t
Xbit_r227_c88 bl[88] br[88] wl[227] vdd gnd cell_6t
Xbit_r228_c88 bl[88] br[88] wl[228] vdd gnd cell_6t
Xbit_r229_c88 bl[88] br[88] wl[229] vdd gnd cell_6t
Xbit_r230_c88 bl[88] br[88] wl[230] vdd gnd cell_6t
Xbit_r231_c88 bl[88] br[88] wl[231] vdd gnd cell_6t
Xbit_r232_c88 bl[88] br[88] wl[232] vdd gnd cell_6t
Xbit_r233_c88 bl[88] br[88] wl[233] vdd gnd cell_6t
Xbit_r234_c88 bl[88] br[88] wl[234] vdd gnd cell_6t
Xbit_r235_c88 bl[88] br[88] wl[235] vdd gnd cell_6t
Xbit_r236_c88 bl[88] br[88] wl[236] vdd gnd cell_6t
Xbit_r237_c88 bl[88] br[88] wl[237] vdd gnd cell_6t
Xbit_r238_c88 bl[88] br[88] wl[238] vdd gnd cell_6t
Xbit_r239_c88 bl[88] br[88] wl[239] vdd gnd cell_6t
Xbit_r240_c88 bl[88] br[88] wl[240] vdd gnd cell_6t
Xbit_r241_c88 bl[88] br[88] wl[241] vdd gnd cell_6t
Xbit_r242_c88 bl[88] br[88] wl[242] vdd gnd cell_6t
Xbit_r243_c88 bl[88] br[88] wl[243] vdd gnd cell_6t
Xbit_r244_c88 bl[88] br[88] wl[244] vdd gnd cell_6t
Xbit_r245_c88 bl[88] br[88] wl[245] vdd gnd cell_6t
Xbit_r246_c88 bl[88] br[88] wl[246] vdd gnd cell_6t
Xbit_r247_c88 bl[88] br[88] wl[247] vdd gnd cell_6t
Xbit_r248_c88 bl[88] br[88] wl[248] vdd gnd cell_6t
Xbit_r249_c88 bl[88] br[88] wl[249] vdd gnd cell_6t
Xbit_r250_c88 bl[88] br[88] wl[250] vdd gnd cell_6t
Xbit_r251_c88 bl[88] br[88] wl[251] vdd gnd cell_6t
Xbit_r252_c88 bl[88] br[88] wl[252] vdd gnd cell_6t
Xbit_r253_c88 bl[88] br[88] wl[253] vdd gnd cell_6t
Xbit_r254_c88 bl[88] br[88] wl[254] vdd gnd cell_6t
Xbit_r255_c88 bl[88] br[88] wl[255] vdd gnd cell_6t
Xbit_r0_c89 bl[89] br[89] wl[0] vdd gnd cell_6t
Xbit_r1_c89 bl[89] br[89] wl[1] vdd gnd cell_6t
Xbit_r2_c89 bl[89] br[89] wl[2] vdd gnd cell_6t
Xbit_r3_c89 bl[89] br[89] wl[3] vdd gnd cell_6t
Xbit_r4_c89 bl[89] br[89] wl[4] vdd gnd cell_6t
Xbit_r5_c89 bl[89] br[89] wl[5] vdd gnd cell_6t
Xbit_r6_c89 bl[89] br[89] wl[6] vdd gnd cell_6t
Xbit_r7_c89 bl[89] br[89] wl[7] vdd gnd cell_6t
Xbit_r8_c89 bl[89] br[89] wl[8] vdd gnd cell_6t
Xbit_r9_c89 bl[89] br[89] wl[9] vdd gnd cell_6t
Xbit_r10_c89 bl[89] br[89] wl[10] vdd gnd cell_6t
Xbit_r11_c89 bl[89] br[89] wl[11] vdd gnd cell_6t
Xbit_r12_c89 bl[89] br[89] wl[12] vdd gnd cell_6t
Xbit_r13_c89 bl[89] br[89] wl[13] vdd gnd cell_6t
Xbit_r14_c89 bl[89] br[89] wl[14] vdd gnd cell_6t
Xbit_r15_c89 bl[89] br[89] wl[15] vdd gnd cell_6t
Xbit_r16_c89 bl[89] br[89] wl[16] vdd gnd cell_6t
Xbit_r17_c89 bl[89] br[89] wl[17] vdd gnd cell_6t
Xbit_r18_c89 bl[89] br[89] wl[18] vdd gnd cell_6t
Xbit_r19_c89 bl[89] br[89] wl[19] vdd gnd cell_6t
Xbit_r20_c89 bl[89] br[89] wl[20] vdd gnd cell_6t
Xbit_r21_c89 bl[89] br[89] wl[21] vdd gnd cell_6t
Xbit_r22_c89 bl[89] br[89] wl[22] vdd gnd cell_6t
Xbit_r23_c89 bl[89] br[89] wl[23] vdd gnd cell_6t
Xbit_r24_c89 bl[89] br[89] wl[24] vdd gnd cell_6t
Xbit_r25_c89 bl[89] br[89] wl[25] vdd gnd cell_6t
Xbit_r26_c89 bl[89] br[89] wl[26] vdd gnd cell_6t
Xbit_r27_c89 bl[89] br[89] wl[27] vdd gnd cell_6t
Xbit_r28_c89 bl[89] br[89] wl[28] vdd gnd cell_6t
Xbit_r29_c89 bl[89] br[89] wl[29] vdd gnd cell_6t
Xbit_r30_c89 bl[89] br[89] wl[30] vdd gnd cell_6t
Xbit_r31_c89 bl[89] br[89] wl[31] vdd gnd cell_6t
Xbit_r32_c89 bl[89] br[89] wl[32] vdd gnd cell_6t
Xbit_r33_c89 bl[89] br[89] wl[33] vdd gnd cell_6t
Xbit_r34_c89 bl[89] br[89] wl[34] vdd gnd cell_6t
Xbit_r35_c89 bl[89] br[89] wl[35] vdd gnd cell_6t
Xbit_r36_c89 bl[89] br[89] wl[36] vdd gnd cell_6t
Xbit_r37_c89 bl[89] br[89] wl[37] vdd gnd cell_6t
Xbit_r38_c89 bl[89] br[89] wl[38] vdd gnd cell_6t
Xbit_r39_c89 bl[89] br[89] wl[39] vdd gnd cell_6t
Xbit_r40_c89 bl[89] br[89] wl[40] vdd gnd cell_6t
Xbit_r41_c89 bl[89] br[89] wl[41] vdd gnd cell_6t
Xbit_r42_c89 bl[89] br[89] wl[42] vdd gnd cell_6t
Xbit_r43_c89 bl[89] br[89] wl[43] vdd gnd cell_6t
Xbit_r44_c89 bl[89] br[89] wl[44] vdd gnd cell_6t
Xbit_r45_c89 bl[89] br[89] wl[45] vdd gnd cell_6t
Xbit_r46_c89 bl[89] br[89] wl[46] vdd gnd cell_6t
Xbit_r47_c89 bl[89] br[89] wl[47] vdd gnd cell_6t
Xbit_r48_c89 bl[89] br[89] wl[48] vdd gnd cell_6t
Xbit_r49_c89 bl[89] br[89] wl[49] vdd gnd cell_6t
Xbit_r50_c89 bl[89] br[89] wl[50] vdd gnd cell_6t
Xbit_r51_c89 bl[89] br[89] wl[51] vdd gnd cell_6t
Xbit_r52_c89 bl[89] br[89] wl[52] vdd gnd cell_6t
Xbit_r53_c89 bl[89] br[89] wl[53] vdd gnd cell_6t
Xbit_r54_c89 bl[89] br[89] wl[54] vdd gnd cell_6t
Xbit_r55_c89 bl[89] br[89] wl[55] vdd gnd cell_6t
Xbit_r56_c89 bl[89] br[89] wl[56] vdd gnd cell_6t
Xbit_r57_c89 bl[89] br[89] wl[57] vdd gnd cell_6t
Xbit_r58_c89 bl[89] br[89] wl[58] vdd gnd cell_6t
Xbit_r59_c89 bl[89] br[89] wl[59] vdd gnd cell_6t
Xbit_r60_c89 bl[89] br[89] wl[60] vdd gnd cell_6t
Xbit_r61_c89 bl[89] br[89] wl[61] vdd gnd cell_6t
Xbit_r62_c89 bl[89] br[89] wl[62] vdd gnd cell_6t
Xbit_r63_c89 bl[89] br[89] wl[63] vdd gnd cell_6t
Xbit_r64_c89 bl[89] br[89] wl[64] vdd gnd cell_6t
Xbit_r65_c89 bl[89] br[89] wl[65] vdd gnd cell_6t
Xbit_r66_c89 bl[89] br[89] wl[66] vdd gnd cell_6t
Xbit_r67_c89 bl[89] br[89] wl[67] vdd gnd cell_6t
Xbit_r68_c89 bl[89] br[89] wl[68] vdd gnd cell_6t
Xbit_r69_c89 bl[89] br[89] wl[69] vdd gnd cell_6t
Xbit_r70_c89 bl[89] br[89] wl[70] vdd gnd cell_6t
Xbit_r71_c89 bl[89] br[89] wl[71] vdd gnd cell_6t
Xbit_r72_c89 bl[89] br[89] wl[72] vdd gnd cell_6t
Xbit_r73_c89 bl[89] br[89] wl[73] vdd gnd cell_6t
Xbit_r74_c89 bl[89] br[89] wl[74] vdd gnd cell_6t
Xbit_r75_c89 bl[89] br[89] wl[75] vdd gnd cell_6t
Xbit_r76_c89 bl[89] br[89] wl[76] vdd gnd cell_6t
Xbit_r77_c89 bl[89] br[89] wl[77] vdd gnd cell_6t
Xbit_r78_c89 bl[89] br[89] wl[78] vdd gnd cell_6t
Xbit_r79_c89 bl[89] br[89] wl[79] vdd gnd cell_6t
Xbit_r80_c89 bl[89] br[89] wl[80] vdd gnd cell_6t
Xbit_r81_c89 bl[89] br[89] wl[81] vdd gnd cell_6t
Xbit_r82_c89 bl[89] br[89] wl[82] vdd gnd cell_6t
Xbit_r83_c89 bl[89] br[89] wl[83] vdd gnd cell_6t
Xbit_r84_c89 bl[89] br[89] wl[84] vdd gnd cell_6t
Xbit_r85_c89 bl[89] br[89] wl[85] vdd gnd cell_6t
Xbit_r86_c89 bl[89] br[89] wl[86] vdd gnd cell_6t
Xbit_r87_c89 bl[89] br[89] wl[87] vdd gnd cell_6t
Xbit_r88_c89 bl[89] br[89] wl[88] vdd gnd cell_6t
Xbit_r89_c89 bl[89] br[89] wl[89] vdd gnd cell_6t
Xbit_r90_c89 bl[89] br[89] wl[90] vdd gnd cell_6t
Xbit_r91_c89 bl[89] br[89] wl[91] vdd gnd cell_6t
Xbit_r92_c89 bl[89] br[89] wl[92] vdd gnd cell_6t
Xbit_r93_c89 bl[89] br[89] wl[93] vdd gnd cell_6t
Xbit_r94_c89 bl[89] br[89] wl[94] vdd gnd cell_6t
Xbit_r95_c89 bl[89] br[89] wl[95] vdd gnd cell_6t
Xbit_r96_c89 bl[89] br[89] wl[96] vdd gnd cell_6t
Xbit_r97_c89 bl[89] br[89] wl[97] vdd gnd cell_6t
Xbit_r98_c89 bl[89] br[89] wl[98] vdd gnd cell_6t
Xbit_r99_c89 bl[89] br[89] wl[99] vdd gnd cell_6t
Xbit_r100_c89 bl[89] br[89] wl[100] vdd gnd cell_6t
Xbit_r101_c89 bl[89] br[89] wl[101] vdd gnd cell_6t
Xbit_r102_c89 bl[89] br[89] wl[102] vdd gnd cell_6t
Xbit_r103_c89 bl[89] br[89] wl[103] vdd gnd cell_6t
Xbit_r104_c89 bl[89] br[89] wl[104] vdd gnd cell_6t
Xbit_r105_c89 bl[89] br[89] wl[105] vdd gnd cell_6t
Xbit_r106_c89 bl[89] br[89] wl[106] vdd gnd cell_6t
Xbit_r107_c89 bl[89] br[89] wl[107] vdd gnd cell_6t
Xbit_r108_c89 bl[89] br[89] wl[108] vdd gnd cell_6t
Xbit_r109_c89 bl[89] br[89] wl[109] vdd gnd cell_6t
Xbit_r110_c89 bl[89] br[89] wl[110] vdd gnd cell_6t
Xbit_r111_c89 bl[89] br[89] wl[111] vdd gnd cell_6t
Xbit_r112_c89 bl[89] br[89] wl[112] vdd gnd cell_6t
Xbit_r113_c89 bl[89] br[89] wl[113] vdd gnd cell_6t
Xbit_r114_c89 bl[89] br[89] wl[114] vdd gnd cell_6t
Xbit_r115_c89 bl[89] br[89] wl[115] vdd gnd cell_6t
Xbit_r116_c89 bl[89] br[89] wl[116] vdd gnd cell_6t
Xbit_r117_c89 bl[89] br[89] wl[117] vdd gnd cell_6t
Xbit_r118_c89 bl[89] br[89] wl[118] vdd gnd cell_6t
Xbit_r119_c89 bl[89] br[89] wl[119] vdd gnd cell_6t
Xbit_r120_c89 bl[89] br[89] wl[120] vdd gnd cell_6t
Xbit_r121_c89 bl[89] br[89] wl[121] vdd gnd cell_6t
Xbit_r122_c89 bl[89] br[89] wl[122] vdd gnd cell_6t
Xbit_r123_c89 bl[89] br[89] wl[123] vdd gnd cell_6t
Xbit_r124_c89 bl[89] br[89] wl[124] vdd gnd cell_6t
Xbit_r125_c89 bl[89] br[89] wl[125] vdd gnd cell_6t
Xbit_r126_c89 bl[89] br[89] wl[126] vdd gnd cell_6t
Xbit_r127_c89 bl[89] br[89] wl[127] vdd gnd cell_6t
Xbit_r128_c89 bl[89] br[89] wl[128] vdd gnd cell_6t
Xbit_r129_c89 bl[89] br[89] wl[129] vdd gnd cell_6t
Xbit_r130_c89 bl[89] br[89] wl[130] vdd gnd cell_6t
Xbit_r131_c89 bl[89] br[89] wl[131] vdd gnd cell_6t
Xbit_r132_c89 bl[89] br[89] wl[132] vdd gnd cell_6t
Xbit_r133_c89 bl[89] br[89] wl[133] vdd gnd cell_6t
Xbit_r134_c89 bl[89] br[89] wl[134] vdd gnd cell_6t
Xbit_r135_c89 bl[89] br[89] wl[135] vdd gnd cell_6t
Xbit_r136_c89 bl[89] br[89] wl[136] vdd gnd cell_6t
Xbit_r137_c89 bl[89] br[89] wl[137] vdd gnd cell_6t
Xbit_r138_c89 bl[89] br[89] wl[138] vdd gnd cell_6t
Xbit_r139_c89 bl[89] br[89] wl[139] vdd gnd cell_6t
Xbit_r140_c89 bl[89] br[89] wl[140] vdd gnd cell_6t
Xbit_r141_c89 bl[89] br[89] wl[141] vdd gnd cell_6t
Xbit_r142_c89 bl[89] br[89] wl[142] vdd gnd cell_6t
Xbit_r143_c89 bl[89] br[89] wl[143] vdd gnd cell_6t
Xbit_r144_c89 bl[89] br[89] wl[144] vdd gnd cell_6t
Xbit_r145_c89 bl[89] br[89] wl[145] vdd gnd cell_6t
Xbit_r146_c89 bl[89] br[89] wl[146] vdd gnd cell_6t
Xbit_r147_c89 bl[89] br[89] wl[147] vdd gnd cell_6t
Xbit_r148_c89 bl[89] br[89] wl[148] vdd gnd cell_6t
Xbit_r149_c89 bl[89] br[89] wl[149] vdd gnd cell_6t
Xbit_r150_c89 bl[89] br[89] wl[150] vdd gnd cell_6t
Xbit_r151_c89 bl[89] br[89] wl[151] vdd gnd cell_6t
Xbit_r152_c89 bl[89] br[89] wl[152] vdd gnd cell_6t
Xbit_r153_c89 bl[89] br[89] wl[153] vdd gnd cell_6t
Xbit_r154_c89 bl[89] br[89] wl[154] vdd gnd cell_6t
Xbit_r155_c89 bl[89] br[89] wl[155] vdd gnd cell_6t
Xbit_r156_c89 bl[89] br[89] wl[156] vdd gnd cell_6t
Xbit_r157_c89 bl[89] br[89] wl[157] vdd gnd cell_6t
Xbit_r158_c89 bl[89] br[89] wl[158] vdd gnd cell_6t
Xbit_r159_c89 bl[89] br[89] wl[159] vdd gnd cell_6t
Xbit_r160_c89 bl[89] br[89] wl[160] vdd gnd cell_6t
Xbit_r161_c89 bl[89] br[89] wl[161] vdd gnd cell_6t
Xbit_r162_c89 bl[89] br[89] wl[162] vdd gnd cell_6t
Xbit_r163_c89 bl[89] br[89] wl[163] vdd gnd cell_6t
Xbit_r164_c89 bl[89] br[89] wl[164] vdd gnd cell_6t
Xbit_r165_c89 bl[89] br[89] wl[165] vdd gnd cell_6t
Xbit_r166_c89 bl[89] br[89] wl[166] vdd gnd cell_6t
Xbit_r167_c89 bl[89] br[89] wl[167] vdd gnd cell_6t
Xbit_r168_c89 bl[89] br[89] wl[168] vdd gnd cell_6t
Xbit_r169_c89 bl[89] br[89] wl[169] vdd gnd cell_6t
Xbit_r170_c89 bl[89] br[89] wl[170] vdd gnd cell_6t
Xbit_r171_c89 bl[89] br[89] wl[171] vdd gnd cell_6t
Xbit_r172_c89 bl[89] br[89] wl[172] vdd gnd cell_6t
Xbit_r173_c89 bl[89] br[89] wl[173] vdd gnd cell_6t
Xbit_r174_c89 bl[89] br[89] wl[174] vdd gnd cell_6t
Xbit_r175_c89 bl[89] br[89] wl[175] vdd gnd cell_6t
Xbit_r176_c89 bl[89] br[89] wl[176] vdd gnd cell_6t
Xbit_r177_c89 bl[89] br[89] wl[177] vdd gnd cell_6t
Xbit_r178_c89 bl[89] br[89] wl[178] vdd gnd cell_6t
Xbit_r179_c89 bl[89] br[89] wl[179] vdd gnd cell_6t
Xbit_r180_c89 bl[89] br[89] wl[180] vdd gnd cell_6t
Xbit_r181_c89 bl[89] br[89] wl[181] vdd gnd cell_6t
Xbit_r182_c89 bl[89] br[89] wl[182] vdd gnd cell_6t
Xbit_r183_c89 bl[89] br[89] wl[183] vdd gnd cell_6t
Xbit_r184_c89 bl[89] br[89] wl[184] vdd gnd cell_6t
Xbit_r185_c89 bl[89] br[89] wl[185] vdd gnd cell_6t
Xbit_r186_c89 bl[89] br[89] wl[186] vdd gnd cell_6t
Xbit_r187_c89 bl[89] br[89] wl[187] vdd gnd cell_6t
Xbit_r188_c89 bl[89] br[89] wl[188] vdd gnd cell_6t
Xbit_r189_c89 bl[89] br[89] wl[189] vdd gnd cell_6t
Xbit_r190_c89 bl[89] br[89] wl[190] vdd gnd cell_6t
Xbit_r191_c89 bl[89] br[89] wl[191] vdd gnd cell_6t
Xbit_r192_c89 bl[89] br[89] wl[192] vdd gnd cell_6t
Xbit_r193_c89 bl[89] br[89] wl[193] vdd gnd cell_6t
Xbit_r194_c89 bl[89] br[89] wl[194] vdd gnd cell_6t
Xbit_r195_c89 bl[89] br[89] wl[195] vdd gnd cell_6t
Xbit_r196_c89 bl[89] br[89] wl[196] vdd gnd cell_6t
Xbit_r197_c89 bl[89] br[89] wl[197] vdd gnd cell_6t
Xbit_r198_c89 bl[89] br[89] wl[198] vdd gnd cell_6t
Xbit_r199_c89 bl[89] br[89] wl[199] vdd gnd cell_6t
Xbit_r200_c89 bl[89] br[89] wl[200] vdd gnd cell_6t
Xbit_r201_c89 bl[89] br[89] wl[201] vdd gnd cell_6t
Xbit_r202_c89 bl[89] br[89] wl[202] vdd gnd cell_6t
Xbit_r203_c89 bl[89] br[89] wl[203] vdd gnd cell_6t
Xbit_r204_c89 bl[89] br[89] wl[204] vdd gnd cell_6t
Xbit_r205_c89 bl[89] br[89] wl[205] vdd gnd cell_6t
Xbit_r206_c89 bl[89] br[89] wl[206] vdd gnd cell_6t
Xbit_r207_c89 bl[89] br[89] wl[207] vdd gnd cell_6t
Xbit_r208_c89 bl[89] br[89] wl[208] vdd gnd cell_6t
Xbit_r209_c89 bl[89] br[89] wl[209] vdd gnd cell_6t
Xbit_r210_c89 bl[89] br[89] wl[210] vdd gnd cell_6t
Xbit_r211_c89 bl[89] br[89] wl[211] vdd gnd cell_6t
Xbit_r212_c89 bl[89] br[89] wl[212] vdd gnd cell_6t
Xbit_r213_c89 bl[89] br[89] wl[213] vdd gnd cell_6t
Xbit_r214_c89 bl[89] br[89] wl[214] vdd gnd cell_6t
Xbit_r215_c89 bl[89] br[89] wl[215] vdd gnd cell_6t
Xbit_r216_c89 bl[89] br[89] wl[216] vdd gnd cell_6t
Xbit_r217_c89 bl[89] br[89] wl[217] vdd gnd cell_6t
Xbit_r218_c89 bl[89] br[89] wl[218] vdd gnd cell_6t
Xbit_r219_c89 bl[89] br[89] wl[219] vdd gnd cell_6t
Xbit_r220_c89 bl[89] br[89] wl[220] vdd gnd cell_6t
Xbit_r221_c89 bl[89] br[89] wl[221] vdd gnd cell_6t
Xbit_r222_c89 bl[89] br[89] wl[222] vdd gnd cell_6t
Xbit_r223_c89 bl[89] br[89] wl[223] vdd gnd cell_6t
Xbit_r224_c89 bl[89] br[89] wl[224] vdd gnd cell_6t
Xbit_r225_c89 bl[89] br[89] wl[225] vdd gnd cell_6t
Xbit_r226_c89 bl[89] br[89] wl[226] vdd gnd cell_6t
Xbit_r227_c89 bl[89] br[89] wl[227] vdd gnd cell_6t
Xbit_r228_c89 bl[89] br[89] wl[228] vdd gnd cell_6t
Xbit_r229_c89 bl[89] br[89] wl[229] vdd gnd cell_6t
Xbit_r230_c89 bl[89] br[89] wl[230] vdd gnd cell_6t
Xbit_r231_c89 bl[89] br[89] wl[231] vdd gnd cell_6t
Xbit_r232_c89 bl[89] br[89] wl[232] vdd gnd cell_6t
Xbit_r233_c89 bl[89] br[89] wl[233] vdd gnd cell_6t
Xbit_r234_c89 bl[89] br[89] wl[234] vdd gnd cell_6t
Xbit_r235_c89 bl[89] br[89] wl[235] vdd gnd cell_6t
Xbit_r236_c89 bl[89] br[89] wl[236] vdd gnd cell_6t
Xbit_r237_c89 bl[89] br[89] wl[237] vdd gnd cell_6t
Xbit_r238_c89 bl[89] br[89] wl[238] vdd gnd cell_6t
Xbit_r239_c89 bl[89] br[89] wl[239] vdd gnd cell_6t
Xbit_r240_c89 bl[89] br[89] wl[240] vdd gnd cell_6t
Xbit_r241_c89 bl[89] br[89] wl[241] vdd gnd cell_6t
Xbit_r242_c89 bl[89] br[89] wl[242] vdd gnd cell_6t
Xbit_r243_c89 bl[89] br[89] wl[243] vdd gnd cell_6t
Xbit_r244_c89 bl[89] br[89] wl[244] vdd gnd cell_6t
Xbit_r245_c89 bl[89] br[89] wl[245] vdd gnd cell_6t
Xbit_r246_c89 bl[89] br[89] wl[246] vdd gnd cell_6t
Xbit_r247_c89 bl[89] br[89] wl[247] vdd gnd cell_6t
Xbit_r248_c89 bl[89] br[89] wl[248] vdd gnd cell_6t
Xbit_r249_c89 bl[89] br[89] wl[249] vdd gnd cell_6t
Xbit_r250_c89 bl[89] br[89] wl[250] vdd gnd cell_6t
Xbit_r251_c89 bl[89] br[89] wl[251] vdd gnd cell_6t
Xbit_r252_c89 bl[89] br[89] wl[252] vdd gnd cell_6t
Xbit_r253_c89 bl[89] br[89] wl[253] vdd gnd cell_6t
Xbit_r254_c89 bl[89] br[89] wl[254] vdd gnd cell_6t
Xbit_r255_c89 bl[89] br[89] wl[255] vdd gnd cell_6t
Xbit_r0_c90 bl[90] br[90] wl[0] vdd gnd cell_6t
Xbit_r1_c90 bl[90] br[90] wl[1] vdd gnd cell_6t
Xbit_r2_c90 bl[90] br[90] wl[2] vdd gnd cell_6t
Xbit_r3_c90 bl[90] br[90] wl[3] vdd gnd cell_6t
Xbit_r4_c90 bl[90] br[90] wl[4] vdd gnd cell_6t
Xbit_r5_c90 bl[90] br[90] wl[5] vdd gnd cell_6t
Xbit_r6_c90 bl[90] br[90] wl[6] vdd gnd cell_6t
Xbit_r7_c90 bl[90] br[90] wl[7] vdd gnd cell_6t
Xbit_r8_c90 bl[90] br[90] wl[8] vdd gnd cell_6t
Xbit_r9_c90 bl[90] br[90] wl[9] vdd gnd cell_6t
Xbit_r10_c90 bl[90] br[90] wl[10] vdd gnd cell_6t
Xbit_r11_c90 bl[90] br[90] wl[11] vdd gnd cell_6t
Xbit_r12_c90 bl[90] br[90] wl[12] vdd gnd cell_6t
Xbit_r13_c90 bl[90] br[90] wl[13] vdd gnd cell_6t
Xbit_r14_c90 bl[90] br[90] wl[14] vdd gnd cell_6t
Xbit_r15_c90 bl[90] br[90] wl[15] vdd gnd cell_6t
Xbit_r16_c90 bl[90] br[90] wl[16] vdd gnd cell_6t
Xbit_r17_c90 bl[90] br[90] wl[17] vdd gnd cell_6t
Xbit_r18_c90 bl[90] br[90] wl[18] vdd gnd cell_6t
Xbit_r19_c90 bl[90] br[90] wl[19] vdd gnd cell_6t
Xbit_r20_c90 bl[90] br[90] wl[20] vdd gnd cell_6t
Xbit_r21_c90 bl[90] br[90] wl[21] vdd gnd cell_6t
Xbit_r22_c90 bl[90] br[90] wl[22] vdd gnd cell_6t
Xbit_r23_c90 bl[90] br[90] wl[23] vdd gnd cell_6t
Xbit_r24_c90 bl[90] br[90] wl[24] vdd gnd cell_6t
Xbit_r25_c90 bl[90] br[90] wl[25] vdd gnd cell_6t
Xbit_r26_c90 bl[90] br[90] wl[26] vdd gnd cell_6t
Xbit_r27_c90 bl[90] br[90] wl[27] vdd gnd cell_6t
Xbit_r28_c90 bl[90] br[90] wl[28] vdd gnd cell_6t
Xbit_r29_c90 bl[90] br[90] wl[29] vdd gnd cell_6t
Xbit_r30_c90 bl[90] br[90] wl[30] vdd gnd cell_6t
Xbit_r31_c90 bl[90] br[90] wl[31] vdd gnd cell_6t
Xbit_r32_c90 bl[90] br[90] wl[32] vdd gnd cell_6t
Xbit_r33_c90 bl[90] br[90] wl[33] vdd gnd cell_6t
Xbit_r34_c90 bl[90] br[90] wl[34] vdd gnd cell_6t
Xbit_r35_c90 bl[90] br[90] wl[35] vdd gnd cell_6t
Xbit_r36_c90 bl[90] br[90] wl[36] vdd gnd cell_6t
Xbit_r37_c90 bl[90] br[90] wl[37] vdd gnd cell_6t
Xbit_r38_c90 bl[90] br[90] wl[38] vdd gnd cell_6t
Xbit_r39_c90 bl[90] br[90] wl[39] vdd gnd cell_6t
Xbit_r40_c90 bl[90] br[90] wl[40] vdd gnd cell_6t
Xbit_r41_c90 bl[90] br[90] wl[41] vdd gnd cell_6t
Xbit_r42_c90 bl[90] br[90] wl[42] vdd gnd cell_6t
Xbit_r43_c90 bl[90] br[90] wl[43] vdd gnd cell_6t
Xbit_r44_c90 bl[90] br[90] wl[44] vdd gnd cell_6t
Xbit_r45_c90 bl[90] br[90] wl[45] vdd gnd cell_6t
Xbit_r46_c90 bl[90] br[90] wl[46] vdd gnd cell_6t
Xbit_r47_c90 bl[90] br[90] wl[47] vdd gnd cell_6t
Xbit_r48_c90 bl[90] br[90] wl[48] vdd gnd cell_6t
Xbit_r49_c90 bl[90] br[90] wl[49] vdd gnd cell_6t
Xbit_r50_c90 bl[90] br[90] wl[50] vdd gnd cell_6t
Xbit_r51_c90 bl[90] br[90] wl[51] vdd gnd cell_6t
Xbit_r52_c90 bl[90] br[90] wl[52] vdd gnd cell_6t
Xbit_r53_c90 bl[90] br[90] wl[53] vdd gnd cell_6t
Xbit_r54_c90 bl[90] br[90] wl[54] vdd gnd cell_6t
Xbit_r55_c90 bl[90] br[90] wl[55] vdd gnd cell_6t
Xbit_r56_c90 bl[90] br[90] wl[56] vdd gnd cell_6t
Xbit_r57_c90 bl[90] br[90] wl[57] vdd gnd cell_6t
Xbit_r58_c90 bl[90] br[90] wl[58] vdd gnd cell_6t
Xbit_r59_c90 bl[90] br[90] wl[59] vdd gnd cell_6t
Xbit_r60_c90 bl[90] br[90] wl[60] vdd gnd cell_6t
Xbit_r61_c90 bl[90] br[90] wl[61] vdd gnd cell_6t
Xbit_r62_c90 bl[90] br[90] wl[62] vdd gnd cell_6t
Xbit_r63_c90 bl[90] br[90] wl[63] vdd gnd cell_6t
Xbit_r64_c90 bl[90] br[90] wl[64] vdd gnd cell_6t
Xbit_r65_c90 bl[90] br[90] wl[65] vdd gnd cell_6t
Xbit_r66_c90 bl[90] br[90] wl[66] vdd gnd cell_6t
Xbit_r67_c90 bl[90] br[90] wl[67] vdd gnd cell_6t
Xbit_r68_c90 bl[90] br[90] wl[68] vdd gnd cell_6t
Xbit_r69_c90 bl[90] br[90] wl[69] vdd gnd cell_6t
Xbit_r70_c90 bl[90] br[90] wl[70] vdd gnd cell_6t
Xbit_r71_c90 bl[90] br[90] wl[71] vdd gnd cell_6t
Xbit_r72_c90 bl[90] br[90] wl[72] vdd gnd cell_6t
Xbit_r73_c90 bl[90] br[90] wl[73] vdd gnd cell_6t
Xbit_r74_c90 bl[90] br[90] wl[74] vdd gnd cell_6t
Xbit_r75_c90 bl[90] br[90] wl[75] vdd gnd cell_6t
Xbit_r76_c90 bl[90] br[90] wl[76] vdd gnd cell_6t
Xbit_r77_c90 bl[90] br[90] wl[77] vdd gnd cell_6t
Xbit_r78_c90 bl[90] br[90] wl[78] vdd gnd cell_6t
Xbit_r79_c90 bl[90] br[90] wl[79] vdd gnd cell_6t
Xbit_r80_c90 bl[90] br[90] wl[80] vdd gnd cell_6t
Xbit_r81_c90 bl[90] br[90] wl[81] vdd gnd cell_6t
Xbit_r82_c90 bl[90] br[90] wl[82] vdd gnd cell_6t
Xbit_r83_c90 bl[90] br[90] wl[83] vdd gnd cell_6t
Xbit_r84_c90 bl[90] br[90] wl[84] vdd gnd cell_6t
Xbit_r85_c90 bl[90] br[90] wl[85] vdd gnd cell_6t
Xbit_r86_c90 bl[90] br[90] wl[86] vdd gnd cell_6t
Xbit_r87_c90 bl[90] br[90] wl[87] vdd gnd cell_6t
Xbit_r88_c90 bl[90] br[90] wl[88] vdd gnd cell_6t
Xbit_r89_c90 bl[90] br[90] wl[89] vdd gnd cell_6t
Xbit_r90_c90 bl[90] br[90] wl[90] vdd gnd cell_6t
Xbit_r91_c90 bl[90] br[90] wl[91] vdd gnd cell_6t
Xbit_r92_c90 bl[90] br[90] wl[92] vdd gnd cell_6t
Xbit_r93_c90 bl[90] br[90] wl[93] vdd gnd cell_6t
Xbit_r94_c90 bl[90] br[90] wl[94] vdd gnd cell_6t
Xbit_r95_c90 bl[90] br[90] wl[95] vdd gnd cell_6t
Xbit_r96_c90 bl[90] br[90] wl[96] vdd gnd cell_6t
Xbit_r97_c90 bl[90] br[90] wl[97] vdd gnd cell_6t
Xbit_r98_c90 bl[90] br[90] wl[98] vdd gnd cell_6t
Xbit_r99_c90 bl[90] br[90] wl[99] vdd gnd cell_6t
Xbit_r100_c90 bl[90] br[90] wl[100] vdd gnd cell_6t
Xbit_r101_c90 bl[90] br[90] wl[101] vdd gnd cell_6t
Xbit_r102_c90 bl[90] br[90] wl[102] vdd gnd cell_6t
Xbit_r103_c90 bl[90] br[90] wl[103] vdd gnd cell_6t
Xbit_r104_c90 bl[90] br[90] wl[104] vdd gnd cell_6t
Xbit_r105_c90 bl[90] br[90] wl[105] vdd gnd cell_6t
Xbit_r106_c90 bl[90] br[90] wl[106] vdd gnd cell_6t
Xbit_r107_c90 bl[90] br[90] wl[107] vdd gnd cell_6t
Xbit_r108_c90 bl[90] br[90] wl[108] vdd gnd cell_6t
Xbit_r109_c90 bl[90] br[90] wl[109] vdd gnd cell_6t
Xbit_r110_c90 bl[90] br[90] wl[110] vdd gnd cell_6t
Xbit_r111_c90 bl[90] br[90] wl[111] vdd gnd cell_6t
Xbit_r112_c90 bl[90] br[90] wl[112] vdd gnd cell_6t
Xbit_r113_c90 bl[90] br[90] wl[113] vdd gnd cell_6t
Xbit_r114_c90 bl[90] br[90] wl[114] vdd gnd cell_6t
Xbit_r115_c90 bl[90] br[90] wl[115] vdd gnd cell_6t
Xbit_r116_c90 bl[90] br[90] wl[116] vdd gnd cell_6t
Xbit_r117_c90 bl[90] br[90] wl[117] vdd gnd cell_6t
Xbit_r118_c90 bl[90] br[90] wl[118] vdd gnd cell_6t
Xbit_r119_c90 bl[90] br[90] wl[119] vdd gnd cell_6t
Xbit_r120_c90 bl[90] br[90] wl[120] vdd gnd cell_6t
Xbit_r121_c90 bl[90] br[90] wl[121] vdd gnd cell_6t
Xbit_r122_c90 bl[90] br[90] wl[122] vdd gnd cell_6t
Xbit_r123_c90 bl[90] br[90] wl[123] vdd gnd cell_6t
Xbit_r124_c90 bl[90] br[90] wl[124] vdd gnd cell_6t
Xbit_r125_c90 bl[90] br[90] wl[125] vdd gnd cell_6t
Xbit_r126_c90 bl[90] br[90] wl[126] vdd gnd cell_6t
Xbit_r127_c90 bl[90] br[90] wl[127] vdd gnd cell_6t
Xbit_r128_c90 bl[90] br[90] wl[128] vdd gnd cell_6t
Xbit_r129_c90 bl[90] br[90] wl[129] vdd gnd cell_6t
Xbit_r130_c90 bl[90] br[90] wl[130] vdd gnd cell_6t
Xbit_r131_c90 bl[90] br[90] wl[131] vdd gnd cell_6t
Xbit_r132_c90 bl[90] br[90] wl[132] vdd gnd cell_6t
Xbit_r133_c90 bl[90] br[90] wl[133] vdd gnd cell_6t
Xbit_r134_c90 bl[90] br[90] wl[134] vdd gnd cell_6t
Xbit_r135_c90 bl[90] br[90] wl[135] vdd gnd cell_6t
Xbit_r136_c90 bl[90] br[90] wl[136] vdd gnd cell_6t
Xbit_r137_c90 bl[90] br[90] wl[137] vdd gnd cell_6t
Xbit_r138_c90 bl[90] br[90] wl[138] vdd gnd cell_6t
Xbit_r139_c90 bl[90] br[90] wl[139] vdd gnd cell_6t
Xbit_r140_c90 bl[90] br[90] wl[140] vdd gnd cell_6t
Xbit_r141_c90 bl[90] br[90] wl[141] vdd gnd cell_6t
Xbit_r142_c90 bl[90] br[90] wl[142] vdd gnd cell_6t
Xbit_r143_c90 bl[90] br[90] wl[143] vdd gnd cell_6t
Xbit_r144_c90 bl[90] br[90] wl[144] vdd gnd cell_6t
Xbit_r145_c90 bl[90] br[90] wl[145] vdd gnd cell_6t
Xbit_r146_c90 bl[90] br[90] wl[146] vdd gnd cell_6t
Xbit_r147_c90 bl[90] br[90] wl[147] vdd gnd cell_6t
Xbit_r148_c90 bl[90] br[90] wl[148] vdd gnd cell_6t
Xbit_r149_c90 bl[90] br[90] wl[149] vdd gnd cell_6t
Xbit_r150_c90 bl[90] br[90] wl[150] vdd gnd cell_6t
Xbit_r151_c90 bl[90] br[90] wl[151] vdd gnd cell_6t
Xbit_r152_c90 bl[90] br[90] wl[152] vdd gnd cell_6t
Xbit_r153_c90 bl[90] br[90] wl[153] vdd gnd cell_6t
Xbit_r154_c90 bl[90] br[90] wl[154] vdd gnd cell_6t
Xbit_r155_c90 bl[90] br[90] wl[155] vdd gnd cell_6t
Xbit_r156_c90 bl[90] br[90] wl[156] vdd gnd cell_6t
Xbit_r157_c90 bl[90] br[90] wl[157] vdd gnd cell_6t
Xbit_r158_c90 bl[90] br[90] wl[158] vdd gnd cell_6t
Xbit_r159_c90 bl[90] br[90] wl[159] vdd gnd cell_6t
Xbit_r160_c90 bl[90] br[90] wl[160] vdd gnd cell_6t
Xbit_r161_c90 bl[90] br[90] wl[161] vdd gnd cell_6t
Xbit_r162_c90 bl[90] br[90] wl[162] vdd gnd cell_6t
Xbit_r163_c90 bl[90] br[90] wl[163] vdd gnd cell_6t
Xbit_r164_c90 bl[90] br[90] wl[164] vdd gnd cell_6t
Xbit_r165_c90 bl[90] br[90] wl[165] vdd gnd cell_6t
Xbit_r166_c90 bl[90] br[90] wl[166] vdd gnd cell_6t
Xbit_r167_c90 bl[90] br[90] wl[167] vdd gnd cell_6t
Xbit_r168_c90 bl[90] br[90] wl[168] vdd gnd cell_6t
Xbit_r169_c90 bl[90] br[90] wl[169] vdd gnd cell_6t
Xbit_r170_c90 bl[90] br[90] wl[170] vdd gnd cell_6t
Xbit_r171_c90 bl[90] br[90] wl[171] vdd gnd cell_6t
Xbit_r172_c90 bl[90] br[90] wl[172] vdd gnd cell_6t
Xbit_r173_c90 bl[90] br[90] wl[173] vdd gnd cell_6t
Xbit_r174_c90 bl[90] br[90] wl[174] vdd gnd cell_6t
Xbit_r175_c90 bl[90] br[90] wl[175] vdd gnd cell_6t
Xbit_r176_c90 bl[90] br[90] wl[176] vdd gnd cell_6t
Xbit_r177_c90 bl[90] br[90] wl[177] vdd gnd cell_6t
Xbit_r178_c90 bl[90] br[90] wl[178] vdd gnd cell_6t
Xbit_r179_c90 bl[90] br[90] wl[179] vdd gnd cell_6t
Xbit_r180_c90 bl[90] br[90] wl[180] vdd gnd cell_6t
Xbit_r181_c90 bl[90] br[90] wl[181] vdd gnd cell_6t
Xbit_r182_c90 bl[90] br[90] wl[182] vdd gnd cell_6t
Xbit_r183_c90 bl[90] br[90] wl[183] vdd gnd cell_6t
Xbit_r184_c90 bl[90] br[90] wl[184] vdd gnd cell_6t
Xbit_r185_c90 bl[90] br[90] wl[185] vdd gnd cell_6t
Xbit_r186_c90 bl[90] br[90] wl[186] vdd gnd cell_6t
Xbit_r187_c90 bl[90] br[90] wl[187] vdd gnd cell_6t
Xbit_r188_c90 bl[90] br[90] wl[188] vdd gnd cell_6t
Xbit_r189_c90 bl[90] br[90] wl[189] vdd gnd cell_6t
Xbit_r190_c90 bl[90] br[90] wl[190] vdd gnd cell_6t
Xbit_r191_c90 bl[90] br[90] wl[191] vdd gnd cell_6t
Xbit_r192_c90 bl[90] br[90] wl[192] vdd gnd cell_6t
Xbit_r193_c90 bl[90] br[90] wl[193] vdd gnd cell_6t
Xbit_r194_c90 bl[90] br[90] wl[194] vdd gnd cell_6t
Xbit_r195_c90 bl[90] br[90] wl[195] vdd gnd cell_6t
Xbit_r196_c90 bl[90] br[90] wl[196] vdd gnd cell_6t
Xbit_r197_c90 bl[90] br[90] wl[197] vdd gnd cell_6t
Xbit_r198_c90 bl[90] br[90] wl[198] vdd gnd cell_6t
Xbit_r199_c90 bl[90] br[90] wl[199] vdd gnd cell_6t
Xbit_r200_c90 bl[90] br[90] wl[200] vdd gnd cell_6t
Xbit_r201_c90 bl[90] br[90] wl[201] vdd gnd cell_6t
Xbit_r202_c90 bl[90] br[90] wl[202] vdd gnd cell_6t
Xbit_r203_c90 bl[90] br[90] wl[203] vdd gnd cell_6t
Xbit_r204_c90 bl[90] br[90] wl[204] vdd gnd cell_6t
Xbit_r205_c90 bl[90] br[90] wl[205] vdd gnd cell_6t
Xbit_r206_c90 bl[90] br[90] wl[206] vdd gnd cell_6t
Xbit_r207_c90 bl[90] br[90] wl[207] vdd gnd cell_6t
Xbit_r208_c90 bl[90] br[90] wl[208] vdd gnd cell_6t
Xbit_r209_c90 bl[90] br[90] wl[209] vdd gnd cell_6t
Xbit_r210_c90 bl[90] br[90] wl[210] vdd gnd cell_6t
Xbit_r211_c90 bl[90] br[90] wl[211] vdd gnd cell_6t
Xbit_r212_c90 bl[90] br[90] wl[212] vdd gnd cell_6t
Xbit_r213_c90 bl[90] br[90] wl[213] vdd gnd cell_6t
Xbit_r214_c90 bl[90] br[90] wl[214] vdd gnd cell_6t
Xbit_r215_c90 bl[90] br[90] wl[215] vdd gnd cell_6t
Xbit_r216_c90 bl[90] br[90] wl[216] vdd gnd cell_6t
Xbit_r217_c90 bl[90] br[90] wl[217] vdd gnd cell_6t
Xbit_r218_c90 bl[90] br[90] wl[218] vdd gnd cell_6t
Xbit_r219_c90 bl[90] br[90] wl[219] vdd gnd cell_6t
Xbit_r220_c90 bl[90] br[90] wl[220] vdd gnd cell_6t
Xbit_r221_c90 bl[90] br[90] wl[221] vdd gnd cell_6t
Xbit_r222_c90 bl[90] br[90] wl[222] vdd gnd cell_6t
Xbit_r223_c90 bl[90] br[90] wl[223] vdd gnd cell_6t
Xbit_r224_c90 bl[90] br[90] wl[224] vdd gnd cell_6t
Xbit_r225_c90 bl[90] br[90] wl[225] vdd gnd cell_6t
Xbit_r226_c90 bl[90] br[90] wl[226] vdd gnd cell_6t
Xbit_r227_c90 bl[90] br[90] wl[227] vdd gnd cell_6t
Xbit_r228_c90 bl[90] br[90] wl[228] vdd gnd cell_6t
Xbit_r229_c90 bl[90] br[90] wl[229] vdd gnd cell_6t
Xbit_r230_c90 bl[90] br[90] wl[230] vdd gnd cell_6t
Xbit_r231_c90 bl[90] br[90] wl[231] vdd gnd cell_6t
Xbit_r232_c90 bl[90] br[90] wl[232] vdd gnd cell_6t
Xbit_r233_c90 bl[90] br[90] wl[233] vdd gnd cell_6t
Xbit_r234_c90 bl[90] br[90] wl[234] vdd gnd cell_6t
Xbit_r235_c90 bl[90] br[90] wl[235] vdd gnd cell_6t
Xbit_r236_c90 bl[90] br[90] wl[236] vdd gnd cell_6t
Xbit_r237_c90 bl[90] br[90] wl[237] vdd gnd cell_6t
Xbit_r238_c90 bl[90] br[90] wl[238] vdd gnd cell_6t
Xbit_r239_c90 bl[90] br[90] wl[239] vdd gnd cell_6t
Xbit_r240_c90 bl[90] br[90] wl[240] vdd gnd cell_6t
Xbit_r241_c90 bl[90] br[90] wl[241] vdd gnd cell_6t
Xbit_r242_c90 bl[90] br[90] wl[242] vdd gnd cell_6t
Xbit_r243_c90 bl[90] br[90] wl[243] vdd gnd cell_6t
Xbit_r244_c90 bl[90] br[90] wl[244] vdd gnd cell_6t
Xbit_r245_c90 bl[90] br[90] wl[245] vdd gnd cell_6t
Xbit_r246_c90 bl[90] br[90] wl[246] vdd gnd cell_6t
Xbit_r247_c90 bl[90] br[90] wl[247] vdd gnd cell_6t
Xbit_r248_c90 bl[90] br[90] wl[248] vdd gnd cell_6t
Xbit_r249_c90 bl[90] br[90] wl[249] vdd gnd cell_6t
Xbit_r250_c90 bl[90] br[90] wl[250] vdd gnd cell_6t
Xbit_r251_c90 bl[90] br[90] wl[251] vdd gnd cell_6t
Xbit_r252_c90 bl[90] br[90] wl[252] vdd gnd cell_6t
Xbit_r253_c90 bl[90] br[90] wl[253] vdd gnd cell_6t
Xbit_r254_c90 bl[90] br[90] wl[254] vdd gnd cell_6t
Xbit_r255_c90 bl[90] br[90] wl[255] vdd gnd cell_6t
Xbit_r0_c91 bl[91] br[91] wl[0] vdd gnd cell_6t
Xbit_r1_c91 bl[91] br[91] wl[1] vdd gnd cell_6t
Xbit_r2_c91 bl[91] br[91] wl[2] vdd gnd cell_6t
Xbit_r3_c91 bl[91] br[91] wl[3] vdd gnd cell_6t
Xbit_r4_c91 bl[91] br[91] wl[4] vdd gnd cell_6t
Xbit_r5_c91 bl[91] br[91] wl[5] vdd gnd cell_6t
Xbit_r6_c91 bl[91] br[91] wl[6] vdd gnd cell_6t
Xbit_r7_c91 bl[91] br[91] wl[7] vdd gnd cell_6t
Xbit_r8_c91 bl[91] br[91] wl[8] vdd gnd cell_6t
Xbit_r9_c91 bl[91] br[91] wl[9] vdd gnd cell_6t
Xbit_r10_c91 bl[91] br[91] wl[10] vdd gnd cell_6t
Xbit_r11_c91 bl[91] br[91] wl[11] vdd gnd cell_6t
Xbit_r12_c91 bl[91] br[91] wl[12] vdd gnd cell_6t
Xbit_r13_c91 bl[91] br[91] wl[13] vdd gnd cell_6t
Xbit_r14_c91 bl[91] br[91] wl[14] vdd gnd cell_6t
Xbit_r15_c91 bl[91] br[91] wl[15] vdd gnd cell_6t
Xbit_r16_c91 bl[91] br[91] wl[16] vdd gnd cell_6t
Xbit_r17_c91 bl[91] br[91] wl[17] vdd gnd cell_6t
Xbit_r18_c91 bl[91] br[91] wl[18] vdd gnd cell_6t
Xbit_r19_c91 bl[91] br[91] wl[19] vdd gnd cell_6t
Xbit_r20_c91 bl[91] br[91] wl[20] vdd gnd cell_6t
Xbit_r21_c91 bl[91] br[91] wl[21] vdd gnd cell_6t
Xbit_r22_c91 bl[91] br[91] wl[22] vdd gnd cell_6t
Xbit_r23_c91 bl[91] br[91] wl[23] vdd gnd cell_6t
Xbit_r24_c91 bl[91] br[91] wl[24] vdd gnd cell_6t
Xbit_r25_c91 bl[91] br[91] wl[25] vdd gnd cell_6t
Xbit_r26_c91 bl[91] br[91] wl[26] vdd gnd cell_6t
Xbit_r27_c91 bl[91] br[91] wl[27] vdd gnd cell_6t
Xbit_r28_c91 bl[91] br[91] wl[28] vdd gnd cell_6t
Xbit_r29_c91 bl[91] br[91] wl[29] vdd gnd cell_6t
Xbit_r30_c91 bl[91] br[91] wl[30] vdd gnd cell_6t
Xbit_r31_c91 bl[91] br[91] wl[31] vdd gnd cell_6t
Xbit_r32_c91 bl[91] br[91] wl[32] vdd gnd cell_6t
Xbit_r33_c91 bl[91] br[91] wl[33] vdd gnd cell_6t
Xbit_r34_c91 bl[91] br[91] wl[34] vdd gnd cell_6t
Xbit_r35_c91 bl[91] br[91] wl[35] vdd gnd cell_6t
Xbit_r36_c91 bl[91] br[91] wl[36] vdd gnd cell_6t
Xbit_r37_c91 bl[91] br[91] wl[37] vdd gnd cell_6t
Xbit_r38_c91 bl[91] br[91] wl[38] vdd gnd cell_6t
Xbit_r39_c91 bl[91] br[91] wl[39] vdd gnd cell_6t
Xbit_r40_c91 bl[91] br[91] wl[40] vdd gnd cell_6t
Xbit_r41_c91 bl[91] br[91] wl[41] vdd gnd cell_6t
Xbit_r42_c91 bl[91] br[91] wl[42] vdd gnd cell_6t
Xbit_r43_c91 bl[91] br[91] wl[43] vdd gnd cell_6t
Xbit_r44_c91 bl[91] br[91] wl[44] vdd gnd cell_6t
Xbit_r45_c91 bl[91] br[91] wl[45] vdd gnd cell_6t
Xbit_r46_c91 bl[91] br[91] wl[46] vdd gnd cell_6t
Xbit_r47_c91 bl[91] br[91] wl[47] vdd gnd cell_6t
Xbit_r48_c91 bl[91] br[91] wl[48] vdd gnd cell_6t
Xbit_r49_c91 bl[91] br[91] wl[49] vdd gnd cell_6t
Xbit_r50_c91 bl[91] br[91] wl[50] vdd gnd cell_6t
Xbit_r51_c91 bl[91] br[91] wl[51] vdd gnd cell_6t
Xbit_r52_c91 bl[91] br[91] wl[52] vdd gnd cell_6t
Xbit_r53_c91 bl[91] br[91] wl[53] vdd gnd cell_6t
Xbit_r54_c91 bl[91] br[91] wl[54] vdd gnd cell_6t
Xbit_r55_c91 bl[91] br[91] wl[55] vdd gnd cell_6t
Xbit_r56_c91 bl[91] br[91] wl[56] vdd gnd cell_6t
Xbit_r57_c91 bl[91] br[91] wl[57] vdd gnd cell_6t
Xbit_r58_c91 bl[91] br[91] wl[58] vdd gnd cell_6t
Xbit_r59_c91 bl[91] br[91] wl[59] vdd gnd cell_6t
Xbit_r60_c91 bl[91] br[91] wl[60] vdd gnd cell_6t
Xbit_r61_c91 bl[91] br[91] wl[61] vdd gnd cell_6t
Xbit_r62_c91 bl[91] br[91] wl[62] vdd gnd cell_6t
Xbit_r63_c91 bl[91] br[91] wl[63] vdd gnd cell_6t
Xbit_r64_c91 bl[91] br[91] wl[64] vdd gnd cell_6t
Xbit_r65_c91 bl[91] br[91] wl[65] vdd gnd cell_6t
Xbit_r66_c91 bl[91] br[91] wl[66] vdd gnd cell_6t
Xbit_r67_c91 bl[91] br[91] wl[67] vdd gnd cell_6t
Xbit_r68_c91 bl[91] br[91] wl[68] vdd gnd cell_6t
Xbit_r69_c91 bl[91] br[91] wl[69] vdd gnd cell_6t
Xbit_r70_c91 bl[91] br[91] wl[70] vdd gnd cell_6t
Xbit_r71_c91 bl[91] br[91] wl[71] vdd gnd cell_6t
Xbit_r72_c91 bl[91] br[91] wl[72] vdd gnd cell_6t
Xbit_r73_c91 bl[91] br[91] wl[73] vdd gnd cell_6t
Xbit_r74_c91 bl[91] br[91] wl[74] vdd gnd cell_6t
Xbit_r75_c91 bl[91] br[91] wl[75] vdd gnd cell_6t
Xbit_r76_c91 bl[91] br[91] wl[76] vdd gnd cell_6t
Xbit_r77_c91 bl[91] br[91] wl[77] vdd gnd cell_6t
Xbit_r78_c91 bl[91] br[91] wl[78] vdd gnd cell_6t
Xbit_r79_c91 bl[91] br[91] wl[79] vdd gnd cell_6t
Xbit_r80_c91 bl[91] br[91] wl[80] vdd gnd cell_6t
Xbit_r81_c91 bl[91] br[91] wl[81] vdd gnd cell_6t
Xbit_r82_c91 bl[91] br[91] wl[82] vdd gnd cell_6t
Xbit_r83_c91 bl[91] br[91] wl[83] vdd gnd cell_6t
Xbit_r84_c91 bl[91] br[91] wl[84] vdd gnd cell_6t
Xbit_r85_c91 bl[91] br[91] wl[85] vdd gnd cell_6t
Xbit_r86_c91 bl[91] br[91] wl[86] vdd gnd cell_6t
Xbit_r87_c91 bl[91] br[91] wl[87] vdd gnd cell_6t
Xbit_r88_c91 bl[91] br[91] wl[88] vdd gnd cell_6t
Xbit_r89_c91 bl[91] br[91] wl[89] vdd gnd cell_6t
Xbit_r90_c91 bl[91] br[91] wl[90] vdd gnd cell_6t
Xbit_r91_c91 bl[91] br[91] wl[91] vdd gnd cell_6t
Xbit_r92_c91 bl[91] br[91] wl[92] vdd gnd cell_6t
Xbit_r93_c91 bl[91] br[91] wl[93] vdd gnd cell_6t
Xbit_r94_c91 bl[91] br[91] wl[94] vdd gnd cell_6t
Xbit_r95_c91 bl[91] br[91] wl[95] vdd gnd cell_6t
Xbit_r96_c91 bl[91] br[91] wl[96] vdd gnd cell_6t
Xbit_r97_c91 bl[91] br[91] wl[97] vdd gnd cell_6t
Xbit_r98_c91 bl[91] br[91] wl[98] vdd gnd cell_6t
Xbit_r99_c91 bl[91] br[91] wl[99] vdd gnd cell_6t
Xbit_r100_c91 bl[91] br[91] wl[100] vdd gnd cell_6t
Xbit_r101_c91 bl[91] br[91] wl[101] vdd gnd cell_6t
Xbit_r102_c91 bl[91] br[91] wl[102] vdd gnd cell_6t
Xbit_r103_c91 bl[91] br[91] wl[103] vdd gnd cell_6t
Xbit_r104_c91 bl[91] br[91] wl[104] vdd gnd cell_6t
Xbit_r105_c91 bl[91] br[91] wl[105] vdd gnd cell_6t
Xbit_r106_c91 bl[91] br[91] wl[106] vdd gnd cell_6t
Xbit_r107_c91 bl[91] br[91] wl[107] vdd gnd cell_6t
Xbit_r108_c91 bl[91] br[91] wl[108] vdd gnd cell_6t
Xbit_r109_c91 bl[91] br[91] wl[109] vdd gnd cell_6t
Xbit_r110_c91 bl[91] br[91] wl[110] vdd gnd cell_6t
Xbit_r111_c91 bl[91] br[91] wl[111] vdd gnd cell_6t
Xbit_r112_c91 bl[91] br[91] wl[112] vdd gnd cell_6t
Xbit_r113_c91 bl[91] br[91] wl[113] vdd gnd cell_6t
Xbit_r114_c91 bl[91] br[91] wl[114] vdd gnd cell_6t
Xbit_r115_c91 bl[91] br[91] wl[115] vdd gnd cell_6t
Xbit_r116_c91 bl[91] br[91] wl[116] vdd gnd cell_6t
Xbit_r117_c91 bl[91] br[91] wl[117] vdd gnd cell_6t
Xbit_r118_c91 bl[91] br[91] wl[118] vdd gnd cell_6t
Xbit_r119_c91 bl[91] br[91] wl[119] vdd gnd cell_6t
Xbit_r120_c91 bl[91] br[91] wl[120] vdd gnd cell_6t
Xbit_r121_c91 bl[91] br[91] wl[121] vdd gnd cell_6t
Xbit_r122_c91 bl[91] br[91] wl[122] vdd gnd cell_6t
Xbit_r123_c91 bl[91] br[91] wl[123] vdd gnd cell_6t
Xbit_r124_c91 bl[91] br[91] wl[124] vdd gnd cell_6t
Xbit_r125_c91 bl[91] br[91] wl[125] vdd gnd cell_6t
Xbit_r126_c91 bl[91] br[91] wl[126] vdd gnd cell_6t
Xbit_r127_c91 bl[91] br[91] wl[127] vdd gnd cell_6t
Xbit_r128_c91 bl[91] br[91] wl[128] vdd gnd cell_6t
Xbit_r129_c91 bl[91] br[91] wl[129] vdd gnd cell_6t
Xbit_r130_c91 bl[91] br[91] wl[130] vdd gnd cell_6t
Xbit_r131_c91 bl[91] br[91] wl[131] vdd gnd cell_6t
Xbit_r132_c91 bl[91] br[91] wl[132] vdd gnd cell_6t
Xbit_r133_c91 bl[91] br[91] wl[133] vdd gnd cell_6t
Xbit_r134_c91 bl[91] br[91] wl[134] vdd gnd cell_6t
Xbit_r135_c91 bl[91] br[91] wl[135] vdd gnd cell_6t
Xbit_r136_c91 bl[91] br[91] wl[136] vdd gnd cell_6t
Xbit_r137_c91 bl[91] br[91] wl[137] vdd gnd cell_6t
Xbit_r138_c91 bl[91] br[91] wl[138] vdd gnd cell_6t
Xbit_r139_c91 bl[91] br[91] wl[139] vdd gnd cell_6t
Xbit_r140_c91 bl[91] br[91] wl[140] vdd gnd cell_6t
Xbit_r141_c91 bl[91] br[91] wl[141] vdd gnd cell_6t
Xbit_r142_c91 bl[91] br[91] wl[142] vdd gnd cell_6t
Xbit_r143_c91 bl[91] br[91] wl[143] vdd gnd cell_6t
Xbit_r144_c91 bl[91] br[91] wl[144] vdd gnd cell_6t
Xbit_r145_c91 bl[91] br[91] wl[145] vdd gnd cell_6t
Xbit_r146_c91 bl[91] br[91] wl[146] vdd gnd cell_6t
Xbit_r147_c91 bl[91] br[91] wl[147] vdd gnd cell_6t
Xbit_r148_c91 bl[91] br[91] wl[148] vdd gnd cell_6t
Xbit_r149_c91 bl[91] br[91] wl[149] vdd gnd cell_6t
Xbit_r150_c91 bl[91] br[91] wl[150] vdd gnd cell_6t
Xbit_r151_c91 bl[91] br[91] wl[151] vdd gnd cell_6t
Xbit_r152_c91 bl[91] br[91] wl[152] vdd gnd cell_6t
Xbit_r153_c91 bl[91] br[91] wl[153] vdd gnd cell_6t
Xbit_r154_c91 bl[91] br[91] wl[154] vdd gnd cell_6t
Xbit_r155_c91 bl[91] br[91] wl[155] vdd gnd cell_6t
Xbit_r156_c91 bl[91] br[91] wl[156] vdd gnd cell_6t
Xbit_r157_c91 bl[91] br[91] wl[157] vdd gnd cell_6t
Xbit_r158_c91 bl[91] br[91] wl[158] vdd gnd cell_6t
Xbit_r159_c91 bl[91] br[91] wl[159] vdd gnd cell_6t
Xbit_r160_c91 bl[91] br[91] wl[160] vdd gnd cell_6t
Xbit_r161_c91 bl[91] br[91] wl[161] vdd gnd cell_6t
Xbit_r162_c91 bl[91] br[91] wl[162] vdd gnd cell_6t
Xbit_r163_c91 bl[91] br[91] wl[163] vdd gnd cell_6t
Xbit_r164_c91 bl[91] br[91] wl[164] vdd gnd cell_6t
Xbit_r165_c91 bl[91] br[91] wl[165] vdd gnd cell_6t
Xbit_r166_c91 bl[91] br[91] wl[166] vdd gnd cell_6t
Xbit_r167_c91 bl[91] br[91] wl[167] vdd gnd cell_6t
Xbit_r168_c91 bl[91] br[91] wl[168] vdd gnd cell_6t
Xbit_r169_c91 bl[91] br[91] wl[169] vdd gnd cell_6t
Xbit_r170_c91 bl[91] br[91] wl[170] vdd gnd cell_6t
Xbit_r171_c91 bl[91] br[91] wl[171] vdd gnd cell_6t
Xbit_r172_c91 bl[91] br[91] wl[172] vdd gnd cell_6t
Xbit_r173_c91 bl[91] br[91] wl[173] vdd gnd cell_6t
Xbit_r174_c91 bl[91] br[91] wl[174] vdd gnd cell_6t
Xbit_r175_c91 bl[91] br[91] wl[175] vdd gnd cell_6t
Xbit_r176_c91 bl[91] br[91] wl[176] vdd gnd cell_6t
Xbit_r177_c91 bl[91] br[91] wl[177] vdd gnd cell_6t
Xbit_r178_c91 bl[91] br[91] wl[178] vdd gnd cell_6t
Xbit_r179_c91 bl[91] br[91] wl[179] vdd gnd cell_6t
Xbit_r180_c91 bl[91] br[91] wl[180] vdd gnd cell_6t
Xbit_r181_c91 bl[91] br[91] wl[181] vdd gnd cell_6t
Xbit_r182_c91 bl[91] br[91] wl[182] vdd gnd cell_6t
Xbit_r183_c91 bl[91] br[91] wl[183] vdd gnd cell_6t
Xbit_r184_c91 bl[91] br[91] wl[184] vdd gnd cell_6t
Xbit_r185_c91 bl[91] br[91] wl[185] vdd gnd cell_6t
Xbit_r186_c91 bl[91] br[91] wl[186] vdd gnd cell_6t
Xbit_r187_c91 bl[91] br[91] wl[187] vdd gnd cell_6t
Xbit_r188_c91 bl[91] br[91] wl[188] vdd gnd cell_6t
Xbit_r189_c91 bl[91] br[91] wl[189] vdd gnd cell_6t
Xbit_r190_c91 bl[91] br[91] wl[190] vdd gnd cell_6t
Xbit_r191_c91 bl[91] br[91] wl[191] vdd gnd cell_6t
Xbit_r192_c91 bl[91] br[91] wl[192] vdd gnd cell_6t
Xbit_r193_c91 bl[91] br[91] wl[193] vdd gnd cell_6t
Xbit_r194_c91 bl[91] br[91] wl[194] vdd gnd cell_6t
Xbit_r195_c91 bl[91] br[91] wl[195] vdd gnd cell_6t
Xbit_r196_c91 bl[91] br[91] wl[196] vdd gnd cell_6t
Xbit_r197_c91 bl[91] br[91] wl[197] vdd gnd cell_6t
Xbit_r198_c91 bl[91] br[91] wl[198] vdd gnd cell_6t
Xbit_r199_c91 bl[91] br[91] wl[199] vdd gnd cell_6t
Xbit_r200_c91 bl[91] br[91] wl[200] vdd gnd cell_6t
Xbit_r201_c91 bl[91] br[91] wl[201] vdd gnd cell_6t
Xbit_r202_c91 bl[91] br[91] wl[202] vdd gnd cell_6t
Xbit_r203_c91 bl[91] br[91] wl[203] vdd gnd cell_6t
Xbit_r204_c91 bl[91] br[91] wl[204] vdd gnd cell_6t
Xbit_r205_c91 bl[91] br[91] wl[205] vdd gnd cell_6t
Xbit_r206_c91 bl[91] br[91] wl[206] vdd gnd cell_6t
Xbit_r207_c91 bl[91] br[91] wl[207] vdd gnd cell_6t
Xbit_r208_c91 bl[91] br[91] wl[208] vdd gnd cell_6t
Xbit_r209_c91 bl[91] br[91] wl[209] vdd gnd cell_6t
Xbit_r210_c91 bl[91] br[91] wl[210] vdd gnd cell_6t
Xbit_r211_c91 bl[91] br[91] wl[211] vdd gnd cell_6t
Xbit_r212_c91 bl[91] br[91] wl[212] vdd gnd cell_6t
Xbit_r213_c91 bl[91] br[91] wl[213] vdd gnd cell_6t
Xbit_r214_c91 bl[91] br[91] wl[214] vdd gnd cell_6t
Xbit_r215_c91 bl[91] br[91] wl[215] vdd gnd cell_6t
Xbit_r216_c91 bl[91] br[91] wl[216] vdd gnd cell_6t
Xbit_r217_c91 bl[91] br[91] wl[217] vdd gnd cell_6t
Xbit_r218_c91 bl[91] br[91] wl[218] vdd gnd cell_6t
Xbit_r219_c91 bl[91] br[91] wl[219] vdd gnd cell_6t
Xbit_r220_c91 bl[91] br[91] wl[220] vdd gnd cell_6t
Xbit_r221_c91 bl[91] br[91] wl[221] vdd gnd cell_6t
Xbit_r222_c91 bl[91] br[91] wl[222] vdd gnd cell_6t
Xbit_r223_c91 bl[91] br[91] wl[223] vdd gnd cell_6t
Xbit_r224_c91 bl[91] br[91] wl[224] vdd gnd cell_6t
Xbit_r225_c91 bl[91] br[91] wl[225] vdd gnd cell_6t
Xbit_r226_c91 bl[91] br[91] wl[226] vdd gnd cell_6t
Xbit_r227_c91 bl[91] br[91] wl[227] vdd gnd cell_6t
Xbit_r228_c91 bl[91] br[91] wl[228] vdd gnd cell_6t
Xbit_r229_c91 bl[91] br[91] wl[229] vdd gnd cell_6t
Xbit_r230_c91 bl[91] br[91] wl[230] vdd gnd cell_6t
Xbit_r231_c91 bl[91] br[91] wl[231] vdd gnd cell_6t
Xbit_r232_c91 bl[91] br[91] wl[232] vdd gnd cell_6t
Xbit_r233_c91 bl[91] br[91] wl[233] vdd gnd cell_6t
Xbit_r234_c91 bl[91] br[91] wl[234] vdd gnd cell_6t
Xbit_r235_c91 bl[91] br[91] wl[235] vdd gnd cell_6t
Xbit_r236_c91 bl[91] br[91] wl[236] vdd gnd cell_6t
Xbit_r237_c91 bl[91] br[91] wl[237] vdd gnd cell_6t
Xbit_r238_c91 bl[91] br[91] wl[238] vdd gnd cell_6t
Xbit_r239_c91 bl[91] br[91] wl[239] vdd gnd cell_6t
Xbit_r240_c91 bl[91] br[91] wl[240] vdd gnd cell_6t
Xbit_r241_c91 bl[91] br[91] wl[241] vdd gnd cell_6t
Xbit_r242_c91 bl[91] br[91] wl[242] vdd gnd cell_6t
Xbit_r243_c91 bl[91] br[91] wl[243] vdd gnd cell_6t
Xbit_r244_c91 bl[91] br[91] wl[244] vdd gnd cell_6t
Xbit_r245_c91 bl[91] br[91] wl[245] vdd gnd cell_6t
Xbit_r246_c91 bl[91] br[91] wl[246] vdd gnd cell_6t
Xbit_r247_c91 bl[91] br[91] wl[247] vdd gnd cell_6t
Xbit_r248_c91 bl[91] br[91] wl[248] vdd gnd cell_6t
Xbit_r249_c91 bl[91] br[91] wl[249] vdd gnd cell_6t
Xbit_r250_c91 bl[91] br[91] wl[250] vdd gnd cell_6t
Xbit_r251_c91 bl[91] br[91] wl[251] vdd gnd cell_6t
Xbit_r252_c91 bl[91] br[91] wl[252] vdd gnd cell_6t
Xbit_r253_c91 bl[91] br[91] wl[253] vdd gnd cell_6t
Xbit_r254_c91 bl[91] br[91] wl[254] vdd gnd cell_6t
Xbit_r255_c91 bl[91] br[91] wl[255] vdd gnd cell_6t
Xbit_r0_c92 bl[92] br[92] wl[0] vdd gnd cell_6t
Xbit_r1_c92 bl[92] br[92] wl[1] vdd gnd cell_6t
Xbit_r2_c92 bl[92] br[92] wl[2] vdd gnd cell_6t
Xbit_r3_c92 bl[92] br[92] wl[3] vdd gnd cell_6t
Xbit_r4_c92 bl[92] br[92] wl[4] vdd gnd cell_6t
Xbit_r5_c92 bl[92] br[92] wl[5] vdd gnd cell_6t
Xbit_r6_c92 bl[92] br[92] wl[6] vdd gnd cell_6t
Xbit_r7_c92 bl[92] br[92] wl[7] vdd gnd cell_6t
Xbit_r8_c92 bl[92] br[92] wl[8] vdd gnd cell_6t
Xbit_r9_c92 bl[92] br[92] wl[9] vdd gnd cell_6t
Xbit_r10_c92 bl[92] br[92] wl[10] vdd gnd cell_6t
Xbit_r11_c92 bl[92] br[92] wl[11] vdd gnd cell_6t
Xbit_r12_c92 bl[92] br[92] wl[12] vdd gnd cell_6t
Xbit_r13_c92 bl[92] br[92] wl[13] vdd gnd cell_6t
Xbit_r14_c92 bl[92] br[92] wl[14] vdd gnd cell_6t
Xbit_r15_c92 bl[92] br[92] wl[15] vdd gnd cell_6t
Xbit_r16_c92 bl[92] br[92] wl[16] vdd gnd cell_6t
Xbit_r17_c92 bl[92] br[92] wl[17] vdd gnd cell_6t
Xbit_r18_c92 bl[92] br[92] wl[18] vdd gnd cell_6t
Xbit_r19_c92 bl[92] br[92] wl[19] vdd gnd cell_6t
Xbit_r20_c92 bl[92] br[92] wl[20] vdd gnd cell_6t
Xbit_r21_c92 bl[92] br[92] wl[21] vdd gnd cell_6t
Xbit_r22_c92 bl[92] br[92] wl[22] vdd gnd cell_6t
Xbit_r23_c92 bl[92] br[92] wl[23] vdd gnd cell_6t
Xbit_r24_c92 bl[92] br[92] wl[24] vdd gnd cell_6t
Xbit_r25_c92 bl[92] br[92] wl[25] vdd gnd cell_6t
Xbit_r26_c92 bl[92] br[92] wl[26] vdd gnd cell_6t
Xbit_r27_c92 bl[92] br[92] wl[27] vdd gnd cell_6t
Xbit_r28_c92 bl[92] br[92] wl[28] vdd gnd cell_6t
Xbit_r29_c92 bl[92] br[92] wl[29] vdd gnd cell_6t
Xbit_r30_c92 bl[92] br[92] wl[30] vdd gnd cell_6t
Xbit_r31_c92 bl[92] br[92] wl[31] vdd gnd cell_6t
Xbit_r32_c92 bl[92] br[92] wl[32] vdd gnd cell_6t
Xbit_r33_c92 bl[92] br[92] wl[33] vdd gnd cell_6t
Xbit_r34_c92 bl[92] br[92] wl[34] vdd gnd cell_6t
Xbit_r35_c92 bl[92] br[92] wl[35] vdd gnd cell_6t
Xbit_r36_c92 bl[92] br[92] wl[36] vdd gnd cell_6t
Xbit_r37_c92 bl[92] br[92] wl[37] vdd gnd cell_6t
Xbit_r38_c92 bl[92] br[92] wl[38] vdd gnd cell_6t
Xbit_r39_c92 bl[92] br[92] wl[39] vdd gnd cell_6t
Xbit_r40_c92 bl[92] br[92] wl[40] vdd gnd cell_6t
Xbit_r41_c92 bl[92] br[92] wl[41] vdd gnd cell_6t
Xbit_r42_c92 bl[92] br[92] wl[42] vdd gnd cell_6t
Xbit_r43_c92 bl[92] br[92] wl[43] vdd gnd cell_6t
Xbit_r44_c92 bl[92] br[92] wl[44] vdd gnd cell_6t
Xbit_r45_c92 bl[92] br[92] wl[45] vdd gnd cell_6t
Xbit_r46_c92 bl[92] br[92] wl[46] vdd gnd cell_6t
Xbit_r47_c92 bl[92] br[92] wl[47] vdd gnd cell_6t
Xbit_r48_c92 bl[92] br[92] wl[48] vdd gnd cell_6t
Xbit_r49_c92 bl[92] br[92] wl[49] vdd gnd cell_6t
Xbit_r50_c92 bl[92] br[92] wl[50] vdd gnd cell_6t
Xbit_r51_c92 bl[92] br[92] wl[51] vdd gnd cell_6t
Xbit_r52_c92 bl[92] br[92] wl[52] vdd gnd cell_6t
Xbit_r53_c92 bl[92] br[92] wl[53] vdd gnd cell_6t
Xbit_r54_c92 bl[92] br[92] wl[54] vdd gnd cell_6t
Xbit_r55_c92 bl[92] br[92] wl[55] vdd gnd cell_6t
Xbit_r56_c92 bl[92] br[92] wl[56] vdd gnd cell_6t
Xbit_r57_c92 bl[92] br[92] wl[57] vdd gnd cell_6t
Xbit_r58_c92 bl[92] br[92] wl[58] vdd gnd cell_6t
Xbit_r59_c92 bl[92] br[92] wl[59] vdd gnd cell_6t
Xbit_r60_c92 bl[92] br[92] wl[60] vdd gnd cell_6t
Xbit_r61_c92 bl[92] br[92] wl[61] vdd gnd cell_6t
Xbit_r62_c92 bl[92] br[92] wl[62] vdd gnd cell_6t
Xbit_r63_c92 bl[92] br[92] wl[63] vdd gnd cell_6t
Xbit_r64_c92 bl[92] br[92] wl[64] vdd gnd cell_6t
Xbit_r65_c92 bl[92] br[92] wl[65] vdd gnd cell_6t
Xbit_r66_c92 bl[92] br[92] wl[66] vdd gnd cell_6t
Xbit_r67_c92 bl[92] br[92] wl[67] vdd gnd cell_6t
Xbit_r68_c92 bl[92] br[92] wl[68] vdd gnd cell_6t
Xbit_r69_c92 bl[92] br[92] wl[69] vdd gnd cell_6t
Xbit_r70_c92 bl[92] br[92] wl[70] vdd gnd cell_6t
Xbit_r71_c92 bl[92] br[92] wl[71] vdd gnd cell_6t
Xbit_r72_c92 bl[92] br[92] wl[72] vdd gnd cell_6t
Xbit_r73_c92 bl[92] br[92] wl[73] vdd gnd cell_6t
Xbit_r74_c92 bl[92] br[92] wl[74] vdd gnd cell_6t
Xbit_r75_c92 bl[92] br[92] wl[75] vdd gnd cell_6t
Xbit_r76_c92 bl[92] br[92] wl[76] vdd gnd cell_6t
Xbit_r77_c92 bl[92] br[92] wl[77] vdd gnd cell_6t
Xbit_r78_c92 bl[92] br[92] wl[78] vdd gnd cell_6t
Xbit_r79_c92 bl[92] br[92] wl[79] vdd gnd cell_6t
Xbit_r80_c92 bl[92] br[92] wl[80] vdd gnd cell_6t
Xbit_r81_c92 bl[92] br[92] wl[81] vdd gnd cell_6t
Xbit_r82_c92 bl[92] br[92] wl[82] vdd gnd cell_6t
Xbit_r83_c92 bl[92] br[92] wl[83] vdd gnd cell_6t
Xbit_r84_c92 bl[92] br[92] wl[84] vdd gnd cell_6t
Xbit_r85_c92 bl[92] br[92] wl[85] vdd gnd cell_6t
Xbit_r86_c92 bl[92] br[92] wl[86] vdd gnd cell_6t
Xbit_r87_c92 bl[92] br[92] wl[87] vdd gnd cell_6t
Xbit_r88_c92 bl[92] br[92] wl[88] vdd gnd cell_6t
Xbit_r89_c92 bl[92] br[92] wl[89] vdd gnd cell_6t
Xbit_r90_c92 bl[92] br[92] wl[90] vdd gnd cell_6t
Xbit_r91_c92 bl[92] br[92] wl[91] vdd gnd cell_6t
Xbit_r92_c92 bl[92] br[92] wl[92] vdd gnd cell_6t
Xbit_r93_c92 bl[92] br[92] wl[93] vdd gnd cell_6t
Xbit_r94_c92 bl[92] br[92] wl[94] vdd gnd cell_6t
Xbit_r95_c92 bl[92] br[92] wl[95] vdd gnd cell_6t
Xbit_r96_c92 bl[92] br[92] wl[96] vdd gnd cell_6t
Xbit_r97_c92 bl[92] br[92] wl[97] vdd gnd cell_6t
Xbit_r98_c92 bl[92] br[92] wl[98] vdd gnd cell_6t
Xbit_r99_c92 bl[92] br[92] wl[99] vdd gnd cell_6t
Xbit_r100_c92 bl[92] br[92] wl[100] vdd gnd cell_6t
Xbit_r101_c92 bl[92] br[92] wl[101] vdd gnd cell_6t
Xbit_r102_c92 bl[92] br[92] wl[102] vdd gnd cell_6t
Xbit_r103_c92 bl[92] br[92] wl[103] vdd gnd cell_6t
Xbit_r104_c92 bl[92] br[92] wl[104] vdd gnd cell_6t
Xbit_r105_c92 bl[92] br[92] wl[105] vdd gnd cell_6t
Xbit_r106_c92 bl[92] br[92] wl[106] vdd gnd cell_6t
Xbit_r107_c92 bl[92] br[92] wl[107] vdd gnd cell_6t
Xbit_r108_c92 bl[92] br[92] wl[108] vdd gnd cell_6t
Xbit_r109_c92 bl[92] br[92] wl[109] vdd gnd cell_6t
Xbit_r110_c92 bl[92] br[92] wl[110] vdd gnd cell_6t
Xbit_r111_c92 bl[92] br[92] wl[111] vdd gnd cell_6t
Xbit_r112_c92 bl[92] br[92] wl[112] vdd gnd cell_6t
Xbit_r113_c92 bl[92] br[92] wl[113] vdd gnd cell_6t
Xbit_r114_c92 bl[92] br[92] wl[114] vdd gnd cell_6t
Xbit_r115_c92 bl[92] br[92] wl[115] vdd gnd cell_6t
Xbit_r116_c92 bl[92] br[92] wl[116] vdd gnd cell_6t
Xbit_r117_c92 bl[92] br[92] wl[117] vdd gnd cell_6t
Xbit_r118_c92 bl[92] br[92] wl[118] vdd gnd cell_6t
Xbit_r119_c92 bl[92] br[92] wl[119] vdd gnd cell_6t
Xbit_r120_c92 bl[92] br[92] wl[120] vdd gnd cell_6t
Xbit_r121_c92 bl[92] br[92] wl[121] vdd gnd cell_6t
Xbit_r122_c92 bl[92] br[92] wl[122] vdd gnd cell_6t
Xbit_r123_c92 bl[92] br[92] wl[123] vdd gnd cell_6t
Xbit_r124_c92 bl[92] br[92] wl[124] vdd gnd cell_6t
Xbit_r125_c92 bl[92] br[92] wl[125] vdd gnd cell_6t
Xbit_r126_c92 bl[92] br[92] wl[126] vdd gnd cell_6t
Xbit_r127_c92 bl[92] br[92] wl[127] vdd gnd cell_6t
Xbit_r128_c92 bl[92] br[92] wl[128] vdd gnd cell_6t
Xbit_r129_c92 bl[92] br[92] wl[129] vdd gnd cell_6t
Xbit_r130_c92 bl[92] br[92] wl[130] vdd gnd cell_6t
Xbit_r131_c92 bl[92] br[92] wl[131] vdd gnd cell_6t
Xbit_r132_c92 bl[92] br[92] wl[132] vdd gnd cell_6t
Xbit_r133_c92 bl[92] br[92] wl[133] vdd gnd cell_6t
Xbit_r134_c92 bl[92] br[92] wl[134] vdd gnd cell_6t
Xbit_r135_c92 bl[92] br[92] wl[135] vdd gnd cell_6t
Xbit_r136_c92 bl[92] br[92] wl[136] vdd gnd cell_6t
Xbit_r137_c92 bl[92] br[92] wl[137] vdd gnd cell_6t
Xbit_r138_c92 bl[92] br[92] wl[138] vdd gnd cell_6t
Xbit_r139_c92 bl[92] br[92] wl[139] vdd gnd cell_6t
Xbit_r140_c92 bl[92] br[92] wl[140] vdd gnd cell_6t
Xbit_r141_c92 bl[92] br[92] wl[141] vdd gnd cell_6t
Xbit_r142_c92 bl[92] br[92] wl[142] vdd gnd cell_6t
Xbit_r143_c92 bl[92] br[92] wl[143] vdd gnd cell_6t
Xbit_r144_c92 bl[92] br[92] wl[144] vdd gnd cell_6t
Xbit_r145_c92 bl[92] br[92] wl[145] vdd gnd cell_6t
Xbit_r146_c92 bl[92] br[92] wl[146] vdd gnd cell_6t
Xbit_r147_c92 bl[92] br[92] wl[147] vdd gnd cell_6t
Xbit_r148_c92 bl[92] br[92] wl[148] vdd gnd cell_6t
Xbit_r149_c92 bl[92] br[92] wl[149] vdd gnd cell_6t
Xbit_r150_c92 bl[92] br[92] wl[150] vdd gnd cell_6t
Xbit_r151_c92 bl[92] br[92] wl[151] vdd gnd cell_6t
Xbit_r152_c92 bl[92] br[92] wl[152] vdd gnd cell_6t
Xbit_r153_c92 bl[92] br[92] wl[153] vdd gnd cell_6t
Xbit_r154_c92 bl[92] br[92] wl[154] vdd gnd cell_6t
Xbit_r155_c92 bl[92] br[92] wl[155] vdd gnd cell_6t
Xbit_r156_c92 bl[92] br[92] wl[156] vdd gnd cell_6t
Xbit_r157_c92 bl[92] br[92] wl[157] vdd gnd cell_6t
Xbit_r158_c92 bl[92] br[92] wl[158] vdd gnd cell_6t
Xbit_r159_c92 bl[92] br[92] wl[159] vdd gnd cell_6t
Xbit_r160_c92 bl[92] br[92] wl[160] vdd gnd cell_6t
Xbit_r161_c92 bl[92] br[92] wl[161] vdd gnd cell_6t
Xbit_r162_c92 bl[92] br[92] wl[162] vdd gnd cell_6t
Xbit_r163_c92 bl[92] br[92] wl[163] vdd gnd cell_6t
Xbit_r164_c92 bl[92] br[92] wl[164] vdd gnd cell_6t
Xbit_r165_c92 bl[92] br[92] wl[165] vdd gnd cell_6t
Xbit_r166_c92 bl[92] br[92] wl[166] vdd gnd cell_6t
Xbit_r167_c92 bl[92] br[92] wl[167] vdd gnd cell_6t
Xbit_r168_c92 bl[92] br[92] wl[168] vdd gnd cell_6t
Xbit_r169_c92 bl[92] br[92] wl[169] vdd gnd cell_6t
Xbit_r170_c92 bl[92] br[92] wl[170] vdd gnd cell_6t
Xbit_r171_c92 bl[92] br[92] wl[171] vdd gnd cell_6t
Xbit_r172_c92 bl[92] br[92] wl[172] vdd gnd cell_6t
Xbit_r173_c92 bl[92] br[92] wl[173] vdd gnd cell_6t
Xbit_r174_c92 bl[92] br[92] wl[174] vdd gnd cell_6t
Xbit_r175_c92 bl[92] br[92] wl[175] vdd gnd cell_6t
Xbit_r176_c92 bl[92] br[92] wl[176] vdd gnd cell_6t
Xbit_r177_c92 bl[92] br[92] wl[177] vdd gnd cell_6t
Xbit_r178_c92 bl[92] br[92] wl[178] vdd gnd cell_6t
Xbit_r179_c92 bl[92] br[92] wl[179] vdd gnd cell_6t
Xbit_r180_c92 bl[92] br[92] wl[180] vdd gnd cell_6t
Xbit_r181_c92 bl[92] br[92] wl[181] vdd gnd cell_6t
Xbit_r182_c92 bl[92] br[92] wl[182] vdd gnd cell_6t
Xbit_r183_c92 bl[92] br[92] wl[183] vdd gnd cell_6t
Xbit_r184_c92 bl[92] br[92] wl[184] vdd gnd cell_6t
Xbit_r185_c92 bl[92] br[92] wl[185] vdd gnd cell_6t
Xbit_r186_c92 bl[92] br[92] wl[186] vdd gnd cell_6t
Xbit_r187_c92 bl[92] br[92] wl[187] vdd gnd cell_6t
Xbit_r188_c92 bl[92] br[92] wl[188] vdd gnd cell_6t
Xbit_r189_c92 bl[92] br[92] wl[189] vdd gnd cell_6t
Xbit_r190_c92 bl[92] br[92] wl[190] vdd gnd cell_6t
Xbit_r191_c92 bl[92] br[92] wl[191] vdd gnd cell_6t
Xbit_r192_c92 bl[92] br[92] wl[192] vdd gnd cell_6t
Xbit_r193_c92 bl[92] br[92] wl[193] vdd gnd cell_6t
Xbit_r194_c92 bl[92] br[92] wl[194] vdd gnd cell_6t
Xbit_r195_c92 bl[92] br[92] wl[195] vdd gnd cell_6t
Xbit_r196_c92 bl[92] br[92] wl[196] vdd gnd cell_6t
Xbit_r197_c92 bl[92] br[92] wl[197] vdd gnd cell_6t
Xbit_r198_c92 bl[92] br[92] wl[198] vdd gnd cell_6t
Xbit_r199_c92 bl[92] br[92] wl[199] vdd gnd cell_6t
Xbit_r200_c92 bl[92] br[92] wl[200] vdd gnd cell_6t
Xbit_r201_c92 bl[92] br[92] wl[201] vdd gnd cell_6t
Xbit_r202_c92 bl[92] br[92] wl[202] vdd gnd cell_6t
Xbit_r203_c92 bl[92] br[92] wl[203] vdd gnd cell_6t
Xbit_r204_c92 bl[92] br[92] wl[204] vdd gnd cell_6t
Xbit_r205_c92 bl[92] br[92] wl[205] vdd gnd cell_6t
Xbit_r206_c92 bl[92] br[92] wl[206] vdd gnd cell_6t
Xbit_r207_c92 bl[92] br[92] wl[207] vdd gnd cell_6t
Xbit_r208_c92 bl[92] br[92] wl[208] vdd gnd cell_6t
Xbit_r209_c92 bl[92] br[92] wl[209] vdd gnd cell_6t
Xbit_r210_c92 bl[92] br[92] wl[210] vdd gnd cell_6t
Xbit_r211_c92 bl[92] br[92] wl[211] vdd gnd cell_6t
Xbit_r212_c92 bl[92] br[92] wl[212] vdd gnd cell_6t
Xbit_r213_c92 bl[92] br[92] wl[213] vdd gnd cell_6t
Xbit_r214_c92 bl[92] br[92] wl[214] vdd gnd cell_6t
Xbit_r215_c92 bl[92] br[92] wl[215] vdd gnd cell_6t
Xbit_r216_c92 bl[92] br[92] wl[216] vdd gnd cell_6t
Xbit_r217_c92 bl[92] br[92] wl[217] vdd gnd cell_6t
Xbit_r218_c92 bl[92] br[92] wl[218] vdd gnd cell_6t
Xbit_r219_c92 bl[92] br[92] wl[219] vdd gnd cell_6t
Xbit_r220_c92 bl[92] br[92] wl[220] vdd gnd cell_6t
Xbit_r221_c92 bl[92] br[92] wl[221] vdd gnd cell_6t
Xbit_r222_c92 bl[92] br[92] wl[222] vdd gnd cell_6t
Xbit_r223_c92 bl[92] br[92] wl[223] vdd gnd cell_6t
Xbit_r224_c92 bl[92] br[92] wl[224] vdd gnd cell_6t
Xbit_r225_c92 bl[92] br[92] wl[225] vdd gnd cell_6t
Xbit_r226_c92 bl[92] br[92] wl[226] vdd gnd cell_6t
Xbit_r227_c92 bl[92] br[92] wl[227] vdd gnd cell_6t
Xbit_r228_c92 bl[92] br[92] wl[228] vdd gnd cell_6t
Xbit_r229_c92 bl[92] br[92] wl[229] vdd gnd cell_6t
Xbit_r230_c92 bl[92] br[92] wl[230] vdd gnd cell_6t
Xbit_r231_c92 bl[92] br[92] wl[231] vdd gnd cell_6t
Xbit_r232_c92 bl[92] br[92] wl[232] vdd gnd cell_6t
Xbit_r233_c92 bl[92] br[92] wl[233] vdd gnd cell_6t
Xbit_r234_c92 bl[92] br[92] wl[234] vdd gnd cell_6t
Xbit_r235_c92 bl[92] br[92] wl[235] vdd gnd cell_6t
Xbit_r236_c92 bl[92] br[92] wl[236] vdd gnd cell_6t
Xbit_r237_c92 bl[92] br[92] wl[237] vdd gnd cell_6t
Xbit_r238_c92 bl[92] br[92] wl[238] vdd gnd cell_6t
Xbit_r239_c92 bl[92] br[92] wl[239] vdd gnd cell_6t
Xbit_r240_c92 bl[92] br[92] wl[240] vdd gnd cell_6t
Xbit_r241_c92 bl[92] br[92] wl[241] vdd gnd cell_6t
Xbit_r242_c92 bl[92] br[92] wl[242] vdd gnd cell_6t
Xbit_r243_c92 bl[92] br[92] wl[243] vdd gnd cell_6t
Xbit_r244_c92 bl[92] br[92] wl[244] vdd gnd cell_6t
Xbit_r245_c92 bl[92] br[92] wl[245] vdd gnd cell_6t
Xbit_r246_c92 bl[92] br[92] wl[246] vdd gnd cell_6t
Xbit_r247_c92 bl[92] br[92] wl[247] vdd gnd cell_6t
Xbit_r248_c92 bl[92] br[92] wl[248] vdd gnd cell_6t
Xbit_r249_c92 bl[92] br[92] wl[249] vdd gnd cell_6t
Xbit_r250_c92 bl[92] br[92] wl[250] vdd gnd cell_6t
Xbit_r251_c92 bl[92] br[92] wl[251] vdd gnd cell_6t
Xbit_r252_c92 bl[92] br[92] wl[252] vdd gnd cell_6t
Xbit_r253_c92 bl[92] br[92] wl[253] vdd gnd cell_6t
Xbit_r254_c92 bl[92] br[92] wl[254] vdd gnd cell_6t
Xbit_r255_c92 bl[92] br[92] wl[255] vdd gnd cell_6t
Xbit_r0_c93 bl[93] br[93] wl[0] vdd gnd cell_6t
Xbit_r1_c93 bl[93] br[93] wl[1] vdd gnd cell_6t
Xbit_r2_c93 bl[93] br[93] wl[2] vdd gnd cell_6t
Xbit_r3_c93 bl[93] br[93] wl[3] vdd gnd cell_6t
Xbit_r4_c93 bl[93] br[93] wl[4] vdd gnd cell_6t
Xbit_r5_c93 bl[93] br[93] wl[5] vdd gnd cell_6t
Xbit_r6_c93 bl[93] br[93] wl[6] vdd gnd cell_6t
Xbit_r7_c93 bl[93] br[93] wl[7] vdd gnd cell_6t
Xbit_r8_c93 bl[93] br[93] wl[8] vdd gnd cell_6t
Xbit_r9_c93 bl[93] br[93] wl[9] vdd gnd cell_6t
Xbit_r10_c93 bl[93] br[93] wl[10] vdd gnd cell_6t
Xbit_r11_c93 bl[93] br[93] wl[11] vdd gnd cell_6t
Xbit_r12_c93 bl[93] br[93] wl[12] vdd gnd cell_6t
Xbit_r13_c93 bl[93] br[93] wl[13] vdd gnd cell_6t
Xbit_r14_c93 bl[93] br[93] wl[14] vdd gnd cell_6t
Xbit_r15_c93 bl[93] br[93] wl[15] vdd gnd cell_6t
Xbit_r16_c93 bl[93] br[93] wl[16] vdd gnd cell_6t
Xbit_r17_c93 bl[93] br[93] wl[17] vdd gnd cell_6t
Xbit_r18_c93 bl[93] br[93] wl[18] vdd gnd cell_6t
Xbit_r19_c93 bl[93] br[93] wl[19] vdd gnd cell_6t
Xbit_r20_c93 bl[93] br[93] wl[20] vdd gnd cell_6t
Xbit_r21_c93 bl[93] br[93] wl[21] vdd gnd cell_6t
Xbit_r22_c93 bl[93] br[93] wl[22] vdd gnd cell_6t
Xbit_r23_c93 bl[93] br[93] wl[23] vdd gnd cell_6t
Xbit_r24_c93 bl[93] br[93] wl[24] vdd gnd cell_6t
Xbit_r25_c93 bl[93] br[93] wl[25] vdd gnd cell_6t
Xbit_r26_c93 bl[93] br[93] wl[26] vdd gnd cell_6t
Xbit_r27_c93 bl[93] br[93] wl[27] vdd gnd cell_6t
Xbit_r28_c93 bl[93] br[93] wl[28] vdd gnd cell_6t
Xbit_r29_c93 bl[93] br[93] wl[29] vdd gnd cell_6t
Xbit_r30_c93 bl[93] br[93] wl[30] vdd gnd cell_6t
Xbit_r31_c93 bl[93] br[93] wl[31] vdd gnd cell_6t
Xbit_r32_c93 bl[93] br[93] wl[32] vdd gnd cell_6t
Xbit_r33_c93 bl[93] br[93] wl[33] vdd gnd cell_6t
Xbit_r34_c93 bl[93] br[93] wl[34] vdd gnd cell_6t
Xbit_r35_c93 bl[93] br[93] wl[35] vdd gnd cell_6t
Xbit_r36_c93 bl[93] br[93] wl[36] vdd gnd cell_6t
Xbit_r37_c93 bl[93] br[93] wl[37] vdd gnd cell_6t
Xbit_r38_c93 bl[93] br[93] wl[38] vdd gnd cell_6t
Xbit_r39_c93 bl[93] br[93] wl[39] vdd gnd cell_6t
Xbit_r40_c93 bl[93] br[93] wl[40] vdd gnd cell_6t
Xbit_r41_c93 bl[93] br[93] wl[41] vdd gnd cell_6t
Xbit_r42_c93 bl[93] br[93] wl[42] vdd gnd cell_6t
Xbit_r43_c93 bl[93] br[93] wl[43] vdd gnd cell_6t
Xbit_r44_c93 bl[93] br[93] wl[44] vdd gnd cell_6t
Xbit_r45_c93 bl[93] br[93] wl[45] vdd gnd cell_6t
Xbit_r46_c93 bl[93] br[93] wl[46] vdd gnd cell_6t
Xbit_r47_c93 bl[93] br[93] wl[47] vdd gnd cell_6t
Xbit_r48_c93 bl[93] br[93] wl[48] vdd gnd cell_6t
Xbit_r49_c93 bl[93] br[93] wl[49] vdd gnd cell_6t
Xbit_r50_c93 bl[93] br[93] wl[50] vdd gnd cell_6t
Xbit_r51_c93 bl[93] br[93] wl[51] vdd gnd cell_6t
Xbit_r52_c93 bl[93] br[93] wl[52] vdd gnd cell_6t
Xbit_r53_c93 bl[93] br[93] wl[53] vdd gnd cell_6t
Xbit_r54_c93 bl[93] br[93] wl[54] vdd gnd cell_6t
Xbit_r55_c93 bl[93] br[93] wl[55] vdd gnd cell_6t
Xbit_r56_c93 bl[93] br[93] wl[56] vdd gnd cell_6t
Xbit_r57_c93 bl[93] br[93] wl[57] vdd gnd cell_6t
Xbit_r58_c93 bl[93] br[93] wl[58] vdd gnd cell_6t
Xbit_r59_c93 bl[93] br[93] wl[59] vdd gnd cell_6t
Xbit_r60_c93 bl[93] br[93] wl[60] vdd gnd cell_6t
Xbit_r61_c93 bl[93] br[93] wl[61] vdd gnd cell_6t
Xbit_r62_c93 bl[93] br[93] wl[62] vdd gnd cell_6t
Xbit_r63_c93 bl[93] br[93] wl[63] vdd gnd cell_6t
Xbit_r64_c93 bl[93] br[93] wl[64] vdd gnd cell_6t
Xbit_r65_c93 bl[93] br[93] wl[65] vdd gnd cell_6t
Xbit_r66_c93 bl[93] br[93] wl[66] vdd gnd cell_6t
Xbit_r67_c93 bl[93] br[93] wl[67] vdd gnd cell_6t
Xbit_r68_c93 bl[93] br[93] wl[68] vdd gnd cell_6t
Xbit_r69_c93 bl[93] br[93] wl[69] vdd gnd cell_6t
Xbit_r70_c93 bl[93] br[93] wl[70] vdd gnd cell_6t
Xbit_r71_c93 bl[93] br[93] wl[71] vdd gnd cell_6t
Xbit_r72_c93 bl[93] br[93] wl[72] vdd gnd cell_6t
Xbit_r73_c93 bl[93] br[93] wl[73] vdd gnd cell_6t
Xbit_r74_c93 bl[93] br[93] wl[74] vdd gnd cell_6t
Xbit_r75_c93 bl[93] br[93] wl[75] vdd gnd cell_6t
Xbit_r76_c93 bl[93] br[93] wl[76] vdd gnd cell_6t
Xbit_r77_c93 bl[93] br[93] wl[77] vdd gnd cell_6t
Xbit_r78_c93 bl[93] br[93] wl[78] vdd gnd cell_6t
Xbit_r79_c93 bl[93] br[93] wl[79] vdd gnd cell_6t
Xbit_r80_c93 bl[93] br[93] wl[80] vdd gnd cell_6t
Xbit_r81_c93 bl[93] br[93] wl[81] vdd gnd cell_6t
Xbit_r82_c93 bl[93] br[93] wl[82] vdd gnd cell_6t
Xbit_r83_c93 bl[93] br[93] wl[83] vdd gnd cell_6t
Xbit_r84_c93 bl[93] br[93] wl[84] vdd gnd cell_6t
Xbit_r85_c93 bl[93] br[93] wl[85] vdd gnd cell_6t
Xbit_r86_c93 bl[93] br[93] wl[86] vdd gnd cell_6t
Xbit_r87_c93 bl[93] br[93] wl[87] vdd gnd cell_6t
Xbit_r88_c93 bl[93] br[93] wl[88] vdd gnd cell_6t
Xbit_r89_c93 bl[93] br[93] wl[89] vdd gnd cell_6t
Xbit_r90_c93 bl[93] br[93] wl[90] vdd gnd cell_6t
Xbit_r91_c93 bl[93] br[93] wl[91] vdd gnd cell_6t
Xbit_r92_c93 bl[93] br[93] wl[92] vdd gnd cell_6t
Xbit_r93_c93 bl[93] br[93] wl[93] vdd gnd cell_6t
Xbit_r94_c93 bl[93] br[93] wl[94] vdd gnd cell_6t
Xbit_r95_c93 bl[93] br[93] wl[95] vdd gnd cell_6t
Xbit_r96_c93 bl[93] br[93] wl[96] vdd gnd cell_6t
Xbit_r97_c93 bl[93] br[93] wl[97] vdd gnd cell_6t
Xbit_r98_c93 bl[93] br[93] wl[98] vdd gnd cell_6t
Xbit_r99_c93 bl[93] br[93] wl[99] vdd gnd cell_6t
Xbit_r100_c93 bl[93] br[93] wl[100] vdd gnd cell_6t
Xbit_r101_c93 bl[93] br[93] wl[101] vdd gnd cell_6t
Xbit_r102_c93 bl[93] br[93] wl[102] vdd gnd cell_6t
Xbit_r103_c93 bl[93] br[93] wl[103] vdd gnd cell_6t
Xbit_r104_c93 bl[93] br[93] wl[104] vdd gnd cell_6t
Xbit_r105_c93 bl[93] br[93] wl[105] vdd gnd cell_6t
Xbit_r106_c93 bl[93] br[93] wl[106] vdd gnd cell_6t
Xbit_r107_c93 bl[93] br[93] wl[107] vdd gnd cell_6t
Xbit_r108_c93 bl[93] br[93] wl[108] vdd gnd cell_6t
Xbit_r109_c93 bl[93] br[93] wl[109] vdd gnd cell_6t
Xbit_r110_c93 bl[93] br[93] wl[110] vdd gnd cell_6t
Xbit_r111_c93 bl[93] br[93] wl[111] vdd gnd cell_6t
Xbit_r112_c93 bl[93] br[93] wl[112] vdd gnd cell_6t
Xbit_r113_c93 bl[93] br[93] wl[113] vdd gnd cell_6t
Xbit_r114_c93 bl[93] br[93] wl[114] vdd gnd cell_6t
Xbit_r115_c93 bl[93] br[93] wl[115] vdd gnd cell_6t
Xbit_r116_c93 bl[93] br[93] wl[116] vdd gnd cell_6t
Xbit_r117_c93 bl[93] br[93] wl[117] vdd gnd cell_6t
Xbit_r118_c93 bl[93] br[93] wl[118] vdd gnd cell_6t
Xbit_r119_c93 bl[93] br[93] wl[119] vdd gnd cell_6t
Xbit_r120_c93 bl[93] br[93] wl[120] vdd gnd cell_6t
Xbit_r121_c93 bl[93] br[93] wl[121] vdd gnd cell_6t
Xbit_r122_c93 bl[93] br[93] wl[122] vdd gnd cell_6t
Xbit_r123_c93 bl[93] br[93] wl[123] vdd gnd cell_6t
Xbit_r124_c93 bl[93] br[93] wl[124] vdd gnd cell_6t
Xbit_r125_c93 bl[93] br[93] wl[125] vdd gnd cell_6t
Xbit_r126_c93 bl[93] br[93] wl[126] vdd gnd cell_6t
Xbit_r127_c93 bl[93] br[93] wl[127] vdd gnd cell_6t
Xbit_r128_c93 bl[93] br[93] wl[128] vdd gnd cell_6t
Xbit_r129_c93 bl[93] br[93] wl[129] vdd gnd cell_6t
Xbit_r130_c93 bl[93] br[93] wl[130] vdd gnd cell_6t
Xbit_r131_c93 bl[93] br[93] wl[131] vdd gnd cell_6t
Xbit_r132_c93 bl[93] br[93] wl[132] vdd gnd cell_6t
Xbit_r133_c93 bl[93] br[93] wl[133] vdd gnd cell_6t
Xbit_r134_c93 bl[93] br[93] wl[134] vdd gnd cell_6t
Xbit_r135_c93 bl[93] br[93] wl[135] vdd gnd cell_6t
Xbit_r136_c93 bl[93] br[93] wl[136] vdd gnd cell_6t
Xbit_r137_c93 bl[93] br[93] wl[137] vdd gnd cell_6t
Xbit_r138_c93 bl[93] br[93] wl[138] vdd gnd cell_6t
Xbit_r139_c93 bl[93] br[93] wl[139] vdd gnd cell_6t
Xbit_r140_c93 bl[93] br[93] wl[140] vdd gnd cell_6t
Xbit_r141_c93 bl[93] br[93] wl[141] vdd gnd cell_6t
Xbit_r142_c93 bl[93] br[93] wl[142] vdd gnd cell_6t
Xbit_r143_c93 bl[93] br[93] wl[143] vdd gnd cell_6t
Xbit_r144_c93 bl[93] br[93] wl[144] vdd gnd cell_6t
Xbit_r145_c93 bl[93] br[93] wl[145] vdd gnd cell_6t
Xbit_r146_c93 bl[93] br[93] wl[146] vdd gnd cell_6t
Xbit_r147_c93 bl[93] br[93] wl[147] vdd gnd cell_6t
Xbit_r148_c93 bl[93] br[93] wl[148] vdd gnd cell_6t
Xbit_r149_c93 bl[93] br[93] wl[149] vdd gnd cell_6t
Xbit_r150_c93 bl[93] br[93] wl[150] vdd gnd cell_6t
Xbit_r151_c93 bl[93] br[93] wl[151] vdd gnd cell_6t
Xbit_r152_c93 bl[93] br[93] wl[152] vdd gnd cell_6t
Xbit_r153_c93 bl[93] br[93] wl[153] vdd gnd cell_6t
Xbit_r154_c93 bl[93] br[93] wl[154] vdd gnd cell_6t
Xbit_r155_c93 bl[93] br[93] wl[155] vdd gnd cell_6t
Xbit_r156_c93 bl[93] br[93] wl[156] vdd gnd cell_6t
Xbit_r157_c93 bl[93] br[93] wl[157] vdd gnd cell_6t
Xbit_r158_c93 bl[93] br[93] wl[158] vdd gnd cell_6t
Xbit_r159_c93 bl[93] br[93] wl[159] vdd gnd cell_6t
Xbit_r160_c93 bl[93] br[93] wl[160] vdd gnd cell_6t
Xbit_r161_c93 bl[93] br[93] wl[161] vdd gnd cell_6t
Xbit_r162_c93 bl[93] br[93] wl[162] vdd gnd cell_6t
Xbit_r163_c93 bl[93] br[93] wl[163] vdd gnd cell_6t
Xbit_r164_c93 bl[93] br[93] wl[164] vdd gnd cell_6t
Xbit_r165_c93 bl[93] br[93] wl[165] vdd gnd cell_6t
Xbit_r166_c93 bl[93] br[93] wl[166] vdd gnd cell_6t
Xbit_r167_c93 bl[93] br[93] wl[167] vdd gnd cell_6t
Xbit_r168_c93 bl[93] br[93] wl[168] vdd gnd cell_6t
Xbit_r169_c93 bl[93] br[93] wl[169] vdd gnd cell_6t
Xbit_r170_c93 bl[93] br[93] wl[170] vdd gnd cell_6t
Xbit_r171_c93 bl[93] br[93] wl[171] vdd gnd cell_6t
Xbit_r172_c93 bl[93] br[93] wl[172] vdd gnd cell_6t
Xbit_r173_c93 bl[93] br[93] wl[173] vdd gnd cell_6t
Xbit_r174_c93 bl[93] br[93] wl[174] vdd gnd cell_6t
Xbit_r175_c93 bl[93] br[93] wl[175] vdd gnd cell_6t
Xbit_r176_c93 bl[93] br[93] wl[176] vdd gnd cell_6t
Xbit_r177_c93 bl[93] br[93] wl[177] vdd gnd cell_6t
Xbit_r178_c93 bl[93] br[93] wl[178] vdd gnd cell_6t
Xbit_r179_c93 bl[93] br[93] wl[179] vdd gnd cell_6t
Xbit_r180_c93 bl[93] br[93] wl[180] vdd gnd cell_6t
Xbit_r181_c93 bl[93] br[93] wl[181] vdd gnd cell_6t
Xbit_r182_c93 bl[93] br[93] wl[182] vdd gnd cell_6t
Xbit_r183_c93 bl[93] br[93] wl[183] vdd gnd cell_6t
Xbit_r184_c93 bl[93] br[93] wl[184] vdd gnd cell_6t
Xbit_r185_c93 bl[93] br[93] wl[185] vdd gnd cell_6t
Xbit_r186_c93 bl[93] br[93] wl[186] vdd gnd cell_6t
Xbit_r187_c93 bl[93] br[93] wl[187] vdd gnd cell_6t
Xbit_r188_c93 bl[93] br[93] wl[188] vdd gnd cell_6t
Xbit_r189_c93 bl[93] br[93] wl[189] vdd gnd cell_6t
Xbit_r190_c93 bl[93] br[93] wl[190] vdd gnd cell_6t
Xbit_r191_c93 bl[93] br[93] wl[191] vdd gnd cell_6t
Xbit_r192_c93 bl[93] br[93] wl[192] vdd gnd cell_6t
Xbit_r193_c93 bl[93] br[93] wl[193] vdd gnd cell_6t
Xbit_r194_c93 bl[93] br[93] wl[194] vdd gnd cell_6t
Xbit_r195_c93 bl[93] br[93] wl[195] vdd gnd cell_6t
Xbit_r196_c93 bl[93] br[93] wl[196] vdd gnd cell_6t
Xbit_r197_c93 bl[93] br[93] wl[197] vdd gnd cell_6t
Xbit_r198_c93 bl[93] br[93] wl[198] vdd gnd cell_6t
Xbit_r199_c93 bl[93] br[93] wl[199] vdd gnd cell_6t
Xbit_r200_c93 bl[93] br[93] wl[200] vdd gnd cell_6t
Xbit_r201_c93 bl[93] br[93] wl[201] vdd gnd cell_6t
Xbit_r202_c93 bl[93] br[93] wl[202] vdd gnd cell_6t
Xbit_r203_c93 bl[93] br[93] wl[203] vdd gnd cell_6t
Xbit_r204_c93 bl[93] br[93] wl[204] vdd gnd cell_6t
Xbit_r205_c93 bl[93] br[93] wl[205] vdd gnd cell_6t
Xbit_r206_c93 bl[93] br[93] wl[206] vdd gnd cell_6t
Xbit_r207_c93 bl[93] br[93] wl[207] vdd gnd cell_6t
Xbit_r208_c93 bl[93] br[93] wl[208] vdd gnd cell_6t
Xbit_r209_c93 bl[93] br[93] wl[209] vdd gnd cell_6t
Xbit_r210_c93 bl[93] br[93] wl[210] vdd gnd cell_6t
Xbit_r211_c93 bl[93] br[93] wl[211] vdd gnd cell_6t
Xbit_r212_c93 bl[93] br[93] wl[212] vdd gnd cell_6t
Xbit_r213_c93 bl[93] br[93] wl[213] vdd gnd cell_6t
Xbit_r214_c93 bl[93] br[93] wl[214] vdd gnd cell_6t
Xbit_r215_c93 bl[93] br[93] wl[215] vdd gnd cell_6t
Xbit_r216_c93 bl[93] br[93] wl[216] vdd gnd cell_6t
Xbit_r217_c93 bl[93] br[93] wl[217] vdd gnd cell_6t
Xbit_r218_c93 bl[93] br[93] wl[218] vdd gnd cell_6t
Xbit_r219_c93 bl[93] br[93] wl[219] vdd gnd cell_6t
Xbit_r220_c93 bl[93] br[93] wl[220] vdd gnd cell_6t
Xbit_r221_c93 bl[93] br[93] wl[221] vdd gnd cell_6t
Xbit_r222_c93 bl[93] br[93] wl[222] vdd gnd cell_6t
Xbit_r223_c93 bl[93] br[93] wl[223] vdd gnd cell_6t
Xbit_r224_c93 bl[93] br[93] wl[224] vdd gnd cell_6t
Xbit_r225_c93 bl[93] br[93] wl[225] vdd gnd cell_6t
Xbit_r226_c93 bl[93] br[93] wl[226] vdd gnd cell_6t
Xbit_r227_c93 bl[93] br[93] wl[227] vdd gnd cell_6t
Xbit_r228_c93 bl[93] br[93] wl[228] vdd gnd cell_6t
Xbit_r229_c93 bl[93] br[93] wl[229] vdd gnd cell_6t
Xbit_r230_c93 bl[93] br[93] wl[230] vdd gnd cell_6t
Xbit_r231_c93 bl[93] br[93] wl[231] vdd gnd cell_6t
Xbit_r232_c93 bl[93] br[93] wl[232] vdd gnd cell_6t
Xbit_r233_c93 bl[93] br[93] wl[233] vdd gnd cell_6t
Xbit_r234_c93 bl[93] br[93] wl[234] vdd gnd cell_6t
Xbit_r235_c93 bl[93] br[93] wl[235] vdd gnd cell_6t
Xbit_r236_c93 bl[93] br[93] wl[236] vdd gnd cell_6t
Xbit_r237_c93 bl[93] br[93] wl[237] vdd gnd cell_6t
Xbit_r238_c93 bl[93] br[93] wl[238] vdd gnd cell_6t
Xbit_r239_c93 bl[93] br[93] wl[239] vdd gnd cell_6t
Xbit_r240_c93 bl[93] br[93] wl[240] vdd gnd cell_6t
Xbit_r241_c93 bl[93] br[93] wl[241] vdd gnd cell_6t
Xbit_r242_c93 bl[93] br[93] wl[242] vdd gnd cell_6t
Xbit_r243_c93 bl[93] br[93] wl[243] vdd gnd cell_6t
Xbit_r244_c93 bl[93] br[93] wl[244] vdd gnd cell_6t
Xbit_r245_c93 bl[93] br[93] wl[245] vdd gnd cell_6t
Xbit_r246_c93 bl[93] br[93] wl[246] vdd gnd cell_6t
Xbit_r247_c93 bl[93] br[93] wl[247] vdd gnd cell_6t
Xbit_r248_c93 bl[93] br[93] wl[248] vdd gnd cell_6t
Xbit_r249_c93 bl[93] br[93] wl[249] vdd gnd cell_6t
Xbit_r250_c93 bl[93] br[93] wl[250] vdd gnd cell_6t
Xbit_r251_c93 bl[93] br[93] wl[251] vdd gnd cell_6t
Xbit_r252_c93 bl[93] br[93] wl[252] vdd gnd cell_6t
Xbit_r253_c93 bl[93] br[93] wl[253] vdd gnd cell_6t
Xbit_r254_c93 bl[93] br[93] wl[254] vdd gnd cell_6t
Xbit_r255_c93 bl[93] br[93] wl[255] vdd gnd cell_6t
Xbit_r0_c94 bl[94] br[94] wl[0] vdd gnd cell_6t
Xbit_r1_c94 bl[94] br[94] wl[1] vdd gnd cell_6t
Xbit_r2_c94 bl[94] br[94] wl[2] vdd gnd cell_6t
Xbit_r3_c94 bl[94] br[94] wl[3] vdd gnd cell_6t
Xbit_r4_c94 bl[94] br[94] wl[4] vdd gnd cell_6t
Xbit_r5_c94 bl[94] br[94] wl[5] vdd gnd cell_6t
Xbit_r6_c94 bl[94] br[94] wl[6] vdd gnd cell_6t
Xbit_r7_c94 bl[94] br[94] wl[7] vdd gnd cell_6t
Xbit_r8_c94 bl[94] br[94] wl[8] vdd gnd cell_6t
Xbit_r9_c94 bl[94] br[94] wl[9] vdd gnd cell_6t
Xbit_r10_c94 bl[94] br[94] wl[10] vdd gnd cell_6t
Xbit_r11_c94 bl[94] br[94] wl[11] vdd gnd cell_6t
Xbit_r12_c94 bl[94] br[94] wl[12] vdd gnd cell_6t
Xbit_r13_c94 bl[94] br[94] wl[13] vdd gnd cell_6t
Xbit_r14_c94 bl[94] br[94] wl[14] vdd gnd cell_6t
Xbit_r15_c94 bl[94] br[94] wl[15] vdd gnd cell_6t
Xbit_r16_c94 bl[94] br[94] wl[16] vdd gnd cell_6t
Xbit_r17_c94 bl[94] br[94] wl[17] vdd gnd cell_6t
Xbit_r18_c94 bl[94] br[94] wl[18] vdd gnd cell_6t
Xbit_r19_c94 bl[94] br[94] wl[19] vdd gnd cell_6t
Xbit_r20_c94 bl[94] br[94] wl[20] vdd gnd cell_6t
Xbit_r21_c94 bl[94] br[94] wl[21] vdd gnd cell_6t
Xbit_r22_c94 bl[94] br[94] wl[22] vdd gnd cell_6t
Xbit_r23_c94 bl[94] br[94] wl[23] vdd gnd cell_6t
Xbit_r24_c94 bl[94] br[94] wl[24] vdd gnd cell_6t
Xbit_r25_c94 bl[94] br[94] wl[25] vdd gnd cell_6t
Xbit_r26_c94 bl[94] br[94] wl[26] vdd gnd cell_6t
Xbit_r27_c94 bl[94] br[94] wl[27] vdd gnd cell_6t
Xbit_r28_c94 bl[94] br[94] wl[28] vdd gnd cell_6t
Xbit_r29_c94 bl[94] br[94] wl[29] vdd gnd cell_6t
Xbit_r30_c94 bl[94] br[94] wl[30] vdd gnd cell_6t
Xbit_r31_c94 bl[94] br[94] wl[31] vdd gnd cell_6t
Xbit_r32_c94 bl[94] br[94] wl[32] vdd gnd cell_6t
Xbit_r33_c94 bl[94] br[94] wl[33] vdd gnd cell_6t
Xbit_r34_c94 bl[94] br[94] wl[34] vdd gnd cell_6t
Xbit_r35_c94 bl[94] br[94] wl[35] vdd gnd cell_6t
Xbit_r36_c94 bl[94] br[94] wl[36] vdd gnd cell_6t
Xbit_r37_c94 bl[94] br[94] wl[37] vdd gnd cell_6t
Xbit_r38_c94 bl[94] br[94] wl[38] vdd gnd cell_6t
Xbit_r39_c94 bl[94] br[94] wl[39] vdd gnd cell_6t
Xbit_r40_c94 bl[94] br[94] wl[40] vdd gnd cell_6t
Xbit_r41_c94 bl[94] br[94] wl[41] vdd gnd cell_6t
Xbit_r42_c94 bl[94] br[94] wl[42] vdd gnd cell_6t
Xbit_r43_c94 bl[94] br[94] wl[43] vdd gnd cell_6t
Xbit_r44_c94 bl[94] br[94] wl[44] vdd gnd cell_6t
Xbit_r45_c94 bl[94] br[94] wl[45] vdd gnd cell_6t
Xbit_r46_c94 bl[94] br[94] wl[46] vdd gnd cell_6t
Xbit_r47_c94 bl[94] br[94] wl[47] vdd gnd cell_6t
Xbit_r48_c94 bl[94] br[94] wl[48] vdd gnd cell_6t
Xbit_r49_c94 bl[94] br[94] wl[49] vdd gnd cell_6t
Xbit_r50_c94 bl[94] br[94] wl[50] vdd gnd cell_6t
Xbit_r51_c94 bl[94] br[94] wl[51] vdd gnd cell_6t
Xbit_r52_c94 bl[94] br[94] wl[52] vdd gnd cell_6t
Xbit_r53_c94 bl[94] br[94] wl[53] vdd gnd cell_6t
Xbit_r54_c94 bl[94] br[94] wl[54] vdd gnd cell_6t
Xbit_r55_c94 bl[94] br[94] wl[55] vdd gnd cell_6t
Xbit_r56_c94 bl[94] br[94] wl[56] vdd gnd cell_6t
Xbit_r57_c94 bl[94] br[94] wl[57] vdd gnd cell_6t
Xbit_r58_c94 bl[94] br[94] wl[58] vdd gnd cell_6t
Xbit_r59_c94 bl[94] br[94] wl[59] vdd gnd cell_6t
Xbit_r60_c94 bl[94] br[94] wl[60] vdd gnd cell_6t
Xbit_r61_c94 bl[94] br[94] wl[61] vdd gnd cell_6t
Xbit_r62_c94 bl[94] br[94] wl[62] vdd gnd cell_6t
Xbit_r63_c94 bl[94] br[94] wl[63] vdd gnd cell_6t
Xbit_r64_c94 bl[94] br[94] wl[64] vdd gnd cell_6t
Xbit_r65_c94 bl[94] br[94] wl[65] vdd gnd cell_6t
Xbit_r66_c94 bl[94] br[94] wl[66] vdd gnd cell_6t
Xbit_r67_c94 bl[94] br[94] wl[67] vdd gnd cell_6t
Xbit_r68_c94 bl[94] br[94] wl[68] vdd gnd cell_6t
Xbit_r69_c94 bl[94] br[94] wl[69] vdd gnd cell_6t
Xbit_r70_c94 bl[94] br[94] wl[70] vdd gnd cell_6t
Xbit_r71_c94 bl[94] br[94] wl[71] vdd gnd cell_6t
Xbit_r72_c94 bl[94] br[94] wl[72] vdd gnd cell_6t
Xbit_r73_c94 bl[94] br[94] wl[73] vdd gnd cell_6t
Xbit_r74_c94 bl[94] br[94] wl[74] vdd gnd cell_6t
Xbit_r75_c94 bl[94] br[94] wl[75] vdd gnd cell_6t
Xbit_r76_c94 bl[94] br[94] wl[76] vdd gnd cell_6t
Xbit_r77_c94 bl[94] br[94] wl[77] vdd gnd cell_6t
Xbit_r78_c94 bl[94] br[94] wl[78] vdd gnd cell_6t
Xbit_r79_c94 bl[94] br[94] wl[79] vdd gnd cell_6t
Xbit_r80_c94 bl[94] br[94] wl[80] vdd gnd cell_6t
Xbit_r81_c94 bl[94] br[94] wl[81] vdd gnd cell_6t
Xbit_r82_c94 bl[94] br[94] wl[82] vdd gnd cell_6t
Xbit_r83_c94 bl[94] br[94] wl[83] vdd gnd cell_6t
Xbit_r84_c94 bl[94] br[94] wl[84] vdd gnd cell_6t
Xbit_r85_c94 bl[94] br[94] wl[85] vdd gnd cell_6t
Xbit_r86_c94 bl[94] br[94] wl[86] vdd gnd cell_6t
Xbit_r87_c94 bl[94] br[94] wl[87] vdd gnd cell_6t
Xbit_r88_c94 bl[94] br[94] wl[88] vdd gnd cell_6t
Xbit_r89_c94 bl[94] br[94] wl[89] vdd gnd cell_6t
Xbit_r90_c94 bl[94] br[94] wl[90] vdd gnd cell_6t
Xbit_r91_c94 bl[94] br[94] wl[91] vdd gnd cell_6t
Xbit_r92_c94 bl[94] br[94] wl[92] vdd gnd cell_6t
Xbit_r93_c94 bl[94] br[94] wl[93] vdd gnd cell_6t
Xbit_r94_c94 bl[94] br[94] wl[94] vdd gnd cell_6t
Xbit_r95_c94 bl[94] br[94] wl[95] vdd gnd cell_6t
Xbit_r96_c94 bl[94] br[94] wl[96] vdd gnd cell_6t
Xbit_r97_c94 bl[94] br[94] wl[97] vdd gnd cell_6t
Xbit_r98_c94 bl[94] br[94] wl[98] vdd gnd cell_6t
Xbit_r99_c94 bl[94] br[94] wl[99] vdd gnd cell_6t
Xbit_r100_c94 bl[94] br[94] wl[100] vdd gnd cell_6t
Xbit_r101_c94 bl[94] br[94] wl[101] vdd gnd cell_6t
Xbit_r102_c94 bl[94] br[94] wl[102] vdd gnd cell_6t
Xbit_r103_c94 bl[94] br[94] wl[103] vdd gnd cell_6t
Xbit_r104_c94 bl[94] br[94] wl[104] vdd gnd cell_6t
Xbit_r105_c94 bl[94] br[94] wl[105] vdd gnd cell_6t
Xbit_r106_c94 bl[94] br[94] wl[106] vdd gnd cell_6t
Xbit_r107_c94 bl[94] br[94] wl[107] vdd gnd cell_6t
Xbit_r108_c94 bl[94] br[94] wl[108] vdd gnd cell_6t
Xbit_r109_c94 bl[94] br[94] wl[109] vdd gnd cell_6t
Xbit_r110_c94 bl[94] br[94] wl[110] vdd gnd cell_6t
Xbit_r111_c94 bl[94] br[94] wl[111] vdd gnd cell_6t
Xbit_r112_c94 bl[94] br[94] wl[112] vdd gnd cell_6t
Xbit_r113_c94 bl[94] br[94] wl[113] vdd gnd cell_6t
Xbit_r114_c94 bl[94] br[94] wl[114] vdd gnd cell_6t
Xbit_r115_c94 bl[94] br[94] wl[115] vdd gnd cell_6t
Xbit_r116_c94 bl[94] br[94] wl[116] vdd gnd cell_6t
Xbit_r117_c94 bl[94] br[94] wl[117] vdd gnd cell_6t
Xbit_r118_c94 bl[94] br[94] wl[118] vdd gnd cell_6t
Xbit_r119_c94 bl[94] br[94] wl[119] vdd gnd cell_6t
Xbit_r120_c94 bl[94] br[94] wl[120] vdd gnd cell_6t
Xbit_r121_c94 bl[94] br[94] wl[121] vdd gnd cell_6t
Xbit_r122_c94 bl[94] br[94] wl[122] vdd gnd cell_6t
Xbit_r123_c94 bl[94] br[94] wl[123] vdd gnd cell_6t
Xbit_r124_c94 bl[94] br[94] wl[124] vdd gnd cell_6t
Xbit_r125_c94 bl[94] br[94] wl[125] vdd gnd cell_6t
Xbit_r126_c94 bl[94] br[94] wl[126] vdd gnd cell_6t
Xbit_r127_c94 bl[94] br[94] wl[127] vdd gnd cell_6t
Xbit_r128_c94 bl[94] br[94] wl[128] vdd gnd cell_6t
Xbit_r129_c94 bl[94] br[94] wl[129] vdd gnd cell_6t
Xbit_r130_c94 bl[94] br[94] wl[130] vdd gnd cell_6t
Xbit_r131_c94 bl[94] br[94] wl[131] vdd gnd cell_6t
Xbit_r132_c94 bl[94] br[94] wl[132] vdd gnd cell_6t
Xbit_r133_c94 bl[94] br[94] wl[133] vdd gnd cell_6t
Xbit_r134_c94 bl[94] br[94] wl[134] vdd gnd cell_6t
Xbit_r135_c94 bl[94] br[94] wl[135] vdd gnd cell_6t
Xbit_r136_c94 bl[94] br[94] wl[136] vdd gnd cell_6t
Xbit_r137_c94 bl[94] br[94] wl[137] vdd gnd cell_6t
Xbit_r138_c94 bl[94] br[94] wl[138] vdd gnd cell_6t
Xbit_r139_c94 bl[94] br[94] wl[139] vdd gnd cell_6t
Xbit_r140_c94 bl[94] br[94] wl[140] vdd gnd cell_6t
Xbit_r141_c94 bl[94] br[94] wl[141] vdd gnd cell_6t
Xbit_r142_c94 bl[94] br[94] wl[142] vdd gnd cell_6t
Xbit_r143_c94 bl[94] br[94] wl[143] vdd gnd cell_6t
Xbit_r144_c94 bl[94] br[94] wl[144] vdd gnd cell_6t
Xbit_r145_c94 bl[94] br[94] wl[145] vdd gnd cell_6t
Xbit_r146_c94 bl[94] br[94] wl[146] vdd gnd cell_6t
Xbit_r147_c94 bl[94] br[94] wl[147] vdd gnd cell_6t
Xbit_r148_c94 bl[94] br[94] wl[148] vdd gnd cell_6t
Xbit_r149_c94 bl[94] br[94] wl[149] vdd gnd cell_6t
Xbit_r150_c94 bl[94] br[94] wl[150] vdd gnd cell_6t
Xbit_r151_c94 bl[94] br[94] wl[151] vdd gnd cell_6t
Xbit_r152_c94 bl[94] br[94] wl[152] vdd gnd cell_6t
Xbit_r153_c94 bl[94] br[94] wl[153] vdd gnd cell_6t
Xbit_r154_c94 bl[94] br[94] wl[154] vdd gnd cell_6t
Xbit_r155_c94 bl[94] br[94] wl[155] vdd gnd cell_6t
Xbit_r156_c94 bl[94] br[94] wl[156] vdd gnd cell_6t
Xbit_r157_c94 bl[94] br[94] wl[157] vdd gnd cell_6t
Xbit_r158_c94 bl[94] br[94] wl[158] vdd gnd cell_6t
Xbit_r159_c94 bl[94] br[94] wl[159] vdd gnd cell_6t
Xbit_r160_c94 bl[94] br[94] wl[160] vdd gnd cell_6t
Xbit_r161_c94 bl[94] br[94] wl[161] vdd gnd cell_6t
Xbit_r162_c94 bl[94] br[94] wl[162] vdd gnd cell_6t
Xbit_r163_c94 bl[94] br[94] wl[163] vdd gnd cell_6t
Xbit_r164_c94 bl[94] br[94] wl[164] vdd gnd cell_6t
Xbit_r165_c94 bl[94] br[94] wl[165] vdd gnd cell_6t
Xbit_r166_c94 bl[94] br[94] wl[166] vdd gnd cell_6t
Xbit_r167_c94 bl[94] br[94] wl[167] vdd gnd cell_6t
Xbit_r168_c94 bl[94] br[94] wl[168] vdd gnd cell_6t
Xbit_r169_c94 bl[94] br[94] wl[169] vdd gnd cell_6t
Xbit_r170_c94 bl[94] br[94] wl[170] vdd gnd cell_6t
Xbit_r171_c94 bl[94] br[94] wl[171] vdd gnd cell_6t
Xbit_r172_c94 bl[94] br[94] wl[172] vdd gnd cell_6t
Xbit_r173_c94 bl[94] br[94] wl[173] vdd gnd cell_6t
Xbit_r174_c94 bl[94] br[94] wl[174] vdd gnd cell_6t
Xbit_r175_c94 bl[94] br[94] wl[175] vdd gnd cell_6t
Xbit_r176_c94 bl[94] br[94] wl[176] vdd gnd cell_6t
Xbit_r177_c94 bl[94] br[94] wl[177] vdd gnd cell_6t
Xbit_r178_c94 bl[94] br[94] wl[178] vdd gnd cell_6t
Xbit_r179_c94 bl[94] br[94] wl[179] vdd gnd cell_6t
Xbit_r180_c94 bl[94] br[94] wl[180] vdd gnd cell_6t
Xbit_r181_c94 bl[94] br[94] wl[181] vdd gnd cell_6t
Xbit_r182_c94 bl[94] br[94] wl[182] vdd gnd cell_6t
Xbit_r183_c94 bl[94] br[94] wl[183] vdd gnd cell_6t
Xbit_r184_c94 bl[94] br[94] wl[184] vdd gnd cell_6t
Xbit_r185_c94 bl[94] br[94] wl[185] vdd gnd cell_6t
Xbit_r186_c94 bl[94] br[94] wl[186] vdd gnd cell_6t
Xbit_r187_c94 bl[94] br[94] wl[187] vdd gnd cell_6t
Xbit_r188_c94 bl[94] br[94] wl[188] vdd gnd cell_6t
Xbit_r189_c94 bl[94] br[94] wl[189] vdd gnd cell_6t
Xbit_r190_c94 bl[94] br[94] wl[190] vdd gnd cell_6t
Xbit_r191_c94 bl[94] br[94] wl[191] vdd gnd cell_6t
Xbit_r192_c94 bl[94] br[94] wl[192] vdd gnd cell_6t
Xbit_r193_c94 bl[94] br[94] wl[193] vdd gnd cell_6t
Xbit_r194_c94 bl[94] br[94] wl[194] vdd gnd cell_6t
Xbit_r195_c94 bl[94] br[94] wl[195] vdd gnd cell_6t
Xbit_r196_c94 bl[94] br[94] wl[196] vdd gnd cell_6t
Xbit_r197_c94 bl[94] br[94] wl[197] vdd gnd cell_6t
Xbit_r198_c94 bl[94] br[94] wl[198] vdd gnd cell_6t
Xbit_r199_c94 bl[94] br[94] wl[199] vdd gnd cell_6t
Xbit_r200_c94 bl[94] br[94] wl[200] vdd gnd cell_6t
Xbit_r201_c94 bl[94] br[94] wl[201] vdd gnd cell_6t
Xbit_r202_c94 bl[94] br[94] wl[202] vdd gnd cell_6t
Xbit_r203_c94 bl[94] br[94] wl[203] vdd gnd cell_6t
Xbit_r204_c94 bl[94] br[94] wl[204] vdd gnd cell_6t
Xbit_r205_c94 bl[94] br[94] wl[205] vdd gnd cell_6t
Xbit_r206_c94 bl[94] br[94] wl[206] vdd gnd cell_6t
Xbit_r207_c94 bl[94] br[94] wl[207] vdd gnd cell_6t
Xbit_r208_c94 bl[94] br[94] wl[208] vdd gnd cell_6t
Xbit_r209_c94 bl[94] br[94] wl[209] vdd gnd cell_6t
Xbit_r210_c94 bl[94] br[94] wl[210] vdd gnd cell_6t
Xbit_r211_c94 bl[94] br[94] wl[211] vdd gnd cell_6t
Xbit_r212_c94 bl[94] br[94] wl[212] vdd gnd cell_6t
Xbit_r213_c94 bl[94] br[94] wl[213] vdd gnd cell_6t
Xbit_r214_c94 bl[94] br[94] wl[214] vdd gnd cell_6t
Xbit_r215_c94 bl[94] br[94] wl[215] vdd gnd cell_6t
Xbit_r216_c94 bl[94] br[94] wl[216] vdd gnd cell_6t
Xbit_r217_c94 bl[94] br[94] wl[217] vdd gnd cell_6t
Xbit_r218_c94 bl[94] br[94] wl[218] vdd gnd cell_6t
Xbit_r219_c94 bl[94] br[94] wl[219] vdd gnd cell_6t
Xbit_r220_c94 bl[94] br[94] wl[220] vdd gnd cell_6t
Xbit_r221_c94 bl[94] br[94] wl[221] vdd gnd cell_6t
Xbit_r222_c94 bl[94] br[94] wl[222] vdd gnd cell_6t
Xbit_r223_c94 bl[94] br[94] wl[223] vdd gnd cell_6t
Xbit_r224_c94 bl[94] br[94] wl[224] vdd gnd cell_6t
Xbit_r225_c94 bl[94] br[94] wl[225] vdd gnd cell_6t
Xbit_r226_c94 bl[94] br[94] wl[226] vdd gnd cell_6t
Xbit_r227_c94 bl[94] br[94] wl[227] vdd gnd cell_6t
Xbit_r228_c94 bl[94] br[94] wl[228] vdd gnd cell_6t
Xbit_r229_c94 bl[94] br[94] wl[229] vdd gnd cell_6t
Xbit_r230_c94 bl[94] br[94] wl[230] vdd gnd cell_6t
Xbit_r231_c94 bl[94] br[94] wl[231] vdd gnd cell_6t
Xbit_r232_c94 bl[94] br[94] wl[232] vdd gnd cell_6t
Xbit_r233_c94 bl[94] br[94] wl[233] vdd gnd cell_6t
Xbit_r234_c94 bl[94] br[94] wl[234] vdd gnd cell_6t
Xbit_r235_c94 bl[94] br[94] wl[235] vdd gnd cell_6t
Xbit_r236_c94 bl[94] br[94] wl[236] vdd gnd cell_6t
Xbit_r237_c94 bl[94] br[94] wl[237] vdd gnd cell_6t
Xbit_r238_c94 bl[94] br[94] wl[238] vdd gnd cell_6t
Xbit_r239_c94 bl[94] br[94] wl[239] vdd gnd cell_6t
Xbit_r240_c94 bl[94] br[94] wl[240] vdd gnd cell_6t
Xbit_r241_c94 bl[94] br[94] wl[241] vdd gnd cell_6t
Xbit_r242_c94 bl[94] br[94] wl[242] vdd gnd cell_6t
Xbit_r243_c94 bl[94] br[94] wl[243] vdd gnd cell_6t
Xbit_r244_c94 bl[94] br[94] wl[244] vdd gnd cell_6t
Xbit_r245_c94 bl[94] br[94] wl[245] vdd gnd cell_6t
Xbit_r246_c94 bl[94] br[94] wl[246] vdd gnd cell_6t
Xbit_r247_c94 bl[94] br[94] wl[247] vdd gnd cell_6t
Xbit_r248_c94 bl[94] br[94] wl[248] vdd gnd cell_6t
Xbit_r249_c94 bl[94] br[94] wl[249] vdd gnd cell_6t
Xbit_r250_c94 bl[94] br[94] wl[250] vdd gnd cell_6t
Xbit_r251_c94 bl[94] br[94] wl[251] vdd gnd cell_6t
Xbit_r252_c94 bl[94] br[94] wl[252] vdd gnd cell_6t
Xbit_r253_c94 bl[94] br[94] wl[253] vdd gnd cell_6t
Xbit_r254_c94 bl[94] br[94] wl[254] vdd gnd cell_6t
Xbit_r255_c94 bl[94] br[94] wl[255] vdd gnd cell_6t
Xbit_r0_c95 bl[95] br[95] wl[0] vdd gnd cell_6t
Xbit_r1_c95 bl[95] br[95] wl[1] vdd gnd cell_6t
Xbit_r2_c95 bl[95] br[95] wl[2] vdd gnd cell_6t
Xbit_r3_c95 bl[95] br[95] wl[3] vdd gnd cell_6t
Xbit_r4_c95 bl[95] br[95] wl[4] vdd gnd cell_6t
Xbit_r5_c95 bl[95] br[95] wl[5] vdd gnd cell_6t
Xbit_r6_c95 bl[95] br[95] wl[6] vdd gnd cell_6t
Xbit_r7_c95 bl[95] br[95] wl[7] vdd gnd cell_6t
Xbit_r8_c95 bl[95] br[95] wl[8] vdd gnd cell_6t
Xbit_r9_c95 bl[95] br[95] wl[9] vdd gnd cell_6t
Xbit_r10_c95 bl[95] br[95] wl[10] vdd gnd cell_6t
Xbit_r11_c95 bl[95] br[95] wl[11] vdd gnd cell_6t
Xbit_r12_c95 bl[95] br[95] wl[12] vdd gnd cell_6t
Xbit_r13_c95 bl[95] br[95] wl[13] vdd gnd cell_6t
Xbit_r14_c95 bl[95] br[95] wl[14] vdd gnd cell_6t
Xbit_r15_c95 bl[95] br[95] wl[15] vdd gnd cell_6t
Xbit_r16_c95 bl[95] br[95] wl[16] vdd gnd cell_6t
Xbit_r17_c95 bl[95] br[95] wl[17] vdd gnd cell_6t
Xbit_r18_c95 bl[95] br[95] wl[18] vdd gnd cell_6t
Xbit_r19_c95 bl[95] br[95] wl[19] vdd gnd cell_6t
Xbit_r20_c95 bl[95] br[95] wl[20] vdd gnd cell_6t
Xbit_r21_c95 bl[95] br[95] wl[21] vdd gnd cell_6t
Xbit_r22_c95 bl[95] br[95] wl[22] vdd gnd cell_6t
Xbit_r23_c95 bl[95] br[95] wl[23] vdd gnd cell_6t
Xbit_r24_c95 bl[95] br[95] wl[24] vdd gnd cell_6t
Xbit_r25_c95 bl[95] br[95] wl[25] vdd gnd cell_6t
Xbit_r26_c95 bl[95] br[95] wl[26] vdd gnd cell_6t
Xbit_r27_c95 bl[95] br[95] wl[27] vdd gnd cell_6t
Xbit_r28_c95 bl[95] br[95] wl[28] vdd gnd cell_6t
Xbit_r29_c95 bl[95] br[95] wl[29] vdd gnd cell_6t
Xbit_r30_c95 bl[95] br[95] wl[30] vdd gnd cell_6t
Xbit_r31_c95 bl[95] br[95] wl[31] vdd gnd cell_6t
Xbit_r32_c95 bl[95] br[95] wl[32] vdd gnd cell_6t
Xbit_r33_c95 bl[95] br[95] wl[33] vdd gnd cell_6t
Xbit_r34_c95 bl[95] br[95] wl[34] vdd gnd cell_6t
Xbit_r35_c95 bl[95] br[95] wl[35] vdd gnd cell_6t
Xbit_r36_c95 bl[95] br[95] wl[36] vdd gnd cell_6t
Xbit_r37_c95 bl[95] br[95] wl[37] vdd gnd cell_6t
Xbit_r38_c95 bl[95] br[95] wl[38] vdd gnd cell_6t
Xbit_r39_c95 bl[95] br[95] wl[39] vdd gnd cell_6t
Xbit_r40_c95 bl[95] br[95] wl[40] vdd gnd cell_6t
Xbit_r41_c95 bl[95] br[95] wl[41] vdd gnd cell_6t
Xbit_r42_c95 bl[95] br[95] wl[42] vdd gnd cell_6t
Xbit_r43_c95 bl[95] br[95] wl[43] vdd gnd cell_6t
Xbit_r44_c95 bl[95] br[95] wl[44] vdd gnd cell_6t
Xbit_r45_c95 bl[95] br[95] wl[45] vdd gnd cell_6t
Xbit_r46_c95 bl[95] br[95] wl[46] vdd gnd cell_6t
Xbit_r47_c95 bl[95] br[95] wl[47] vdd gnd cell_6t
Xbit_r48_c95 bl[95] br[95] wl[48] vdd gnd cell_6t
Xbit_r49_c95 bl[95] br[95] wl[49] vdd gnd cell_6t
Xbit_r50_c95 bl[95] br[95] wl[50] vdd gnd cell_6t
Xbit_r51_c95 bl[95] br[95] wl[51] vdd gnd cell_6t
Xbit_r52_c95 bl[95] br[95] wl[52] vdd gnd cell_6t
Xbit_r53_c95 bl[95] br[95] wl[53] vdd gnd cell_6t
Xbit_r54_c95 bl[95] br[95] wl[54] vdd gnd cell_6t
Xbit_r55_c95 bl[95] br[95] wl[55] vdd gnd cell_6t
Xbit_r56_c95 bl[95] br[95] wl[56] vdd gnd cell_6t
Xbit_r57_c95 bl[95] br[95] wl[57] vdd gnd cell_6t
Xbit_r58_c95 bl[95] br[95] wl[58] vdd gnd cell_6t
Xbit_r59_c95 bl[95] br[95] wl[59] vdd gnd cell_6t
Xbit_r60_c95 bl[95] br[95] wl[60] vdd gnd cell_6t
Xbit_r61_c95 bl[95] br[95] wl[61] vdd gnd cell_6t
Xbit_r62_c95 bl[95] br[95] wl[62] vdd gnd cell_6t
Xbit_r63_c95 bl[95] br[95] wl[63] vdd gnd cell_6t
Xbit_r64_c95 bl[95] br[95] wl[64] vdd gnd cell_6t
Xbit_r65_c95 bl[95] br[95] wl[65] vdd gnd cell_6t
Xbit_r66_c95 bl[95] br[95] wl[66] vdd gnd cell_6t
Xbit_r67_c95 bl[95] br[95] wl[67] vdd gnd cell_6t
Xbit_r68_c95 bl[95] br[95] wl[68] vdd gnd cell_6t
Xbit_r69_c95 bl[95] br[95] wl[69] vdd gnd cell_6t
Xbit_r70_c95 bl[95] br[95] wl[70] vdd gnd cell_6t
Xbit_r71_c95 bl[95] br[95] wl[71] vdd gnd cell_6t
Xbit_r72_c95 bl[95] br[95] wl[72] vdd gnd cell_6t
Xbit_r73_c95 bl[95] br[95] wl[73] vdd gnd cell_6t
Xbit_r74_c95 bl[95] br[95] wl[74] vdd gnd cell_6t
Xbit_r75_c95 bl[95] br[95] wl[75] vdd gnd cell_6t
Xbit_r76_c95 bl[95] br[95] wl[76] vdd gnd cell_6t
Xbit_r77_c95 bl[95] br[95] wl[77] vdd gnd cell_6t
Xbit_r78_c95 bl[95] br[95] wl[78] vdd gnd cell_6t
Xbit_r79_c95 bl[95] br[95] wl[79] vdd gnd cell_6t
Xbit_r80_c95 bl[95] br[95] wl[80] vdd gnd cell_6t
Xbit_r81_c95 bl[95] br[95] wl[81] vdd gnd cell_6t
Xbit_r82_c95 bl[95] br[95] wl[82] vdd gnd cell_6t
Xbit_r83_c95 bl[95] br[95] wl[83] vdd gnd cell_6t
Xbit_r84_c95 bl[95] br[95] wl[84] vdd gnd cell_6t
Xbit_r85_c95 bl[95] br[95] wl[85] vdd gnd cell_6t
Xbit_r86_c95 bl[95] br[95] wl[86] vdd gnd cell_6t
Xbit_r87_c95 bl[95] br[95] wl[87] vdd gnd cell_6t
Xbit_r88_c95 bl[95] br[95] wl[88] vdd gnd cell_6t
Xbit_r89_c95 bl[95] br[95] wl[89] vdd gnd cell_6t
Xbit_r90_c95 bl[95] br[95] wl[90] vdd gnd cell_6t
Xbit_r91_c95 bl[95] br[95] wl[91] vdd gnd cell_6t
Xbit_r92_c95 bl[95] br[95] wl[92] vdd gnd cell_6t
Xbit_r93_c95 bl[95] br[95] wl[93] vdd gnd cell_6t
Xbit_r94_c95 bl[95] br[95] wl[94] vdd gnd cell_6t
Xbit_r95_c95 bl[95] br[95] wl[95] vdd gnd cell_6t
Xbit_r96_c95 bl[95] br[95] wl[96] vdd gnd cell_6t
Xbit_r97_c95 bl[95] br[95] wl[97] vdd gnd cell_6t
Xbit_r98_c95 bl[95] br[95] wl[98] vdd gnd cell_6t
Xbit_r99_c95 bl[95] br[95] wl[99] vdd gnd cell_6t
Xbit_r100_c95 bl[95] br[95] wl[100] vdd gnd cell_6t
Xbit_r101_c95 bl[95] br[95] wl[101] vdd gnd cell_6t
Xbit_r102_c95 bl[95] br[95] wl[102] vdd gnd cell_6t
Xbit_r103_c95 bl[95] br[95] wl[103] vdd gnd cell_6t
Xbit_r104_c95 bl[95] br[95] wl[104] vdd gnd cell_6t
Xbit_r105_c95 bl[95] br[95] wl[105] vdd gnd cell_6t
Xbit_r106_c95 bl[95] br[95] wl[106] vdd gnd cell_6t
Xbit_r107_c95 bl[95] br[95] wl[107] vdd gnd cell_6t
Xbit_r108_c95 bl[95] br[95] wl[108] vdd gnd cell_6t
Xbit_r109_c95 bl[95] br[95] wl[109] vdd gnd cell_6t
Xbit_r110_c95 bl[95] br[95] wl[110] vdd gnd cell_6t
Xbit_r111_c95 bl[95] br[95] wl[111] vdd gnd cell_6t
Xbit_r112_c95 bl[95] br[95] wl[112] vdd gnd cell_6t
Xbit_r113_c95 bl[95] br[95] wl[113] vdd gnd cell_6t
Xbit_r114_c95 bl[95] br[95] wl[114] vdd gnd cell_6t
Xbit_r115_c95 bl[95] br[95] wl[115] vdd gnd cell_6t
Xbit_r116_c95 bl[95] br[95] wl[116] vdd gnd cell_6t
Xbit_r117_c95 bl[95] br[95] wl[117] vdd gnd cell_6t
Xbit_r118_c95 bl[95] br[95] wl[118] vdd gnd cell_6t
Xbit_r119_c95 bl[95] br[95] wl[119] vdd gnd cell_6t
Xbit_r120_c95 bl[95] br[95] wl[120] vdd gnd cell_6t
Xbit_r121_c95 bl[95] br[95] wl[121] vdd gnd cell_6t
Xbit_r122_c95 bl[95] br[95] wl[122] vdd gnd cell_6t
Xbit_r123_c95 bl[95] br[95] wl[123] vdd gnd cell_6t
Xbit_r124_c95 bl[95] br[95] wl[124] vdd gnd cell_6t
Xbit_r125_c95 bl[95] br[95] wl[125] vdd gnd cell_6t
Xbit_r126_c95 bl[95] br[95] wl[126] vdd gnd cell_6t
Xbit_r127_c95 bl[95] br[95] wl[127] vdd gnd cell_6t
Xbit_r128_c95 bl[95] br[95] wl[128] vdd gnd cell_6t
Xbit_r129_c95 bl[95] br[95] wl[129] vdd gnd cell_6t
Xbit_r130_c95 bl[95] br[95] wl[130] vdd gnd cell_6t
Xbit_r131_c95 bl[95] br[95] wl[131] vdd gnd cell_6t
Xbit_r132_c95 bl[95] br[95] wl[132] vdd gnd cell_6t
Xbit_r133_c95 bl[95] br[95] wl[133] vdd gnd cell_6t
Xbit_r134_c95 bl[95] br[95] wl[134] vdd gnd cell_6t
Xbit_r135_c95 bl[95] br[95] wl[135] vdd gnd cell_6t
Xbit_r136_c95 bl[95] br[95] wl[136] vdd gnd cell_6t
Xbit_r137_c95 bl[95] br[95] wl[137] vdd gnd cell_6t
Xbit_r138_c95 bl[95] br[95] wl[138] vdd gnd cell_6t
Xbit_r139_c95 bl[95] br[95] wl[139] vdd gnd cell_6t
Xbit_r140_c95 bl[95] br[95] wl[140] vdd gnd cell_6t
Xbit_r141_c95 bl[95] br[95] wl[141] vdd gnd cell_6t
Xbit_r142_c95 bl[95] br[95] wl[142] vdd gnd cell_6t
Xbit_r143_c95 bl[95] br[95] wl[143] vdd gnd cell_6t
Xbit_r144_c95 bl[95] br[95] wl[144] vdd gnd cell_6t
Xbit_r145_c95 bl[95] br[95] wl[145] vdd gnd cell_6t
Xbit_r146_c95 bl[95] br[95] wl[146] vdd gnd cell_6t
Xbit_r147_c95 bl[95] br[95] wl[147] vdd gnd cell_6t
Xbit_r148_c95 bl[95] br[95] wl[148] vdd gnd cell_6t
Xbit_r149_c95 bl[95] br[95] wl[149] vdd gnd cell_6t
Xbit_r150_c95 bl[95] br[95] wl[150] vdd gnd cell_6t
Xbit_r151_c95 bl[95] br[95] wl[151] vdd gnd cell_6t
Xbit_r152_c95 bl[95] br[95] wl[152] vdd gnd cell_6t
Xbit_r153_c95 bl[95] br[95] wl[153] vdd gnd cell_6t
Xbit_r154_c95 bl[95] br[95] wl[154] vdd gnd cell_6t
Xbit_r155_c95 bl[95] br[95] wl[155] vdd gnd cell_6t
Xbit_r156_c95 bl[95] br[95] wl[156] vdd gnd cell_6t
Xbit_r157_c95 bl[95] br[95] wl[157] vdd gnd cell_6t
Xbit_r158_c95 bl[95] br[95] wl[158] vdd gnd cell_6t
Xbit_r159_c95 bl[95] br[95] wl[159] vdd gnd cell_6t
Xbit_r160_c95 bl[95] br[95] wl[160] vdd gnd cell_6t
Xbit_r161_c95 bl[95] br[95] wl[161] vdd gnd cell_6t
Xbit_r162_c95 bl[95] br[95] wl[162] vdd gnd cell_6t
Xbit_r163_c95 bl[95] br[95] wl[163] vdd gnd cell_6t
Xbit_r164_c95 bl[95] br[95] wl[164] vdd gnd cell_6t
Xbit_r165_c95 bl[95] br[95] wl[165] vdd gnd cell_6t
Xbit_r166_c95 bl[95] br[95] wl[166] vdd gnd cell_6t
Xbit_r167_c95 bl[95] br[95] wl[167] vdd gnd cell_6t
Xbit_r168_c95 bl[95] br[95] wl[168] vdd gnd cell_6t
Xbit_r169_c95 bl[95] br[95] wl[169] vdd gnd cell_6t
Xbit_r170_c95 bl[95] br[95] wl[170] vdd gnd cell_6t
Xbit_r171_c95 bl[95] br[95] wl[171] vdd gnd cell_6t
Xbit_r172_c95 bl[95] br[95] wl[172] vdd gnd cell_6t
Xbit_r173_c95 bl[95] br[95] wl[173] vdd gnd cell_6t
Xbit_r174_c95 bl[95] br[95] wl[174] vdd gnd cell_6t
Xbit_r175_c95 bl[95] br[95] wl[175] vdd gnd cell_6t
Xbit_r176_c95 bl[95] br[95] wl[176] vdd gnd cell_6t
Xbit_r177_c95 bl[95] br[95] wl[177] vdd gnd cell_6t
Xbit_r178_c95 bl[95] br[95] wl[178] vdd gnd cell_6t
Xbit_r179_c95 bl[95] br[95] wl[179] vdd gnd cell_6t
Xbit_r180_c95 bl[95] br[95] wl[180] vdd gnd cell_6t
Xbit_r181_c95 bl[95] br[95] wl[181] vdd gnd cell_6t
Xbit_r182_c95 bl[95] br[95] wl[182] vdd gnd cell_6t
Xbit_r183_c95 bl[95] br[95] wl[183] vdd gnd cell_6t
Xbit_r184_c95 bl[95] br[95] wl[184] vdd gnd cell_6t
Xbit_r185_c95 bl[95] br[95] wl[185] vdd gnd cell_6t
Xbit_r186_c95 bl[95] br[95] wl[186] vdd gnd cell_6t
Xbit_r187_c95 bl[95] br[95] wl[187] vdd gnd cell_6t
Xbit_r188_c95 bl[95] br[95] wl[188] vdd gnd cell_6t
Xbit_r189_c95 bl[95] br[95] wl[189] vdd gnd cell_6t
Xbit_r190_c95 bl[95] br[95] wl[190] vdd gnd cell_6t
Xbit_r191_c95 bl[95] br[95] wl[191] vdd gnd cell_6t
Xbit_r192_c95 bl[95] br[95] wl[192] vdd gnd cell_6t
Xbit_r193_c95 bl[95] br[95] wl[193] vdd gnd cell_6t
Xbit_r194_c95 bl[95] br[95] wl[194] vdd gnd cell_6t
Xbit_r195_c95 bl[95] br[95] wl[195] vdd gnd cell_6t
Xbit_r196_c95 bl[95] br[95] wl[196] vdd gnd cell_6t
Xbit_r197_c95 bl[95] br[95] wl[197] vdd gnd cell_6t
Xbit_r198_c95 bl[95] br[95] wl[198] vdd gnd cell_6t
Xbit_r199_c95 bl[95] br[95] wl[199] vdd gnd cell_6t
Xbit_r200_c95 bl[95] br[95] wl[200] vdd gnd cell_6t
Xbit_r201_c95 bl[95] br[95] wl[201] vdd gnd cell_6t
Xbit_r202_c95 bl[95] br[95] wl[202] vdd gnd cell_6t
Xbit_r203_c95 bl[95] br[95] wl[203] vdd gnd cell_6t
Xbit_r204_c95 bl[95] br[95] wl[204] vdd gnd cell_6t
Xbit_r205_c95 bl[95] br[95] wl[205] vdd gnd cell_6t
Xbit_r206_c95 bl[95] br[95] wl[206] vdd gnd cell_6t
Xbit_r207_c95 bl[95] br[95] wl[207] vdd gnd cell_6t
Xbit_r208_c95 bl[95] br[95] wl[208] vdd gnd cell_6t
Xbit_r209_c95 bl[95] br[95] wl[209] vdd gnd cell_6t
Xbit_r210_c95 bl[95] br[95] wl[210] vdd gnd cell_6t
Xbit_r211_c95 bl[95] br[95] wl[211] vdd gnd cell_6t
Xbit_r212_c95 bl[95] br[95] wl[212] vdd gnd cell_6t
Xbit_r213_c95 bl[95] br[95] wl[213] vdd gnd cell_6t
Xbit_r214_c95 bl[95] br[95] wl[214] vdd gnd cell_6t
Xbit_r215_c95 bl[95] br[95] wl[215] vdd gnd cell_6t
Xbit_r216_c95 bl[95] br[95] wl[216] vdd gnd cell_6t
Xbit_r217_c95 bl[95] br[95] wl[217] vdd gnd cell_6t
Xbit_r218_c95 bl[95] br[95] wl[218] vdd gnd cell_6t
Xbit_r219_c95 bl[95] br[95] wl[219] vdd gnd cell_6t
Xbit_r220_c95 bl[95] br[95] wl[220] vdd gnd cell_6t
Xbit_r221_c95 bl[95] br[95] wl[221] vdd gnd cell_6t
Xbit_r222_c95 bl[95] br[95] wl[222] vdd gnd cell_6t
Xbit_r223_c95 bl[95] br[95] wl[223] vdd gnd cell_6t
Xbit_r224_c95 bl[95] br[95] wl[224] vdd gnd cell_6t
Xbit_r225_c95 bl[95] br[95] wl[225] vdd gnd cell_6t
Xbit_r226_c95 bl[95] br[95] wl[226] vdd gnd cell_6t
Xbit_r227_c95 bl[95] br[95] wl[227] vdd gnd cell_6t
Xbit_r228_c95 bl[95] br[95] wl[228] vdd gnd cell_6t
Xbit_r229_c95 bl[95] br[95] wl[229] vdd gnd cell_6t
Xbit_r230_c95 bl[95] br[95] wl[230] vdd gnd cell_6t
Xbit_r231_c95 bl[95] br[95] wl[231] vdd gnd cell_6t
Xbit_r232_c95 bl[95] br[95] wl[232] vdd gnd cell_6t
Xbit_r233_c95 bl[95] br[95] wl[233] vdd gnd cell_6t
Xbit_r234_c95 bl[95] br[95] wl[234] vdd gnd cell_6t
Xbit_r235_c95 bl[95] br[95] wl[235] vdd gnd cell_6t
Xbit_r236_c95 bl[95] br[95] wl[236] vdd gnd cell_6t
Xbit_r237_c95 bl[95] br[95] wl[237] vdd gnd cell_6t
Xbit_r238_c95 bl[95] br[95] wl[238] vdd gnd cell_6t
Xbit_r239_c95 bl[95] br[95] wl[239] vdd gnd cell_6t
Xbit_r240_c95 bl[95] br[95] wl[240] vdd gnd cell_6t
Xbit_r241_c95 bl[95] br[95] wl[241] vdd gnd cell_6t
Xbit_r242_c95 bl[95] br[95] wl[242] vdd gnd cell_6t
Xbit_r243_c95 bl[95] br[95] wl[243] vdd gnd cell_6t
Xbit_r244_c95 bl[95] br[95] wl[244] vdd gnd cell_6t
Xbit_r245_c95 bl[95] br[95] wl[245] vdd gnd cell_6t
Xbit_r246_c95 bl[95] br[95] wl[246] vdd gnd cell_6t
Xbit_r247_c95 bl[95] br[95] wl[247] vdd gnd cell_6t
Xbit_r248_c95 bl[95] br[95] wl[248] vdd gnd cell_6t
Xbit_r249_c95 bl[95] br[95] wl[249] vdd gnd cell_6t
Xbit_r250_c95 bl[95] br[95] wl[250] vdd gnd cell_6t
Xbit_r251_c95 bl[95] br[95] wl[251] vdd gnd cell_6t
Xbit_r252_c95 bl[95] br[95] wl[252] vdd gnd cell_6t
Xbit_r253_c95 bl[95] br[95] wl[253] vdd gnd cell_6t
Xbit_r254_c95 bl[95] br[95] wl[254] vdd gnd cell_6t
Xbit_r255_c95 bl[95] br[95] wl[255] vdd gnd cell_6t
Xbit_r0_c96 bl[96] br[96] wl[0] vdd gnd cell_6t
Xbit_r1_c96 bl[96] br[96] wl[1] vdd gnd cell_6t
Xbit_r2_c96 bl[96] br[96] wl[2] vdd gnd cell_6t
Xbit_r3_c96 bl[96] br[96] wl[3] vdd gnd cell_6t
Xbit_r4_c96 bl[96] br[96] wl[4] vdd gnd cell_6t
Xbit_r5_c96 bl[96] br[96] wl[5] vdd gnd cell_6t
Xbit_r6_c96 bl[96] br[96] wl[6] vdd gnd cell_6t
Xbit_r7_c96 bl[96] br[96] wl[7] vdd gnd cell_6t
Xbit_r8_c96 bl[96] br[96] wl[8] vdd gnd cell_6t
Xbit_r9_c96 bl[96] br[96] wl[9] vdd gnd cell_6t
Xbit_r10_c96 bl[96] br[96] wl[10] vdd gnd cell_6t
Xbit_r11_c96 bl[96] br[96] wl[11] vdd gnd cell_6t
Xbit_r12_c96 bl[96] br[96] wl[12] vdd gnd cell_6t
Xbit_r13_c96 bl[96] br[96] wl[13] vdd gnd cell_6t
Xbit_r14_c96 bl[96] br[96] wl[14] vdd gnd cell_6t
Xbit_r15_c96 bl[96] br[96] wl[15] vdd gnd cell_6t
Xbit_r16_c96 bl[96] br[96] wl[16] vdd gnd cell_6t
Xbit_r17_c96 bl[96] br[96] wl[17] vdd gnd cell_6t
Xbit_r18_c96 bl[96] br[96] wl[18] vdd gnd cell_6t
Xbit_r19_c96 bl[96] br[96] wl[19] vdd gnd cell_6t
Xbit_r20_c96 bl[96] br[96] wl[20] vdd gnd cell_6t
Xbit_r21_c96 bl[96] br[96] wl[21] vdd gnd cell_6t
Xbit_r22_c96 bl[96] br[96] wl[22] vdd gnd cell_6t
Xbit_r23_c96 bl[96] br[96] wl[23] vdd gnd cell_6t
Xbit_r24_c96 bl[96] br[96] wl[24] vdd gnd cell_6t
Xbit_r25_c96 bl[96] br[96] wl[25] vdd gnd cell_6t
Xbit_r26_c96 bl[96] br[96] wl[26] vdd gnd cell_6t
Xbit_r27_c96 bl[96] br[96] wl[27] vdd gnd cell_6t
Xbit_r28_c96 bl[96] br[96] wl[28] vdd gnd cell_6t
Xbit_r29_c96 bl[96] br[96] wl[29] vdd gnd cell_6t
Xbit_r30_c96 bl[96] br[96] wl[30] vdd gnd cell_6t
Xbit_r31_c96 bl[96] br[96] wl[31] vdd gnd cell_6t
Xbit_r32_c96 bl[96] br[96] wl[32] vdd gnd cell_6t
Xbit_r33_c96 bl[96] br[96] wl[33] vdd gnd cell_6t
Xbit_r34_c96 bl[96] br[96] wl[34] vdd gnd cell_6t
Xbit_r35_c96 bl[96] br[96] wl[35] vdd gnd cell_6t
Xbit_r36_c96 bl[96] br[96] wl[36] vdd gnd cell_6t
Xbit_r37_c96 bl[96] br[96] wl[37] vdd gnd cell_6t
Xbit_r38_c96 bl[96] br[96] wl[38] vdd gnd cell_6t
Xbit_r39_c96 bl[96] br[96] wl[39] vdd gnd cell_6t
Xbit_r40_c96 bl[96] br[96] wl[40] vdd gnd cell_6t
Xbit_r41_c96 bl[96] br[96] wl[41] vdd gnd cell_6t
Xbit_r42_c96 bl[96] br[96] wl[42] vdd gnd cell_6t
Xbit_r43_c96 bl[96] br[96] wl[43] vdd gnd cell_6t
Xbit_r44_c96 bl[96] br[96] wl[44] vdd gnd cell_6t
Xbit_r45_c96 bl[96] br[96] wl[45] vdd gnd cell_6t
Xbit_r46_c96 bl[96] br[96] wl[46] vdd gnd cell_6t
Xbit_r47_c96 bl[96] br[96] wl[47] vdd gnd cell_6t
Xbit_r48_c96 bl[96] br[96] wl[48] vdd gnd cell_6t
Xbit_r49_c96 bl[96] br[96] wl[49] vdd gnd cell_6t
Xbit_r50_c96 bl[96] br[96] wl[50] vdd gnd cell_6t
Xbit_r51_c96 bl[96] br[96] wl[51] vdd gnd cell_6t
Xbit_r52_c96 bl[96] br[96] wl[52] vdd gnd cell_6t
Xbit_r53_c96 bl[96] br[96] wl[53] vdd gnd cell_6t
Xbit_r54_c96 bl[96] br[96] wl[54] vdd gnd cell_6t
Xbit_r55_c96 bl[96] br[96] wl[55] vdd gnd cell_6t
Xbit_r56_c96 bl[96] br[96] wl[56] vdd gnd cell_6t
Xbit_r57_c96 bl[96] br[96] wl[57] vdd gnd cell_6t
Xbit_r58_c96 bl[96] br[96] wl[58] vdd gnd cell_6t
Xbit_r59_c96 bl[96] br[96] wl[59] vdd gnd cell_6t
Xbit_r60_c96 bl[96] br[96] wl[60] vdd gnd cell_6t
Xbit_r61_c96 bl[96] br[96] wl[61] vdd gnd cell_6t
Xbit_r62_c96 bl[96] br[96] wl[62] vdd gnd cell_6t
Xbit_r63_c96 bl[96] br[96] wl[63] vdd gnd cell_6t
Xbit_r64_c96 bl[96] br[96] wl[64] vdd gnd cell_6t
Xbit_r65_c96 bl[96] br[96] wl[65] vdd gnd cell_6t
Xbit_r66_c96 bl[96] br[96] wl[66] vdd gnd cell_6t
Xbit_r67_c96 bl[96] br[96] wl[67] vdd gnd cell_6t
Xbit_r68_c96 bl[96] br[96] wl[68] vdd gnd cell_6t
Xbit_r69_c96 bl[96] br[96] wl[69] vdd gnd cell_6t
Xbit_r70_c96 bl[96] br[96] wl[70] vdd gnd cell_6t
Xbit_r71_c96 bl[96] br[96] wl[71] vdd gnd cell_6t
Xbit_r72_c96 bl[96] br[96] wl[72] vdd gnd cell_6t
Xbit_r73_c96 bl[96] br[96] wl[73] vdd gnd cell_6t
Xbit_r74_c96 bl[96] br[96] wl[74] vdd gnd cell_6t
Xbit_r75_c96 bl[96] br[96] wl[75] vdd gnd cell_6t
Xbit_r76_c96 bl[96] br[96] wl[76] vdd gnd cell_6t
Xbit_r77_c96 bl[96] br[96] wl[77] vdd gnd cell_6t
Xbit_r78_c96 bl[96] br[96] wl[78] vdd gnd cell_6t
Xbit_r79_c96 bl[96] br[96] wl[79] vdd gnd cell_6t
Xbit_r80_c96 bl[96] br[96] wl[80] vdd gnd cell_6t
Xbit_r81_c96 bl[96] br[96] wl[81] vdd gnd cell_6t
Xbit_r82_c96 bl[96] br[96] wl[82] vdd gnd cell_6t
Xbit_r83_c96 bl[96] br[96] wl[83] vdd gnd cell_6t
Xbit_r84_c96 bl[96] br[96] wl[84] vdd gnd cell_6t
Xbit_r85_c96 bl[96] br[96] wl[85] vdd gnd cell_6t
Xbit_r86_c96 bl[96] br[96] wl[86] vdd gnd cell_6t
Xbit_r87_c96 bl[96] br[96] wl[87] vdd gnd cell_6t
Xbit_r88_c96 bl[96] br[96] wl[88] vdd gnd cell_6t
Xbit_r89_c96 bl[96] br[96] wl[89] vdd gnd cell_6t
Xbit_r90_c96 bl[96] br[96] wl[90] vdd gnd cell_6t
Xbit_r91_c96 bl[96] br[96] wl[91] vdd gnd cell_6t
Xbit_r92_c96 bl[96] br[96] wl[92] vdd gnd cell_6t
Xbit_r93_c96 bl[96] br[96] wl[93] vdd gnd cell_6t
Xbit_r94_c96 bl[96] br[96] wl[94] vdd gnd cell_6t
Xbit_r95_c96 bl[96] br[96] wl[95] vdd gnd cell_6t
Xbit_r96_c96 bl[96] br[96] wl[96] vdd gnd cell_6t
Xbit_r97_c96 bl[96] br[96] wl[97] vdd gnd cell_6t
Xbit_r98_c96 bl[96] br[96] wl[98] vdd gnd cell_6t
Xbit_r99_c96 bl[96] br[96] wl[99] vdd gnd cell_6t
Xbit_r100_c96 bl[96] br[96] wl[100] vdd gnd cell_6t
Xbit_r101_c96 bl[96] br[96] wl[101] vdd gnd cell_6t
Xbit_r102_c96 bl[96] br[96] wl[102] vdd gnd cell_6t
Xbit_r103_c96 bl[96] br[96] wl[103] vdd gnd cell_6t
Xbit_r104_c96 bl[96] br[96] wl[104] vdd gnd cell_6t
Xbit_r105_c96 bl[96] br[96] wl[105] vdd gnd cell_6t
Xbit_r106_c96 bl[96] br[96] wl[106] vdd gnd cell_6t
Xbit_r107_c96 bl[96] br[96] wl[107] vdd gnd cell_6t
Xbit_r108_c96 bl[96] br[96] wl[108] vdd gnd cell_6t
Xbit_r109_c96 bl[96] br[96] wl[109] vdd gnd cell_6t
Xbit_r110_c96 bl[96] br[96] wl[110] vdd gnd cell_6t
Xbit_r111_c96 bl[96] br[96] wl[111] vdd gnd cell_6t
Xbit_r112_c96 bl[96] br[96] wl[112] vdd gnd cell_6t
Xbit_r113_c96 bl[96] br[96] wl[113] vdd gnd cell_6t
Xbit_r114_c96 bl[96] br[96] wl[114] vdd gnd cell_6t
Xbit_r115_c96 bl[96] br[96] wl[115] vdd gnd cell_6t
Xbit_r116_c96 bl[96] br[96] wl[116] vdd gnd cell_6t
Xbit_r117_c96 bl[96] br[96] wl[117] vdd gnd cell_6t
Xbit_r118_c96 bl[96] br[96] wl[118] vdd gnd cell_6t
Xbit_r119_c96 bl[96] br[96] wl[119] vdd gnd cell_6t
Xbit_r120_c96 bl[96] br[96] wl[120] vdd gnd cell_6t
Xbit_r121_c96 bl[96] br[96] wl[121] vdd gnd cell_6t
Xbit_r122_c96 bl[96] br[96] wl[122] vdd gnd cell_6t
Xbit_r123_c96 bl[96] br[96] wl[123] vdd gnd cell_6t
Xbit_r124_c96 bl[96] br[96] wl[124] vdd gnd cell_6t
Xbit_r125_c96 bl[96] br[96] wl[125] vdd gnd cell_6t
Xbit_r126_c96 bl[96] br[96] wl[126] vdd gnd cell_6t
Xbit_r127_c96 bl[96] br[96] wl[127] vdd gnd cell_6t
Xbit_r128_c96 bl[96] br[96] wl[128] vdd gnd cell_6t
Xbit_r129_c96 bl[96] br[96] wl[129] vdd gnd cell_6t
Xbit_r130_c96 bl[96] br[96] wl[130] vdd gnd cell_6t
Xbit_r131_c96 bl[96] br[96] wl[131] vdd gnd cell_6t
Xbit_r132_c96 bl[96] br[96] wl[132] vdd gnd cell_6t
Xbit_r133_c96 bl[96] br[96] wl[133] vdd gnd cell_6t
Xbit_r134_c96 bl[96] br[96] wl[134] vdd gnd cell_6t
Xbit_r135_c96 bl[96] br[96] wl[135] vdd gnd cell_6t
Xbit_r136_c96 bl[96] br[96] wl[136] vdd gnd cell_6t
Xbit_r137_c96 bl[96] br[96] wl[137] vdd gnd cell_6t
Xbit_r138_c96 bl[96] br[96] wl[138] vdd gnd cell_6t
Xbit_r139_c96 bl[96] br[96] wl[139] vdd gnd cell_6t
Xbit_r140_c96 bl[96] br[96] wl[140] vdd gnd cell_6t
Xbit_r141_c96 bl[96] br[96] wl[141] vdd gnd cell_6t
Xbit_r142_c96 bl[96] br[96] wl[142] vdd gnd cell_6t
Xbit_r143_c96 bl[96] br[96] wl[143] vdd gnd cell_6t
Xbit_r144_c96 bl[96] br[96] wl[144] vdd gnd cell_6t
Xbit_r145_c96 bl[96] br[96] wl[145] vdd gnd cell_6t
Xbit_r146_c96 bl[96] br[96] wl[146] vdd gnd cell_6t
Xbit_r147_c96 bl[96] br[96] wl[147] vdd gnd cell_6t
Xbit_r148_c96 bl[96] br[96] wl[148] vdd gnd cell_6t
Xbit_r149_c96 bl[96] br[96] wl[149] vdd gnd cell_6t
Xbit_r150_c96 bl[96] br[96] wl[150] vdd gnd cell_6t
Xbit_r151_c96 bl[96] br[96] wl[151] vdd gnd cell_6t
Xbit_r152_c96 bl[96] br[96] wl[152] vdd gnd cell_6t
Xbit_r153_c96 bl[96] br[96] wl[153] vdd gnd cell_6t
Xbit_r154_c96 bl[96] br[96] wl[154] vdd gnd cell_6t
Xbit_r155_c96 bl[96] br[96] wl[155] vdd gnd cell_6t
Xbit_r156_c96 bl[96] br[96] wl[156] vdd gnd cell_6t
Xbit_r157_c96 bl[96] br[96] wl[157] vdd gnd cell_6t
Xbit_r158_c96 bl[96] br[96] wl[158] vdd gnd cell_6t
Xbit_r159_c96 bl[96] br[96] wl[159] vdd gnd cell_6t
Xbit_r160_c96 bl[96] br[96] wl[160] vdd gnd cell_6t
Xbit_r161_c96 bl[96] br[96] wl[161] vdd gnd cell_6t
Xbit_r162_c96 bl[96] br[96] wl[162] vdd gnd cell_6t
Xbit_r163_c96 bl[96] br[96] wl[163] vdd gnd cell_6t
Xbit_r164_c96 bl[96] br[96] wl[164] vdd gnd cell_6t
Xbit_r165_c96 bl[96] br[96] wl[165] vdd gnd cell_6t
Xbit_r166_c96 bl[96] br[96] wl[166] vdd gnd cell_6t
Xbit_r167_c96 bl[96] br[96] wl[167] vdd gnd cell_6t
Xbit_r168_c96 bl[96] br[96] wl[168] vdd gnd cell_6t
Xbit_r169_c96 bl[96] br[96] wl[169] vdd gnd cell_6t
Xbit_r170_c96 bl[96] br[96] wl[170] vdd gnd cell_6t
Xbit_r171_c96 bl[96] br[96] wl[171] vdd gnd cell_6t
Xbit_r172_c96 bl[96] br[96] wl[172] vdd gnd cell_6t
Xbit_r173_c96 bl[96] br[96] wl[173] vdd gnd cell_6t
Xbit_r174_c96 bl[96] br[96] wl[174] vdd gnd cell_6t
Xbit_r175_c96 bl[96] br[96] wl[175] vdd gnd cell_6t
Xbit_r176_c96 bl[96] br[96] wl[176] vdd gnd cell_6t
Xbit_r177_c96 bl[96] br[96] wl[177] vdd gnd cell_6t
Xbit_r178_c96 bl[96] br[96] wl[178] vdd gnd cell_6t
Xbit_r179_c96 bl[96] br[96] wl[179] vdd gnd cell_6t
Xbit_r180_c96 bl[96] br[96] wl[180] vdd gnd cell_6t
Xbit_r181_c96 bl[96] br[96] wl[181] vdd gnd cell_6t
Xbit_r182_c96 bl[96] br[96] wl[182] vdd gnd cell_6t
Xbit_r183_c96 bl[96] br[96] wl[183] vdd gnd cell_6t
Xbit_r184_c96 bl[96] br[96] wl[184] vdd gnd cell_6t
Xbit_r185_c96 bl[96] br[96] wl[185] vdd gnd cell_6t
Xbit_r186_c96 bl[96] br[96] wl[186] vdd gnd cell_6t
Xbit_r187_c96 bl[96] br[96] wl[187] vdd gnd cell_6t
Xbit_r188_c96 bl[96] br[96] wl[188] vdd gnd cell_6t
Xbit_r189_c96 bl[96] br[96] wl[189] vdd gnd cell_6t
Xbit_r190_c96 bl[96] br[96] wl[190] vdd gnd cell_6t
Xbit_r191_c96 bl[96] br[96] wl[191] vdd gnd cell_6t
Xbit_r192_c96 bl[96] br[96] wl[192] vdd gnd cell_6t
Xbit_r193_c96 bl[96] br[96] wl[193] vdd gnd cell_6t
Xbit_r194_c96 bl[96] br[96] wl[194] vdd gnd cell_6t
Xbit_r195_c96 bl[96] br[96] wl[195] vdd gnd cell_6t
Xbit_r196_c96 bl[96] br[96] wl[196] vdd gnd cell_6t
Xbit_r197_c96 bl[96] br[96] wl[197] vdd gnd cell_6t
Xbit_r198_c96 bl[96] br[96] wl[198] vdd gnd cell_6t
Xbit_r199_c96 bl[96] br[96] wl[199] vdd gnd cell_6t
Xbit_r200_c96 bl[96] br[96] wl[200] vdd gnd cell_6t
Xbit_r201_c96 bl[96] br[96] wl[201] vdd gnd cell_6t
Xbit_r202_c96 bl[96] br[96] wl[202] vdd gnd cell_6t
Xbit_r203_c96 bl[96] br[96] wl[203] vdd gnd cell_6t
Xbit_r204_c96 bl[96] br[96] wl[204] vdd gnd cell_6t
Xbit_r205_c96 bl[96] br[96] wl[205] vdd gnd cell_6t
Xbit_r206_c96 bl[96] br[96] wl[206] vdd gnd cell_6t
Xbit_r207_c96 bl[96] br[96] wl[207] vdd gnd cell_6t
Xbit_r208_c96 bl[96] br[96] wl[208] vdd gnd cell_6t
Xbit_r209_c96 bl[96] br[96] wl[209] vdd gnd cell_6t
Xbit_r210_c96 bl[96] br[96] wl[210] vdd gnd cell_6t
Xbit_r211_c96 bl[96] br[96] wl[211] vdd gnd cell_6t
Xbit_r212_c96 bl[96] br[96] wl[212] vdd gnd cell_6t
Xbit_r213_c96 bl[96] br[96] wl[213] vdd gnd cell_6t
Xbit_r214_c96 bl[96] br[96] wl[214] vdd gnd cell_6t
Xbit_r215_c96 bl[96] br[96] wl[215] vdd gnd cell_6t
Xbit_r216_c96 bl[96] br[96] wl[216] vdd gnd cell_6t
Xbit_r217_c96 bl[96] br[96] wl[217] vdd gnd cell_6t
Xbit_r218_c96 bl[96] br[96] wl[218] vdd gnd cell_6t
Xbit_r219_c96 bl[96] br[96] wl[219] vdd gnd cell_6t
Xbit_r220_c96 bl[96] br[96] wl[220] vdd gnd cell_6t
Xbit_r221_c96 bl[96] br[96] wl[221] vdd gnd cell_6t
Xbit_r222_c96 bl[96] br[96] wl[222] vdd gnd cell_6t
Xbit_r223_c96 bl[96] br[96] wl[223] vdd gnd cell_6t
Xbit_r224_c96 bl[96] br[96] wl[224] vdd gnd cell_6t
Xbit_r225_c96 bl[96] br[96] wl[225] vdd gnd cell_6t
Xbit_r226_c96 bl[96] br[96] wl[226] vdd gnd cell_6t
Xbit_r227_c96 bl[96] br[96] wl[227] vdd gnd cell_6t
Xbit_r228_c96 bl[96] br[96] wl[228] vdd gnd cell_6t
Xbit_r229_c96 bl[96] br[96] wl[229] vdd gnd cell_6t
Xbit_r230_c96 bl[96] br[96] wl[230] vdd gnd cell_6t
Xbit_r231_c96 bl[96] br[96] wl[231] vdd gnd cell_6t
Xbit_r232_c96 bl[96] br[96] wl[232] vdd gnd cell_6t
Xbit_r233_c96 bl[96] br[96] wl[233] vdd gnd cell_6t
Xbit_r234_c96 bl[96] br[96] wl[234] vdd gnd cell_6t
Xbit_r235_c96 bl[96] br[96] wl[235] vdd gnd cell_6t
Xbit_r236_c96 bl[96] br[96] wl[236] vdd gnd cell_6t
Xbit_r237_c96 bl[96] br[96] wl[237] vdd gnd cell_6t
Xbit_r238_c96 bl[96] br[96] wl[238] vdd gnd cell_6t
Xbit_r239_c96 bl[96] br[96] wl[239] vdd gnd cell_6t
Xbit_r240_c96 bl[96] br[96] wl[240] vdd gnd cell_6t
Xbit_r241_c96 bl[96] br[96] wl[241] vdd gnd cell_6t
Xbit_r242_c96 bl[96] br[96] wl[242] vdd gnd cell_6t
Xbit_r243_c96 bl[96] br[96] wl[243] vdd gnd cell_6t
Xbit_r244_c96 bl[96] br[96] wl[244] vdd gnd cell_6t
Xbit_r245_c96 bl[96] br[96] wl[245] vdd gnd cell_6t
Xbit_r246_c96 bl[96] br[96] wl[246] vdd gnd cell_6t
Xbit_r247_c96 bl[96] br[96] wl[247] vdd gnd cell_6t
Xbit_r248_c96 bl[96] br[96] wl[248] vdd gnd cell_6t
Xbit_r249_c96 bl[96] br[96] wl[249] vdd gnd cell_6t
Xbit_r250_c96 bl[96] br[96] wl[250] vdd gnd cell_6t
Xbit_r251_c96 bl[96] br[96] wl[251] vdd gnd cell_6t
Xbit_r252_c96 bl[96] br[96] wl[252] vdd gnd cell_6t
Xbit_r253_c96 bl[96] br[96] wl[253] vdd gnd cell_6t
Xbit_r254_c96 bl[96] br[96] wl[254] vdd gnd cell_6t
Xbit_r255_c96 bl[96] br[96] wl[255] vdd gnd cell_6t
Xbit_r0_c97 bl[97] br[97] wl[0] vdd gnd cell_6t
Xbit_r1_c97 bl[97] br[97] wl[1] vdd gnd cell_6t
Xbit_r2_c97 bl[97] br[97] wl[2] vdd gnd cell_6t
Xbit_r3_c97 bl[97] br[97] wl[3] vdd gnd cell_6t
Xbit_r4_c97 bl[97] br[97] wl[4] vdd gnd cell_6t
Xbit_r5_c97 bl[97] br[97] wl[5] vdd gnd cell_6t
Xbit_r6_c97 bl[97] br[97] wl[6] vdd gnd cell_6t
Xbit_r7_c97 bl[97] br[97] wl[7] vdd gnd cell_6t
Xbit_r8_c97 bl[97] br[97] wl[8] vdd gnd cell_6t
Xbit_r9_c97 bl[97] br[97] wl[9] vdd gnd cell_6t
Xbit_r10_c97 bl[97] br[97] wl[10] vdd gnd cell_6t
Xbit_r11_c97 bl[97] br[97] wl[11] vdd gnd cell_6t
Xbit_r12_c97 bl[97] br[97] wl[12] vdd gnd cell_6t
Xbit_r13_c97 bl[97] br[97] wl[13] vdd gnd cell_6t
Xbit_r14_c97 bl[97] br[97] wl[14] vdd gnd cell_6t
Xbit_r15_c97 bl[97] br[97] wl[15] vdd gnd cell_6t
Xbit_r16_c97 bl[97] br[97] wl[16] vdd gnd cell_6t
Xbit_r17_c97 bl[97] br[97] wl[17] vdd gnd cell_6t
Xbit_r18_c97 bl[97] br[97] wl[18] vdd gnd cell_6t
Xbit_r19_c97 bl[97] br[97] wl[19] vdd gnd cell_6t
Xbit_r20_c97 bl[97] br[97] wl[20] vdd gnd cell_6t
Xbit_r21_c97 bl[97] br[97] wl[21] vdd gnd cell_6t
Xbit_r22_c97 bl[97] br[97] wl[22] vdd gnd cell_6t
Xbit_r23_c97 bl[97] br[97] wl[23] vdd gnd cell_6t
Xbit_r24_c97 bl[97] br[97] wl[24] vdd gnd cell_6t
Xbit_r25_c97 bl[97] br[97] wl[25] vdd gnd cell_6t
Xbit_r26_c97 bl[97] br[97] wl[26] vdd gnd cell_6t
Xbit_r27_c97 bl[97] br[97] wl[27] vdd gnd cell_6t
Xbit_r28_c97 bl[97] br[97] wl[28] vdd gnd cell_6t
Xbit_r29_c97 bl[97] br[97] wl[29] vdd gnd cell_6t
Xbit_r30_c97 bl[97] br[97] wl[30] vdd gnd cell_6t
Xbit_r31_c97 bl[97] br[97] wl[31] vdd gnd cell_6t
Xbit_r32_c97 bl[97] br[97] wl[32] vdd gnd cell_6t
Xbit_r33_c97 bl[97] br[97] wl[33] vdd gnd cell_6t
Xbit_r34_c97 bl[97] br[97] wl[34] vdd gnd cell_6t
Xbit_r35_c97 bl[97] br[97] wl[35] vdd gnd cell_6t
Xbit_r36_c97 bl[97] br[97] wl[36] vdd gnd cell_6t
Xbit_r37_c97 bl[97] br[97] wl[37] vdd gnd cell_6t
Xbit_r38_c97 bl[97] br[97] wl[38] vdd gnd cell_6t
Xbit_r39_c97 bl[97] br[97] wl[39] vdd gnd cell_6t
Xbit_r40_c97 bl[97] br[97] wl[40] vdd gnd cell_6t
Xbit_r41_c97 bl[97] br[97] wl[41] vdd gnd cell_6t
Xbit_r42_c97 bl[97] br[97] wl[42] vdd gnd cell_6t
Xbit_r43_c97 bl[97] br[97] wl[43] vdd gnd cell_6t
Xbit_r44_c97 bl[97] br[97] wl[44] vdd gnd cell_6t
Xbit_r45_c97 bl[97] br[97] wl[45] vdd gnd cell_6t
Xbit_r46_c97 bl[97] br[97] wl[46] vdd gnd cell_6t
Xbit_r47_c97 bl[97] br[97] wl[47] vdd gnd cell_6t
Xbit_r48_c97 bl[97] br[97] wl[48] vdd gnd cell_6t
Xbit_r49_c97 bl[97] br[97] wl[49] vdd gnd cell_6t
Xbit_r50_c97 bl[97] br[97] wl[50] vdd gnd cell_6t
Xbit_r51_c97 bl[97] br[97] wl[51] vdd gnd cell_6t
Xbit_r52_c97 bl[97] br[97] wl[52] vdd gnd cell_6t
Xbit_r53_c97 bl[97] br[97] wl[53] vdd gnd cell_6t
Xbit_r54_c97 bl[97] br[97] wl[54] vdd gnd cell_6t
Xbit_r55_c97 bl[97] br[97] wl[55] vdd gnd cell_6t
Xbit_r56_c97 bl[97] br[97] wl[56] vdd gnd cell_6t
Xbit_r57_c97 bl[97] br[97] wl[57] vdd gnd cell_6t
Xbit_r58_c97 bl[97] br[97] wl[58] vdd gnd cell_6t
Xbit_r59_c97 bl[97] br[97] wl[59] vdd gnd cell_6t
Xbit_r60_c97 bl[97] br[97] wl[60] vdd gnd cell_6t
Xbit_r61_c97 bl[97] br[97] wl[61] vdd gnd cell_6t
Xbit_r62_c97 bl[97] br[97] wl[62] vdd gnd cell_6t
Xbit_r63_c97 bl[97] br[97] wl[63] vdd gnd cell_6t
Xbit_r64_c97 bl[97] br[97] wl[64] vdd gnd cell_6t
Xbit_r65_c97 bl[97] br[97] wl[65] vdd gnd cell_6t
Xbit_r66_c97 bl[97] br[97] wl[66] vdd gnd cell_6t
Xbit_r67_c97 bl[97] br[97] wl[67] vdd gnd cell_6t
Xbit_r68_c97 bl[97] br[97] wl[68] vdd gnd cell_6t
Xbit_r69_c97 bl[97] br[97] wl[69] vdd gnd cell_6t
Xbit_r70_c97 bl[97] br[97] wl[70] vdd gnd cell_6t
Xbit_r71_c97 bl[97] br[97] wl[71] vdd gnd cell_6t
Xbit_r72_c97 bl[97] br[97] wl[72] vdd gnd cell_6t
Xbit_r73_c97 bl[97] br[97] wl[73] vdd gnd cell_6t
Xbit_r74_c97 bl[97] br[97] wl[74] vdd gnd cell_6t
Xbit_r75_c97 bl[97] br[97] wl[75] vdd gnd cell_6t
Xbit_r76_c97 bl[97] br[97] wl[76] vdd gnd cell_6t
Xbit_r77_c97 bl[97] br[97] wl[77] vdd gnd cell_6t
Xbit_r78_c97 bl[97] br[97] wl[78] vdd gnd cell_6t
Xbit_r79_c97 bl[97] br[97] wl[79] vdd gnd cell_6t
Xbit_r80_c97 bl[97] br[97] wl[80] vdd gnd cell_6t
Xbit_r81_c97 bl[97] br[97] wl[81] vdd gnd cell_6t
Xbit_r82_c97 bl[97] br[97] wl[82] vdd gnd cell_6t
Xbit_r83_c97 bl[97] br[97] wl[83] vdd gnd cell_6t
Xbit_r84_c97 bl[97] br[97] wl[84] vdd gnd cell_6t
Xbit_r85_c97 bl[97] br[97] wl[85] vdd gnd cell_6t
Xbit_r86_c97 bl[97] br[97] wl[86] vdd gnd cell_6t
Xbit_r87_c97 bl[97] br[97] wl[87] vdd gnd cell_6t
Xbit_r88_c97 bl[97] br[97] wl[88] vdd gnd cell_6t
Xbit_r89_c97 bl[97] br[97] wl[89] vdd gnd cell_6t
Xbit_r90_c97 bl[97] br[97] wl[90] vdd gnd cell_6t
Xbit_r91_c97 bl[97] br[97] wl[91] vdd gnd cell_6t
Xbit_r92_c97 bl[97] br[97] wl[92] vdd gnd cell_6t
Xbit_r93_c97 bl[97] br[97] wl[93] vdd gnd cell_6t
Xbit_r94_c97 bl[97] br[97] wl[94] vdd gnd cell_6t
Xbit_r95_c97 bl[97] br[97] wl[95] vdd gnd cell_6t
Xbit_r96_c97 bl[97] br[97] wl[96] vdd gnd cell_6t
Xbit_r97_c97 bl[97] br[97] wl[97] vdd gnd cell_6t
Xbit_r98_c97 bl[97] br[97] wl[98] vdd gnd cell_6t
Xbit_r99_c97 bl[97] br[97] wl[99] vdd gnd cell_6t
Xbit_r100_c97 bl[97] br[97] wl[100] vdd gnd cell_6t
Xbit_r101_c97 bl[97] br[97] wl[101] vdd gnd cell_6t
Xbit_r102_c97 bl[97] br[97] wl[102] vdd gnd cell_6t
Xbit_r103_c97 bl[97] br[97] wl[103] vdd gnd cell_6t
Xbit_r104_c97 bl[97] br[97] wl[104] vdd gnd cell_6t
Xbit_r105_c97 bl[97] br[97] wl[105] vdd gnd cell_6t
Xbit_r106_c97 bl[97] br[97] wl[106] vdd gnd cell_6t
Xbit_r107_c97 bl[97] br[97] wl[107] vdd gnd cell_6t
Xbit_r108_c97 bl[97] br[97] wl[108] vdd gnd cell_6t
Xbit_r109_c97 bl[97] br[97] wl[109] vdd gnd cell_6t
Xbit_r110_c97 bl[97] br[97] wl[110] vdd gnd cell_6t
Xbit_r111_c97 bl[97] br[97] wl[111] vdd gnd cell_6t
Xbit_r112_c97 bl[97] br[97] wl[112] vdd gnd cell_6t
Xbit_r113_c97 bl[97] br[97] wl[113] vdd gnd cell_6t
Xbit_r114_c97 bl[97] br[97] wl[114] vdd gnd cell_6t
Xbit_r115_c97 bl[97] br[97] wl[115] vdd gnd cell_6t
Xbit_r116_c97 bl[97] br[97] wl[116] vdd gnd cell_6t
Xbit_r117_c97 bl[97] br[97] wl[117] vdd gnd cell_6t
Xbit_r118_c97 bl[97] br[97] wl[118] vdd gnd cell_6t
Xbit_r119_c97 bl[97] br[97] wl[119] vdd gnd cell_6t
Xbit_r120_c97 bl[97] br[97] wl[120] vdd gnd cell_6t
Xbit_r121_c97 bl[97] br[97] wl[121] vdd gnd cell_6t
Xbit_r122_c97 bl[97] br[97] wl[122] vdd gnd cell_6t
Xbit_r123_c97 bl[97] br[97] wl[123] vdd gnd cell_6t
Xbit_r124_c97 bl[97] br[97] wl[124] vdd gnd cell_6t
Xbit_r125_c97 bl[97] br[97] wl[125] vdd gnd cell_6t
Xbit_r126_c97 bl[97] br[97] wl[126] vdd gnd cell_6t
Xbit_r127_c97 bl[97] br[97] wl[127] vdd gnd cell_6t
Xbit_r128_c97 bl[97] br[97] wl[128] vdd gnd cell_6t
Xbit_r129_c97 bl[97] br[97] wl[129] vdd gnd cell_6t
Xbit_r130_c97 bl[97] br[97] wl[130] vdd gnd cell_6t
Xbit_r131_c97 bl[97] br[97] wl[131] vdd gnd cell_6t
Xbit_r132_c97 bl[97] br[97] wl[132] vdd gnd cell_6t
Xbit_r133_c97 bl[97] br[97] wl[133] vdd gnd cell_6t
Xbit_r134_c97 bl[97] br[97] wl[134] vdd gnd cell_6t
Xbit_r135_c97 bl[97] br[97] wl[135] vdd gnd cell_6t
Xbit_r136_c97 bl[97] br[97] wl[136] vdd gnd cell_6t
Xbit_r137_c97 bl[97] br[97] wl[137] vdd gnd cell_6t
Xbit_r138_c97 bl[97] br[97] wl[138] vdd gnd cell_6t
Xbit_r139_c97 bl[97] br[97] wl[139] vdd gnd cell_6t
Xbit_r140_c97 bl[97] br[97] wl[140] vdd gnd cell_6t
Xbit_r141_c97 bl[97] br[97] wl[141] vdd gnd cell_6t
Xbit_r142_c97 bl[97] br[97] wl[142] vdd gnd cell_6t
Xbit_r143_c97 bl[97] br[97] wl[143] vdd gnd cell_6t
Xbit_r144_c97 bl[97] br[97] wl[144] vdd gnd cell_6t
Xbit_r145_c97 bl[97] br[97] wl[145] vdd gnd cell_6t
Xbit_r146_c97 bl[97] br[97] wl[146] vdd gnd cell_6t
Xbit_r147_c97 bl[97] br[97] wl[147] vdd gnd cell_6t
Xbit_r148_c97 bl[97] br[97] wl[148] vdd gnd cell_6t
Xbit_r149_c97 bl[97] br[97] wl[149] vdd gnd cell_6t
Xbit_r150_c97 bl[97] br[97] wl[150] vdd gnd cell_6t
Xbit_r151_c97 bl[97] br[97] wl[151] vdd gnd cell_6t
Xbit_r152_c97 bl[97] br[97] wl[152] vdd gnd cell_6t
Xbit_r153_c97 bl[97] br[97] wl[153] vdd gnd cell_6t
Xbit_r154_c97 bl[97] br[97] wl[154] vdd gnd cell_6t
Xbit_r155_c97 bl[97] br[97] wl[155] vdd gnd cell_6t
Xbit_r156_c97 bl[97] br[97] wl[156] vdd gnd cell_6t
Xbit_r157_c97 bl[97] br[97] wl[157] vdd gnd cell_6t
Xbit_r158_c97 bl[97] br[97] wl[158] vdd gnd cell_6t
Xbit_r159_c97 bl[97] br[97] wl[159] vdd gnd cell_6t
Xbit_r160_c97 bl[97] br[97] wl[160] vdd gnd cell_6t
Xbit_r161_c97 bl[97] br[97] wl[161] vdd gnd cell_6t
Xbit_r162_c97 bl[97] br[97] wl[162] vdd gnd cell_6t
Xbit_r163_c97 bl[97] br[97] wl[163] vdd gnd cell_6t
Xbit_r164_c97 bl[97] br[97] wl[164] vdd gnd cell_6t
Xbit_r165_c97 bl[97] br[97] wl[165] vdd gnd cell_6t
Xbit_r166_c97 bl[97] br[97] wl[166] vdd gnd cell_6t
Xbit_r167_c97 bl[97] br[97] wl[167] vdd gnd cell_6t
Xbit_r168_c97 bl[97] br[97] wl[168] vdd gnd cell_6t
Xbit_r169_c97 bl[97] br[97] wl[169] vdd gnd cell_6t
Xbit_r170_c97 bl[97] br[97] wl[170] vdd gnd cell_6t
Xbit_r171_c97 bl[97] br[97] wl[171] vdd gnd cell_6t
Xbit_r172_c97 bl[97] br[97] wl[172] vdd gnd cell_6t
Xbit_r173_c97 bl[97] br[97] wl[173] vdd gnd cell_6t
Xbit_r174_c97 bl[97] br[97] wl[174] vdd gnd cell_6t
Xbit_r175_c97 bl[97] br[97] wl[175] vdd gnd cell_6t
Xbit_r176_c97 bl[97] br[97] wl[176] vdd gnd cell_6t
Xbit_r177_c97 bl[97] br[97] wl[177] vdd gnd cell_6t
Xbit_r178_c97 bl[97] br[97] wl[178] vdd gnd cell_6t
Xbit_r179_c97 bl[97] br[97] wl[179] vdd gnd cell_6t
Xbit_r180_c97 bl[97] br[97] wl[180] vdd gnd cell_6t
Xbit_r181_c97 bl[97] br[97] wl[181] vdd gnd cell_6t
Xbit_r182_c97 bl[97] br[97] wl[182] vdd gnd cell_6t
Xbit_r183_c97 bl[97] br[97] wl[183] vdd gnd cell_6t
Xbit_r184_c97 bl[97] br[97] wl[184] vdd gnd cell_6t
Xbit_r185_c97 bl[97] br[97] wl[185] vdd gnd cell_6t
Xbit_r186_c97 bl[97] br[97] wl[186] vdd gnd cell_6t
Xbit_r187_c97 bl[97] br[97] wl[187] vdd gnd cell_6t
Xbit_r188_c97 bl[97] br[97] wl[188] vdd gnd cell_6t
Xbit_r189_c97 bl[97] br[97] wl[189] vdd gnd cell_6t
Xbit_r190_c97 bl[97] br[97] wl[190] vdd gnd cell_6t
Xbit_r191_c97 bl[97] br[97] wl[191] vdd gnd cell_6t
Xbit_r192_c97 bl[97] br[97] wl[192] vdd gnd cell_6t
Xbit_r193_c97 bl[97] br[97] wl[193] vdd gnd cell_6t
Xbit_r194_c97 bl[97] br[97] wl[194] vdd gnd cell_6t
Xbit_r195_c97 bl[97] br[97] wl[195] vdd gnd cell_6t
Xbit_r196_c97 bl[97] br[97] wl[196] vdd gnd cell_6t
Xbit_r197_c97 bl[97] br[97] wl[197] vdd gnd cell_6t
Xbit_r198_c97 bl[97] br[97] wl[198] vdd gnd cell_6t
Xbit_r199_c97 bl[97] br[97] wl[199] vdd gnd cell_6t
Xbit_r200_c97 bl[97] br[97] wl[200] vdd gnd cell_6t
Xbit_r201_c97 bl[97] br[97] wl[201] vdd gnd cell_6t
Xbit_r202_c97 bl[97] br[97] wl[202] vdd gnd cell_6t
Xbit_r203_c97 bl[97] br[97] wl[203] vdd gnd cell_6t
Xbit_r204_c97 bl[97] br[97] wl[204] vdd gnd cell_6t
Xbit_r205_c97 bl[97] br[97] wl[205] vdd gnd cell_6t
Xbit_r206_c97 bl[97] br[97] wl[206] vdd gnd cell_6t
Xbit_r207_c97 bl[97] br[97] wl[207] vdd gnd cell_6t
Xbit_r208_c97 bl[97] br[97] wl[208] vdd gnd cell_6t
Xbit_r209_c97 bl[97] br[97] wl[209] vdd gnd cell_6t
Xbit_r210_c97 bl[97] br[97] wl[210] vdd gnd cell_6t
Xbit_r211_c97 bl[97] br[97] wl[211] vdd gnd cell_6t
Xbit_r212_c97 bl[97] br[97] wl[212] vdd gnd cell_6t
Xbit_r213_c97 bl[97] br[97] wl[213] vdd gnd cell_6t
Xbit_r214_c97 bl[97] br[97] wl[214] vdd gnd cell_6t
Xbit_r215_c97 bl[97] br[97] wl[215] vdd gnd cell_6t
Xbit_r216_c97 bl[97] br[97] wl[216] vdd gnd cell_6t
Xbit_r217_c97 bl[97] br[97] wl[217] vdd gnd cell_6t
Xbit_r218_c97 bl[97] br[97] wl[218] vdd gnd cell_6t
Xbit_r219_c97 bl[97] br[97] wl[219] vdd gnd cell_6t
Xbit_r220_c97 bl[97] br[97] wl[220] vdd gnd cell_6t
Xbit_r221_c97 bl[97] br[97] wl[221] vdd gnd cell_6t
Xbit_r222_c97 bl[97] br[97] wl[222] vdd gnd cell_6t
Xbit_r223_c97 bl[97] br[97] wl[223] vdd gnd cell_6t
Xbit_r224_c97 bl[97] br[97] wl[224] vdd gnd cell_6t
Xbit_r225_c97 bl[97] br[97] wl[225] vdd gnd cell_6t
Xbit_r226_c97 bl[97] br[97] wl[226] vdd gnd cell_6t
Xbit_r227_c97 bl[97] br[97] wl[227] vdd gnd cell_6t
Xbit_r228_c97 bl[97] br[97] wl[228] vdd gnd cell_6t
Xbit_r229_c97 bl[97] br[97] wl[229] vdd gnd cell_6t
Xbit_r230_c97 bl[97] br[97] wl[230] vdd gnd cell_6t
Xbit_r231_c97 bl[97] br[97] wl[231] vdd gnd cell_6t
Xbit_r232_c97 bl[97] br[97] wl[232] vdd gnd cell_6t
Xbit_r233_c97 bl[97] br[97] wl[233] vdd gnd cell_6t
Xbit_r234_c97 bl[97] br[97] wl[234] vdd gnd cell_6t
Xbit_r235_c97 bl[97] br[97] wl[235] vdd gnd cell_6t
Xbit_r236_c97 bl[97] br[97] wl[236] vdd gnd cell_6t
Xbit_r237_c97 bl[97] br[97] wl[237] vdd gnd cell_6t
Xbit_r238_c97 bl[97] br[97] wl[238] vdd gnd cell_6t
Xbit_r239_c97 bl[97] br[97] wl[239] vdd gnd cell_6t
Xbit_r240_c97 bl[97] br[97] wl[240] vdd gnd cell_6t
Xbit_r241_c97 bl[97] br[97] wl[241] vdd gnd cell_6t
Xbit_r242_c97 bl[97] br[97] wl[242] vdd gnd cell_6t
Xbit_r243_c97 bl[97] br[97] wl[243] vdd gnd cell_6t
Xbit_r244_c97 bl[97] br[97] wl[244] vdd gnd cell_6t
Xbit_r245_c97 bl[97] br[97] wl[245] vdd gnd cell_6t
Xbit_r246_c97 bl[97] br[97] wl[246] vdd gnd cell_6t
Xbit_r247_c97 bl[97] br[97] wl[247] vdd gnd cell_6t
Xbit_r248_c97 bl[97] br[97] wl[248] vdd gnd cell_6t
Xbit_r249_c97 bl[97] br[97] wl[249] vdd gnd cell_6t
Xbit_r250_c97 bl[97] br[97] wl[250] vdd gnd cell_6t
Xbit_r251_c97 bl[97] br[97] wl[251] vdd gnd cell_6t
Xbit_r252_c97 bl[97] br[97] wl[252] vdd gnd cell_6t
Xbit_r253_c97 bl[97] br[97] wl[253] vdd gnd cell_6t
Xbit_r254_c97 bl[97] br[97] wl[254] vdd gnd cell_6t
Xbit_r255_c97 bl[97] br[97] wl[255] vdd gnd cell_6t
Xbit_r0_c98 bl[98] br[98] wl[0] vdd gnd cell_6t
Xbit_r1_c98 bl[98] br[98] wl[1] vdd gnd cell_6t
Xbit_r2_c98 bl[98] br[98] wl[2] vdd gnd cell_6t
Xbit_r3_c98 bl[98] br[98] wl[3] vdd gnd cell_6t
Xbit_r4_c98 bl[98] br[98] wl[4] vdd gnd cell_6t
Xbit_r5_c98 bl[98] br[98] wl[5] vdd gnd cell_6t
Xbit_r6_c98 bl[98] br[98] wl[6] vdd gnd cell_6t
Xbit_r7_c98 bl[98] br[98] wl[7] vdd gnd cell_6t
Xbit_r8_c98 bl[98] br[98] wl[8] vdd gnd cell_6t
Xbit_r9_c98 bl[98] br[98] wl[9] vdd gnd cell_6t
Xbit_r10_c98 bl[98] br[98] wl[10] vdd gnd cell_6t
Xbit_r11_c98 bl[98] br[98] wl[11] vdd gnd cell_6t
Xbit_r12_c98 bl[98] br[98] wl[12] vdd gnd cell_6t
Xbit_r13_c98 bl[98] br[98] wl[13] vdd gnd cell_6t
Xbit_r14_c98 bl[98] br[98] wl[14] vdd gnd cell_6t
Xbit_r15_c98 bl[98] br[98] wl[15] vdd gnd cell_6t
Xbit_r16_c98 bl[98] br[98] wl[16] vdd gnd cell_6t
Xbit_r17_c98 bl[98] br[98] wl[17] vdd gnd cell_6t
Xbit_r18_c98 bl[98] br[98] wl[18] vdd gnd cell_6t
Xbit_r19_c98 bl[98] br[98] wl[19] vdd gnd cell_6t
Xbit_r20_c98 bl[98] br[98] wl[20] vdd gnd cell_6t
Xbit_r21_c98 bl[98] br[98] wl[21] vdd gnd cell_6t
Xbit_r22_c98 bl[98] br[98] wl[22] vdd gnd cell_6t
Xbit_r23_c98 bl[98] br[98] wl[23] vdd gnd cell_6t
Xbit_r24_c98 bl[98] br[98] wl[24] vdd gnd cell_6t
Xbit_r25_c98 bl[98] br[98] wl[25] vdd gnd cell_6t
Xbit_r26_c98 bl[98] br[98] wl[26] vdd gnd cell_6t
Xbit_r27_c98 bl[98] br[98] wl[27] vdd gnd cell_6t
Xbit_r28_c98 bl[98] br[98] wl[28] vdd gnd cell_6t
Xbit_r29_c98 bl[98] br[98] wl[29] vdd gnd cell_6t
Xbit_r30_c98 bl[98] br[98] wl[30] vdd gnd cell_6t
Xbit_r31_c98 bl[98] br[98] wl[31] vdd gnd cell_6t
Xbit_r32_c98 bl[98] br[98] wl[32] vdd gnd cell_6t
Xbit_r33_c98 bl[98] br[98] wl[33] vdd gnd cell_6t
Xbit_r34_c98 bl[98] br[98] wl[34] vdd gnd cell_6t
Xbit_r35_c98 bl[98] br[98] wl[35] vdd gnd cell_6t
Xbit_r36_c98 bl[98] br[98] wl[36] vdd gnd cell_6t
Xbit_r37_c98 bl[98] br[98] wl[37] vdd gnd cell_6t
Xbit_r38_c98 bl[98] br[98] wl[38] vdd gnd cell_6t
Xbit_r39_c98 bl[98] br[98] wl[39] vdd gnd cell_6t
Xbit_r40_c98 bl[98] br[98] wl[40] vdd gnd cell_6t
Xbit_r41_c98 bl[98] br[98] wl[41] vdd gnd cell_6t
Xbit_r42_c98 bl[98] br[98] wl[42] vdd gnd cell_6t
Xbit_r43_c98 bl[98] br[98] wl[43] vdd gnd cell_6t
Xbit_r44_c98 bl[98] br[98] wl[44] vdd gnd cell_6t
Xbit_r45_c98 bl[98] br[98] wl[45] vdd gnd cell_6t
Xbit_r46_c98 bl[98] br[98] wl[46] vdd gnd cell_6t
Xbit_r47_c98 bl[98] br[98] wl[47] vdd gnd cell_6t
Xbit_r48_c98 bl[98] br[98] wl[48] vdd gnd cell_6t
Xbit_r49_c98 bl[98] br[98] wl[49] vdd gnd cell_6t
Xbit_r50_c98 bl[98] br[98] wl[50] vdd gnd cell_6t
Xbit_r51_c98 bl[98] br[98] wl[51] vdd gnd cell_6t
Xbit_r52_c98 bl[98] br[98] wl[52] vdd gnd cell_6t
Xbit_r53_c98 bl[98] br[98] wl[53] vdd gnd cell_6t
Xbit_r54_c98 bl[98] br[98] wl[54] vdd gnd cell_6t
Xbit_r55_c98 bl[98] br[98] wl[55] vdd gnd cell_6t
Xbit_r56_c98 bl[98] br[98] wl[56] vdd gnd cell_6t
Xbit_r57_c98 bl[98] br[98] wl[57] vdd gnd cell_6t
Xbit_r58_c98 bl[98] br[98] wl[58] vdd gnd cell_6t
Xbit_r59_c98 bl[98] br[98] wl[59] vdd gnd cell_6t
Xbit_r60_c98 bl[98] br[98] wl[60] vdd gnd cell_6t
Xbit_r61_c98 bl[98] br[98] wl[61] vdd gnd cell_6t
Xbit_r62_c98 bl[98] br[98] wl[62] vdd gnd cell_6t
Xbit_r63_c98 bl[98] br[98] wl[63] vdd gnd cell_6t
Xbit_r64_c98 bl[98] br[98] wl[64] vdd gnd cell_6t
Xbit_r65_c98 bl[98] br[98] wl[65] vdd gnd cell_6t
Xbit_r66_c98 bl[98] br[98] wl[66] vdd gnd cell_6t
Xbit_r67_c98 bl[98] br[98] wl[67] vdd gnd cell_6t
Xbit_r68_c98 bl[98] br[98] wl[68] vdd gnd cell_6t
Xbit_r69_c98 bl[98] br[98] wl[69] vdd gnd cell_6t
Xbit_r70_c98 bl[98] br[98] wl[70] vdd gnd cell_6t
Xbit_r71_c98 bl[98] br[98] wl[71] vdd gnd cell_6t
Xbit_r72_c98 bl[98] br[98] wl[72] vdd gnd cell_6t
Xbit_r73_c98 bl[98] br[98] wl[73] vdd gnd cell_6t
Xbit_r74_c98 bl[98] br[98] wl[74] vdd gnd cell_6t
Xbit_r75_c98 bl[98] br[98] wl[75] vdd gnd cell_6t
Xbit_r76_c98 bl[98] br[98] wl[76] vdd gnd cell_6t
Xbit_r77_c98 bl[98] br[98] wl[77] vdd gnd cell_6t
Xbit_r78_c98 bl[98] br[98] wl[78] vdd gnd cell_6t
Xbit_r79_c98 bl[98] br[98] wl[79] vdd gnd cell_6t
Xbit_r80_c98 bl[98] br[98] wl[80] vdd gnd cell_6t
Xbit_r81_c98 bl[98] br[98] wl[81] vdd gnd cell_6t
Xbit_r82_c98 bl[98] br[98] wl[82] vdd gnd cell_6t
Xbit_r83_c98 bl[98] br[98] wl[83] vdd gnd cell_6t
Xbit_r84_c98 bl[98] br[98] wl[84] vdd gnd cell_6t
Xbit_r85_c98 bl[98] br[98] wl[85] vdd gnd cell_6t
Xbit_r86_c98 bl[98] br[98] wl[86] vdd gnd cell_6t
Xbit_r87_c98 bl[98] br[98] wl[87] vdd gnd cell_6t
Xbit_r88_c98 bl[98] br[98] wl[88] vdd gnd cell_6t
Xbit_r89_c98 bl[98] br[98] wl[89] vdd gnd cell_6t
Xbit_r90_c98 bl[98] br[98] wl[90] vdd gnd cell_6t
Xbit_r91_c98 bl[98] br[98] wl[91] vdd gnd cell_6t
Xbit_r92_c98 bl[98] br[98] wl[92] vdd gnd cell_6t
Xbit_r93_c98 bl[98] br[98] wl[93] vdd gnd cell_6t
Xbit_r94_c98 bl[98] br[98] wl[94] vdd gnd cell_6t
Xbit_r95_c98 bl[98] br[98] wl[95] vdd gnd cell_6t
Xbit_r96_c98 bl[98] br[98] wl[96] vdd gnd cell_6t
Xbit_r97_c98 bl[98] br[98] wl[97] vdd gnd cell_6t
Xbit_r98_c98 bl[98] br[98] wl[98] vdd gnd cell_6t
Xbit_r99_c98 bl[98] br[98] wl[99] vdd gnd cell_6t
Xbit_r100_c98 bl[98] br[98] wl[100] vdd gnd cell_6t
Xbit_r101_c98 bl[98] br[98] wl[101] vdd gnd cell_6t
Xbit_r102_c98 bl[98] br[98] wl[102] vdd gnd cell_6t
Xbit_r103_c98 bl[98] br[98] wl[103] vdd gnd cell_6t
Xbit_r104_c98 bl[98] br[98] wl[104] vdd gnd cell_6t
Xbit_r105_c98 bl[98] br[98] wl[105] vdd gnd cell_6t
Xbit_r106_c98 bl[98] br[98] wl[106] vdd gnd cell_6t
Xbit_r107_c98 bl[98] br[98] wl[107] vdd gnd cell_6t
Xbit_r108_c98 bl[98] br[98] wl[108] vdd gnd cell_6t
Xbit_r109_c98 bl[98] br[98] wl[109] vdd gnd cell_6t
Xbit_r110_c98 bl[98] br[98] wl[110] vdd gnd cell_6t
Xbit_r111_c98 bl[98] br[98] wl[111] vdd gnd cell_6t
Xbit_r112_c98 bl[98] br[98] wl[112] vdd gnd cell_6t
Xbit_r113_c98 bl[98] br[98] wl[113] vdd gnd cell_6t
Xbit_r114_c98 bl[98] br[98] wl[114] vdd gnd cell_6t
Xbit_r115_c98 bl[98] br[98] wl[115] vdd gnd cell_6t
Xbit_r116_c98 bl[98] br[98] wl[116] vdd gnd cell_6t
Xbit_r117_c98 bl[98] br[98] wl[117] vdd gnd cell_6t
Xbit_r118_c98 bl[98] br[98] wl[118] vdd gnd cell_6t
Xbit_r119_c98 bl[98] br[98] wl[119] vdd gnd cell_6t
Xbit_r120_c98 bl[98] br[98] wl[120] vdd gnd cell_6t
Xbit_r121_c98 bl[98] br[98] wl[121] vdd gnd cell_6t
Xbit_r122_c98 bl[98] br[98] wl[122] vdd gnd cell_6t
Xbit_r123_c98 bl[98] br[98] wl[123] vdd gnd cell_6t
Xbit_r124_c98 bl[98] br[98] wl[124] vdd gnd cell_6t
Xbit_r125_c98 bl[98] br[98] wl[125] vdd gnd cell_6t
Xbit_r126_c98 bl[98] br[98] wl[126] vdd gnd cell_6t
Xbit_r127_c98 bl[98] br[98] wl[127] vdd gnd cell_6t
Xbit_r128_c98 bl[98] br[98] wl[128] vdd gnd cell_6t
Xbit_r129_c98 bl[98] br[98] wl[129] vdd gnd cell_6t
Xbit_r130_c98 bl[98] br[98] wl[130] vdd gnd cell_6t
Xbit_r131_c98 bl[98] br[98] wl[131] vdd gnd cell_6t
Xbit_r132_c98 bl[98] br[98] wl[132] vdd gnd cell_6t
Xbit_r133_c98 bl[98] br[98] wl[133] vdd gnd cell_6t
Xbit_r134_c98 bl[98] br[98] wl[134] vdd gnd cell_6t
Xbit_r135_c98 bl[98] br[98] wl[135] vdd gnd cell_6t
Xbit_r136_c98 bl[98] br[98] wl[136] vdd gnd cell_6t
Xbit_r137_c98 bl[98] br[98] wl[137] vdd gnd cell_6t
Xbit_r138_c98 bl[98] br[98] wl[138] vdd gnd cell_6t
Xbit_r139_c98 bl[98] br[98] wl[139] vdd gnd cell_6t
Xbit_r140_c98 bl[98] br[98] wl[140] vdd gnd cell_6t
Xbit_r141_c98 bl[98] br[98] wl[141] vdd gnd cell_6t
Xbit_r142_c98 bl[98] br[98] wl[142] vdd gnd cell_6t
Xbit_r143_c98 bl[98] br[98] wl[143] vdd gnd cell_6t
Xbit_r144_c98 bl[98] br[98] wl[144] vdd gnd cell_6t
Xbit_r145_c98 bl[98] br[98] wl[145] vdd gnd cell_6t
Xbit_r146_c98 bl[98] br[98] wl[146] vdd gnd cell_6t
Xbit_r147_c98 bl[98] br[98] wl[147] vdd gnd cell_6t
Xbit_r148_c98 bl[98] br[98] wl[148] vdd gnd cell_6t
Xbit_r149_c98 bl[98] br[98] wl[149] vdd gnd cell_6t
Xbit_r150_c98 bl[98] br[98] wl[150] vdd gnd cell_6t
Xbit_r151_c98 bl[98] br[98] wl[151] vdd gnd cell_6t
Xbit_r152_c98 bl[98] br[98] wl[152] vdd gnd cell_6t
Xbit_r153_c98 bl[98] br[98] wl[153] vdd gnd cell_6t
Xbit_r154_c98 bl[98] br[98] wl[154] vdd gnd cell_6t
Xbit_r155_c98 bl[98] br[98] wl[155] vdd gnd cell_6t
Xbit_r156_c98 bl[98] br[98] wl[156] vdd gnd cell_6t
Xbit_r157_c98 bl[98] br[98] wl[157] vdd gnd cell_6t
Xbit_r158_c98 bl[98] br[98] wl[158] vdd gnd cell_6t
Xbit_r159_c98 bl[98] br[98] wl[159] vdd gnd cell_6t
Xbit_r160_c98 bl[98] br[98] wl[160] vdd gnd cell_6t
Xbit_r161_c98 bl[98] br[98] wl[161] vdd gnd cell_6t
Xbit_r162_c98 bl[98] br[98] wl[162] vdd gnd cell_6t
Xbit_r163_c98 bl[98] br[98] wl[163] vdd gnd cell_6t
Xbit_r164_c98 bl[98] br[98] wl[164] vdd gnd cell_6t
Xbit_r165_c98 bl[98] br[98] wl[165] vdd gnd cell_6t
Xbit_r166_c98 bl[98] br[98] wl[166] vdd gnd cell_6t
Xbit_r167_c98 bl[98] br[98] wl[167] vdd gnd cell_6t
Xbit_r168_c98 bl[98] br[98] wl[168] vdd gnd cell_6t
Xbit_r169_c98 bl[98] br[98] wl[169] vdd gnd cell_6t
Xbit_r170_c98 bl[98] br[98] wl[170] vdd gnd cell_6t
Xbit_r171_c98 bl[98] br[98] wl[171] vdd gnd cell_6t
Xbit_r172_c98 bl[98] br[98] wl[172] vdd gnd cell_6t
Xbit_r173_c98 bl[98] br[98] wl[173] vdd gnd cell_6t
Xbit_r174_c98 bl[98] br[98] wl[174] vdd gnd cell_6t
Xbit_r175_c98 bl[98] br[98] wl[175] vdd gnd cell_6t
Xbit_r176_c98 bl[98] br[98] wl[176] vdd gnd cell_6t
Xbit_r177_c98 bl[98] br[98] wl[177] vdd gnd cell_6t
Xbit_r178_c98 bl[98] br[98] wl[178] vdd gnd cell_6t
Xbit_r179_c98 bl[98] br[98] wl[179] vdd gnd cell_6t
Xbit_r180_c98 bl[98] br[98] wl[180] vdd gnd cell_6t
Xbit_r181_c98 bl[98] br[98] wl[181] vdd gnd cell_6t
Xbit_r182_c98 bl[98] br[98] wl[182] vdd gnd cell_6t
Xbit_r183_c98 bl[98] br[98] wl[183] vdd gnd cell_6t
Xbit_r184_c98 bl[98] br[98] wl[184] vdd gnd cell_6t
Xbit_r185_c98 bl[98] br[98] wl[185] vdd gnd cell_6t
Xbit_r186_c98 bl[98] br[98] wl[186] vdd gnd cell_6t
Xbit_r187_c98 bl[98] br[98] wl[187] vdd gnd cell_6t
Xbit_r188_c98 bl[98] br[98] wl[188] vdd gnd cell_6t
Xbit_r189_c98 bl[98] br[98] wl[189] vdd gnd cell_6t
Xbit_r190_c98 bl[98] br[98] wl[190] vdd gnd cell_6t
Xbit_r191_c98 bl[98] br[98] wl[191] vdd gnd cell_6t
Xbit_r192_c98 bl[98] br[98] wl[192] vdd gnd cell_6t
Xbit_r193_c98 bl[98] br[98] wl[193] vdd gnd cell_6t
Xbit_r194_c98 bl[98] br[98] wl[194] vdd gnd cell_6t
Xbit_r195_c98 bl[98] br[98] wl[195] vdd gnd cell_6t
Xbit_r196_c98 bl[98] br[98] wl[196] vdd gnd cell_6t
Xbit_r197_c98 bl[98] br[98] wl[197] vdd gnd cell_6t
Xbit_r198_c98 bl[98] br[98] wl[198] vdd gnd cell_6t
Xbit_r199_c98 bl[98] br[98] wl[199] vdd gnd cell_6t
Xbit_r200_c98 bl[98] br[98] wl[200] vdd gnd cell_6t
Xbit_r201_c98 bl[98] br[98] wl[201] vdd gnd cell_6t
Xbit_r202_c98 bl[98] br[98] wl[202] vdd gnd cell_6t
Xbit_r203_c98 bl[98] br[98] wl[203] vdd gnd cell_6t
Xbit_r204_c98 bl[98] br[98] wl[204] vdd gnd cell_6t
Xbit_r205_c98 bl[98] br[98] wl[205] vdd gnd cell_6t
Xbit_r206_c98 bl[98] br[98] wl[206] vdd gnd cell_6t
Xbit_r207_c98 bl[98] br[98] wl[207] vdd gnd cell_6t
Xbit_r208_c98 bl[98] br[98] wl[208] vdd gnd cell_6t
Xbit_r209_c98 bl[98] br[98] wl[209] vdd gnd cell_6t
Xbit_r210_c98 bl[98] br[98] wl[210] vdd gnd cell_6t
Xbit_r211_c98 bl[98] br[98] wl[211] vdd gnd cell_6t
Xbit_r212_c98 bl[98] br[98] wl[212] vdd gnd cell_6t
Xbit_r213_c98 bl[98] br[98] wl[213] vdd gnd cell_6t
Xbit_r214_c98 bl[98] br[98] wl[214] vdd gnd cell_6t
Xbit_r215_c98 bl[98] br[98] wl[215] vdd gnd cell_6t
Xbit_r216_c98 bl[98] br[98] wl[216] vdd gnd cell_6t
Xbit_r217_c98 bl[98] br[98] wl[217] vdd gnd cell_6t
Xbit_r218_c98 bl[98] br[98] wl[218] vdd gnd cell_6t
Xbit_r219_c98 bl[98] br[98] wl[219] vdd gnd cell_6t
Xbit_r220_c98 bl[98] br[98] wl[220] vdd gnd cell_6t
Xbit_r221_c98 bl[98] br[98] wl[221] vdd gnd cell_6t
Xbit_r222_c98 bl[98] br[98] wl[222] vdd gnd cell_6t
Xbit_r223_c98 bl[98] br[98] wl[223] vdd gnd cell_6t
Xbit_r224_c98 bl[98] br[98] wl[224] vdd gnd cell_6t
Xbit_r225_c98 bl[98] br[98] wl[225] vdd gnd cell_6t
Xbit_r226_c98 bl[98] br[98] wl[226] vdd gnd cell_6t
Xbit_r227_c98 bl[98] br[98] wl[227] vdd gnd cell_6t
Xbit_r228_c98 bl[98] br[98] wl[228] vdd gnd cell_6t
Xbit_r229_c98 bl[98] br[98] wl[229] vdd gnd cell_6t
Xbit_r230_c98 bl[98] br[98] wl[230] vdd gnd cell_6t
Xbit_r231_c98 bl[98] br[98] wl[231] vdd gnd cell_6t
Xbit_r232_c98 bl[98] br[98] wl[232] vdd gnd cell_6t
Xbit_r233_c98 bl[98] br[98] wl[233] vdd gnd cell_6t
Xbit_r234_c98 bl[98] br[98] wl[234] vdd gnd cell_6t
Xbit_r235_c98 bl[98] br[98] wl[235] vdd gnd cell_6t
Xbit_r236_c98 bl[98] br[98] wl[236] vdd gnd cell_6t
Xbit_r237_c98 bl[98] br[98] wl[237] vdd gnd cell_6t
Xbit_r238_c98 bl[98] br[98] wl[238] vdd gnd cell_6t
Xbit_r239_c98 bl[98] br[98] wl[239] vdd gnd cell_6t
Xbit_r240_c98 bl[98] br[98] wl[240] vdd gnd cell_6t
Xbit_r241_c98 bl[98] br[98] wl[241] vdd gnd cell_6t
Xbit_r242_c98 bl[98] br[98] wl[242] vdd gnd cell_6t
Xbit_r243_c98 bl[98] br[98] wl[243] vdd gnd cell_6t
Xbit_r244_c98 bl[98] br[98] wl[244] vdd gnd cell_6t
Xbit_r245_c98 bl[98] br[98] wl[245] vdd gnd cell_6t
Xbit_r246_c98 bl[98] br[98] wl[246] vdd gnd cell_6t
Xbit_r247_c98 bl[98] br[98] wl[247] vdd gnd cell_6t
Xbit_r248_c98 bl[98] br[98] wl[248] vdd gnd cell_6t
Xbit_r249_c98 bl[98] br[98] wl[249] vdd gnd cell_6t
Xbit_r250_c98 bl[98] br[98] wl[250] vdd gnd cell_6t
Xbit_r251_c98 bl[98] br[98] wl[251] vdd gnd cell_6t
Xbit_r252_c98 bl[98] br[98] wl[252] vdd gnd cell_6t
Xbit_r253_c98 bl[98] br[98] wl[253] vdd gnd cell_6t
Xbit_r254_c98 bl[98] br[98] wl[254] vdd gnd cell_6t
Xbit_r255_c98 bl[98] br[98] wl[255] vdd gnd cell_6t
Xbit_r0_c99 bl[99] br[99] wl[0] vdd gnd cell_6t
Xbit_r1_c99 bl[99] br[99] wl[1] vdd gnd cell_6t
Xbit_r2_c99 bl[99] br[99] wl[2] vdd gnd cell_6t
Xbit_r3_c99 bl[99] br[99] wl[3] vdd gnd cell_6t
Xbit_r4_c99 bl[99] br[99] wl[4] vdd gnd cell_6t
Xbit_r5_c99 bl[99] br[99] wl[5] vdd gnd cell_6t
Xbit_r6_c99 bl[99] br[99] wl[6] vdd gnd cell_6t
Xbit_r7_c99 bl[99] br[99] wl[7] vdd gnd cell_6t
Xbit_r8_c99 bl[99] br[99] wl[8] vdd gnd cell_6t
Xbit_r9_c99 bl[99] br[99] wl[9] vdd gnd cell_6t
Xbit_r10_c99 bl[99] br[99] wl[10] vdd gnd cell_6t
Xbit_r11_c99 bl[99] br[99] wl[11] vdd gnd cell_6t
Xbit_r12_c99 bl[99] br[99] wl[12] vdd gnd cell_6t
Xbit_r13_c99 bl[99] br[99] wl[13] vdd gnd cell_6t
Xbit_r14_c99 bl[99] br[99] wl[14] vdd gnd cell_6t
Xbit_r15_c99 bl[99] br[99] wl[15] vdd gnd cell_6t
Xbit_r16_c99 bl[99] br[99] wl[16] vdd gnd cell_6t
Xbit_r17_c99 bl[99] br[99] wl[17] vdd gnd cell_6t
Xbit_r18_c99 bl[99] br[99] wl[18] vdd gnd cell_6t
Xbit_r19_c99 bl[99] br[99] wl[19] vdd gnd cell_6t
Xbit_r20_c99 bl[99] br[99] wl[20] vdd gnd cell_6t
Xbit_r21_c99 bl[99] br[99] wl[21] vdd gnd cell_6t
Xbit_r22_c99 bl[99] br[99] wl[22] vdd gnd cell_6t
Xbit_r23_c99 bl[99] br[99] wl[23] vdd gnd cell_6t
Xbit_r24_c99 bl[99] br[99] wl[24] vdd gnd cell_6t
Xbit_r25_c99 bl[99] br[99] wl[25] vdd gnd cell_6t
Xbit_r26_c99 bl[99] br[99] wl[26] vdd gnd cell_6t
Xbit_r27_c99 bl[99] br[99] wl[27] vdd gnd cell_6t
Xbit_r28_c99 bl[99] br[99] wl[28] vdd gnd cell_6t
Xbit_r29_c99 bl[99] br[99] wl[29] vdd gnd cell_6t
Xbit_r30_c99 bl[99] br[99] wl[30] vdd gnd cell_6t
Xbit_r31_c99 bl[99] br[99] wl[31] vdd gnd cell_6t
Xbit_r32_c99 bl[99] br[99] wl[32] vdd gnd cell_6t
Xbit_r33_c99 bl[99] br[99] wl[33] vdd gnd cell_6t
Xbit_r34_c99 bl[99] br[99] wl[34] vdd gnd cell_6t
Xbit_r35_c99 bl[99] br[99] wl[35] vdd gnd cell_6t
Xbit_r36_c99 bl[99] br[99] wl[36] vdd gnd cell_6t
Xbit_r37_c99 bl[99] br[99] wl[37] vdd gnd cell_6t
Xbit_r38_c99 bl[99] br[99] wl[38] vdd gnd cell_6t
Xbit_r39_c99 bl[99] br[99] wl[39] vdd gnd cell_6t
Xbit_r40_c99 bl[99] br[99] wl[40] vdd gnd cell_6t
Xbit_r41_c99 bl[99] br[99] wl[41] vdd gnd cell_6t
Xbit_r42_c99 bl[99] br[99] wl[42] vdd gnd cell_6t
Xbit_r43_c99 bl[99] br[99] wl[43] vdd gnd cell_6t
Xbit_r44_c99 bl[99] br[99] wl[44] vdd gnd cell_6t
Xbit_r45_c99 bl[99] br[99] wl[45] vdd gnd cell_6t
Xbit_r46_c99 bl[99] br[99] wl[46] vdd gnd cell_6t
Xbit_r47_c99 bl[99] br[99] wl[47] vdd gnd cell_6t
Xbit_r48_c99 bl[99] br[99] wl[48] vdd gnd cell_6t
Xbit_r49_c99 bl[99] br[99] wl[49] vdd gnd cell_6t
Xbit_r50_c99 bl[99] br[99] wl[50] vdd gnd cell_6t
Xbit_r51_c99 bl[99] br[99] wl[51] vdd gnd cell_6t
Xbit_r52_c99 bl[99] br[99] wl[52] vdd gnd cell_6t
Xbit_r53_c99 bl[99] br[99] wl[53] vdd gnd cell_6t
Xbit_r54_c99 bl[99] br[99] wl[54] vdd gnd cell_6t
Xbit_r55_c99 bl[99] br[99] wl[55] vdd gnd cell_6t
Xbit_r56_c99 bl[99] br[99] wl[56] vdd gnd cell_6t
Xbit_r57_c99 bl[99] br[99] wl[57] vdd gnd cell_6t
Xbit_r58_c99 bl[99] br[99] wl[58] vdd gnd cell_6t
Xbit_r59_c99 bl[99] br[99] wl[59] vdd gnd cell_6t
Xbit_r60_c99 bl[99] br[99] wl[60] vdd gnd cell_6t
Xbit_r61_c99 bl[99] br[99] wl[61] vdd gnd cell_6t
Xbit_r62_c99 bl[99] br[99] wl[62] vdd gnd cell_6t
Xbit_r63_c99 bl[99] br[99] wl[63] vdd gnd cell_6t
Xbit_r64_c99 bl[99] br[99] wl[64] vdd gnd cell_6t
Xbit_r65_c99 bl[99] br[99] wl[65] vdd gnd cell_6t
Xbit_r66_c99 bl[99] br[99] wl[66] vdd gnd cell_6t
Xbit_r67_c99 bl[99] br[99] wl[67] vdd gnd cell_6t
Xbit_r68_c99 bl[99] br[99] wl[68] vdd gnd cell_6t
Xbit_r69_c99 bl[99] br[99] wl[69] vdd gnd cell_6t
Xbit_r70_c99 bl[99] br[99] wl[70] vdd gnd cell_6t
Xbit_r71_c99 bl[99] br[99] wl[71] vdd gnd cell_6t
Xbit_r72_c99 bl[99] br[99] wl[72] vdd gnd cell_6t
Xbit_r73_c99 bl[99] br[99] wl[73] vdd gnd cell_6t
Xbit_r74_c99 bl[99] br[99] wl[74] vdd gnd cell_6t
Xbit_r75_c99 bl[99] br[99] wl[75] vdd gnd cell_6t
Xbit_r76_c99 bl[99] br[99] wl[76] vdd gnd cell_6t
Xbit_r77_c99 bl[99] br[99] wl[77] vdd gnd cell_6t
Xbit_r78_c99 bl[99] br[99] wl[78] vdd gnd cell_6t
Xbit_r79_c99 bl[99] br[99] wl[79] vdd gnd cell_6t
Xbit_r80_c99 bl[99] br[99] wl[80] vdd gnd cell_6t
Xbit_r81_c99 bl[99] br[99] wl[81] vdd gnd cell_6t
Xbit_r82_c99 bl[99] br[99] wl[82] vdd gnd cell_6t
Xbit_r83_c99 bl[99] br[99] wl[83] vdd gnd cell_6t
Xbit_r84_c99 bl[99] br[99] wl[84] vdd gnd cell_6t
Xbit_r85_c99 bl[99] br[99] wl[85] vdd gnd cell_6t
Xbit_r86_c99 bl[99] br[99] wl[86] vdd gnd cell_6t
Xbit_r87_c99 bl[99] br[99] wl[87] vdd gnd cell_6t
Xbit_r88_c99 bl[99] br[99] wl[88] vdd gnd cell_6t
Xbit_r89_c99 bl[99] br[99] wl[89] vdd gnd cell_6t
Xbit_r90_c99 bl[99] br[99] wl[90] vdd gnd cell_6t
Xbit_r91_c99 bl[99] br[99] wl[91] vdd gnd cell_6t
Xbit_r92_c99 bl[99] br[99] wl[92] vdd gnd cell_6t
Xbit_r93_c99 bl[99] br[99] wl[93] vdd gnd cell_6t
Xbit_r94_c99 bl[99] br[99] wl[94] vdd gnd cell_6t
Xbit_r95_c99 bl[99] br[99] wl[95] vdd gnd cell_6t
Xbit_r96_c99 bl[99] br[99] wl[96] vdd gnd cell_6t
Xbit_r97_c99 bl[99] br[99] wl[97] vdd gnd cell_6t
Xbit_r98_c99 bl[99] br[99] wl[98] vdd gnd cell_6t
Xbit_r99_c99 bl[99] br[99] wl[99] vdd gnd cell_6t
Xbit_r100_c99 bl[99] br[99] wl[100] vdd gnd cell_6t
Xbit_r101_c99 bl[99] br[99] wl[101] vdd gnd cell_6t
Xbit_r102_c99 bl[99] br[99] wl[102] vdd gnd cell_6t
Xbit_r103_c99 bl[99] br[99] wl[103] vdd gnd cell_6t
Xbit_r104_c99 bl[99] br[99] wl[104] vdd gnd cell_6t
Xbit_r105_c99 bl[99] br[99] wl[105] vdd gnd cell_6t
Xbit_r106_c99 bl[99] br[99] wl[106] vdd gnd cell_6t
Xbit_r107_c99 bl[99] br[99] wl[107] vdd gnd cell_6t
Xbit_r108_c99 bl[99] br[99] wl[108] vdd gnd cell_6t
Xbit_r109_c99 bl[99] br[99] wl[109] vdd gnd cell_6t
Xbit_r110_c99 bl[99] br[99] wl[110] vdd gnd cell_6t
Xbit_r111_c99 bl[99] br[99] wl[111] vdd gnd cell_6t
Xbit_r112_c99 bl[99] br[99] wl[112] vdd gnd cell_6t
Xbit_r113_c99 bl[99] br[99] wl[113] vdd gnd cell_6t
Xbit_r114_c99 bl[99] br[99] wl[114] vdd gnd cell_6t
Xbit_r115_c99 bl[99] br[99] wl[115] vdd gnd cell_6t
Xbit_r116_c99 bl[99] br[99] wl[116] vdd gnd cell_6t
Xbit_r117_c99 bl[99] br[99] wl[117] vdd gnd cell_6t
Xbit_r118_c99 bl[99] br[99] wl[118] vdd gnd cell_6t
Xbit_r119_c99 bl[99] br[99] wl[119] vdd gnd cell_6t
Xbit_r120_c99 bl[99] br[99] wl[120] vdd gnd cell_6t
Xbit_r121_c99 bl[99] br[99] wl[121] vdd gnd cell_6t
Xbit_r122_c99 bl[99] br[99] wl[122] vdd gnd cell_6t
Xbit_r123_c99 bl[99] br[99] wl[123] vdd gnd cell_6t
Xbit_r124_c99 bl[99] br[99] wl[124] vdd gnd cell_6t
Xbit_r125_c99 bl[99] br[99] wl[125] vdd gnd cell_6t
Xbit_r126_c99 bl[99] br[99] wl[126] vdd gnd cell_6t
Xbit_r127_c99 bl[99] br[99] wl[127] vdd gnd cell_6t
Xbit_r128_c99 bl[99] br[99] wl[128] vdd gnd cell_6t
Xbit_r129_c99 bl[99] br[99] wl[129] vdd gnd cell_6t
Xbit_r130_c99 bl[99] br[99] wl[130] vdd gnd cell_6t
Xbit_r131_c99 bl[99] br[99] wl[131] vdd gnd cell_6t
Xbit_r132_c99 bl[99] br[99] wl[132] vdd gnd cell_6t
Xbit_r133_c99 bl[99] br[99] wl[133] vdd gnd cell_6t
Xbit_r134_c99 bl[99] br[99] wl[134] vdd gnd cell_6t
Xbit_r135_c99 bl[99] br[99] wl[135] vdd gnd cell_6t
Xbit_r136_c99 bl[99] br[99] wl[136] vdd gnd cell_6t
Xbit_r137_c99 bl[99] br[99] wl[137] vdd gnd cell_6t
Xbit_r138_c99 bl[99] br[99] wl[138] vdd gnd cell_6t
Xbit_r139_c99 bl[99] br[99] wl[139] vdd gnd cell_6t
Xbit_r140_c99 bl[99] br[99] wl[140] vdd gnd cell_6t
Xbit_r141_c99 bl[99] br[99] wl[141] vdd gnd cell_6t
Xbit_r142_c99 bl[99] br[99] wl[142] vdd gnd cell_6t
Xbit_r143_c99 bl[99] br[99] wl[143] vdd gnd cell_6t
Xbit_r144_c99 bl[99] br[99] wl[144] vdd gnd cell_6t
Xbit_r145_c99 bl[99] br[99] wl[145] vdd gnd cell_6t
Xbit_r146_c99 bl[99] br[99] wl[146] vdd gnd cell_6t
Xbit_r147_c99 bl[99] br[99] wl[147] vdd gnd cell_6t
Xbit_r148_c99 bl[99] br[99] wl[148] vdd gnd cell_6t
Xbit_r149_c99 bl[99] br[99] wl[149] vdd gnd cell_6t
Xbit_r150_c99 bl[99] br[99] wl[150] vdd gnd cell_6t
Xbit_r151_c99 bl[99] br[99] wl[151] vdd gnd cell_6t
Xbit_r152_c99 bl[99] br[99] wl[152] vdd gnd cell_6t
Xbit_r153_c99 bl[99] br[99] wl[153] vdd gnd cell_6t
Xbit_r154_c99 bl[99] br[99] wl[154] vdd gnd cell_6t
Xbit_r155_c99 bl[99] br[99] wl[155] vdd gnd cell_6t
Xbit_r156_c99 bl[99] br[99] wl[156] vdd gnd cell_6t
Xbit_r157_c99 bl[99] br[99] wl[157] vdd gnd cell_6t
Xbit_r158_c99 bl[99] br[99] wl[158] vdd gnd cell_6t
Xbit_r159_c99 bl[99] br[99] wl[159] vdd gnd cell_6t
Xbit_r160_c99 bl[99] br[99] wl[160] vdd gnd cell_6t
Xbit_r161_c99 bl[99] br[99] wl[161] vdd gnd cell_6t
Xbit_r162_c99 bl[99] br[99] wl[162] vdd gnd cell_6t
Xbit_r163_c99 bl[99] br[99] wl[163] vdd gnd cell_6t
Xbit_r164_c99 bl[99] br[99] wl[164] vdd gnd cell_6t
Xbit_r165_c99 bl[99] br[99] wl[165] vdd gnd cell_6t
Xbit_r166_c99 bl[99] br[99] wl[166] vdd gnd cell_6t
Xbit_r167_c99 bl[99] br[99] wl[167] vdd gnd cell_6t
Xbit_r168_c99 bl[99] br[99] wl[168] vdd gnd cell_6t
Xbit_r169_c99 bl[99] br[99] wl[169] vdd gnd cell_6t
Xbit_r170_c99 bl[99] br[99] wl[170] vdd gnd cell_6t
Xbit_r171_c99 bl[99] br[99] wl[171] vdd gnd cell_6t
Xbit_r172_c99 bl[99] br[99] wl[172] vdd gnd cell_6t
Xbit_r173_c99 bl[99] br[99] wl[173] vdd gnd cell_6t
Xbit_r174_c99 bl[99] br[99] wl[174] vdd gnd cell_6t
Xbit_r175_c99 bl[99] br[99] wl[175] vdd gnd cell_6t
Xbit_r176_c99 bl[99] br[99] wl[176] vdd gnd cell_6t
Xbit_r177_c99 bl[99] br[99] wl[177] vdd gnd cell_6t
Xbit_r178_c99 bl[99] br[99] wl[178] vdd gnd cell_6t
Xbit_r179_c99 bl[99] br[99] wl[179] vdd gnd cell_6t
Xbit_r180_c99 bl[99] br[99] wl[180] vdd gnd cell_6t
Xbit_r181_c99 bl[99] br[99] wl[181] vdd gnd cell_6t
Xbit_r182_c99 bl[99] br[99] wl[182] vdd gnd cell_6t
Xbit_r183_c99 bl[99] br[99] wl[183] vdd gnd cell_6t
Xbit_r184_c99 bl[99] br[99] wl[184] vdd gnd cell_6t
Xbit_r185_c99 bl[99] br[99] wl[185] vdd gnd cell_6t
Xbit_r186_c99 bl[99] br[99] wl[186] vdd gnd cell_6t
Xbit_r187_c99 bl[99] br[99] wl[187] vdd gnd cell_6t
Xbit_r188_c99 bl[99] br[99] wl[188] vdd gnd cell_6t
Xbit_r189_c99 bl[99] br[99] wl[189] vdd gnd cell_6t
Xbit_r190_c99 bl[99] br[99] wl[190] vdd gnd cell_6t
Xbit_r191_c99 bl[99] br[99] wl[191] vdd gnd cell_6t
Xbit_r192_c99 bl[99] br[99] wl[192] vdd gnd cell_6t
Xbit_r193_c99 bl[99] br[99] wl[193] vdd gnd cell_6t
Xbit_r194_c99 bl[99] br[99] wl[194] vdd gnd cell_6t
Xbit_r195_c99 bl[99] br[99] wl[195] vdd gnd cell_6t
Xbit_r196_c99 bl[99] br[99] wl[196] vdd gnd cell_6t
Xbit_r197_c99 bl[99] br[99] wl[197] vdd gnd cell_6t
Xbit_r198_c99 bl[99] br[99] wl[198] vdd gnd cell_6t
Xbit_r199_c99 bl[99] br[99] wl[199] vdd gnd cell_6t
Xbit_r200_c99 bl[99] br[99] wl[200] vdd gnd cell_6t
Xbit_r201_c99 bl[99] br[99] wl[201] vdd gnd cell_6t
Xbit_r202_c99 bl[99] br[99] wl[202] vdd gnd cell_6t
Xbit_r203_c99 bl[99] br[99] wl[203] vdd gnd cell_6t
Xbit_r204_c99 bl[99] br[99] wl[204] vdd gnd cell_6t
Xbit_r205_c99 bl[99] br[99] wl[205] vdd gnd cell_6t
Xbit_r206_c99 bl[99] br[99] wl[206] vdd gnd cell_6t
Xbit_r207_c99 bl[99] br[99] wl[207] vdd gnd cell_6t
Xbit_r208_c99 bl[99] br[99] wl[208] vdd gnd cell_6t
Xbit_r209_c99 bl[99] br[99] wl[209] vdd gnd cell_6t
Xbit_r210_c99 bl[99] br[99] wl[210] vdd gnd cell_6t
Xbit_r211_c99 bl[99] br[99] wl[211] vdd gnd cell_6t
Xbit_r212_c99 bl[99] br[99] wl[212] vdd gnd cell_6t
Xbit_r213_c99 bl[99] br[99] wl[213] vdd gnd cell_6t
Xbit_r214_c99 bl[99] br[99] wl[214] vdd gnd cell_6t
Xbit_r215_c99 bl[99] br[99] wl[215] vdd gnd cell_6t
Xbit_r216_c99 bl[99] br[99] wl[216] vdd gnd cell_6t
Xbit_r217_c99 bl[99] br[99] wl[217] vdd gnd cell_6t
Xbit_r218_c99 bl[99] br[99] wl[218] vdd gnd cell_6t
Xbit_r219_c99 bl[99] br[99] wl[219] vdd gnd cell_6t
Xbit_r220_c99 bl[99] br[99] wl[220] vdd gnd cell_6t
Xbit_r221_c99 bl[99] br[99] wl[221] vdd gnd cell_6t
Xbit_r222_c99 bl[99] br[99] wl[222] vdd gnd cell_6t
Xbit_r223_c99 bl[99] br[99] wl[223] vdd gnd cell_6t
Xbit_r224_c99 bl[99] br[99] wl[224] vdd gnd cell_6t
Xbit_r225_c99 bl[99] br[99] wl[225] vdd gnd cell_6t
Xbit_r226_c99 bl[99] br[99] wl[226] vdd gnd cell_6t
Xbit_r227_c99 bl[99] br[99] wl[227] vdd gnd cell_6t
Xbit_r228_c99 bl[99] br[99] wl[228] vdd gnd cell_6t
Xbit_r229_c99 bl[99] br[99] wl[229] vdd gnd cell_6t
Xbit_r230_c99 bl[99] br[99] wl[230] vdd gnd cell_6t
Xbit_r231_c99 bl[99] br[99] wl[231] vdd gnd cell_6t
Xbit_r232_c99 bl[99] br[99] wl[232] vdd gnd cell_6t
Xbit_r233_c99 bl[99] br[99] wl[233] vdd gnd cell_6t
Xbit_r234_c99 bl[99] br[99] wl[234] vdd gnd cell_6t
Xbit_r235_c99 bl[99] br[99] wl[235] vdd gnd cell_6t
Xbit_r236_c99 bl[99] br[99] wl[236] vdd gnd cell_6t
Xbit_r237_c99 bl[99] br[99] wl[237] vdd gnd cell_6t
Xbit_r238_c99 bl[99] br[99] wl[238] vdd gnd cell_6t
Xbit_r239_c99 bl[99] br[99] wl[239] vdd gnd cell_6t
Xbit_r240_c99 bl[99] br[99] wl[240] vdd gnd cell_6t
Xbit_r241_c99 bl[99] br[99] wl[241] vdd gnd cell_6t
Xbit_r242_c99 bl[99] br[99] wl[242] vdd gnd cell_6t
Xbit_r243_c99 bl[99] br[99] wl[243] vdd gnd cell_6t
Xbit_r244_c99 bl[99] br[99] wl[244] vdd gnd cell_6t
Xbit_r245_c99 bl[99] br[99] wl[245] vdd gnd cell_6t
Xbit_r246_c99 bl[99] br[99] wl[246] vdd gnd cell_6t
Xbit_r247_c99 bl[99] br[99] wl[247] vdd gnd cell_6t
Xbit_r248_c99 bl[99] br[99] wl[248] vdd gnd cell_6t
Xbit_r249_c99 bl[99] br[99] wl[249] vdd gnd cell_6t
Xbit_r250_c99 bl[99] br[99] wl[250] vdd gnd cell_6t
Xbit_r251_c99 bl[99] br[99] wl[251] vdd gnd cell_6t
Xbit_r252_c99 bl[99] br[99] wl[252] vdd gnd cell_6t
Xbit_r253_c99 bl[99] br[99] wl[253] vdd gnd cell_6t
Xbit_r254_c99 bl[99] br[99] wl[254] vdd gnd cell_6t
Xbit_r255_c99 bl[99] br[99] wl[255] vdd gnd cell_6t
Xbit_r0_c100 bl[100] br[100] wl[0] vdd gnd cell_6t
Xbit_r1_c100 bl[100] br[100] wl[1] vdd gnd cell_6t
Xbit_r2_c100 bl[100] br[100] wl[2] vdd gnd cell_6t
Xbit_r3_c100 bl[100] br[100] wl[3] vdd gnd cell_6t
Xbit_r4_c100 bl[100] br[100] wl[4] vdd gnd cell_6t
Xbit_r5_c100 bl[100] br[100] wl[5] vdd gnd cell_6t
Xbit_r6_c100 bl[100] br[100] wl[6] vdd gnd cell_6t
Xbit_r7_c100 bl[100] br[100] wl[7] vdd gnd cell_6t
Xbit_r8_c100 bl[100] br[100] wl[8] vdd gnd cell_6t
Xbit_r9_c100 bl[100] br[100] wl[9] vdd gnd cell_6t
Xbit_r10_c100 bl[100] br[100] wl[10] vdd gnd cell_6t
Xbit_r11_c100 bl[100] br[100] wl[11] vdd gnd cell_6t
Xbit_r12_c100 bl[100] br[100] wl[12] vdd gnd cell_6t
Xbit_r13_c100 bl[100] br[100] wl[13] vdd gnd cell_6t
Xbit_r14_c100 bl[100] br[100] wl[14] vdd gnd cell_6t
Xbit_r15_c100 bl[100] br[100] wl[15] vdd gnd cell_6t
Xbit_r16_c100 bl[100] br[100] wl[16] vdd gnd cell_6t
Xbit_r17_c100 bl[100] br[100] wl[17] vdd gnd cell_6t
Xbit_r18_c100 bl[100] br[100] wl[18] vdd gnd cell_6t
Xbit_r19_c100 bl[100] br[100] wl[19] vdd gnd cell_6t
Xbit_r20_c100 bl[100] br[100] wl[20] vdd gnd cell_6t
Xbit_r21_c100 bl[100] br[100] wl[21] vdd gnd cell_6t
Xbit_r22_c100 bl[100] br[100] wl[22] vdd gnd cell_6t
Xbit_r23_c100 bl[100] br[100] wl[23] vdd gnd cell_6t
Xbit_r24_c100 bl[100] br[100] wl[24] vdd gnd cell_6t
Xbit_r25_c100 bl[100] br[100] wl[25] vdd gnd cell_6t
Xbit_r26_c100 bl[100] br[100] wl[26] vdd gnd cell_6t
Xbit_r27_c100 bl[100] br[100] wl[27] vdd gnd cell_6t
Xbit_r28_c100 bl[100] br[100] wl[28] vdd gnd cell_6t
Xbit_r29_c100 bl[100] br[100] wl[29] vdd gnd cell_6t
Xbit_r30_c100 bl[100] br[100] wl[30] vdd gnd cell_6t
Xbit_r31_c100 bl[100] br[100] wl[31] vdd gnd cell_6t
Xbit_r32_c100 bl[100] br[100] wl[32] vdd gnd cell_6t
Xbit_r33_c100 bl[100] br[100] wl[33] vdd gnd cell_6t
Xbit_r34_c100 bl[100] br[100] wl[34] vdd gnd cell_6t
Xbit_r35_c100 bl[100] br[100] wl[35] vdd gnd cell_6t
Xbit_r36_c100 bl[100] br[100] wl[36] vdd gnd cell_6t
Xbit_r37_c100 bl[100] br[100] wl[37] vdd gnd cell_6t
Xbit_r38_c100 bl[100] br[100] wl[38] vdd gnd cell_6t
Xbit_r39_c100 bl[100] br[100] wl[39] vdd gnd cell_6t
Xbit_r40_c100 bl[100] br[100] wl[40] vdd gnd cell_6t
Xbit_r41_c100 bl[100] br[100] wl[41] vdd gnd cell_6t
Xbit_r42_c100 bl[100] br[100] wl[42] vdd gnd cell_6t
Xbit_r43_c100 bl[100] br[100] wl[43] vdd gnd cell_6t
Xbit_r44_c100 bl[100] br[100] wl[44] vdd gnd cell_6t
Xbit_r45_c100 bl[100] br[100] wl[45] vdd gnd cell_6t
Xbit_r46_c100 bl[100] br[100] wl[46] vdd gnd cell_6t
Xbit_r47_c100 bl[100] br[100] wl[47] vdd gnd cell_6t
Xbit_r48_c100 bl[100] br[100] wl[48] vdd gnd cell_6t
Xbit_r49_c100 bl[100] br[100] wl[49] vdd gnd cell_6t
Xbit_r50_c100 bl[100] br[100] wl[50] vdd gnd cell_6t
Xbit_r51_c100 bl[100] br[100] wl[51] vdd gnd cell_6t
Xbit_r52_c100 bl[100] br[100] wl[52] vdd gnd cell_6t
Xbit_r53_c100 bl[100] br[100] wl[53] vdd gnd cell_6t
Xbit_r54_c100 bl[100] br[100] wl[54] vdd gnd cell_6t
Xbit_r55_c100 bl[100] br[100] wl[55] vdd gnd cell_6t
Xbit_r56_c100 bl[100] br[100] wl[56] vdd gnd cell_6t
Xbit_r57_c100 bl[100] br[100] wl[57] vdd gnd cell_6t
Xbit_r58_c100 bl[100] br[100] wl[58] vdd gnd cell_6t
Xbit_r59_c100 bl[100] br[100] wl[59] vdd gnd cell_6t
Xbit_r60_c100 bl[100] br[100] wl[60] vdd gnd cell_6t
Xbit_r61_c100 bl[100] br[100] wl[61] vdd gnd cell_6t
Xbit_r62_c100 bl[100] br[100] wl[62] vdd gnd cell_6t
Xbit_r63_c100 bl[100] br[100] wl[63] vdd gnd cell_6t
Xbit_r64_c100 bl[100] br[100] wl[64] vdd gnd cell_6t
Xbit_r65_c100 bl[100] br[100] wl[65] vdd gnd cell_6t
Xbit_r66_c100 bl[100] br[100] wl[66] vdd gnd cell_6t
Xbit_r67_c100 bl[100] br[100] wl[67] vdd gnd cell_6t
Xbit_r68_c100 bl[100] br[100] wl[68] vdd gnd cell_6t
Xbit_r69_c100 bl[100] br[100] wl[69] vdd gnd cell_6t
Xbit_r70_c100 bl[100] br[100] wl[70] vdd gnd cell_6t
Xbit_r71_c100 bl[100] br[100] wl[71] vdd gnd cell_6t
Xbit_r72_c100 bl[100] br[100] wl[72] vdd gnd cell_6t
Xbit_r73_c100 bl[100] br[100] wl[73] vdd gnd cell_6t
Xbit_r74_c100 bl[100] br[100] wl[74] vdd gnd cell_6t
Xbit_r75_c100 bl[100] br[100] wl[75] vdd gnd cell_6t
Xbit_r76_c100 bl[100] br[100] wl[76] vdd gnd cell_6t
Xbit_r77_c100 bl[100] br[100] wl[77] vdd gnd cell_6t
Xbit_r78_c100 bl[100] br[100] wl[78] vdd gnd cell_6t
Xbit_r79_c100 bl[100] br[100] wl[79] vdd gnd cell_6t
Xbit_r80_c100 bl[100] br[100] wl[80] vdd gnd cell_6t
Xbit_r81_c100 bl[100] br[100] wl[81] vdd gnd cell_6t
Xbit_r82_c100 bl[100] br[100] wl[82] vdd gnd cell_6t
Xbit_r83_c100 bl[100] br[100] wl[83] vdd gnd cell_6t
Xbit_r84_c100 bl[100] br[100] wl[84] vdd gnd cell_6t
Xbit_r85_c100 bl[100] br[100] wl[85] vdd gnd cell_6t
Xbit_r86_c100 bl[100] br[100] wl[86] vdd gnd cell_6t
Xbit_r87_c100 bl[100] br[100] wl[87] vdd gnd cell_6t
Xbit_r88_c100 bl[100] br[100] wl[88] vdd gnd cell_6t
Xbit_r89_c100 bl[100] br[100] wl[89] vdd gnd cell_6t
Xbit_r90_c100 bl[100] br[100] wl[90] vdd gnd cell_6t
Xbit_r91_c100 bl[100] br[100] wl[91] vdd gnd cell_6t
Xbit_r92_c100 bl[100] br[100] wl[92] vdd gnd cell_6t
Xbit_r93_c100 bl[100] br[100] wl[93] vdd gnd cell_6t
Xbit_r94_c100 bl[100] br[100] wl[94] vdd gnd cell_6t
Xbit_r95_c100 bl[100] br[100] wl[95] vdd gnd cell_6t
Xbit_r96_c100 bl[100] br[100] wl[96] vdd gnd cell_6t
Xbit_r97_c100 bl[100] br[100] wl[97] vdd gnd cell_6t
Xbit_r98_c100 bl[100] br[100] wl[98] vdd gnd cell_6t
Xbit_r99_c100 bl[100] br[100] wl[99] vdd gnd cell_6t
Xbit_r100_c100 bl[100] br[100] wl[100] vdd gnd cell_6t
Xbit_r101_c100 bl[100] br[100] wl[101] vdd gnd cell_6t
Xbit_r102_c100 bl[100] br[100] wl[102] vdd gnd cell_6t
Xbit_r103_c100 bl[100] br[100] wl[103] vdd gnd cell_6t
Xbit_r104_c100 bl[100] br[100] wl[104] vdd gnd cell_6t
Xbit_r105_c100 bl[100] br[100] wl[105] vdd gnd cell_6t
Xbit_r106_c100 bl[100] br[100] wl[106] vdd gnd cell_6t
Xbit_r107_c100 bl[100] br[100] wl[107] vdd gnd cell_6t
Xbit_r108_c100 bl[100] br[100] wl[108] vdd gnd cell_6t
Xbit_r109_c100 bl[100] br[100] wl[109] vdd gnd cell_6t
Xbit_r110_c100 bl[100] br[100] wl[110] vdd gnd cell_6t
Xbit_r111_c100 bl[100] br[100] wl[111] vdd gnd cell_6t
Xbit_r112_c100 bl[100] br[100] wl[112] vdd gnd cell_6t
Xbit_r113_c100 bl[100] br[100] wl[113] vdd gnd cell_6t
Xbit_r114_c100 bl[100] br[100] wl[114] vdd gnd cell_6t
Xbit_r115_c100 bl[100] br[100] wl[115] vdd gnd cell_6t
Xbit_r116_c100 bl[100] br[100] wl[116] vdd gnd cell_6t
Xbit_r117_c100 bl[100] br[100] wl[117] vdd gnd cell_6t
Xbit_r118_c100 bl[100] br[100] wl[118] vdd gnd cell_6t
Xbit_r119_c100 bl[100] br[100] wl[119] vdd gnd cell_6t
Xbit_r120_c100 bl[100] br[100] wl[120] vdd gnd cell_6t
Xbit_r121_c100 bl[100] br[100] wl[121] vdd gnd cell_6t
Xbit_r122_c100 bl[100] br[100] wl[122] vdd gnd cell_6t
Xbit_r123_c100 bl[100] br[100] wl[123] vdd gnd cell_6t
Xbit_r124_c100 bl[100] br[100] wl[124] vdd gnd cell_6t
Xbit_r125_c100 bl[100] br[100] wl[125] vdd gnd cell_6t
Xbit_r126_c100 bl[100] br[100] wl[126] vdd gnd cell_6t
Xbit_r127_c100 bl[100] br[100] wl[127] vdd gnd cell_6t
Xbit_r128_c100 bl[100] br[100] wl[128] vdd gnd cell_6t
Xbit_r129_c100 bl[100] br[100] wl[129] vdd gnd cell_6t
Xbit_r130_c100 bl[100] br[100] wl[130] vdd gnd cell_6t
Xbit_r131_c100 bl[100] br[100] wl[131] vdd gnd cell_6t
Xbit_r132_c100 bl[100] br[100] wl[132] vdd gnd cell_6t
Xbit_r133_c100 bl[100] br[100] wl[133] vdd gnd cell_6t
Xbit_r134_c100 bl[100] br[100] wl[134] vdd gnd cell_6t
Xbit_r135_c100 bl[100] br[100] wl[135] vdd gnd cell_6t
Xbit_r136_c100 bl[100] br[100] wl[136] vdd gnd cell_6t
Xbit_r137_c100 bl[100] br[100] wl[137] vdd gnd cell_6t
Xbit_r138_c100 bl[100] br[100] wl[138] vdd gnd cell_6t
Xbit_r139_c100 bl[100] br[100] wl[139] vdd gnd cell_6t
Xbit_r140_c100 bl[100] br[100] wl[140] vdd gnd cell_6t
Xbit_r141_c100 bl[100] br[100] wl[141] vdd gnd cell_6t
Xbit_r142_c100 bl[100] br[100] wl[142] vdd gnd cell_6t
Xbit_r143_c100 bl[100] br[100] wl[143] vdd gnd cell_6t
Xbit_r144_c100 bl[100] br[100] wl[144] vdd gnd cell_6t
Xbit_r145_c100 bl[100] br[100] wl[145] vdd gnd cell_6t
Xbit_r146_c100 bl[100] br[100] wl[146] vdd gnd cell_6t
Xbit_r147_c100 bl[100] br[100] wl[147] vdd gnd cell_6t
Xbit_r148_c100 bl[100] br[100] wl[148] vdd gnd cell_6t
Xbit_r149_c100 bl[100] br[100] wl[149] vdd gnd cell_6t
Xbit_r150_c100 bl[100] br[100] wl[150] vdd gnd cell_6t
Xbit_r151_c100 bl[100] br[100] wl[151] vdd gnd cell_6t
Xbit_r152_c100 bl[100] br[100] wl[152] vdd gnd cell_6t
Xbit_r153_c100 bl[100] br[100] wl[153] vdd gnd cell_6t
Xbit_r154_c100 bl[100] br[100] wl[154] vdd gnd cell_6t
Xbit_r155_c100 bl[100] br[100] wl[155] vdd gnd cell_6t
Xbit_r156_c100 bl[100] br[100] wl[156] vdd gnd cell_6t
Xbit_r157_c100 bl[100] br[100] wl[157] vdd gnd cell_6t
Xbit_r158_c100 bl[100] br[100] wl[158] vdd gnd cell_6t
Xbit_r159_c100 bl[100] br[100] wl[159] vdd gnd cell_6t
Xbit_r160_c100 bl[100] br[100] wl[160] vdd gnd cell_6t
Xbit_r161_c100 bl[100] br[100] wl[161] vdd gnd cell_6t
Xbit_r162_c100 bl[100] br[100] wl[162] vdd gnd cell_6t
Xbit_r163_c100 bl[100] br[100] wl[163] vdd gnd cell_6t
Xbit_r164_c100 bl[100] br[100] wl[164] vdd gnd cell_6t
Xbit_r165_c100 bl[100] br[100] wl[165] vdd gnd cell_6t
Xbit_r166_c100 bl[100] br[100] wl[166] vdd gnd cell_6t
Xbit_r167_c100 bl[100] br[100] wl[167] vdd gnd cell_6t
Xbit_r168_c100 bl[100] br[100] wl[168] vdd gnd cell_6t
Xbit_r169_c100 bl[100] br[100] wl[169] vdd gnd cell_6t
Xbit_r170_c100 bl[100] br[100] wl[170] vdd gnd cell_6t
Xbit_r171_c100 bl[100] br[100] wl[171] vdd gnd cell_6t
Xbit_r172_c100 bl[100] br[100] wl[172] vdd gnd cell_6t
Xbit_r173_c100 bl[100] br[100] wl[173] vdd gnd cell_6t
Xbit_r174_c100 bl[100] br[100] wl[174] vdd gnd cell_6t
Xbit_r175_c100 bl[100] br[100] wl[175] vdd gnd cell_6t
Xbit_r176_c100 bl[100] br[100] wl[176] vdd gnd cell_6t
Xbit_r177_c100 bl[100] br[100] wl[177] vdd gnd cell_6t
Xbit_r178_c100 bl[100] br[100] wl[178] vdd gnd cell_6t
Xbit_r179_c100 bl[100] br[100] wl[179] vdd gnd cell_6t
Xbit_r180_c100 bl[100] br[100] wl[180] vdd gnd cell_6t
Xbit_r181_c100 bl[100] br[100] wl[181] vdd gnd cell_6t
Xbit_r182_c100 bl[100] br[100] wl[182] vdd gnd cell_6t
Xbit_r183_c100 bl[100] br[100] wl[183] vdd gnd cell_6t
Xbit_r184_c100 bl[100] br[100] wl[184] vdd gnd cell_6t
Xbit_r185_c100 bl[100] br[100] wl[185] vdd gnd cell_6t
Xbit_r186_c100 bl[100] br[100] wl[186] vdd gnd cell_6t
Xbit_r187_c100 bl[100] br[100] wl[187] vdd gnd cell_6t
Xbit_r188_c100 bl[100] br[100] wl[188] vdd gnd cell_6t
Xbit_r189_c100 bl[100] br[100] wl[189] vdd gnd cell_6t
Xbit_r190_c100 bl[100] br[100] wl[190] vdd gnd cell_6t
Xbit_r191_c100 bl[100] br[100] wl[191] vdd gnd cell_6t
Xbit_r192_c100 bl[100] br[100] wl[192] vdd gnd cell_6t
Xbit_r193_c100 bl[100] br[100] wl[193] vdd gnd cell_6t
Xbit_r194_c100 bl[100] br[100] wl[194] vdd gnd cell_6t
Xbit_r195_c100 bl[100] br[100] wl[195] vdd gnd cell_6t
Xbit_r196_c100 bl[100] br[100] wl[196] vdd gnd cell_6t
Xbit_r197_c100 bl[100] br[100] wl[197] vdd gnd cell_6t
Xbit_r198_c100 bl[100] br[100] wl[198] vdd gnd cell_6t
Xbit_r199_c100 bl[100] br[100] wl[199] vdd gnd cell_6t
Xbit_r200_c100 bl[100] br[100] wl[200] vdd gnd cell_6t
Xbit_r201_c100 bl[100] br[100] wl[201] vdd gnd cell_6t
Xbit_r202_c100 bl[100] br[100] wl[202] vdd gnd cell_6t
Xbit_r203_c100 bl[100] br[100] wl[203] vdd gnd cell_6t
Xbit_r204_c100 bl[100] br[100] wl[204] vdd gnd cell_6t
Xbit_r205_c100 bl[100] br[100] wl[205] vdd gnd cell_6t
Xbit_r206_c100 bl[100] br[100] wl[206] vdd gnd cell_6t
Xbit_r207_c100 bl[100] br[100] wl[207] vdd gnd cell_6t
Xbit_r208_c100 bl[100] br[100] wl[208] vdd gnd cell_6t
Xbit_r209_c100 bl[100] br[100] wl[209] vdd gnd cell_6t
Xbit_r210_c100 bl[100] br[100] wl[210] vdd gnd cell_6t
Xbit_r211_c100 bl[100] br[100] wl[211] vdd gnd cell_6t
Xbit_r212_c100 bl[100] br[100] wl[212] vdd gnd cell_6t
Xbit_r213_c100 bl[100] br[100] wl[213] vdd gnd cell_6t
Xbit_r214_c100 bl[100] br[100] wl[214] vdd gnd cell_6t
Xbit_r215_c100 bl[100] br[100] wl[215] vdd gnd cell_6t
Xbit_r216_c100 bl[100] br[100] wl[216] vdd gnd cell_6t
Xbit_r217_c100 bl[100] br[100] wl[217] vdd gnd cell_6t
Xbit_r218_c100 bl[100] br[100] wl[218] vdd gnd cell_6t
Xbit_r219_c100 bl[100] br[100] wl[219] vdd gnd cell_6t
Xbit_r220_c100 bl[100] br[100] wl[220] vdd gnd cell_6t
Xbit_r221_c100 bl[100] br[100] wl[221] vdd gnd cell_6t
Xbit_r222_c100 bl[100] br[100] wl[222] vdd gnd cell_6t
Xbit_r223_c100 bl[100] br[100] wl[223] vdd gnd cell_6t
Xbit_r224_c100 bl[100] br[100] wl[224] vdd gnd cell_6t
Xbit_r225_c100 bl[100] br[100] wl[225] vdd gnd cell_6t
Xbit_r226_c100 bl[100] br[100] wl[226] vdd gnd cell_6t
Xbit_r227_c100 bl[100] br[100] wl[227] vdd gnd cell_6t
Xbit_r228_c100 bl[100] br[100] wl[228] vdd gnd cell_6t
Xbit_r229_c100 bl[100] br[100] wl[229] vdd gnd cell_6t
Xbit_r230_c100 bl[100] br[100] wl[230] vdd gnd cell_6t
Xbit_r231_c100 bl[100] br[100] wl[231] vdd gnd cell_6t
Xbit_r232_c100 bl[100] br[100] wl[232] vdd gnd cell_6t
Xbit_r233_c100 bl[100] br[100] wl[233] vdd gnd cell_6t
Xbit_r234_c100 bl[100] br[100] wl[234] vdd gnd cell_6t
Xbit_r235_c100 bl[100] br[100] wl[235] vdd gnd cell_6t
Xbit_r236_c100 bl[100] br[100] wl[236] vdd gnd cell_6t
Xbit_r237_c100 bl[100] br[100] wl[237] vdd gnd cell_6t
Xbit_r238_c100 bl[100] br[100] wl[238] vdd gnd cell_6t
Xbit_r239_c100 bl[100] br[100] wl[239] vdd gnd cell_6t
Xbit_r240_c100 bl[100] br[100] wl[240] vdd gnd cell_6t
Xbit_r241_c100 bl[100] br[100] wl[241] vdd gnd cell_6t
Xbit_r242_c100 bl[100] br[100] wl[242] vdd gnd cell_6t
Xbit_r243_c100 bl[100] br[100] wl[243] vdd gnd cell_6t
Xbit_r244_c100 bl[100] br[100] wl[244] vdd gnd cell_6t
Xbit_r245_c100 bl[100] br[100] wl[245] vdd gnd cell_6t
Xbit_r246_c100 bl[100] br[100] wl[246] vdd gnd cell_6t
Xbit_r247_c100 bl[100] br[100] wl[247] vdd gnd cell_6t
Xbit_r248_c100 bl[100] br[100] wl[248] vdd gnd cell_6t
Xbit_r249_c100 bl[100] br[100] wl[249] vdd gnd cell_6t
Xbit_r250_c100 bl[100] br[100] wl[250] vdd gnd cell_6t
Xbit_r251_c100 bl[100] br[100] wl[251] vdd gnd cell_6t
Xbit_r252_c100 bl[100] br[100] wl[252] vdd gnd cell_6t
Xbit_r253_c100 bl[100] br[100] wl[253] vdd gnd cell_6t
Xbit_r254_c100 bl[100] br[100] wl[254] vdd gnd cell_6t
Xbit_r255_c100 bl[100] br[100] wl[255] vdd gnd cell_6t
Xbit_r0_c101 bl[101] br[101] wl[0] vdd gnd cell_6t
Xbit_r1_c101 bl[101] br[101] wl[1] vdd gnd cell_6t
Xbit_r2_c101 bl[101] br[101] wl[2] vdd gnd cell_6t
Xbit_r3_c101 bl[101] br[101] wl[3] vdd gnd cell_6t
Xbit_r4_c101 bl[101] br[101] wl[4] vdd gnd cell_6t
Xbit_r5_c101 bl[101] br[101] wl[5] vdd gnd cell_6t
Xbit_r6_c101 bl[101] br[101] wl[6] vdd gnd cell_6t
Xbit_r7_c101 bl[101] br[101] wl[7] vdd gnd cell_6t
Xbit_r8_c101 bl[101] br[101] wl[8] vdd gnd cell_6t
Xbit_r9_c101 bl[101] br[101] wl[9] vdd gnd cell_6t
Xbit_r10_c101 bl[101] br[101] wl[10] vdd gnd cell_6t
Xbit_r11_c101 bl[101] br[101] wl[11] vdd gnd cell_6t
Xbit_r12_c101 bl[101] br[101] wl[12] vdd gnd cell_6t
Xbit_r13_c101 bl[101] br[101] wl[13] vdd gnd cell_6t
Xbit_r14_c101 bl[101] br[101] wl[14] vdd gnd cell_6t
Xbit_r15_c101 bl[101] br[101] wl[15] vdd gnd cell_6t
Xbit_r16_c101 bl[101] br[101] wl[16] vdd gnd cell_6t
Xbit_r17_c101 bl[101] br[101] wl[17] vdd gnd cell_6t
Xbit_r18_c101 bl[101] br[101] wl[18] vdd gnd cell_6t
Xbit_r19_c101 bl[101] br[101] wl[19] vdd gnd cell_6t
Xbit_r20_c101 bl[101] br[101] wl[20] vdd gnd cell_6t
Xbit_r21_c101 bl[101] br[101] wl[21] vdd gnd cell_6t
Xbit_r22_c101 bl[101] br[101] wl[22] vdd gnd cell_6t
Xbit_r23_c101 bl[101] br[101] wl[23] vdd gnd cell_6t
Xbit_r24_c101 bl[101] br[101] wl[24] vdd gnd cell_6t
Xbit_r25_c101 bl[101] br[101] wl[25] vdd gnd cell_6t
Xbit_r26_c101 bl[101] br[101] wl[26] vdd gnd cell_6t
Xbit_r27_c101 bl[101] br[101] wl[27] vdd gnd cell_6t
Xbit_r28_c101 bl[101] br[101] wl[28] vdd gnd cell_6t
Xbit_r29_c101 bl[101] br[101] wl[29] vdd gnd cell_6t
Xbit_r30_c101 bl[101] br[101] wl[30] vdd gnd cell_6t
Xbit_r31_c101 bl[101] br[101] wl[31] vdd gnd cell_6t
Xbit_r32_c101 bl[101] br[101] wl[32] vdd gnd cell_6t
Xbit_r33_c101 bl[101] br[101] wl[33] vdd gnd cell_6t
Xbit_r34_c101 bl[101] br[101] wl[34] vdd gnd cell_6t
Xbit_r35_c101 bl[101] br[101] wl[35] vdd gnd cell_6t
Xbit_r36_c101 bl[101] br[101] wl[36] vdd gnd cell_6t
Xbit_r37_c101 bl[101] br[101] wl[37] vdd gnd cell_6t
Xbit_r38_c101 bl[101] br[101] wl[38] vdd gnd cell_6t
Xbit_r39_c101 bl[101] br[101] wl[39] vdd gnd cell_6t
Xbit_r40_c101 bl[101] br[101] wl[40] vdd gnd cell_6t
Xbit_r41_c101 bl[101] br[101] wl[41] vdd gnd cell_6t
Xbit_r42_c101 bl[101] br[101] wl[42] vdd gnd cell_6t
Xbit_r43_c101 bl[101] br[101] wl[43] vdd gnd cell_6t
Xbit_r44_c101 bl[101] br[101] wl[44] vdd gnd cell_6t
Xbit_r45_c101 bl[101] br[101] wl[45] vdd gnd cell_6t
Xbit_r46_c101 bl[101] br[101] wl[46] vdd gnd cell_6t
Xbit_r47_c101 bl[101] br[101] wl[47] vdd gnd cell_6t
Xbit_r48_c101 bl[101] br[101] wl[48] vdd gnd cell_6t
Xbit_r49_c101 bl[101] br[101] wl[49] vdd gnd cell_6t
Xbit_r50_c101 bl[101] br[101] wl[50] vdd gnd cell_6t
Xbit_r51_c101 bl[101] br[101] wl[51] vdd gnd cell_6t
Xbit_r52_c101 bl[101] br[101] wl[52] vdd gnd cell_6t
Xbit_r53_c101 bl[101] br[101] wl[53] vdd gnd cell_6t
Xbit_r54_c101 bl[101] br[101] wl[54] vdd gnd cell_6t
Xbit_r55_c101 bl[101] br[101] wl[55] vdd gnd cell_6t
Xbit_r56_c101 bl[101] br[101] wl[56] vdd gnd cell_6t
Xbit_r57_c101 bl[101] br[101] wl[57] vdd gnd cell_6t
Xbit_r58_c101 bl[101] br[101] wl[58] vdd gnd cell_6t
Xbit_r59_c101 bl[101] br[101] wl[59] vdd gnd cell_6t
Xbit_r60_c101 bl[101] br[101] wl[60] vdd gnd cell_6t
Xbit_r61_c101 bl[101] br[101] wl[61] vdd gnd cell_6t
Xbit_r62_c101 bl[101] br[101] wl[62] vdd gnd cell_6t
Xbit_r63_c101 bl[101] br[101] wl[63] vdd gnd cell_6t
Xbit_r64_c101 bl[101] br[101] wl[64] vdd gnd cell_6t
Xbit_r65_c101 bl[101] br[101] wl[65] vdd gnd cell_6t
Xbit_r66_c101 bl[101] br[101] wl[66] vdd gnd cell_6t
Xbit_r67_c101 bl[101] br[101] wl[67] vdd gnd cell_6t
Xbit_r68_c101 bl[101] br[101] wl[68] vdd gnd cell_6t
Xbit_r69_c101 bl[101] br[101] wl[69] vdd gnd cell_6t
Xbit_r70_c101 bl[101] br[101] wl[70] vdd gnd cell_6t
Xbit_r71_c101 bl[101] br[101] wl[71] vdd gnd cell_6t
Xbit_r72_c101 bl[101] br[101] wl[72] vdd gnd cell_6t
Xbit_r73_c101 bl[101] br[101] wl[73] vdd gnd cell_6t
Xbit_r74_c101 bl[101] br[101] wl[74] vdd gnd cell_6t
Xbit_r75_c101 bl[101] br[101] wl[75] vdd gnd cell_6t
Xbit_r76_c101 bl[101] br[101] wl[76] vdd gnd cell_6t
Xbit_r77_c101 bl[101] br[101] wl[77] vdd gnd cell_6t
Xbit_r78_c101 bl[101] br[101] wl[78] vdd gnd cell_6t
Xbit_r79_c101 bl[101] br[101] wl[79] vdd gnd cell_6t
Xbit_r80_c101 bl[101] br[101] wl[80] vdd gnd cell_6t
Xbit_r81_c101 bl[101] br[101] wl[81] vdd gnd cell_6t
Xbit_r82_c101 bl[101] br[101] wl[82] vdd gnd cell_6t
Xbit_r83_c101 bl[101] br[101] wl[83] vdd gnd cell_6t
Xbit_r84_c101 bl[101] br[101] wl[84] vdd gnd cell_6t
Xbit_r85_c101 bl[101] br[101] wl[85] vdd gnd cell_6t
Xbit_r86_c101 bl[101] br[101] wl[86] vdd gnd cell_6t
Xbit_r87_c101 bl[101] br[101] wl[87] vdd gnd cell_6t
Xbit_r88_c101 bl[101] br[101] wl[88] vdd gnd cell_6t
Xbit_r89_c101 bl[101] br[101] wl[89] vdd gnd cell_6t
Xbit_r90_c101 bl[101] br[101] wl[90] vdd gnd cell_6t
Xbit_r91_c101 bl[101] br[101] wl[91] vdd gnd cell_6t
Xbit_r92_c101 bl[101] br[101] wl[92] vdd gnd cell_6t
Xbit_r93_c101 bl[101] br[101] wl[93] vdd gnd cell_6t
Xbit_r94_c101 bl[101] br[101] wl[94] vdd gnd cell_6t
Xbit_r95_c101 bl[101] br[101] wl[95] vdd gnd cell_6t
Xbit_r96_c101 bl[101] br[101] wl[96] vdd gnd cell_6t
Xbit_r97_c101 bl[101] br[101] wl[97] vdd gnd cell_6t
Xbit_r98_c101 bl[101] br[101] wl[98] vdd gnd cell_6t
Xbit_r99_c101 bl[101] br[101] wl[99] vdd gnd cell_6t
Xbit_r100_c101 bl[101] br[101] wl[100] vdd gnd cell_6t
Xbit_r101_c101 bl[101] br[101] wl[101] vdd gnd cell_6t
Xbit_r102_c101 bl[101] br[101] wl[102] vdd gnd cell_6t
Xbit_r103_c101 bl[101] br[101] wl[103] vdd gnd cell_6t
Xbit_r104_c101 bl[101] br[101] wl[104] vdd gnd cell_6t
Xbit_r105_c101 bl[101] br[101] wl[105] vdd gnd cell_6t
Xbit_r106_c101 bl[101] br[101] wl[106] vdd gnd cell_6t
Xbit_r107_c101 bl[101] br[101] wl[107] vdd gnd cell_6t
Xbit_r108_c101 bl[101] br[101] wl[108] vdd gnd cell_6t
Xbit_r109_c101 bl[101] br[101] wl[109] vdd gnd cell_6t
Xbit_r110_c101 bl[101] br[101] wl[110] vdd gnd cell_6t
Xbit_r111_c101 bl[101] br[101] wl[111] vdd gnd cell_6t
Xbit_r112_c101 bl[101] br[101] wl[112] vdd gnd cell_6t
Xbit_r113_c101 bl[101] br[101] wl[113] vdd gnd cell_6t
Xbit_r114_c101 bl[101] br[101] wl[114] vdd gnd cell_6t
Xbit_r115_c101 bl[101] br[101] wl[115] vdd gnd cell_6t
Xbit_r116_c101 bl[101] br[101] wl[116] vdd gnd cell_6t
Xbit_r117_c101 bl[101] br[101] wl[117] vdd gnd cell_6t
Xbit_r118_c101 bl[101] br[101] wl[118] vdd gnd cell_6t
Xbit_r119_c101 bl[101] br[101] wl[119] vdd gnd cell_6t
Xbit_r120_c101 bl[101] br[101] wl[120] vdd gnd cell_6t
Xbit_r121_c101 bl[101] br[101] wl[121] vdd gnd cell_6t
Xbit_r122_c101 bl[101] br[101] wl[122] vdd gnd cell_6t
Xbit_r123_c101 bl[101] br[101] wl[123] vdd gnd cell_6t
Xbit_r124_c101 bl[101] br[101] wl[124] vdd gnd cell_6t
Xbit_r125_c101 bl[101] br[101] wl[125] vdd gnd cell_6t
Xbit_r126_c101 bl[101] br[101] wl[126] vdd gnd cell_6t
Xbit_r127_c101 bl[101] br[101] wl[127] vdd gnd cell_6t
Xbit_r128_c101 bl[101] br[101] wl[128] vdd gnd cell_6t
Xbit_r129_c101 bl[101] br[101] wl[129] vdd gnd cell_6t
Xbit_r130_c101 bl[101] br[101] wl[130] vdd gnd cell_6t
Xbit_r131_c101 bl[101] br[101] wl[131] vdd gnd cell_6t
Xbit_r132_c101 bl[101] br[101] wl[132] vdd gnd cell_6t
Xbit_r133_c101 bl[101] br[101] wl[133] vdd gnd cell_6t
Xbit_r134_c101 bl[101] br[101] wl[134] vdd gnd cell_6t
Xbit_r135_c101 bl[101] br[101] wl[135] vdd gnd cell_6t
Xbit_r136_c101 bl[101] br[101] wl[136] vdd gnd cell_6t
Xbit_r137_c101 bl[101] br[101] wl[137] vdd gnd cell_6t
Xbit_r138_c101 bl[101] br[101] wl[138] vdd gnd cell_6t
Xbit_r139_c101 bl[101] br[101] wl[139] vdd gnd cell_6t
Xbit_r140_c101 bl[101] br[101] wl[140] vdd gnd cell_6t
Xbit_r141_c101 bl[101] br[101] wl[141] vdd gnd cell_6t
Xbit_r142_c101 bl[101] br[101] wl[142] vdd gnd cell_6t
Xbit_r143_c101 bl[101] br[101] wl[143] vdd gnd cell_6t
Xbit_r144_c101 bl[101] br[101] wl[144] vdd gnd cell_6t
Xbit_r145_c101 bl[101] br[101] wl[145] vdd gnd cell_6t
Xbit_r146_c101 bl[101] br[101] wl[146] vdd gnd cell_6t
Xbit_r147_c101 bl[101] br[101] wl[147] vdd gnd cell_6t
Xbit_r148_c101 bl[101] br[101] wl[148] vdd gnd cell_6t
Xbit_r149_c101 bl[101] br[101] wl[149] vdd gnd cell_6t
Xbit_r150_c101 bl[101] br[101] wl[150] vdd gnd cell_6t
Xbit_r151_c101 bl[101] br[101] wl[151] vdd gnd cell_6t
Xbit_r152_c101 bl[101] br[101] wl[152] vdd gnd cell_6t
Xbit_r153_c101 bl[101] br[101] wl[153] vdd gnd cell_6t
Xbit_r154_c101 bl[101] br[101] wl[154] vdd gnd cell_6t
Xbit_r155_c101 bl[101] br[101] wl[155] vdd gnd cell_6t
Xbit_r156_c101 bl[101] br[101] wl[156] vdd gnd cell_6t
Xbit_r157_c101 bl[101] br[101] wl[157] vdd gnd cell_6t
Xbit_r158_c101 bl[101] br[101] wl[158] vdd gnd cell_6t
Xbit_r159_c101 bl[101] br[101] wl[159] vdd gnd cell_6t
Xbit_r160_c101 bl[101] br[101] wl[160] vdd gnd cell_6t
Xbit_r161_c101 bl[101] br[101] wl[161] vdd gnd cell_6t
Xbit_r162_c101 bl[101] br[101] wl[162] vdd gnd cell_6t
Xbit_r163_c101 bl[101] br[101] wl[163] vdd gnd cell_6t
Xbit_r164_c101 bl[101] br[101] wl[164] vdd gnd cell_6t
Xbit_r165_c101 bl[101] br[101] wl[165] vdd gnd cell_6t
Xbit_r166_c101 bl[101] br[101] wl[166] vdd gnd cell_6t
Xbit_r167_c101 bl[101] br[101] wl[167] vdd gnd cell_6t
Xbit_r168_c101 bl[101] br[101] wl[168] vdd gnd cell_6t
Xbit_r169_c101 bl[101] br[101] wl[169] vdd gnd cell_6t
Xbit_r170_c101 bl[101] br[101] wl[170] vdd gnd cell_6t
Xbit_r171_c101 bl[101] br[101] wl[171] vdd gnd cell_6t
Xbit_r172_c101 bl[101] br[101] wl[172] vdd gnd cell_6t
Xbit_r173_c101 bl[101] br[101] wl[173] vdd gnd cell_6t
Xbit_r174_c101 bl[101] br[101] wl[174] vdd gnd cell_6t
Xbit_r175_c101 bl[101] br[101] wl[175] vdd gnd cell_6t
Xbit_r176_c101 bl[101] br[101] wl[176] vdd gnd cell_6t
Xbit_r177_c101 bl[101] br[101] wl[177] vdd gnd cell_6t
Xbit_r178_c101 bl[101] br[101] wl[178] vdd gnd cell_6t
Xbit_r179_c101 bl[101] br[101] wl[179] vdd gnd cell_6t
Xbit_r180_c101 bl[101] br[101] wl[180] vdd gnd cell_6t
Xbit_r181_c101 bl[101] br[101] wl[181] vdd gnd cell_6t
Xbit_r182_c101 bl[101] br[101] wl[182] vdd gnd cell_6t
Xbit_r183_c101 bl[101] br[101] wl[183] vdd gnd cell_6t
Xbit_r184_c101 bl[101] br[101] wl[184] vdd gnd cell_6t
Xbit_r185_c101 bl[101] br[101] wl[185] vdd gnd cell_6t
Xbit_r186_c101 bl[101] br[101] wl[186] vdd gnd cell_6t
Xbit_r187_c101 bl[101] br[101] wl[187] vdd gnd cell_6t
Xbit_r188_c101 bl[101] br[101] wl[188] vdd gnd cell_6t
Xbit_r189_c101 bl[101] br[101] wl[189] vdd gnd cell_6t
Xbit_r190_c101 bl[101] br[101] wl[190] vdd gnd cell_6t
Xbit_r191_c101 bl[101] br[101] wl[191] vdd gnd cell_6t
Xbit_r192_c101 bl[101] br[101] wl[192] vdd gnd cell_6t
Xbit_r193_c101 bl[101] br[101] wl[193] vdd gnd cell_6t
Xbit_r194_c101 bl[101] br[101] wl[194] vdd gnd cell_6t
Xbit_r195_c101 bl[101] br[101] wl[195] vdd gnd cell_6t
Xbit_r196_c101 bl[101] br[101] wl[196] vdd gnd cell_6t
Xbit_r197_c101 bl[101] br[101] wl[197] vdd gnd cell_6t
Xbit_r198_c101 bl[101] br[101] wl[198] vdd gnd cell_6t
Xbit_r199_c101 bl[101] br[101] wl[199] vdd gnd cell_6t
Xbit_r200_c101 bl[101] br[101] wl[200] vdd gnd cell_6t
Xbit_r201_c101 bl[101] br[101] wl[201] vdd gnd cell_6t
Xbit_r202_c101 bl[101] br[101] wl[202] vdd gnd cell_6t
Xbit_r203_c101 bl[101] br[101] wl[203] vdd gnd cell_6t
Xbit_r204_c101 bl[101] br[101] wl[204] vdd gnd cell_6t
Xbit_r205_c101 bl[101] br[101] wl[205] vdd gnd cell_6t
Xbit_r206_c101 bl[101] br[101] wl[206] vdd gnd cell_6t
Xbit_r207_c101 bl[101] br[101] wl[207] vdd gnd cell_6t
Xbit_r208_c101 bl[101] br[101] wl[208] vdd gnd cell_6t
Xbit_r209_c101 bl[101] br[101] wl[209] vdd gnd cell_6t
Xbit_r210_c101 bl[101] br[101] wl[210] vdd gnd cell_6t
Xbit_r211_c101 bl[101] br[101] wl[211] vdd gnd cell_6t
Xbit_r212_c101 bl[101] br[101] wl[212] vdd gnd cell_6t
Xbit_r213_c101 bl[101] br[101] wl[213] vdd gnd cell_6t
Xbit_r214_c101 bl[101] br[101] wl[214] vdd gnd cell_6t
Xbit_r215_c101 bl[101] br[101] wl[215] vdd gnd cell_6t
Xbit_r216_c101 bl[101] br[101] wl[216] vdd gnd cell_6t
Xbit_r217_c101 bl[101] br[101] wl[217] vdd gnd cell_6t
Xbit_r218_c101 bl[101] br[101] wl[218] vdd gnd cell_6t
Xbit_r219_c101 bl[101] br[101] wl[219] vdd gnd cell_6t
Xbit_r220_c101 bl[101] br[101] wl[220] vdd gnd cell_6t
Xbit_r221_c101 bl[101] br[101] wl[221] vdd gnd cell_6t
Xbit_r222_c101 bl[101] br[101] wl[222] vdd gnd cell_6t
Xbit_r223_c101 bl[101] br[101] wl[223] vdd gnd cell_6t
Xbit_r224_c101 bl[101] br[101] wl[224] vdd gnd cell_6t
Xbit_r225_c101 bl[101] br[101] wl[225] vdd gnd cell_6t
Xbit_r226_c101 bl[101] br[101] wl[226] vdd gnd cell_6t
Xbit_r227_c101 bl[101] br[101] wl[227] vdd gnd cell_6t
Xbit_r228_c101 bl[101] br[101] wl[228] vdd gnd cell_6t
Xbit_r229_c101 bl[101] br[101] wl[229] vdd gnd cell_6t
Xbit_r230_c101 bl[101] br[101] wl[230] vdd gnd cell_6t
Xbit_r231_c101 bl[101] br[101] wl[231] vdd gnd cell_6t
Xbit_r232_c101 bl[101] br[101] wl[232] vdd gnd cell_6t
Xbit_r233_c101 bl[101] br[101] wl[233] vdd gnd cell_6t
Xbit_r234_c101 bl[101] br[101] wl[234] vdd gnd cell_6t
Xbit_r235_c101 bl[101] br[101] wl[235] vdd gnd cell_6t
Xbit_r236_c101 bl[101] br[101] wl[236] vdd gnd cell_6t
Xbit_r237_c101 bl[101] br[101] wl[237] vdd gnd cell_6t
Xbit_r238_c101 bl[101] br[101] wl[238] vdd gnd cell_6t
Xbit_r239_c101 bl[101] br[101] wl[239] vdd gnd cell_6t
Xbit_r240_c101 bl[101] br[101] wl[240] vdd gnd cell_6t
Xbit_r241_c101 bl[101] br[101] wl[241] vdd gnd cell_6t
Xbit_r242_c101 bl[101] br[101] wl[242] vdd gnd cell_6t
Xbit_r243_c101 bl[101] br[101] wl[243] vdd gnd cell_6t
Xbit_r244_c101 bl[101] br[101] wl[244] vdd gnd cell_6t
Xbit_r245_c101 bl[101] br[101] wl[245] vdd gnd cell_6t
Xbit_r246_c101 bl[101] br[101] wl[246] vdd gnd cell_6t
Xbit_r247_c101 bl[101] br[101] wl[247] vdd gnd cell_6t
Xbit_r248_c101 bl[101] br[101] wl[248] vdd gnd cell_6t
Xbit_r249_c101 bl[101] br[101] wl[249] vdd gnd cell_6t
Xbit_r250_c101 bl[101] br[101] wl[250] vdd gnd cell_6t
Xbit_r251_c101 bl[101] br[101] wl[251] vdd gnd cell_6t
Xbit_r252_c101 bl[101] br[101] wl[252] vdd gnd cell_6t
Xbit_r253_c101 bl[101] br[101] wl[253] vdd gnd cell_6t
Xbit_r254_c101 bl[101] br[101] wl[254] vdd gnd cell_6t
Xbit_r255_c101 bl[101] br[101] wl[255] vdd gnd cell_6t
Xbit_r0_c102 bl[102] br[102] wl[0] vdd gnd cell_6t
Xbit_r1_c102 bl[102] br[102] wl[1] vdd gnd cell_6t
Xbit_r2_c102 bl[102] br[102] wl[2] vdd gnd cell_6t
Xbit_r3_c102 bl[102] br[102] wl[3] vdd gnd cell_6t
Xbit_r4_c102 bl[102] br[102] wl[4] vdd gnd cell_6t
Xbit_r5_c102 bl[102] br[102] wl[5] vdd gnd cell_6t
Xbit_r6_c102 bl[102] br[102] wl[6] vdd gnd cell_6t
Xbit_r7_c102 bl[102] br[102] wl[7] vdd gnd cell_6t
Xbit_r8_c102 bl[102] br[102] wl[8] vdd gnd cell_6t
Xbit_r9_c102 bl[102] br[102] wl[9] vdd gnd cell_6t
Xbit_r10_c102 bl[102] br[102] wl[10] vdd gnd cell_6t
Xbit_r11_c102 bl[102] br[102] wl[11] vdd gnd cell_6t
Xbit_r12_c102 bl[102] br[102] wl[12] vdd gnd cell_6t
Xbit_r13_c102 bl[102] br[102] wl[13] vdd gnd cell_6t
Xbit_r14_c102 bl[102] br[102] wl[14] vdd gnd cell_6t
Xbit_r15_c102 bl[102] br[102] wl[15] vdd gnd cell_6t
Xbit_r16_c102 bl[102] br[102] wl[16] vdd gnd cell_6t
Xbit_r17_c102 bl[102] br[102] wl[17] vdd gnd cell_6t
Xbit_r18_c102 bl[102] br[102] wl[18] vdd gnd cell_6t
Xbit_r19_c102 bl[102] br[102] wl[19] vdd gnd cell_6t
Xbit_r20_c102 bl[102] br[102] wl[20] vdd gnd cell_6t
Xbit_r21_c102 bl[102] br[102] wl[21] vdd gnd cell_6t
Xbit_r22_c102 bl[102] br[102] wl[22] vdd gnd cell_6t
Xbit_r23_c102 bl[102] br[102] wl[23] vdd gnd cell_6t
Xbit_r24_c102 bl[102] br[102] wl[24] vdd gnd cell_6t
Xbit_r25_c102 bl[102] br[102] wl[25] vdd gnd cell_6t
Xbit_r26_c102 bl[102] br[102] wl[26] vdd gnd cell_6t
Xbit_r27_c102 bl[102] br[102] wl[27] vdd gnd cell_6t
Xbit_r28_c102 bl[102] br[102] wl[28] vdd gnd cell_6t
Xbit_r29_c102 bl[102] br[102] wl[29] vdd gnd cell_6t
Xbit_r30_c102 bl[102] br[102] wl[30] vdd gnd cell_6t
Xbit_r31_c102 bl[102] br[102] wl[31] vdd gnd cell_6t
Xbit_r32_c102 bl[102] br[102] wl[32] vdd gnd cell_6t
Xbit_r33_c102 bl[102] br[102] wl[33] vdd gnd cell_6t
Xbit_r34_c102 bl[102] br[102] wl[34] vdd gnd cell_6t
Xbit_r35_c102 bl[102] br[102] wl[35] vdd gnd cell_6t
Xbit_r36_c102 bl[102] br[102] wl[36] vdd gnd cell_6t
Xbit_r37_c102 bl[102] br[102] wl[37] vdd gnd cell_6t
Xbit_r38_c102 bl[102] br[102] wl[38] vdd gnd cell_6t
Xbit_r39_c102 bl[102] br[102] wl[39] vdd gnd cell_6t
Xbit_r40_c102 bl[102] br[102] wl[40] vdd gnd cell_6t
Xbit_r41_c102 bl[102] br[102] wl[41] vdd gnd cell_6t
Xbit_r42_c102 bl[102] br[102] wl[42] vdd gnd cell_6t
Xbit_r43_c102 bl[102] br[102] wl[43] vdd gnd cell_6t
Xbit_r44_c102 bl[102] br[102] wl[44] vdd gnd cell_6t
Xbit_r45_c102 bl[102] br[102] wl[45] vdd gnd cell_6t
Xbit_r46_c102 bl[102] br[102] wl[46] vdd gnd cell_6t
Xbit_r47_c102 bl[102] br[102] wl[47] vdd gnd cell_6t
Xbit_r48_c102 bl[102] br[102] wl[48] vdd gnd cell_6t
Xbit_r49_c102 bl[102] br[102] wl[49] vdd gnd cell_6t
Xbit_r50_c102 bl[102] br[102] wl[50] vdd gnd cell_6t
Xbit_r51_c102 bl[102] br[102] wl[51] vdd gnd cell_6t
Xbit_r52_c102 bl[102] br[102] wl[52] vdd gnd cell_6t
Xbit_r53_c102 bl[102] br[102] wl[53] vdd gnd cell_6t
Xbit_r54_c102 bl[102] br[102] wl[54] vdd gnd cell_6t
Xbit_r55_c102 bl[102] br[102] wl[55] vdd gnd cell_6t
Xbit_r56_c102 bl[102] br[102] wl[56] vdd gnd cell_6t
Xbit_r57_c102 bl[102] br[102] wl[57] vdd gnd cell_6t
Xbit_r58_c102 bl[102] br[102] wl[58] vdd gnd cell_6t
Xbit_r59_c102 bl[102] br[102] wl[59] vdd gnd cell_6t
Xbit_r60_c102 bl[102] br[102] wl[60] vdd gnd cell_6t
Xbit_r61_c102 bl[102] br[102] wl[61] vdd gnd cell_6t
Xbit_r62_c102 bl[102] br[102] wl[62] vdd gnd cell_6t
Xbit_r63_c102 bl[102] br[102] wl[63] vdd gnd cell_6t
Xbit_r64_c102 bl[102] br[102] wl[64] vdd gnd cell_6t
Xbit_r65_c102 bl[102] br[102] wl[65] vdd gnd cell_6t
Xbit_r66_c102 bl[102] br[102] wl[66] vdd gnd cell_6t
Xbit_r67_c102 bl[102] br[102] wl[67] vdd gnd cell_6t
Xbit_r68_c102 bl[102] br[102] wl[68] vdd gnd cell_6t
Xbit_r69_c102 bl[102] br[102] wl[69] vdd gnd cell_6t
Xbit_r70_c102 bl[102] br[102] wl[70] vdd gnd cell_6t
Xbit_r71_c102 bl[102] br[102] wl[71] vdd gnd cell_6t
Xbit_r72_c102 bl[102] br[102] wl[72] vdd gnd cell_6t
Xbit_r73_c102 bl[102] br[102] wl[73] vdd gnd cell_6t
Xbit_r74_c102 bl[102] br[102] wl[74] vdd gnd cell_6t
Xbit_r75_c102 bl[102] br[102] wl[75] vdd gnd cell_6t
Xbit_r76_c102 bl[102] br[102] wl[76] vdd gnd cell_6t
Xbit_r77_c102 bl[102] br[102] wl[77] vdd gnd cell_6t
Xbit_r78_c102 bl[102] br[102] wl[78] vdd gnd cell_6t
Xbit_r79_c102 bl[102] br[102] wl[79] vdd gnd cell_6t
Xbit_r80_c102 bl[102] br[102] wl[80] vdd gnd cell_6t
Xbit_r81_c102 bl[102] br[102] wl[81] vdd gnd cell_6t
Xbit_r82_c102 bl[102] br[102] wl[82] vdd gnd cell_6t
Xbit_r83_c102 bl[102] br[102] wl[83] vdd gnd cell_6t
Xbit_r84_c102 bl[102] br[102] wl[84] vdd gnd cell_6t
Xbit_r85_c102 bl[102] br[102] wl[85] vdd gnd cell_6t
Xbit_r86_c102 bl[102] br[102] wl[86] vdd gnd cell_6t
Xbit_r87_c102 bl[102] br[102] wl[87] vdd gnd cell_6t
Xbit_r88_c102 bl[102] br[102] wl[88] vdd gnd cell_6t
Xbit_r89_c102 bl[102] br[102] wl[89] vdd gnd cell_6t
Xbit_r90_c102 bl[102] br[102] wl[90] vdd gnd cell_6t
Xbit_r91_c102 bl[102] br[102] wl[91] vdd gnd cell_6t
Xbit_r92_c102 bl[102] br[102] wl[92] vdd gnd cell_6t
Xbit_r93_c102 bl[102] br[102] wl[93] vdd gnd cell_6t
Xbit_r94_c102 bl[102] br[102] wl[94] vdd gnd cell_6t
Xbit_r95_c102 bl[102] br[102] wl[95] vdd gnd cell_6t
Xbit_r96_c102 bl[102] br[102] wl[96] vdd gnd cell_6t
Xbit_r97_c102 bl[102] br[102] wl[97] vdd gnd cell_6t
Xbit_r98_c102 bl[102] br[102] wl[98] vdd gnd cell_6t
Xbit_r99_c102 bl[102] br[102] wl[99] vdd gnd cell_6t
Xbit_r100_c102 bl[102] br[102] wl[100] vdd gnd cell_6t
Xbit_r101_c102 bl[102] br[102] wl[101] vdd gnd cell_6t
Xbit_r102_c102 bl[102] br[102] wl[102] vdd gnd cell_6t
Xbit_r103_c102 bl[102] br[102] wl[103] vdd gnd cell_6t
Xbit_r104_c102 bl[102] br[102] wl[104] vdd gnd cell_6t
Xbit_r105_c102 bl[102] br[102] wl[105] vdd gnd cell_6t
Xbit_r106_c102 bl[102] br[102] wl[106] vdd gnd cell_6t
Xbit_r107_c102 bl[102] br[102] wl[107] vdd gnd cell_6t
Xbit_r108_c102 bl[102] br[102] wl[108] vdd gnd cell_6t
Xbit_r109_c102 bl[102] br[102] wl[109] vdd gnd cell_6t
Xbit_r110_c102 bl[102] br[102] wl[110] vdd gnd cell_6t
Xbit_r111_c102 bl[102] br[102] wl[111] vdd gnd cell_6t
Xbit_r112_c102 bl[102] br[102] wl[112] vdd gnd cell_6t
Xbit_r113_c102 bl[102] br[102] wl[113] vdd gnd cell_6t
Xbit_r114_c102 bl[102] br[102] wl[114] vdd gnd cell_6t
Xbit_r115_c102 bl[102] br[102] wl[115] vdd gnd cell_6t
Xbit_r116_c102 bl[102] br[102] wl[116] vdd gnd cell_6t
Xbit_r117_c102 bl[102] br[102] wl[117] vdd gnd cell_6t
Xbit_r118_c102 bl[102] br[102] wl[118] vdd gnd cell_6t
Xbit_r119_c102 bl[102] br[102] wl[119] vdd gnd cell_6t
Xbit_r120_c102 bl[102] br[102] wl[120] vdd gnd cell_6t
Xbit_r121_c102 bl[102] br[102] wl[121] vdd gnd cell_6t
Xbit_r122_c102 bl[102] br[102] wl[122] vdd gnd cell_6t
Xbit_r123_c102 bl[102] br[102] wl[123] vdd gnd cell_6t
Xbit_r124_c102 bl[102] br[102] wl[124] vdd gnd cell_6t
Xbit_r125_c102 bl[102] br[102] wl[125] vdd gnd cell_6t
Xbit_r126_c102 bl[102] br[102] wl[126] vdd gnd cell_6t
Xbit_r127_c102 bl[102] br[102] wl[127] vdd gnd cell_6t
Xbit_r128_c102 bl[102] br[102] wl[128] vdd gnd cell_6t
Xbit_r129_c102 bl[102] br[102] wl[129] vdd gnd cell_6t
Xbit_r130_c102 bl[102] br[102] wl[130] vdd gnd cell_6t
Xbit_r131_c102 bl[102] br[102] wl[131] vdd gnd cell_6t
Xbit_r132_c102 bl[102] br[102] wl[132] vdd gnd cell_6t
Xbit_r133_c102 bl[102] br[102] wl[133] vdd gnd cell_6t
Xbit_r134_c102 bl[102] br[102] wl[134] vdd gnd cell_6t
Xbit_r135_c102 bl[102] br[102] wl[135] vdd gnd cell_6t
Xbit_r136_c102 bl[102] br[102] wl[136] vdd gnd cell_6t
Xbit_r137_c102 bl[102] br[102] wl[137] vdd gnd cell_6t
Xbit_r138_c102 bl[102] br[102] wl[138] vdd gnd cell_6t
Xbit_r139_c102 bl[102] br[102] wl[139] vdd gnd cell_6t
Xbit_r140_c102 bl[102] br[102] wl[140] vdd gnd cell_6t
Xbit_r141_c102 bl[102] br[102] wl[141] vdd gnd cell_6t
Xbit_r142_c102 bl[102] br[102] wl[142] vdd gnd cell_6t
Xbit_r143_c102 bl[102] br[102] wl[143] vdd gnd cell_6t
Xbit_r144_c102 bl[102] br[102] wl[144] vdd gnd cell_6t
Xbit_r145_c102 bl[102] br[102] wl[145] vdd gnd cell_6t
Xbit_r146_c102 bl[102] br[102] wl[146] vdd gnd cell_6t
Xbit_r147_c102 bl[102] br[102] wl[147] vdd gnd cell_6t
Xbit_r148_c102 bl[102] br[102] wl[148] vdd gnd cell_6t
Xbit_r149_c102 bl[102] br[102] wl[149] vdd gnd cell_6t
Xbit_r150_c102 bl[102] br[102] wl[150] vdd gnd cell_6t
Xbit_r151_c102 bl[102] br[102] wl[151] vdd gnd cell_6t
Xbit_r152_c102 bl[102] br[102] wl[152] vdd gnd cell_6t
Xbit_r153_c102 bl[102] br[102] wl[153] vdd gnd cell_6t
Xbit_r154_c102 bl[102] br[102] wl[154] vdd gnd cell_6t
Xbit_r155_c102 bl[102] br[102] wl[155] vdd gnd cell_6t
Xbit_r156_c102 bl[102] br[102] wl[156] vdd gnd cell_6t
Xbit_r157_c102 bl[102] br[102] wl[157] vdd gnd cell_6t
Xbit_r158_c102 bl[102] br[102] wl[158] vdd gnd cell_6t
Xbit_r159_c102 bl[102] br[102] wl[159] vdd gnd cell_6t
Xbit_r160_c102 bl[102] br[102] wl[160] vdd gnd cell_6t
Xbit_r161_c102 bl[102] br[102] wl[161] vdd gnd cell_6t
Xbit_r162_c102 bl[102] br[102] wl[162] vdd gnd cell_6t
Xbit_r163_c102 bl[102] br[102] wl[163] vdd gnd cell_6t
Xbit_r164_c102 bl[102] br[102] wl[164] vdd gnd cell_6t
Xbit_r165_c102 bl[102] br[102] wl[165] vdd gnd cell_6t
Xbit_r166_c102 bl[102] br[102] wl[166] vdd gnd cell_6t
Xbit_r167_c102 bl[102] br[102] wl[167] vdd gnd cell_6t
Xbit_r168_c102 bl[102] br[102] wl[168] vdd gnd cell_6t
Xbit_r169_c102 bl[102] br[102] wl[169] vdd gnd cell_6t
Xbit_r170_c102 bl[102] br[102] wl[170] vdd gnd cell_6t
Xbit_r171_c102 bl[102] br[102] wl[171] vdd gnd cell_6t
Xbit_r172_c102 bl[102] br[102] wl[172] vdd gnd cell_6t
Xbit_r173_c102 bl[102] br[102] wl[173] vdd gnd cell_6t
Xbit_r174_c102 bl[102] br[102] wl[174] vdd gnd cell_6t
Xbit_r175_c102 bl[102] br[102] wl[175] vdd gnd cell_6t
Xbit_r176_c102 bl[102] br[102] wl[176] vdd gnd cell_6t
Xbit_r177_c102 bl[102] br[102] wl[177] vdd gnd cell_6t
Xbit_r178_c102 bl[102] br[102] wl[178] vdd gnd cell_6t
Xbit_r179_c102 bl[102] br[102] wl[179] vdd gnd cell_6t
Xbit_r180_c102 bl[102] br[102] wl[180] vdd gnd cell_6t
Xbit_r181_c102 bl[102] br[102] wl[181] vdd gnd cell_6t
Xbit_r182_c102 bl[102] br[102] wl[182] vdd gnd cell_6t
Xbit_r183_c102 bl[102] br[102] wl[183] vdd gnd cell_6t
Xbit_r184_c102 bl[102] br[102] wl[184] vdd gnd cell_6t
Xbit_r185_c102 bl[102] br[102] wl[185] vdd gnd cell_6t
Xbit_r186_c102 bl[102] br[102] wl[186] vdd gnd cell_6t
Xbit_r187_c102 bl[102] br[102] wl[187] vdd gnd cell_6t
Xbit_r188_c102 bl[102] br[102] wl[188] vdd gnd cell_6t
Xbit_r189_c102 bl[102] br[102] wl[189] vdd gnd cell_6t
Xbit_r190_c102 bl[102] br[102] wl[190] vdd gnd cell_6t
Xbit_r191_c102 bl[102] br[102] wl[191] vdd gnd cell_6t
Xbit_r192_c102 bl[102] br[102] wl[192] vdd gnd cell_6t
Xbit_r193_c102 bl[102] br[102] wl[193] vdd gnd cell_6t
Xbit_r194_c102 bl[102] br[102] wl[194] vdd gnd cell_6t
Xbit_r195_c102 bl[102] br[102] wl[195] vdd gnd cell_6t
Xbit_r196_c102 bl[102] br[102] wl[196] vdd gnd cell_6t
Xbit_r197_c102 bl[102] br[102] wl[197] vdd gnd cell_6t
Xbit_r198_c102 bl[102] br[102] wl[198] vdd gnd cell_6t
Xbit_r199_c102 bl[102] br[102] wl[199] vdd gnd cell_6t
Xbit_r200_c102 bl[102] br[102] wl[200] vdd gnd cell_6t
Xbit_r201_c102 bl[102] br[102] wl[201] vdd gnd cell_6t
Xbit_r202_c102 bl[102] br[102] wl[202] vdd gnd cell_6t
Xbit_r203_c102 bl[102] br[102] wl[203] vdd gnd cell_6t
Xbit_r204_c102 bl[102] br[102] wl[204] vdd gnd cell_6t
Xbit_r205_c102 bl[102] br[102] wl[205] vdd gnd cell_6t
Xbit_r206_c102 bl[102] br[102] wl[206] vdd gnd cell_6t
Xbit_r207_c102 bl[102] br[102] wl[207] vdd gnd cell_6t
Xbit_r208_c102 bl[102] br[102] wl[208] vdd gnd cell_6t
Xbit_r209_c102 bl[102] br[102] wl[209] vdd gnd cell_6t
Xbit_r210_c102 bl[102] br[102] wl[210] vdd gnd cell_6t
Xbit_r211_c102 bl[102] br[102] wl[211] vdd gnd cell_6t
Xbit_r212_c102 bl[102] br[102] wl[212] vdd gnd cell_6t
Xbit_r213_c102 bl[102] br[102] wl[213] vdd gnd cell_6t
Xbit_r214_c102 bl[102] br[102] wl[214] vdd gnd cell_6t
Xbit_r215_c102 bl[102] br[102] wl[215] vdd gnd cell_6t
Xbit_r216_c102 bl[102] br[102] wl[216] vdd gnd cell_6t
Xbit_r217_c102 bl[102] br[102] wl[217] vdd gnd cell_6t
Xbit_r218_c102 bl[102] br[102] wl[218] vdd gnd cell_6t
Xbit_r219_c102 bl[102] br[102] wl[219] vdd gnd cell_6t
Xbit_r220_c102 bl[102] br[102] wl[220] vdd gnd cell_6t
Xbit_r221_c102 bl[102] br[102] wl[221] vdd gnd cell_6t
Xbit_r222_c102 bl[102] br[102] wl[222] vdd gnd cell_6t
Xbit_r223_c102 bl[102] br[102] wl[223] vdd gnd cell_6t
Xbit_r224_c102 bl[102] br[102] wl[224] vdd gnd cell_6t
Xbit_r225_c102 bl[102] br[102] wl[225] vdd gnd cell_6t
Xbit_r226_c102 bl[102] br[102] wl[226] vdd gnd cell_6t
Xbit_r227_c102 bl[102] br[102] wl[227] vdd gnd cell_6t
Xbit_r228_c102 bl[102] br[102] wl[228] vdd gnd cell_6t
Xbit_r229_c102 bl[102] br[102] wl[229] vdd gnd cell_6t
Xbit_r230_c102 bl[102] br[102] wl[230] vdd gnd cell_6t
Xbit_r231_c102 bl[102] br[102] wl[231] vdd gnd cell_6t
Xbit_r232_c102 bl[102] br[102] wl[232] vdd gnd cell_6t
Xbit_r233_c102 bl[102] br[102] wl[233] vdd gnd cell_6t
Xbit_r234_c102 bl[102] br[102] wl[234] vdd gnd cell_6t
Xbit_r235_c102 bl[102] br[102] wl[235] vdd gnd cell_6t
Xbit_r236_c102 bl[102] br[102] wl[236] vdd gnd cell_6t
Xbit_r237_c102 bl[102] br[102] wl[237] vdd gnd cell_6t
Xbit_r238_c102 bl[102] br[102] wl[238] vdd gnd cell_6t
Xbit_r239_c102 bl[102] br[102] wl[239] vdd gnd cell_6t
Xbit_r240_c102 bl[102] br[102] wl[240] vdd gnd cell_6t
Xbit_r241_c102 bl[102] br[102] wl[241] vdd gnd cell_6t
Xbit_r242_c102 bl[102] br[102] wl[242] vdd gnd cell_6t
Xbit_r243_c102 bl[102] br[102] wl[243] vdd gnd cell_6t
Xbit_r244_c102 bl[102] br[102] wl[244] vdd gnd cell_6t
Xbit_r245_c102 bl[102] br[102] wl[245] vdd gnd cell_6t
Xbit_r246_c102 bl[102] br[102] wl[246] vdd gnd cell_6t
Xbit_r247_c102 bl[102] br[102] wl[247] vdd gnd cell_6t
Xbit_r248_c102 bl[102] br[102] wl[248] vdd gnd cell_6t
Xbit_r249_c102 bl[102] br[102] wl[249] vdd gnd cell_6t
Xbit_r250_c102 bl[102] br[102] wl[250] vdd gnd cell_6t
Xbit_r251_c102 bl[102] br[102] wl[251] vdd gnd cell_6t
Xbit_r252_c102 bl[102] br[102] wl[252] vdd gnd cell_6t
Xbit_r253_c102 bl[102] br[102] wl[253] vdd gnd cell_6t
Xbit_r254_c102 bl[102] br[102] wl[254] vdd gnd cell_6t
Xbit_r255_c102 bl[102] br[102] wl[255] vdd gnd cell_6t
Xbit_r0_c103 bl[103] br[103] wl[0] vdd gnd cell_6t
Xbit_r1_c103 bl[103] br[103] wl[1] vdd gnd cell_6t
Xbit_r2_c103 bl[103] br[103] wl[2] vdd gnd cell_6t
Xbit_r3_c103 bl[103] br[103] wl[3] vdd gnd cell_6t
Xbit_r4_c103 bl[103] br[103] wl[4] vdd gnd cell_6t
Xbit_r5_c103 bl[103] br[103] wl[5] vdd gnd cell_6t
Xbit_r6_c103 bl[103] br[103] wl[6] vdd gnd cell_6t
Xbit_r7_c103 bl[103] br[103] wl[7] vdd gnd cell_6t
Xbit_r8_c103 bl[103] br[103] wl[8] vdd gnd cell_6t
Xbit_r9_c103 bl[103] br[103] wl[9] vdd gnd cell_6t
Xbit_r10_c103 bl[103] br[103] wl[10] vdd gnd cell_6t
Xbit_r11_c103 bl[103] br[103] wl[11] vdd gnd cell_6t
Xbit_r12_c103 bl[103] br[103] wl[12] vdd gnd cell_6t
Xbit_r13_c103 bl[103] br[103] wl[13] vdd gnd cell_6t
Xbit_r14_c103 bl[103] br[103] wl[14] vdd gnd cell_6t
Xbit_r15_c103 bl[103] br[103] wl[15] vdd gnd cell_6t
Xbit_r16_c103 bl[103] br[103] wl[16] vdd gnd cell_6t
Xbit_r17_c103 bl[103] br[103] wl[17] vdd gnd cell_6t
Xbit_r18_c103 bl[103] br[103] wl[18] vdd gnd cell_6t
Xbit_r19_c103 bl[103] br[103] wl[19] vdd gnd cell_6t
Xbit_r20_c103 bl[103] br[103] wl[20] vdd gnd cell_6t
Xbit_r21_c103 bl[103] br[103] wl[21] vdd gnd cell_6t
Xbit_r22_c103 bl[103] br[103] wl[22] vdd gnd cell_6t
Xbit_r23_c103 bl[103] br[103] wl[23] vdd gnd cell_6t
Xbit_r24_c103 bl[103] br[103] wl[24] vdd gnd cell_6t
Xbit_r25_c103 bl[103] br[103] wl[25] vdd gnd cell_6t
Xbit_r26_c103 bl[103] br[103] wl[26] vdd gnd cell_6t
Xbit_r27_c103 bl[103] br[103] wl[27] vdd gnd cell_6t
Xbit_r28_c103 bl[103] br[103] wl[28] vdd gnd cell_6t
Xbit_r29_c103 bl[103] br[103] wl[29] vdd gnd cell_6t
Xbit_r30_c103 bl[103] br[103] wl[30] vdd gnd cell_6t
Xbit_r31_c103 bl[103] br[103] wl[31] vdd gnd cell_6t
Xbit_r32_c103 bl[103] br[103] wl[32] vdd gnd cell_6t
Xbit_r33_c103 bl[103] br[103] wl[33] vdd gnd cell_6t
Xbit_r34_c103 bl[103] br[103] wl[34] vdd gnd cell_6t
Xbit_r35_c103 bl[103] br[103] wl[35] vdd gnd cell_6t
Xbit_r36_c103 bl[103] br[103] wl[36] vdd gnd cell_6t
Xbit_r37_c103 bl[103] br[103] wl[37] vdd gnd cell_6t
Xbit_r38_c103 bl[103] br[103] wl[38] vdd gnd cell_6t
Xbit_r39_c103 bl[103] br[103] wl[39] vdd gnd cell_6t
Xbit_r40_c103 bl[103] br[103] wl[40] vdd gnd cell_6t
Xbit_r41_c103 bl[103] br[103] wl[41] vdd gnd cell_6t
Xbit_r42_c103 bl[103] br[103] wl[42] vdd gnd cell_6t
Xbit_r43_c103 bl[103] br[103] wl[43] vdd gnd cell_6t
Xbit_r44_c103 bl[103] br[103] wl[44] vdd gnd cell_6t
Xbit_r45_c103 bl[103] br[103] wl[45] vdd gnd cell_6t
Xbit_r46_c103 bl[103] br[103] wl[46] vdd gnd cell_6t
Xbit_r47_c103 bl[103] br[103] wl[47] vdd gnd cell_6t
Xbit_r48_c103 bl[103] br[103] wl[48] vdd gnd cell_6t
Xbit_r49_c103 bl[103] br[103] wl[49] vdd gnd cell_6t
Xbit_r50_c103 bl[103] br[103] wl[50] vdd gnd cell_6t
Xbit_r51_c103 bl[103] br[103] wl[51] vdd gnd cell_6t
Xbit_r52_c103 bl[103] br[103] wl[52] vdd gnd cell_6t
Xbit_r53_c103 bl[103] br[103] wl[53] vdd gnd cell_6t
Xbit_r54_c103 bl[103] br[103] wl[54] vdd gnd cell_6t
Xbit_r55_c103 bl[103] br[103] wl[55] vdd gnd cell_6t
Xbit_r56_c103 bl[103] br[103] wl[56] vdd gnd cell_6t
Xbit_r57_c103 bl[103] br[103] wl[57] vdd gnd cell_6t
Xbit_r58_c103 bl[103] br[103] wl[58] vdd gnd cell_6t
Xbit_r59_c103 bl[103] br[103] wl[59] vdd gnd cell_6t
Xbit_r60_c103 bl[103] br[103] wl[60] vdd gnd cell_6t
Xbit_r61_c103 bl[103] br[103] wl[61] vdd gnd cell_6t
Xbit_r62_c103 bl[103] br[103] wl[62] vdd gnd cell_6t
Xbit_r63_c103 bl[103] br[103] wl[63] vdd gnd cell_6t
Xbit_r64_c103 bl[103] br[103] wl[64] vdd gnd cell_6t
Xbit_r65_c103 bl[103] br[103] wl[65] vdd gnd cell_6t
Xbit_r66_c103 bl[103] br[103] wl[66] vdd gnd cell_6t
Xbit_r67_c103 bl[103] br[103] wl[67] vdd gnd cell_6t
Xbit_r68_c103 bl[103] br[103] wl[68] vdd gnd cell_6t
Xbit_r69_c103 bl[103] br[103] wl[69] vdd gnd cell_6t
Xbit_r70_c103 bl[103] br[103] wl[70] vdd gnd cell_6t
Xbit_r71_c103 bl[103] br[103] wl[71] vdd gnd cell_6t
Xbit_r72_c103 bl[103] br[103] wl[72] vdd gnd cell_6t
Xbit_r73_c103 bl[103] br[103] wl[73] vdd gnd cell_6t
Xbit_r74_c103 bl[103] br[103] wl[74] vdd gnd cell_6t
Xbit_r75_c103 bl[103] br[103] wl[75] vdd gnd cell_6t
Xbit_r76_c103 bl[103] br[103] wl[76] vdd gnd cell_6t
Xbit_r77_c103 bl[103] br[103] wl[77] vdd gnd cell_6t
Xbit_r78_c103 bl[103] br[103] wl[78] vdd gnd cell_6t
Xbit_r79_c103 bl[103] br[103] wl[79] vdd gnd cell_6t
Xbit_r80_c103 bl[103] br[103] wl[80] vdd gnd cell_6t
Xbit_r81_c103 bl[103] br[103] wl[81] vdd gnd cell_6t
Xbit_r82_c103 bl[103] br[103] wl[82] vdd gnd cell_6t
Xbit_r83_c103 bl[103] br[103] wl[83] vdd gnd cell_6t
Xbit_r84_c103 bl[103] br[103] wl[84] vdd gnd cell_6t
Xbit_r85_c103 bl[103] br[103] wl[85] vdd gnd cell_6t
Xbit_r86_c103 bl[103] br[103] wl[86] vdd gnd cell_6t
Xbit_r87_c103 bl[103] br[103] wl[87] vdd gnd cell_6t
Xbit_r88_c103 bl[103] br[103] wl[88] vdd gnd cell_6t
Xbit_r89_c103 bl[103] br[103] wl[89] vdd gnd cell_6t
Xbit_r90_c103 bl[103] br[103] wl[90] vdd gnd cell_6t
Xbit_r91_c103 bl[103] br[103] wl[91] vdd gnd cell_6t
Xbit_r92_c103 bl[103] br[103] wl[92] vdd gnd cell_6t
Xbit_r93_c103 bl[103] br[103] wl[93] vdd gnd cell_6t
Xbit_r94_c103 bl[103] br[103] wl[94] vdd gnd cell_6t
Xbit_r95_c103 bl[103] br[103] wl[95] vdd gnd cell_6t
Xbit_r96_c103 bl[103] br[103] wl[96] vdd gnd cell_6t
Xbit_r97_c103 bl[103] br[103] wl[97] vdd gnd cell_6t
Xbit_r98_c103 bl[103] br[103] wl[98] vdd gnd cell_6t
Xbit_r99_c103 bl[103] br[103] wl[99] vdd gnd cell_6t
Xbit_r100_c103 bl[103] br[103] wl[100] vdd gnd cell_6t
Xbit_r101_c103 bl[103] br[103] wl[101] vdd gnd cell_6t
Xbit_r102_c103 bl[103] br[103] wl[102] vdd gnd cell_6t
Xbit_r103_c103 bl[103] br[103] wl[103] vdd gnd cell_6t
Xbit_r104_c103 bl[103] br[103] wl[104] vdd gnd cell_6t
Xbit_r105_c103 bl[103] br[103] wl[105] vdd gnd cell_6t
Xbit_r106_c103 bl[103] br[103] wl[106] vdd gnd cell_6t
Xbit_r107_c103 bl[103] br[103] wl[107] vdd gnd cell_6t
Xbit_r108_c103 bl[103] br[103] wl[108] vdd gnd cell_6t
Xbit_r109_c103 bl[103] br[103] wl[109] vdd gnd cell_6t
Xbit_r110_c103 bl[103] br[103] wl[110] vdd gnd cell_6t
Xbit_r111_c103 bl[103] br[103] wl[111] vdd gnd cell_6t
Xbit_r112_c103 bl[103] br[103] wl[112] vdd gnd cell_6t
Xbit_r113_c103 bl[103] br[103] wl[113] vdd gnd cell_6t
Xbit_r114_c103 bl[103] br[103] wl[114] vdd gnd cell_6t
Xbit_r115_c103 bl[103] br[103] wl[115] vdd gnd cell_6t
Xbit_r116_c103 bl[103] br[103] wl[116] vdd gnd cell_6t
Xbit_r117_c103 bl[103] br[103] wl[117] vdd gnd cell_6t
Xbit_r118_c103 bl[103] br[103] wl[118] vdd gnd cell_6t
Xbit_r119_c103 bl[103] br[103] wl[119] vdd gnd cell_6t
Xbit_r120_c103 bl[103] br[103] wl[120] vdd gnd cell_6t
Xbit_r121_c103 bl[103] br[103] wl[121] vdd gnd cell_6t
Xbit_r122_c103 bl[103] br[103] wl[122] vdd gnd cell_6t
Xbit_r123_c103 bl[103] br[103] wl[123] vdd gnd cell_6t
Xbit_r124_c103 bl[103] br[103] wl[124] vdd gnd cell_6t
Xbit_r125_c103 bl[103] br[103] wl[125] vdd gnd cell_6t
Xbit_r126_c103 bl[103] br[103] wl[126] vdd gnd cell_6t
Xbit_r127_c103 bl[103] br[103] wl[127] vdd gnd cell_6t
Xbit_r128_c103 bl[103] br[103] wl[128] vdd gnd cell_6t
Xbit_r129_c103 bl[103] br[103] wl[129] vdd gnd cell_6t
Xbit_r130_c103 bl[103] br[103] wl[130] vdd gnd cell_6t
Xbit_r131_c103 bl[103] br[103] wl[131] vdd gnd cell_6t
Xbit_r132_c103 bl[103] br[103] wl[132] vdd gnd cell_6t
Xbit_r133_c103 bl[103] br[103] wl[133] vdd gnd cell_6t
Xbit_r134_c103 bl[103] br[103] wl[134] vdd gnd cell_6t
Xbit_r135_c103 bl[103] br[103] wl[135] vdd gnd cell_6t
Xbit_r136_c103 bl[103] br[103] wl[136] vdd gnd cell_6t
Xbit_r137_c103 bl[103] br[103] wl[137] vdd gnd cell_6t
Xbit_r138_c103 bl[103] br[103] wl[138] vdd gnd cell_6t
Xbit_r139_c103 bl[103] br[103] wl[139] vdd gnd cell_6t
Xbit_r140_c103 bl[103] br[103] wl[140] vdd gnd cell_6t
Xbit_r141_c103 bl[103] br[103] wl[141] vdd gnd cell_6t
Xbit_r142_c103 bl[103] br[103] wl[142] vdd gnd cell_6t
Xbit_r143_c103 bl[103] br[103] wl[143] vdd gnd cell_6t
Xbit_r144_c103 bl[103] br[103] wl[144] vdd gnd cell_6t
Xbit_r145_c103 bl[103] br[103] wl[145] vdd gnd cell_6t
Xbit_r146_c103 bl[103] br[103] wl[146] vdd gnd cell_6t
Xbit_r147_c103 bl[103] br[103] wl[147] vdd gnd cell_6t
Xbit_r148_c103 bl[103] br[103] wl[148] vdd gnd cell_6t
Xbit_r149_c103 bl[103] br[103] wl[149] vdd gnd cell_6t
Xbit_r150_c103 bl[103] br[103] wl[150] vdd gnd cell_6t
Xbit_r151_c103 bl[103] br[103] wl[151] vdd gnd cell_6t
Xbit_r152_c103 bl[103] br[103] wl[152] vdd gnd cell_6t
Xbit_r153_c103 bl[103] br[103] wl[153] vdd gnd cell_6t
Xbit_r154_c103 bl[103] br[103] wl[154] vdd gnd cell_6t
Xbit_r155_c103 bl[103] br[103] wl[155] vdd gnd cell_6t
Xbit_r156_c103 bl[103] br[103] wl[156] vdd gnd cell_6t
Xbit_r157_c103 bl[103] br[103] wl[157] vdd gnd cell_6t
Xbit_r158_c103 bl[103] br[103] wl[158] vdd gnd cell_6t
Xbit_r159_c103 bl[103] br[103] wl[159] vdd gnd cell_6t
Xbit_r160_c103 bl[103] br[103] wl[160] vdd gnd cell_6t
Xbit_r161_c103 bl[103] br[103] wl[161] vdd gnd cell_6t
Xbit_r162_c103 bl[103] br[103] wl[162] vdd gnd cell_6t
Xbit_r163_c103 bl[103] br[103] wl[163] vdd gnd cell_6t
Xbit_r164_c103 bl[103] br[103] wl[164] vdd gnd cell_6t
Xbit_r165_c103 bl[103] br[103] wl[165] vdd gnd cell_6t
Xbit_r166_c103 bl[103] br[103] wl[166] vdd gnd cell_6t
Xbit_r167_c103 bl[103] br[103] wl[167] vdd gnd cell_6t
Xbit_r168_c103 bl[103] br[103] wl[168] vdd gnd cell_6t
Xbit_r169_c103 bl[103] br[103] wl[169] vdd gnd cell_6t
Xbit_r170_c103 bl[103] br[103] wl[170] vdd gnd cell_6t
Xbit_r171_c103 bl[103] br[103] wl[171] vdd gnd cell_6t
Xbit_r172_c103 bl[103] br[103] wl[172] vdd gnd cell_6t
Xbit_r173_c103 bl[103] br[103] wl[173] vdd gnd cell_6t
Xbit_r174_c103 bl[103] br[103] wl[174] vdd gnd cell_6t
Xbit_r175_c103 bl[103] br[103] wl[175] vdd gnd cell_6t
Xbit_r176_c103 bl[103] br[103] wl[176] vdd gnd cell_6t
Xbit_r177_c103 bl[103] br[103] wl[177] vdd gnd cell_6t
Xbit_r178_c103 bl[103] br[103] wl[178] vdd gnd cell_6t
Xbit_r179_c103 bl[103] br[103] wl[179] vdd gnd cell_6t
Xbit_r180_c103 bl[103] br[103] wl[180] vdd gnd cell_6t
Xbit_r181_c103 bl[103] br[103] wl[181] vdd gnd cell_6t
Xbit_r182_c103 bl[103] br[103] wl[182] vdd gnd cell_6t
Xbit_r183_c103 bl[103] br[103] wl[183] vdd gnd cell_6t
Xbit_r184_c103 bl[103] br[103] wl[184] vdd gnd cell_6t
Xbit_r185_c103 bl[103] br[103] wl[185] vdd gnd cell_6t
Xbit_r186_c103 bl[103] br[103] wl[186] vdd gnd cell_6t
Xbit_r187_c103 bl[103] br[103] wl[187] vdd gnd cell_6t
Xbit_r188_c103 bl[103] br[103] wl[188] vdd gnd cell_6t
Xbit_r189_c103 bl[103] br[103] wl[189] vdd gnd cell_6t
Xbit_r190_c103 bl[103] br[103] wl[190] vdd gnd cell_6t
Xbit_r191_c103 bl[103] br[103] wl[191] vdd gnd cell_6t
Xbit_r192_c103 bl[103] br[103] wl[192] vdd gnd cell_6t
Xbit_r193_c103 bl[103] br[103] wl[193] vdd gnd cell_6t
Xbit_r194_c103 bl[103] br[103] wl[194] vdd gnd cell_6t
Xbit_r195_c103 bl[103] br[103] wl[195] vdd gnd cell_6t
Xbit_r196_c103 bl[103] br[103] wl[196] vdd gnd cell_6t
Xbit_r197_c103 bl[103] br[103] wl[197] vdd gnd cell_6t
Xbit_r198_c103 bl[103] br[103] wl[198] vdd gnd cell_6t
Xbit_r199_c103 bl[103] br[103] wl[199] vdd gnd cell_6t
Xbit_r200_c103 bl[103] br[103] wl[200] vdd gnd cell_6t
Xbit_r201_c103 bl[103] br[103] wl[201] vdd gnd cell_6t
Xbit_r202_c103 bl[103] br[103] wl[202] vdd gnd cell_6t
Xbit_r203_c103 bl[103] br[103] wl[203] vdd gnd cell_6t
Xbit_r204_c103 bl[103] br[103] wl[204] vdd gnd cell_6t
Xbit_r205_c103 bl[103] br[103] wl[205] vdd gnd cell_6t
Xbit_r206_c103 bl[103] br[103] wl[206] vdd gnd cell_6t
Xbit_r207_c103 bl[103] br[103] wl[207] vdd gnd cell_6t
Xbit_r208_c103 bl[103] br[103] wl[208] vdd gnd cell_6t
Xbit_r209_c103 bl[103] br[103] wl[209] vdd gnd cell_6t
Xbit_r210_c103 bl[103] br[103] wl[210] vdd gnd cell_6t
Xbit_r211_c103 bl[103] br[103] wl[211] vdd gnd cell_6t
Xbit_r212_c103 bl[103] br[103] wl[212] vdd gnd cell_6t
Xbit_r213_c103 bl[103] br[103] wl[213] vdd gnd cell_6t
Xbit_r214_c103 bl[103] br[103] wl[214] vdd gnd cell_6t
Xbit_r215_c103 bl[103] br[103] wl[215] vdd gnd cell_6t
Xbit_r216_c103 bl[103] br[103] wl[216] vdd gnd cell_6t
Xbit_r217_c103 bl[103] br[103] wl[217] vdd gnd cell_6t
Xbit_r218_c103 bl[103] br[103] wl[218] vdd gnd cell_6t
Xbit_r219_c103 bl[103] br[103] wl[219] vdd gnd cell_6t
Xbit_r220_c103 bl[103] br[103] wl[220] vdd gnd cell_6t
Xbit_r221_c103 bl[103] br[103] wl[221] vdd gnd cell_6t
Xbit_r222_c103 bl[103] br[103] wl[222] vdd gnd cell_6t
Xbit_r223_c103 bl[103] br[103] wl[223] vdd gnd cell_6t
Xbit_r224_c103 bl[103] br[103] wl[224] vdd gnd cell_6t
Xbit_r225_c103 bl[103] br[103] wl[225] vdd gnd cell_6t
Xbit_r226_c103 bl[103] br[103] wl[226] vdd gnd cell_6t
Xbit_r227_c103 bl[103] br[103] wl[227] vdd gnd cell_6t
Xbit_r228_c103 bl[103] br[103] wl[228] vdd gnd cell_6t
Xbit_r229_c103 bl[103] br[103] wl[229] vdd gnd cell_6t
Xbit_r230_c103 bl[103] br[103] wl[230] vdd gnd cell_6t
Xbit_r231_c103 bl[103] br[103] wl[231] vdd gnd cell_6t
Xbit_r232_c103 bl[103] br[103] wl[232] vdd gnd cell_6t
Xbit_r233_c103 bl[103] br[103] wl[233] vdd gnd cell_6t
Xbit_r234_c103 bl[103] br[103] wl[234] vdd gnd cell_6t
Xbit_r235_c103 bl[103] br[103] wl[235] vdd gnd cell_6t
Xbit_r236_c103 bl[103] br[103] wl[236] vdd gnd cell_6t
Xbit_r237_c103 bl[103] br[103] wl[237] vdd gnd cell_6t
Xbit_r238_c103 bl[103] br[103] wl[238] vdd gnd cell_6t
Xbit_r239_c103 bl[103] br[103] wl[239] vdd gnd cell_6t
Xbit_r240_c103 bl[103] br[103] wl[240] vdd gnd cell_6t
Xbit_r241_c103 bl[103] br[103] wl[241] vdd gnd cell_6t
Xbit_r242_c103 bl[103] br[103] wl[242] vdd gnd cell_6t
Xbit_r243_c103 bl[103] br[103] wl[243] vdd gnd cell_6t
Xbit_r244_c103 bl[103] br[103] wl[244] vdd gnd cell_6t
Xbit_r245_c103 bl[103] br[103] wl[245] vdd gnd cell_6t
Xbit_r246_c103 bl[103] br[103] wl[246] vdd gnd cell_6t
Xbit_r247_c103 bl[103] br[103] wl[247] vdd gnd cell_6t
Xbit_r248_c103 bl[103] br[103] wl[248] vdd gnd cell_6t
Xbit_r249_c103 bl[103] br[103] wl[249] vdd gnd cell_6t
Xbit_r250_c103 bl[103] br[103] wl[250] vdd gnd cell_6t
Xbit_r251_c103 bl[103] br[103] wl[251] vdd gnd cell_6t
Xbit_r252_c103 bl[103] br[103] wl[252] vdd gnd cell_6t
Xbit_r253_c103 bl[103] br[103] wl[253] vdd gnd cell_6t
Xbit_r254_c103 bl[103] br[103] wl[254] vdd gnd cell_6t
Xbit_r255_c103 bl[103] br[103] wl[255] vdd gnd cell_6t
Xbit_r0_c104 bl[104] br[104] wl[0] vdd gnd cell_6t
Xbit_r1_c104 bl[104] br[104] wl[1] vdd gnd cell_6t
Xbit_r2_c104 bl[104] br[104] wl[2] vdd gnd cell_6t
Xbit_r3_c104 bl[104] br[104] wl[3] vdd gnd cell_6t
Xbit_r4_c104 bl[104] br[104] wl[4] vdd gnd cell_6t
Xbit_r5_c104 bl[104] br[104] wl[5] vdd gnd cell_6t
Xbit_r6_c104 bl[104] br[104] wl[6] vdd gnd cell_6t
Xbit_r7_c104 bl[104] br[104] wl[7] vdd gnd cell_6t
Xbit_r8_c104 bl[104] br[104] wl[8] vdd gnd cell_6t
Xbit_r9_c104 bl[104] br[104] wl[9] vdd gnd cell_6t
Xbit_r10_c104 bl[104] br[104] wl[10] vdd gnd cell_6t
Xbit_r11_c104 bl[104] br[104] wl[11] vdd gnd cell_6t
Xbit_r12_c104 bl[104] br[104] wl[12] vdd gnd cell_6t
Xbit_r13_c104 bl[104] br[104] wl[13] vdd gnd cell_6t
Xbit_r14_c104 bl[104] br[104] wl[14] vdd gnd cell_6t
Xbit_r15_c104 bl[104] br[104] wl[15] vdd gnd cell_6t
Xbit_r16_c104 bl[104] br[104] wl[16] vdd gnd cell_6t
Xbit_r17_c104 bl[104] br[104] wl[17] vdd gnd cell_6t
Xbit_r18_c104 bl[104] br[104] wl[18] vdd gnd cell_6t
Xbit_r19_c104 bl[104] br[104] wl[19] vdd gnd cell_6t
Xbit_r20_c104 bl[104] br[104] wl[20] vdd gnd cell_6t
Xbit_r21_c104 bl[104] br[104] wl[21] vdd gnd cell_6t
Xbit_r22_c104 bl[104] br[104] wl[22] vdd gnd cell_6t
Xbit_r23_c104 bl[104] br[104] wl[23] vdd gnd cell_6t
Xbit_r24_c104 bl[104] br[104] wl[24] vdd gnd cell_6t
Xbit_r25_c104 bl[104] br[104] wl[25] vdd gnd cell_6t
Xbit_r26_c104 bl[104] br[104] wl[26] vdd gnd cell_6t
Xbit_r27_c104 bl[104] br[104] wl[27] vdd gnd cell_6t
Xbit_r28_c104 bl[104] br[104] wl[28] vdd gnd cell_6t
Xbit_r29_c104 bl[104] br[104] wl[29] vdd gnd cell_6t
Xbit_r30_c104 bl[104] br[104] wl[30] vdd gnd cell_6t
Xbit_r31_c104 bl[104] br[104] wl[31] vdd gnd cell_6t
Xbit_r32_c104 bl[104] br[104] wl[32] vdd gnd cell_6t
Xbit_r33_c104 bl[104] br[104] wl[33] vdd gnd cell_6t
Xbit_r34_c104 bl[104] br[104] wl[34] vdd gnd cell_6t
Xbit_r35_c104 bl[104] br[104] wl[35] vdd gnd cell_6t
Xbit_r36_c104 bl[104] br[104] wl[36] vdd gnd cell_6t
Xbit_r37_c104 bl[104] br[104] wl[37] vdd gnd cell_6t
Xbit_r38_c104 bl[104] br[104] wl[38] vdd gnd cell_6t
Xbit_r39_c104 bl[104] br[104] wl[39] vdd gnd cell_6t
Xbit_r40_c104 bl[104] br[104] wl[40] vdd gnd cell_6t
Xbit_r41_c104 bl[104] br[104] wl[41] vdd gnd cell_6t
Xbit_r42_c104 bl[104] br[104] wl[42] vdd gnd cell_6t
Xbit_r43_c104 bl[104] br[104] wl[43] vdd gnd cell_6t
Xbit_r44_c104 bl[104] br[104] wl[44] vdd gnd cell_6t
Xbit_r45_c104 bl[104] br[104] wl[45] vdd gnd cell_6t
Xbit_r46_c104 bl[104] br[104] wl[46] vdd gnd cell_6t
Xbit_r47_c104 bl[104] br[104] wl[47] vdd gnd cell_6t
Xbit_r48_c104 bl[104] br[104] wl[48] vdd gnd cell_6t
Xbit_r49_c104 bl[104] br[104] wl[49] vdd gnd cell_6t
Xbit_r50_c104 bl[104] br[104] wl[50] vdd gnd cell_6t
Xbit_r51_c104 bl[104] br[104] wl[51] vdd gnd cell_6t
Xbit_r52_c104 bl[104] br[104] wl[52] vdd gnd cell_6t
Xbit_r53_c104 bl[104] br[104] wl[53] vdd gnd cell_6t
Xbit_r54_c104 bl[104] br[104] wl[54] vdd gnd cell_6t
Xbit_r55_c104 bl[104] br[104] wl[55] vdd gnd cell_6t
Xbit_r56_c104 bl[104] br[104] wl[56] vdd gnd cell_6t
Xbit_r57_c104 bl[104] br[104] wl[57] vdd gnd cell_6t
Xbit_r58_c104 bl[104] br[104] wl[58] vdd gnd cell_6t
Xbit_r59_c104 bl[104] br[104] wl[59] vdd gnd cell_6t
Xbit_r60_c104 bl[104] br[104] wl[60] vdd gnd cell_6t
Xbit_r61_c104 bl[104] br[104] wl[61] vdd gnd cell_6t
Xbit_r62_c104 bl[104] br[104] wl[62] vdd gnd cell_6t
Xbit_r63_c104 bl[104] br[104] wl[63] vdd gnd cell_6t
Xbit_r64_c104 bl[104] br[104] wl[64] vdd gnd cell_6t
Xbit_r65_c104 bl[104] br[104] wl[65] vdd gnd cell_6t
Xbit_r66_c104 bl[104] br[104] wl[66] vdd gnd cell_6t
Xbit_r67_c104 bl[104] br[104] wl[67] vdd gnd cell_6t
Xbit_r68_c104 bl[104] br[104] wl[68] vdd gnd cell_6t
Xbit_r69_c104 bl[104] br[104] wl[69] vdd gnd cell_6t
Xbit_r70_c104 bl[104] br[104] wl[70] vdd gnd cell_6t
Xbit_r71_c104 bl[104] br[104] wl[71] vdd gnd cell_6t
Xbit_r72_c104 bl[104] br[104] wl[72] vdd gnd cell_6t
Xbit_r73_c104 bl[104] br[104] wl[73] vdd gnd cell_6t
Xbit_r74_c104 bl[104] br[104] wl[74] vdd gnd cell_6t
Xbit_r75_c104 bl[104] br[104] wl[75] vdd gnd cell_6t
Xbit_r76_c104 bl[104] br[104] wl[76] vdd gnd cell_6t
Xbit_r77_c104 bl[104] br[104] wl[77] vdd gnd cell_6t
Xbit_r78_c104 bl[104] br[104] wl[78] vdd gnd cell_6t
Xbit_r79_c104 bl[104] br[104] wl[79] vdd gnd cell_6t
Xbit_r80_c104 bl[104] br[104] wl[80] vdd gnd cell_6t
Xbit_r81_c104 bl[104] br[104] wl[81] vdd gnd cell_6t
Xbit_r82_c104 bl[104] br[104] wl[82] vdd gnd cell_6t
Xbit_r83_c104 bl[104] br[104] wl[83] vdd gnd cell_6t
Xbit_r84_c104 bl[104] br[104] wl[84] vdd gnd cell_6t
Xbit_r85_c104 bl[104] br[104] wl[85] vdd gnd cell_6t
Xbit_r86_c104 bl[104] br[104] wl[86] vdd gnd cell_6t
Xbit_r87_c104 bl[104] br[104] wl[87] vdd gnd cell_6t
Xbit_r88_c104 bl[104] br[104] wl[88] vdd gnd cell_6t
Xbit_r89_c104 bl[104] br[104] wl[89] vdd gnd cell_6t
Xbit_r90_c104 bl[104] br[104] wl[90] vdd gnd cell_6t
Xbit_r91_c104 bl[104] br[104] wl[91] vdd gnd cell_6t
Xbit_r92_c104 bl[104] br[104] wl[92] vdd gnd cell_6t
Xbit_r93_c104 bl[104] br[104] wl[93] vdd gnd cell_6t
Xbit_r94_c104 bl[104] br[104] wl[94] vdd gnd cell_6t
Xbit_r95_c104 bl[104] br[104] wl[95] vdd gnd cell_6t
Xbit_r96_c104 bl[104] br[104] wl[96] vdd gnd cell_6t
Xbit_r97_c104 bl[104] br[104] wl[97] vdd gnd cell_6t
Xbit_r98_c104 bl[104] br[104] wl[98] vdd gnd cell_6t
Xbit_r99_c104 bl[104] br[104] wl[99] vdd gnd cell_6t
Xbit_r100_c104 bl[104] br[104] wl[100] vdd gnd cell_6t
Xbit_r101_c104 bl[104] br[104] wl[101] vdd gnd cell_6t
Xbit_r102_c104 bl[104] br[104] wl[102] vdd gnd cell_6t
Xbit_r103_c104 bl[104] br[104] wl[103] vdd gnd cell_6t
Xbit_r104_c104 bl[104] br[104] wl[104] vdd gnd cell_6t
Xbit_r105_c104 bl[104] br[104] wl[105] vdd gnd cell_6t
Xbit_r106_c104 bl[104] br[104] wl[106] vdd gnd cell_6t
Xbit_r107_c104 bl[104] br[104] wl[107] vdd gnd cell_6t
Xbit_r108_c104 bl[104] br[104] wl[108] vdd gnd cell_6t
Xbit_r109_c104 bl[104] br[104] wl[109] vdd gnd cell_6t
Xbit_r110_c104 bl[104] br[104] wl[110] vdd gnd cell_6t
Xbit_r111_c104 bl[104] br[104] wl[111] vdd gnd cell_6t
Xbit_r112_c104 bl[104] br[104] wl[112] vdd gnd cell_6t
Xbit_r113_c104 bl[104] br[104] wl[113] vdd gnd cell_6t
Xbit_r114_c104 bl[104] br[104] wl[114] vdd gnd cell_6t
Xbit_r115_c104 bl[104] br[104] wl[115] vdd gnd cell_6t
Xbit_r116_c104 bl[104] br[104] wl[116] vdd gnd cell_6t
Xbit_r117_c104 bl[104] br[104] wl[117] vdd gnd cell_6t
Xbit_r118_c104 bl[104] br[104] wl[118] vdd gnd cell_6t
Xbit_r119_c104 bl[104] br[104] wl[119] vdd gnd cell_6t
Xbit_r120_c104 bl[104] br[104] wl[120] vdd gnd cell_6t
Xbit_r121_c104 bl[104] br[104] wl[121] vdd gnd cell_6t
Xbit_r122_c104 bl[104] br[104] wl[122] vdd gnd cell_6t
Xbit_r123_c104 bl[104] br[104] wl[123] vdd gnd cell_6t
Xbit_r124_c104 bl[104] br[104] wl[124] vdd gnd cell_6t
Xbit_r125_c104 bl[104] br[104] wl[125] vdd gnd cell_6t
Xbit_r126_c104 bl[104] br[104] wl[126] vdd gnd cell_6t
Xbit_r127_c104 bl[104] br[104] wl[127] vdd gnd cell_6t
Xbit_r128_c104 bl[104] br[104] wl[128] vdd gnd cell_6t
Xbit_r129_c104 bl[104] br[104] wl[129] vdd gnd cell_6t
Xbit_r130_c104 bl[104] br[104] wl[130] vdd gnd cell_6t
Xbit_r131_c104 bl[104] br[104] wl[131] vdd gnd cell_6t
Xbit_r132_c104 bl[104] br[104] wl[132] vdd gnd cell_6t
Xbit_r133_c104 bl[104] br[104] wl[133] vdd gnd cell_6t
Xbit_r134_c104 bl[104] br[104] wl[134] vdd gnd cell_6t
Xbit_r135_c104 bl[104] br[104] wl[135] vdd gnd cell_6t
Xbit_r136_c104 bl[104] br[104] wl[136] vdd gnd cell_6t
Xbit_r137_c104 bl[104] br[104] wl[137] vdd gnd cell_6t
Xbit_r138_c104 bl[104] br[104] wl[138] vdd gnd cell_6t
Xbit_r139_c104 bl[104] br[104] wl[139] vdd gnd cell_6t
Xbit_r140_c104 bl[104] br[104] wl[140] vdd gnd cell_6t
Xbit_r141_c104 bl[104] br[104] wl[141] vdd gnd cell_6t
Xbit_r142_c104 bl[104] br[104] wl[142] vdd gnd cell_6t
Xbit_r143_c104 bl[104] br[104] wl[143] vdd gnd cell_6t
Xbit_r144_c104 bl[104] br[104] wl[144] vdd gnd cell_6t
Xbit_r145_c104 bl[104] br[104] wl[145] vdd gnd cell_6t
Xbit_r146_c104 bl[104] br[104] wl[146] vdd gnd cell_6t
Xbit_r147_c104 bl[104] br[104] wl[147] vdd gnd cell_6t
Xbit_r148_c104 bl[104] br[104] wl[148] vdd gnd cell_6t
Xbit_r149_c104 bl[104] br[104] wl[149] vdd gnd cell_6t
Xbit_r150_c104 bl[104] br[104] wl[150] vdd gnd cell_6t
Xbit_r151_c104 bl[104] br[104] wl[151] vdd gnd cell_6t
Xbit_r152_c104 bl[104] br[104] wl[152] vdd gnd cell_6t
Xbit_r153_c104 bl[104] br[104] wl[153] vdd gnd cell_6t
Xbit_r154_c104 bl[104] br[104] wl[154] vdd gnd cell_6t
Xbit_r155_c104 bl[104] br[104] wl[155] vdd gnd cell_6t
Xbit_r156_c104 bl[104] br[104] wl[156] vdd gnd cell_6t
Xbit_r157_c104 bl[104] br[104] wl[157] vdd gnd cell_6t
Xbit_r158_c104 bl[104] br[104] wl[158] vdd gnd cell_6t
Xbit_r159_c104 bl[104] br[104] wl[159] vdd gnd cell_6t
Xbit_r160_c104 bl[104] br[104] wl[160] vdd gnd cell_6t
Xbit_r161_c104 bl[104] br[104] wl[161] vdd gnd cell_6t
Xbit_r162_c104 bl[104] br[104] wl[162] vdd gnd cell_6t
Xbit_r163_c104 bl[104] br[104] wl[163] vdd gnd cell_6t
Xbit_r164_c104 bl[104] br[104] wl[164] vdd gnd cell_6t
Xbit_r165_c104 bl[104] br[104] wl[165] vdd gnd cell_6t
Xbit_r166_c104 bl[104] br[104] wl[166] vdd gnd cell_6t
Xbit_r167_c104 bl[104] br[104] wl[167] vdd gnd cell_6t
Xbit_r168_c104 bl[104] br[104] wl[168] vdd gnd cell_6t
Xbit_r169_c104 bl[104] br[104] wl[169] vdd gnd cell_6t
Xbit_r170_c104 bl[104] br[104] wl[170] vdd gnd cell_6t
Xbit_r171_c104 bl[104] br[104] wl[171] vdd gnd cell_6t
Xbit_r172_c104 bl[104] br[104] wl[172] vdd gnd cell_6t
Xbit_r173_c104 bl[104] br[104] wl[173] vdd gnd cell_6t
Xbit_r174_c104 bl[104] br[104] wl[174] vdd gnd cell_6t
Xbit_r175_c104 bl[104] br[104] wl[175] vdd gnd cell_6t
Xbit_r176_c104 bl[104] br[104] wl[176] vdd gnd cell_6t
Xbit_r177_c104 bl[104] br[104] wl[177] vdd gnd cell_6t
Xbit_r178_c104 bl[104] br[104] wl[178] vdd gnd cell_6t
Xbit_r179_c104 bl[104] br[104] wl[179] vdd gnd cell_6t
Xbit_r180_c104 bl[104] br[104] wl[180] vdd gnd cell_6t
Xbit_r181_c104 bl[104] br[104] wl[181] vdd gnd cell_6t
Xbit_r182_c104 bl[104] br[104] wl[182] vdd gnd cell_6t
Xbit_r183_c104 bl[104] br[104] wl[183] vdd gnd cell_6t
Xbit_r184_c104 bl[104] br[104] wl[184] vdd gnd cell_6t
Xbit_r185_c104 bl[104] br[104] wl[185] vdd gnd cell_6t
Xbit_r186_c104 bl[104] br[104] wl[186] vdd gnd cell_6t
Xbit_r187_c104 bl[104] br[104] wl[187] vdd gnd cell_6t
Xbit_r188_c104 bl[104] br[104] wl[188] vdd gnd cell_6t
Xbit_r189_c104 bl[104] br[104] wl[189] vdd gnd cell_6t
Xbit_r190_c104 bl[104] br[104] wl[190] vdd gnd cell_6t
Xbit_r191_c104 bl[104] br[104] wl[191] vdd gnd cell_6t
Xbit_r192_c104 bl[104] br[104] wl[192] vdd gnd cell_6t
Xbit_r193_c104 bl[104] br[104] wl[193] vdd gnd cell_6t
Xbit_r194_c104 bl[104] br[104] wl[194] vdd gnd cell_6t
Xbit_r195_c104 bl[104] br[104] wl[195] vdd gnd cell_6t
Xbit_r196_c104 bl[104] br[104] wl[196] vdd gnd cell_6t
Xbit_r197_c104 bl[104] br[104] wl[197] vdd gnd cell_6t
Xbit_r198_c104 bl[104] br[104] wl[198] vdd gnd cell_6t
Xbit_r199_c104 bl[104] br[104] wl[199] vdd gnd cell_6t
Xbit_r200_c104 bl[104] br[104] wl[200] vdd gnd cell_6t
Xbit_r201_c104 bl[104] br[104] wl[201] vdd gnd cell_6t
Xbit_r202_c104 bl[104] br[104] wl[202] vdd gnd cell_6t
Xbit_r203_c104 bl[104] br[104] wl[203] vdd gnd cell_6t
Xbit_r204_c104 bl[104] br[104] wl[204] vdd gnd cell_6t
Xbit_r205_c104 bl[104] br[104] wl[205] vdd gnd cell_6t
Xbit_r206_c104 bl[104] br[104] wl[206] vdd gnd cell_6t
Xbit_r207_c104 bl[104] br[104] wl[207] vdd gnd cell_6t
Xbit_r208_c104 bl[104] br[104] wl[208] vdd gnd cell_6t
Xbit_r209_c104 bl[104] br[104] wl[209] vdd gnd cell_6t
Xbit_r210_c104 bl[104] br[104] wl[210] vdd gnd cell_6t
Xbit_r211_c104 bl[104] br[104] wl[211] vdd gnd cell_6t
Xbit_r212_c104 bl[104] br[104] wl[212] vdd gnd cell_6t
Xbit_r213_c104 bl[104] br[104] wl[213] vdd gnd cell_6t
Xbit_r214_c104 bl[104] br[104] wl[214] vdd gnd cell_6t
Xbit_r215_c104 bl[104] br[104] wl[215] vdd gnd cell_6t
Xbit_r216_c104 bl[104] br[104] wl[216] vdd gnd cell_6t
Xbit_r217_c104 bl[104] br[104] wl[217] vdd gnd cell_6t
Xbit_r218_c104 bl[104] br[104] wl[218] vdd gnd cell_6t
Xbit_r219_c104 bl[104] br[104] wl[219] vdd gnd cell_6t
Xbit_r220_c104 bl[104] br[104] wl[220] vdd gnd cell_6t
Xbit_r221_c104 bl[104] br[104] wl[221] vdd gnd cell_6t
Xbit_r222_c104 bl[104] br[104] wl[222] vdd gnd cell_6t
Xbit_r223_c104 bl[104] br[104] wl[223] vdd gnd cell_6t
Xbit_r224_c104 bl[104] br[104] wl[224] vdd gnd cell_6t
Xbit_r225_c104 bl[104] br[104] wl[225] vdd gnd cell_6t
Xbit_r226_c104 bl[104] br[104] wl[226] vdd gnd cell_6t
Xbit_r227_c104 bl[104] br[104] wl[227] vdd gnd cell_6t
Xbit_r228_c104 bl[104] br[104] wl[228] vdd gnd cell_6t
Xbit_r229_c104 bl[104] br[104] wl[229] vdd gnd cell_6t
Xbit_r230_c104 bl[104] br[104] wl[230] vdd gnd cell_6t
Xbit_r231_c104 bl[104] br[104] wl[231] vdd gnd cell_6t
Xbit_r232_c104 bl[104] br[104] wl[232] vdd gnd cell_6t
Xbit_r233_c104 bl[104] br[104] wl[233] vdd gnd cell_6t
Xbit_r234_c104 bl[104] br[104] wl[234] vdd gnd cell_6t
Xbit_r235_c104 bl[104] br[104] wl[235] vdd gnd cell_6t
Xbit_r236_c104 bl[104] br[104] wl[236] vdd gnd cell_6t
Xbit_r237_c104 bl[104] br[104] wl[237] vdd gnd cell_6t
Xbit_r238_c104 bl[104] br[104] wl[238] vdd gnd cell_6t
Xbit_r239_c104 bl[104] br[104] wl[239] vdd gnd cell_6t
Xbit_r240_c104 bl[104] br[104] wl[240] vdd gnd cell_6t
Xbit_r241_c104 bl[104] br[104] wl[241] vdd gnd cell_6t
Xbit_r242_c104 bl[104] br[104] wl[242] vdd gnd cell_6t
Xbit_r243_c104 bl[104] br[104] wl[243] vdd gnd cell_6t
Xbit_r244_c104 bl[104] br[104] wl[244] vdd gnd cell_6t
Xbit_r245_c104 bl[104] br[104] wl[245] vdd gnd cell_6t
Xbit_r246_c104 bl[104] br[104] wl[246] vdd gnd cell_6t
Xbit_r247_c104 bl[104] br[104] wl[247] vdd gnd cell_6t
Xbit_r248_c104 bl[104] br[104] wl[248] vdd gnd cell_6t
Xbit_r249_c104 bl[104] br[104] wl[249] vdd gnd cell_6t
Xbit_r250_c104 bl[104] br[104] wl[250] vdd gnd cell_6t
Xbit_r251_c104 bl[104] br[104] wl[251] vdd gnd cell_6t
Xbit_r252_c104 bl[104] br[104] wl[252] vdd gnd cell_6t
Xbit_r253_c104 bl[104] br[104] wl[253] vdd gnd cell_6t
Xbit_r254_c104 bl[104] br[104] wl[254] vdd gnd cell_6t
Xbit_r255_c104 bl[104] br[104] wl[255] vdd gnd cell_6t
Xbit_r0_c105 bl[105] br[105] wl[0] vdd gnd cell_6t
Xbit_r1_c105 bl[105] br[105] wl[1] vdd gnd cell_6t
Xbit_r2_c105 bl[105] br[105] wl[2] vdd gnd cell_6t
Xbit_r3_c105 bl[105] br[105] wl[3] vdd gnd cell_6t
Xbit_r4_c105 bl[105] br[105] wl[4] vdd gnd cell_6t
Xbit_r5_c105 bl[105] br[105] wl[5] vdd gnd cell_6t
Xbit_r6_c105 bl[105] br[105] wl[6] vdd gnd cell_6t
Xbit_r7_c105 bl[105] br[105] wl[7] vdd gnd cell_6t
Xbit_r8_c105 bl[105] br[105] wl[8] vdd gnd cell_6t
Xbit_r9_c105 bl[105] br[105] wl[9] vdd gnd cell_6t
Xbit_r10_c105 bl[105] br[105] wl[10] vdd gnd cell_6t
Xbit_r11_c105 bl[105] br[105] wl[11] vdd gnd cell_6t
Xbit_r12_c105 bl[105] br[105] wl[12] vdd gnd cell_6t
Xbit_r13_c105 bl[105] br[105] wl[13] vdd gnd cell_6t
Xbit_r14_c105 bl[105] br[105] wl[14] vdd gnd cell_6t
Xbit_r15_c105 bl[105] br[105] wl[15] vdd gnd cell_6t
Xbit_r16_c105 bl[105] br[105] wl[16] vdd gnd cell_6t
Xbit_r17_c105 bl[105] br[105] wl[17] vdd gnd cell_6t
Xbit_r18_c105 bl[105] br[105] wl[18] vdd gnd cell_6t
Xbit_r19_c105 bl[105] br[105] wl[19] vdd gnd cell_6t
Xbit_r20_c105 bl[105] br[105] wl[20] vdd gnd cell_6t
Xbit_r21_c105 bl[105] br[105] wl[21] vdd gnd cell_6t
Xbit_r22_c105 bl[105] br[105] wl[22] vdd gnd cell_6t
Xbit_r23_c105 bl[105] br[105] wl[23] vdd gnd cell_6t
Xbit_r24_c105 bl[105] br[105] wl[24] vdd gnd cell_6t
Xbit_r25_c105 bl[105] br[105] wl[25] vdd gnd cell_6t
Xbit_r26_c105 bl[105] br[105] wl[26] vdd gnd cell_6t
Xbit_r27_c105 bl[105] br[105] wl[27] vdd gnd cell_6t
Xbit_r28_c105 bl[105] br[105] wl[28] vdd gnd cell_6t
Xbit_r29_c105 bl[105] br[105] wl[29] vdd gnd cell_6t
Xbit_r30_c105 bl[105] br[105] wl[30] vdd gnd cell_6t
Xbit_r31_c105 bl[105] br[105] wl[31] vdd gnd cell_6t
Xbit_r32_c105 bl[105] br[105] wl[32] vdd gnd cell_6t
Xbit_r33_c105 bl[105] br[105] wl[33] vdd gnd cell_6t
Xbit_r34_c105 bl[105] br[105] wl[34] vdd gnd cell_6t
Xbit_r35_c105 bl[105] br[105] wl[35] vdd gnd cell_6t
Xbit_r36_c105 bl[105] br[105] wl[36] vdd gnd cell_6t
Xbit_r37_c105 bl[105] br[105] wl[37] vdd gnd cell_6t
Xbit_r38_c105 bl[105] br[105] wl[38] vdd gnd cell_6t
Xbit_r39_c105 bl[105] br[105] wl[39] vdd gnd cell_6t
Xbit_r40_c105 bl[105] br[105] wl[40] vdd gnd cell_6t
Xbit_r41_c105 bl[105] br[105] wl[41] vdd gnd cell_6t
Xbit_r42_c105 bl[105] br[105] wl[42] vdd gnd cell_6t
Xbit_r43_c105 bl[105] br[105] wl[43] vdd gnd cell_6t
Xbit_r44_c105 bl[105] br[105] wl[44] vdd gnd cell_6t
Xbit_r45_c105 bl[105] br[105] wl[45] vdd gnd cell_6t
Xbit_r46_c105 bl[105] br[105] wl[46] vdd gnd cell_6t
Xbit_r47_c105 bl[105] br[105] wl[47] vdd gnd cell_6t
Xbit_r48_c105 bl[105] br[105] wl[48] vdd gnd cell_6t
Xbit_r49_c105 bl[105] br[105] wl[49] vdd gnd cell_6t
Xbit_r50_c105 bl[105] br[105] wl[50] vdd gnd cell_6t
Xbit_r51_c105 bl[105] br[105] wl[51] vdd gnd cell_6t
Xbit_r52_c105 bl[105] br[105] wl[52] vdd gnd cell_6t
Xbit_r53_c105 bl[105] br[105] wl[53] vdd gnd cell_6t
Xbit_r54_c105 bl[105] br[105] wl[54] vdd gnd cell_6t
Xbit_r55_c105 bl[105] br[105] wl[55] vdd gnd cell_6t
Xbit_r56_c105 bl[105] br[105] wl[56] vdd gnd cell_6t
Xbit_r57_c105 bl[105] br[105] wl[57] vdd gnd cell_6t
Xbit_r58_c105 bl[105] br[105] wl[58] vdd gnd cell_6t
Xbit_r59_c105 bl[105] br[105] wl[59] vdd gnd cell_6t
Xbit_r60_c105 bl[105] br[105] wl[60] vdd gnd cell_6t
Xbit_r61_c105 bl[105] br[105] wl[61] vdd gnd cell_6t
Xbit_r62_c105 bl[105] br[105] wl[62] vdd gnd cell_6t
Xbit_r63_c105 bl[105] br[105] wl[63] vdd gnd cell_6t
Xbit_r64_c105 bl[105] br[105] wl[64] vdd gnd cell_6t
Xbit_r65_c105 bl[105] br[105] wl[65] vdd gnd cell_6t
Xbit_r66_c105 bl[105] br[105] wl[66] vdd gnd cell_6t
Xbit_r67_c105 bl[105] br[105] wl[67] vdd gnd cell_6t
Xbit_r68_c105 bl[105] br[105] wl[68] vdd gnd cell_6t
Xbit_r69_c105 bl[105] br[105] wl[69] vdd gnd cell_6t
Xbit_r70_c105 bl[105] br[105] wl[70] vdd gnd cell_6t
Xbit_r71_c105 bl[105] br[105] wl[71] vdd gnd cell_6t
Xbit_r72_c105 bl[105] br[105] wl[72] vdd gnd cell_6t
Xbit_r73_c105 bl[105] br[105] wl[73] vdd gnd cell_6t
Xbit_r74_c105 bl[105] br[105] wl[74] vdd gnd cell_6t
Xbit_r75_c105 bl[105] br[105] wl[75] vdd gnd cell_6t
Xbit_r76_c105 bl[105] br[105] wl[76] vdd gnd cell_6t
Xbit_r77_c105 bl[105] br[105] wl[77] vdd gnd cell_6t
Xbit_r78_c105 bl[105] br[105] wl[78] vdd gnd cell_6t
Xbit_r79_c105 bl[105] br[105] wl[79] vdd gnd cell_6t
Xbit_r80_c105 bl[105] br[105] wl[80] vdd gnd cell_6t
Xbit_r81_c105 bl[105] br[105] wl[81] vdd gnd cell_6t
Xbit_r82_c105 bl[105] br[105] wl[82] vdd gnd cell_6t
Xbit_r83_c105 bl[105] br[105] wl[83] vdd gnd cell_6t
Xbit_r84_c105 bl[105] br[105] wl[84] vdd gnd cell_6t
Xbit_r85_c105 bl[105] br[105] wl[85] vdd gnd cell_6t
Xbit_r86_c105 bl[105] br[105] wl[86] vdd gnd cell_6t
Xbit_r87_c105 bl[105] br[105] wl[87] vdd gnd cell_6t
Xbit_r88_c105 bl[105] br[105] wl[88] vdd gnd cell_6t
Xbit_r89_c105 bl[105] br[105] wl[89] vdd gnd cell_6t
Xbit_r90_c105 bl[105] br[105] wl[90] vdd gnd cell_6t
Xbit_r91_c105 bl[105] br[105] wl[91] vdd gnd cell_6t
Xbit_r92_c105 bl[105] br[105] wl[92] vdd gnd cell_6t
Xbit_r93_c105 bl[105] br[105] wl[93] vdd gnd cell_6t
Xbit_r94_c105 bl[105] br[105] wl[94] vdd gnd cell_6t
Xbit_r95_c105 bl[105] br[105] wl[95] vdd gnd cell_6t
Xbit_r96_c105 bl[105] br[105] wl[96] vdd gnd cell_6t
Xbit_r97_c105 bl[105] br[105] wl[97] vdd gnd cell_6t
Xbit_r98_c105 bl[105] br[105] wl[98] vdd gnd cell_6t
Xbit_r99_c105 bl[105] br[105] wl[99] vdd gnd cell_6t
Xbit_r100_c105 bl[105] br[105] wl[100] vdd gnd cell_6t
Xbit_r101_c105 bl[105] br[105] wl[101] vdd gnd cell_6t
Xbit_r102_c105 bl[105] br[105] wl[102] vdd gnd cell_6t
Xbit_r103_c105 bl[105] br[105] wl[103] vdd gnd cell_6t
Xbit_r104_c105 bl[105] br[105] wl[104] vdd gnd cell_6t
Xbit_r105_c105 bl[105] br[105] wl[105] vdd gnd cell_6t
Xbit_r106_c105 bl[105] br[105] wl[106] vdd gnd cell_6t
Xbit_r107_c105 bl[105] br[105] wl[107] vdd gnd cell_6t
Xbit_r108_c105 bl[105] br[105] wl[108] vdd gnd cell_6t
Xbit_r109_c105 bl[105] br[105] wl[109] vdd gnd cell_6t
Xbit_r110_c105 bl[105] br[105] wl[110] vdd gnd cell_6t
Xbit_r111_c105 bl[105] br[105] wl[111] vdd gnd cell_6t
Xbit_r112_c105 bl[105] br[105] wl[112] vdd gnd cell_6t
Xbit_r113_c105 bl[105] br[105] wl[113] vdd gnd cell_6t
Xbit_r114_c105 bl[105] br[105] wl[114] vdd gnd cell_6t
Xbit_r115_c105 bl[105] br[105] wl[115] vdd gnd cell_6t
Xbit_r116_c105 bl[105] br[105] wl[116] vdd gnd cell_6t
Xbit_r117_c105 bl[105] br[105] wl[117] vdd gnd cell_6t
Xbit_r118_c105 bl[105] br[105] wl[118] vdd gnd cell_6t
Xbit_r119_c105 bl[105] br[105] wl[119] vdd gnd cell_6t
Xbit_r120_c105 bl[105] br[105] wl[120] vdd gnd cell_6t
Xbit_r121_c105 bl[105] br[105] wl[121] vdd gnd cell_6t
Xbit_r122_c105 bl[105] br[105] wl[122] vdd gnd cell_6t
Xbit_r123_c105 bl[105] br[105] wl[123] vdd gnd cell_6t
Xbit_r124_c105 bl[105] br[105] wl[124] vdd gnd cell_6t
Xbit_r125_c105 bl[105] br[105] wl[125] vdd gnd cell_6t
Xbit_r126_c105 bl[105] br[105] wl[126] vdd gnd cell_6t
Xbit_r127_c105 bl[105] br[105] wl[127] vdd gnd cell_6t
Xbit_r128_c105 bl[105] br[105] wl[128] vdd gnd cell_6t
Xbit_r129_c105 bl[105] br[105] wl[129] vdd gnd cell_6t
Xbit_r130_c105 bl[105] br[105] wl[130] vdd gnd cell_6t
Xbit_r131_c105 bl[105] br[105] wl[131] vdd gnd cell_6t
Xbit_r132_c105 bl[105] br[105] wl[132] vdd gnd cell_6t
Xbit_r133_c105 bl[105] br[105] wl[133] vdd gnd cell_6t
Xbit_r134_c105 bl[105] br[105] wl[134] vdd gnd cell_6t
Xbit_r135_c105 bl[105] br[105] wl[135] vdd gnd cell_6t
Xbit_r136_c105 bl[105] br[105] wl[136] vdd gnd cell_6t
Xbit_r137_c105 bl[105] br[105] wl[137] vdd gnd cell_6t
Xbit_r138_c105 bl[105] br[105] wl[138] vdd gnd cell_6t
Xbit_r139_c105 bl[105] br[105] wl[139] vdd gnd cell_6t
Xbit_r140_c105 bl[105] br[105] wl[140] vdd gnd cell_6t
Xbit_r141_c105 bl[105] br[105] wl[141] vdd gnd cell_6t
Xbit_r142_c105 bl[105] br[105] wl[142] vdd gnd cell_6t
Xbit_r143_c105 bl[105] br[105] wl[143] vdd gnd cell_6t
Xbit_r144_c105 bl[105] br[105] wl[144] vdd gnd cell_6t
Xbit_r145_c105 bl[105] br[105] wl[145] vdd gnd cell_6t
Xbit_r146_c105 bl[105] br[105] wl[146] vdd gnd cell_6t
Xbit_r147_c105 bl[105] br[105] wl[147] vdd gnd cell_6t
Xbit_r148_c105 bl[105] br[105] wl[148] vdd gnd cell_6t
Xbit_r149_c105 bl[105] br[105] wl[149] vdd gnd cell_6t
Xbit_r150_c105 bl[105] br[105] wl[150] vdd gnd cell_6t
Xbit_r151_c105 bl[105] br[105] wl[151] vdd gnd cell_6t
Xbit_r152_c105 bl[105] br[105] wl[152] vdd gnd cell_6t
Xbit_r153_c105 bl[105] br[105] wl[153] vdd gnd cell_6t
Xbit_r154_c105 bl[105] br[105] wl[154] vdd gnd cell_6t
Xbit_r155_c105 bl[105] br[105] wl[155] vdd gnd cell_6t
Xbit_r156_c105 bl[105] br[105] wl[156] vdd gnd cell_6t
Xbit_r157_c105 bl[105] br[105] wl[157] vdd gnd cell_6t
Xbit_r158_c105 bl[105] br[105] wl[158] vdd gnd cell_6t
Xbit_r159_c105 bl[105] br[105] wl[159] vdd gnd cell_6t
Xbit_r160_c105 bl[105] br[105] wl[160] vdd gnd cell_6t
Xbit_r161_c105 bl[105] br[105] wl[161] vdd gnd cell_6t
Xbit_r162_c105 bl[105] br[105] wl[162] vdd gnd cell_6t
Xbit_r163_c105 bl[105] br[105] wl[163] vdd gnd cell_6t
Xbit_r164_c105 bl[105] br[105] wl[164] vdd gnd cell_6t
Xbit_r165_c105 bl[105] br[105] wl[165] vdd gnd cell_6t
Xbit_r166_c105 bl[105] br[105] wl[166] vdd gnd cell_6t
Xbit_r167_c105 bl[105] br[105] wl[167] vdd gnd cell_6t
Xbit_r168_c105 bl[105] br[105] wl[168] vdd gnd cell_6t
Xbit_r169_c105 bl[105] br[105] wl[169] vdd gnd cell_6t
Xbit_r170_c105 bl[105] br[105] wl[170] vdd gnd cell_6t
Xbit_r171_c105 bl[105] br[105] wl[171] vdd gnd cell_6t
Xbit_r172_c105 bl[105] br[105] wl[172] vdd gnd cell_6t
Xbit_r173_c105 bl[105] br[105] wl[173] vdd gnd cell_6t
Xbit_r174_c105 bl[105] br[105] wl[174] vdd gnd cell_6t
Xbit_r175_c105 bl[105] br[105] wl[175] vdd gnd cell_6t
Xbit_r176_c105 bl[105] br[105] wl[176] vdd gnd cell_6t
Xbit_r177_c105 bl[105] br[105] wl[177] vdd gnd cell_6t
Xbit_r178_c105 bl[105] br[105] wl[178] vdd gnd cell_6t
Xbit_r179_c105 bl[105] br[105] wl[179] vdd gnd cell_6t
Xbit_r180_c105 bl[105] br[105] wl[180] vdd gnd cell_6t
Xbit_r181_c105 bl[105] br[105] wl[181] vdd gnd cell_6t
Xbit_r182_c105 bl[105] br[105] wl[182] vdd gnd cell_6t
Xbit_r183_c105 bl[105] br[105] wl[183] vdd gnd cell_6t
Xbit_r184_c105 bl[105] br[105] wl[184] vdd gnd cell_6t
Xbit_r185_c105 bl[105] br[105] wl[185] vdd gnd cell_6t
Xbit_r186_c105 bl[105] br[105] wl[186] vdd gnd cell_6t
Xbit_r187_c105 bl[105] br[105] wl[187] vdd gnd cell_6t
Xbit_r188_c105 bl[105] br[105] wl[188] vdd gnd cell_6t
Xbit_r189_c105 bl[105] br[105] wl[189] vdd gnd cell_6t
Xbit_r190_c105 bl[105] br[105] wl[190] vdd gnd cell_6t
Xbit_r191_c105 bl[105] br[105] wl[191] vdd gnd cell_6t
Xbit_r192_c105 bl[105] br[105] wl[192] vdd gnd cell_6t
Xbit_r193_c105 bl[105] br[105] wl[193] vdd gnd cell_6t
Xbit_r194_c105 bl[105] br[105] wl[194] vdd gnd cell_6t
Xbit_r195_c105 bl[105] br[105] wl[195] vdd gnd cell_6t
Xbit_r196_c105 bl[105] br[105] wl[196] vdd gnd cell_6t
Xbit_r197_c105 bl[105] br[105] wl[197] vdd gnd cell_6t
Xbit_r198_c105 bl[105] br[105] wl[198] vdd gnd cell_6t
Xbit_r199_c105 bl[105] br[105] wl[199] vdd gnd cell_6t
Xbit_r200_c105 bl[105] br[105] wl[200] vdd gnd cell_6t
Xbit_r201_c105 bl[105] br[105] wl[201] vdd gnd cell_6t
Xbit_r202_c105 bl[105] br[105] wl[202] vdd gnd cell_6t
Xbit_r203_c105 bl[105] br[105] wl[203] vdd gnd cell_6t
Xbit_r204_c105 bl[105] br[105] wl[204] vdd gnd cell_6t
Xbit_r205_c105 bl[105] br[105] wl[205] vdd gnd cell_6t
Xbit_r206_c105 bl[105] br[105] wl[206] vdd gnd cell_6t
Xbit_r207_c105 bl[105] br[105] wl[207] vdd gnd cell_6t
Xbit_r208_c105 bl[105] br[105] wl[208] vdd gnd cell_6t
Xbit_r209_c105 bl[105] br[105] wl[209] vdd gnd cell_6t
Xbit_r210_c105 bl[105] br[105] wl[210] vdd gnd cell_6t
Xbit_r211_c105 bl[105] br[105] wl[211] vdd gnd cell_6t
Xbit_r212_c105 bl[105] br[105] wl[212] vdd gnd cell_6t
Xbit_r213_c105 bl[105] br[105] wl[213] vdd gnd cell_6t
Xbit_r214_c105 bl[105] br[105] wl[214] vdd gnd cell_6t
Xbit_r215_c105 bl[105] br[105] wl[215] vdd gnd cell_6t
Xbit_r216_c105 bl[105] br[105] wl[216] vdd gnd cell_6t
Xbit_r217_c105 bl[105] br[105] wl[217] vdd gnd cell_6t
Xbit_r218_c105 bl[105] br[105] wl[218] vdd gnd cell_6t
Xbit_r219_c105 bl[105] br[105] wl[219] vdd gnd cell_6t
Xbit_r220_c105 bl[105] br[105] wl[220] vdd gnd cell_6t
Xbit_r221_c105 bl[105] br[105] wl[221] vdd gnd cell_6t
Xbit_r222_c105 bl[105] br[105] wl[222] vdd gnd cell_6t
Xbit_r223_c105 bl[105] br[105] wl[223] vdd gnd cell_6t
Xbit_r224_c105 bl[105] br[105] wl[224] vdd gnd cell_6t
Xbit_r225_c105 bl[105] br[105] wl[225] vdd gnd cell_6t
Xbit_r226_c105 bl[105] br[105] wl[226] vdd gnd cell_6t
Xbit_r227_c105 bl[105] br[105] wl[227] vdd gnd cell_6t
Xbit_r228_c105 bl[105] br[105] wl[228] vdd gnd cell_6t
Xbit_r229_c105 bl[105] br[105] wl[229] vdd gnd cell_6t
Xbit_r230_c105 bl[105] br[105] wl[230] vdd gnd cell_6t
Xbit_r231_c105 bl[105] br[105] wl[231] vdd gnd cell_6t
Xbit_r232_c105 bl[105] br[105] wl[232] vdd gnd cell_6t
Xbit_r233_c105 bl[105] br[105] wl[233] vdd gnd cell_6t
Xbit_r234_c105 bl[105] br[105] wl[234] vdd gnd cell_6t
Xbit_r235_c105 bl[105] br[105] wl[235] vdd gnd cell_6t
Xbit_r236_c105 bl[105] br[105] wl[236] vdd gnd cell_6t
Xbit_r237_c105 bl[105] br[105] wl[237] vdd gnd cell_6t
Xbit_r238_c105 bl[105] br[105] wl[238] vdd gnd cell_6t
Xbit_r239_c105 bl[105] br[105] wl[239] vdd gnd cell_6t
Xbit_r240_c105 bl[105] br[105] wl[240] vdd gnd cell_6t
Xbit_r241_c105 bl[105] br[105] wl[241] vdd gnd cell_6t
Xbit_r242_c105 bl[105] br[105] wl[242] vdd gnd cell_6t
Xbit_r243_c105 bl[105] br[105] wl[243] vdd gnd cell_6t
Xbit_r244_c105 bl[105] br[105] wl[244] vdd gnd cell_6t
Xbit_r245_c105 bl[105] br[105] wl[245] vdd gnd cell_6t
Xbit_r246_c105 bl[105] br[105] wl[246] vdd gnd cell_6t
Xbit_r247_c105 bl[105] br[105] wl[247] vdd gnd cell_6t
Xbit_r248_c105 bl[105] br[105] wl[248] vdd gnd cell_6t
Xbit_r249_c105 bl[105] br[105] wl[249] vdd gnd cell_6t
Xbit_r250_c105 bl[105] br[105] wl[250] vdd gnd cell_6t
Xbit_r251_c105 bl[105] br[105] wl[251] vdd gnd cell_6t
Xbit_r252_c105 bl[105] br[105] wl[252] vdd gnd cell_6t
Xbit_r253_c105 bl[105] br[105] wl[253] vdd gnd cell_6t
Xbit_r254_c105 bl[105] br[105] wl[254] vdd gnd cell_6t
Xbit_r255_c105 bl[105] br[105] wl[255] vdd gnd cell_6t
Xbit_r0_c106 bl[106] br[106] wl[0] vdd gnd cell_6t
Xbit_r1_c106 bl[106] br[106] wl[1] vdd gnd cell_6t
Xbit_r2_c106 bl[106] br[106] wl[2] vdd gnd cell_6t
Xbit_r3_c106 bl[106] br[106] wl[3] vdd gnd cell_6t
Xbit_r4_c106 bl[106] br[106] wl[4] vdd gnd cell_6t
Xbit_r5_c106 bl[106] br[106] wl[5] vdd gnd cell_6t
Xbit_r6_c106 bl[106] br[106] wl[6] vdd gnd cell_6t
Xbit_r7_c106 bl[106] br[106] wl[7] vdd gnd cell_6t
Xbit_r8_c106 bl[106] br[106] wl[8] vdd gnd cell_6t
Xbit_r9_c106 bl[106] br[106] wl[9] vdd gnd cell_6t
Xbit_r10_c106 bl[106] br[106] wl[10] vdd gnd cell_6t
Xbit_r11_c106 bl[106] br[106] wl[11] vdd gnd cell_6t
Xbit_r12_c106 bl[106] br[106] wl[12] vdd gnd cell_6t
Xbit_r13_c106 bl[106] br[106] wl[13] vdd gnd cell_6t
Xbit_r14_c106 bl[106] br[106] wl[14] vdd gnd cell_6t
Xbit_r15_c106 bl[106] br[106] wl[15] vdd gnd cell_6t
Xbit_r16_c106 bl[106] br[106] wl[16] vdd gnd cell_6t
Xbit_r17_c106 bl[106] br[106] wl[17] vdd gnd cell_6t
Xbit_r18_c106 bl[106] br[106] wl[18] vdd gnd cell_6t
Xbit_r19_c106 bl[106] br[106] wl[19] vdd gnd cell_6t
Xbit_r20_c106 bl[106] br[106] wl[20] vdd gnd cell_6t
Xbit_r21_c106 bl[106] br[106] wl[21] vdd gnd cell_6t
Xbit_r22_c106 bl[106] br[106] wl[22] vdd gnd cell_6t
Xbit_r23_c106 bl[106] br[106] wl[23] vdd gnd cell_6t
Xbit_r24_c106 bl[106] br[106] wl[24] vdd gnd cell_6t
Xbit_r25_c106 bl[106] br[106] wl[25] vdd gnd cell_6t
Xbit_r26_c106 bl[106] br[106] wl[26] vdd gnd cell_6t
Xbit_r27_c106 bl[106] br[106] wl[27] vdd gnd cell_6t
Xbit_r28_c106 bl[106] br[106] wl[28] vdd gnd cell_6t
Xbit_r29_c106 bl[106] br[106] wl[29] vdd gnd cell_6t
Xbit_r30_c106 bl[106] br[106] wl[30] vdd gnd cell_6t
Xbit_r31_c106 bl[106] br[106] wl[31] vdd gnd cell_6t
Xbit_r32_c106 bl[106] br[106] wl[32] vdd gnd cell_6t
Xbit_r33_c106 bl[106] br[106] wl[33] vdd gnd cell_6t
Xbit_r34_c106 bl[106] br[106] wl[34] vdd gnd cell_6t
Xbit_r35_c106 bl[106] br[106] wl[35] vdd gnd cell_6t
Xbit_r36_c106 bl[106] br[106] wl[36] vdd gnd cell_6t
Xbit_r37_c106 bl[106] br[106] wl[37] vdd gnd cell_6t
Xbit_r38_c106 bl[106] br[106] wl[38] vdd gnd cell_6t
Xbit_r39_c106 bl[106] br[106] wl[39] vdd gnd cell_6t
Xbit_r40_c106 bl[106] br[106] wl[40] vdd gnd cell_6t
Xbit_r41_c106 bl[106] br[106] wl[41] vdd gnd cell_6t
Xbit_r42_c106 bl[106] br[106] wl[42] vdd gnd cell_6t
Xbit_r43_c106 bl[106] br[106] wl[43] vdd gnd cell_6t
Xbit_r44_c106 bl[106] br[106] wl[44] vdd gnd cell_6t
Xbit_r45_c106 bl[106] br[106] wl[45] vdd gnd cell_6t
Xbit_r46_c106 bl[106] br[106] wl[46] vdd gnd cell_6t
Xbit_r47_c106 bl[106] br[106] wl[47] vdd gnd cell_6t
Xbit_r48_c106 bl[106] br[106] wl[48] vdd gnd cell_6t
Xbit_r49_c106 bl[106] br[106] wl[49] vdd gnd cell_6t
Xbit_r50_c106 bl[106] br[106] wl[50] vdd gnd cell_6t
Xbit_r51_c106 bl[106] br[106] wl[51] vdd gnd cell_6t
Xbit_r52_c106 bl[106] br[106] wl[52] vdd gnd cell_6t
Xbit_r53_c106 bl[106] br[106] wl[53] vdd gnd cell_6t
Xbit_r54_c106 bl[106] br[106] wl[54] vdd gnd cell_6t
Xbit_r55_c106 bl[106] br[106] wl[55] vdd gnd cell_6t
Xbit_r56_c106 bl[106] br[106] wl[56] vdd gnd cell_6t
Xbit_r57_c106 bl[106] br[106] wl[57] vdd gnd cell_6t
Xbit_r58_c106 bl[106] br[106] wl[58] vdd gnd cell_6t
Xbit_r59_c106 bl[106] br[106] wl[59] vdd gnd cell_6t
Xbit_r60_c106 bl[106] br[106] wl[60] vdd gnd cell_6t
Xbit_r61_c106 bl[106] br[106] wl[61] vdd gnd cell_6t
Xbit_r62_c106 bl[106] br[106] wl[62] vdd gnd cell_6t
Xbit_r63_c106 bl[106] br[106] wl[63] vdd gnd cell_6t
Xbit_r64_c106 bl[106] br[106] wl[64] vdd gnd cell_6t
Xbit_r65_c106 bl[106] br[106] wl[65] vdd gnd cell_6t
Xbit_r66_c106 bl[106] br[106] wl[66] vdd gnd cell_6t
Xbit_r67_c106 bl[106] br[106] wl[67] vdd gnd cell_6t
Xbit_r68_c106 bl[106] br[106] wl[68] vdd gnd cell_6t
Xbit_r69_c106 bl[106] br[106] wl[69] vdd gnd cell_6t
Xbit_r70_c106 bl[106] br[106] wl[70] vdd gnd cell_6t
Xbit_r71_c106 bl[106] br[106] wl[71] vdd gnd cell_6t
Xbit_r72_c106 bl[106] br[106] wl[72] vdd gnd cell_6t
Xbit_r73_c106 bl[106] br[106] wl[73] vdd gnd cell_6t
Xbit_r74_c106 bl[106] br[106] wl[74] vdd gnd cell_6t
Xbit_r75_c106 bl[106] br[106] wl[75] vdd gnd cell_6t
Xbit_r76_c106 bl[106] br[106] wl[76] vdd gnd cell_6t
Xbit_r77_c106 bl[106] br[106] wl[77] vdd gnd cell_6t
Xbit_r78_c106 bl[106] br[106] wl[78] vdd gnd cell_6t
Xbit_r79_c106 bl[106] br[106] wl[79] vdd gnd cell_6t
Xbit_r80_c106 bl[106] br[106] wl[80] vdd gnd cell_6t
Xbit_r81_c106 bl[106] br[106] wl[81] vdd gnd cell_6t
Xbit_r82_c106 bl[106] br[106] wl[82] vdd gnd cell_6t
Xbit_r83_c106 bl[106] br[106] wl[83] vdd gnd cell_6t
Xbit_r84_c106 bl[106] br[106] wl[84] vdd gnd cell_6t
Xbit_r85_c106 bl[106] br[106] wl[85] vdd gnd cell_6t
Xbit_r86_c106 bl[106] br[106] wl[86] vdd gnd cell_6t
Xbit_r87_c106 bl[106] br[106] wl[87] vdd gnd cell_6t
Xbit_r88_c106 bl[106] br[106] wl[88] vdd gnd cell_6t
Xbit_r89_c106 bl[106] br[106] wl[89] vdd gnd cell_6t
Xbit_r90_c106 bl[106] br[106] wl[90] vdd gnd cell_6t
Xbit_r91_c106 bl[106] br[106] wl[91] vdd gnd cell_6t
Xbit_r92_c106 bl[106] br[106] wl[92] vdd gnd cell_6t
Xbit_r93_c106 bl[106] br[106] wl[93] vdd gnd cell_6t
Xbit_r94_c106 bl[106] br[106] wl[94] vdd gnd cell_6t
Xbit_r95_c106 bl[106] br[106] wl[95] vdd gnd cell_6t
Xbit_r96_c106 bl[106] br[106] wl[96] vdd gnd cell_6t
Xbit_r97_c106 bl[106] br[106] wl[97] vdd gnd cell_6t
Xbit_r98_c106 bl[106] br[106] wl[98] vdd gnd cell_6t
Xbit_r99_c106 bl[106] br[106] wl[99] vdd gnd cell_6t
Xbit_r100_c106 bl[106] br[106] wl[100] vdd gnd cell_6t
Xbit_r101_c106 bl[106] br[106] wl[101] vdd gnd cell_6t
Xbit_r102_c106 bl[106] br[106] wl[102] vdd gnd cell_6t
Xbit_r103_c106 bl[106] br[106] wl[103] vdd gnd cell_6t
Xbit_r104_c106 bl[106] br[106] wl[104] vdd gnd cell_6t
Xbit_r105_c106 bl[106] br[106] wl[105] vdd gnd cell_6t
Xbit_r106_c106 bl[106] br[106] wl[106] vdd gnd cell_6t
Xbit_r107_c106 bl[106] br[106] wl[107] vdd gnd cell_6t
Xbit_r108_c106 bl[106] br[106] wl[108] vdd gnd cell_6t
Xbit_r109_c106 bl[106] br[106] wl[109] vdd gnd cell_6t
Xbit_r110_c106 bl[106] br[106] wl[110] vdd gnd cell_6t
Xbit_r111_c106 bl[106] br[106] wl[111] vdd gnd cell_6t
Xbit_r112_c106 bl[106] br[106] wl[112] vdd gnd cell_6t
Xbit_r113_c106 bl[106] br[106] wl[113] vdd gnd cell_6t
Xbit_r114_c106 bl[106] br[106] wl[114] vdd gnd cell_6t
Xbit_r115_c106 bl[106] br[106] wl[115] vdd gnd cell_6t
Xbit_r116_c106 bl[106] br[106] wl[116] vdd gnd cell_6t
Xbit_r117_c106 bl[106] br[106] wl[117] vdd gnd cell_6t
Xbit_r118_c106 bl[106] br[106] wl[118] vdd gnd cell_6t
Xbit_r119_c106 bl[106] br[106] wl[119] vdd gnd cell_6t
Xbit_r120_c106 bl[106] br[106] wl[120] vdd gnd cell_6t
Xbit_r121_c106 bl[106] br[106] wl[121] vdd gnd cell_6t
Xbit_r122_c106 bl[106] br[106] wl[122] vdd gnd cell_6t
Xbit_r123_c106 bl[106] br[106] wl[123] vdd gnd cell_6t
Xbit_r124_c106 bl[106] br[106] wl[124] vdd gnd cell_6t
Xbit_r125_c106 bl[106] br[106] wl[125] vdd gnd cell_6t
Xbit_r126_c106 bl[106] br[106] wl[126] vdd gnd cell_6t
Xbit_r127_c106 bl[106] br[106] wl[127] vdd gnd cell_6t
Xbit_r128_c106 bl[106] br[106] wl[128] vdd gnd cell_6t
Xbit_r129_c106 bl[106] br[106] wl[129] vdd gnd cell_6t
Xbit_r130_c106 bl[106] br[106] wl[130] vdd gnd cell_6t
Xbit_r131_c106 bl[106] br[106] wl[131] vdd gnd cell_6t
Xbit_r132_c106 bl[106] br[106] wl[132] vdd gnd cell_6t
Xbit_r133_c106 bl[106] br[106] wl[133] vdd gnd cell_6t
Xbit_r134_c106 bl[106] br[106] wl[134] vdd gnd cell_6t
Xbit_r135_c106 bl[106] br[106] wl[135] vdd gnd cell_6t
Xbit_r136_c106 bl[106] br[106] wl[136] vdd gnd cell_6t
Xbit_r137_c106 bl[106] br[106] wl[137] vdd gnd cell_6t
Xbit_r138_c106 bl[106] br[106] wl[138] vdd gnd cell_6t
Xbit_r139_c106 bl[106] br[106] wl[139] vdd gnd cell_6t
Xbit_r140_c106 bl[106] br[106] wl[140] vdd gnd cell_6t
Xbit_r141_c106 bl[106] br[106] wl[141] vdd gnd cell_6t
Xbit_r142_c106 bl[106] br[106] wl[142] vdd gnd cell_6t
Xbit_r143_c106 bl[106] br[106] wl[143] vdd gnd cell_6t
Xbit_r144_c106 bl[106] br[106] wl[144] vdd gnd cell_6t
Xbit_r145_c106 bl[106] br[106] wl[145] vdd gnd cell_6t
Xbit_r146_c106 bl[106] br[106] wl[146] vdd gnd cell_6t
Xbit_r147_c106 bl[106] br[106] wl[147] vdd gnd cell_6t
Xbit_r148_c106 bl[106] br[106] wl[148] vdd gnd cell_6t
Xbit_r149_c106 bl[106] br[106] wl[149] vdd gnd cell_6t
Xbit_r150_c106 bl[106] br[106] wl[150] vdd gnd cell_6t
Xbit_r151_c106 bl[106] br[106] wl[151] vdd gnd cell_6t
Xbit_r152_c106 bl[106] br[106] wl[152] vdd gnd cell_6t
Xbit_r153_c106 bl[106] br[106] wl[153] vdd gnd cell_6t
Xbit_r154_c106 bl[106] br[106] wl[154] vdd gnd cell_6t
Xbit_r155_c106 bl[106] br[106] wl[155] vdd gnd cell_6t
Xbit_r156_c106 bl[106] br[106] wl[156] vdd gnd cell_6t
Xbit_r157_c106 bl[106] br[106] wl[157] vdd gnd cell_6t
Xbit_r158_c106 bl[106] br[106] wl[158] vdd gnd cell_6t
Xbit_r159_c106 bl[106] br[106] wl[159] vdd gnd cell_6t
Xbit_r160_c106 bl[106] br[106] wl[160] vdd gnd cell_6t
Xbit_r161_c106 bl[106] br[106] wl[161] vdd gnd cell_6t
Xbit_r162_c106 bl[106] br[106] wl[162] vdd gnd cell_6t
Xbit_r163_c106 bl[106] br[106] wl[163] vdd gnd cell_6t
Xbit_r164_c106 bl[106] br[106] wl[164] vdd gnd cell_6t
Xbit_r165_c106 bl[106] br[106] wl[165] vdd gnd cell_6t
Xbit_r166_c106 bl[106] br[106] wl[166] vdd gnd cell_6t
Xbit_r167_c106 bl[106] br[106] wl[167] vdd gnd cell_6t
Xbit_r168_c106 bl[106] br[106] wl[168] vdd gnd cell_6t
Xbit_r169_c106 bl[106] br[106] wl[169] vdd gnd cell_6t
Xbit_r170_c106 bl[106] br[106] wl[170] vdd gnd cell_6t
Xbit_r171_c106 bl[106] br[106] wl[171] vdd gnd cell_6t
Xbit_r172_c106 bl[106] br[106] wl[172] vdd gnd cell_6t
Xbit_r173_c106 bl[106] br[106] wl[173] vdd gnd cell_6t
Xbit_r174_c106 bl[106] br[106] wl[174] vdd gnd cell_6t
Xbit_r175_c106 bl[106] br[106] wl[175] vdd gnd cell_6t
Xbit_r176_c106 bl[106] br[106] wl[176] vdd gnd cell_6t
Xbit_r177_c106 bl[106] br[106] wl[177] vdd gnd cell_6t
Xbit_r178_c106 bl[106] br[106] wl[178] vdd gnd cell_6t
Xbit_r179_c106 bl[106] br[106] wl[179] vdd gnd cell_6t
Xbit_r180_c106 bl[106] br[106] wl[180] vdd gnd cell_6t
Xbit_r181_c106 bl[106] br[106] wl[181] vdd gnd cell_6t
Xbit_r182_c106 bl[106] br[106] wl[182] vdd gnd cell_6t
Xbit_r183_c106 bl[106] br[106] wl[183] vdd gnd cell_6t
Xbit_r184_c106 bl[106] br[106] wl[184] vdd gnd cell_6t
Xbit_r185_c106 bl[106] br[106] wl[185] vdd gnd cell_6t
Xbit_r186_c106 bl[106] br[106] wl[186] vdd gnd cell_6t
Xbit_r187_c106 bl[106] br[106] wl[187] vdd gnd cell_6t
Xbit_r188_c106 bl[106] br[106] wl[188] vdd gnd cell_6t
Xbit_r189_c106 bl[106] br[106] wl[189] vdd gnd cell_6t
Xbit_r190_c106 bl[106] br[106] wl[190] vdd gnd cell_6t
Xbit_r191_c106 bl[106] br[106] wl[191] vdd gnd cell_6t
Xbit_r192_c106 bl[106] br[106] wl[192] vdd gnd cell_6t
Xbit_r193_c106 bl[106] br[106] wl[193] vdd gnd cell_6t
Xbit_r194_c106 bl[106] br[106] wl[194] vdd gnd cell_6t
Xbit_r195_c106 bl[106] br[106] wl[195] vdd gnd cell_6t
Xbit_r196_c106 bl[106] br[106] wl[196] vdd gnd cell_6t
Xbit_r197_c106 bl[106] br[106] wl[197] vdd gnd cell_6t
Xbit_r198_c106 bl[106] br[106] wl[198] vdd gnd cell_6t
Xbit_r199_c106 bl[106] br[106] wl[199] vdd gnd cell_6t
Xbit_r200_c106 bl[106] br[106] wl[200] vdd gnd cell_6t
Xbit_r201_c106 bl[106] br[106] wl[201] vdd gnd cell_6t
Xbit_r202_c106 bl[106] br[106] wl[202] vdd gnd cell_6t
Xbit_r203_c106 bl[106] br[106] wl[203] vdd gnd cell_6t
Xbit_r204_c106 bl[106] br[106] wl[204] vdd gnd cell_6t
Xbit_r205_c106 bl[106] br[106] wl[205] vdd gnd cell_6t
Xbit_r206_c106 bl[106] br[106] wl[206] vdd gnd cell_6t
Xbit_r207_c106 bl[106] br[106] wl[207] vdd gnd cell_6t
Xbit_r208_c106 bl[106] br[106] wl[208] vdd gnd cell_6t
Xbit_r209_c106 bl[106] br[106] wl[209] vdd gnd cell_6t
Xbit_r210_c106 bl[106] br[106] wl[210] vdd gnd cell_6t
Xbit_r211_c106 bl[106] br[106] wl[211] vdd gnd cell_6t
Xbit_r212_c106 bl[106] br[106] wl[212] vdd gnd cell_6t
Xbit_r213_c106 bl[106] br[106] wl[213] vdd gnd cell_6t
Xbit_r214_c106 bl[106] br[106] wl[214] vdd gnd cell_6t
Xbit_r215_c106 bl[106] br[106] wl[215] vdd gnd cell_6t
Xbit_r216_c106 bl[106] br[106] wl[216] vdd gnd cell_6t
Xbit_r217_c106 bl[106] br[106] wl[217] vdd gnd cell_6t
Xbit_r218_c106 bl[106] br[106] wl[218] vdd gnd cell_6t
Xbit_r219_c106 bl[106] br[106] wl[219] vdd gnd cell_6t
Xbit_r220_c106 bl[106] br[106] wl[220] vdd gnd cell_6t
Xbit_r221_c106 bl[106] br[106] wl[221] vdd gnd cell_6t
Xbit_r222_c106 bl[106] br[106] wl[222] vdd gnd cell_6t
Xbit_r223_c106 bl[106] br[106] wl[223] vdd gnd cell_6t
Xbit_r224_c106 bl[106] br[106] wl[224] vdd gnd cell_6t
Xbit_r225_c106 bl[106] br[106] wl[225] vdd gnd cell_6t
Xbit_r226_c106 bl[106] br[106] wl[226] vdd gnd cell_6t
Xbit_r227_c106 bl[106] br[106] wl[227] vdd gnd cell_6t
Xbit_r228_c106 bl[106] br[106] wl[228] vdd gnd cell_6t
Xbit_r229_c106 bl[106] br[106] wl[229] vdd gnd cell_6t
Xbit_r230_c106 bl[106] br[106] wl[230] vdd gnd cell_6t
Xbit_r231_c106 bl[106] br[106] wl[231] vdd gnd cell_6t
Xbit_r232_c106 bl[106] br[106] wl[232] vdd gnd cell_6t
Xbit_r233_c106 bl[106] br[106] wl[233] vdd gnd cell_6t
Xbit_r234_c106 bl[106] br[106] wl[234] vdd gnd cell_6t
Xbit_r235_c106 bl[106] br[106] wl[235] vdd gnd cell_6t
Xbit_r236_c106 bl[106] br[106] wl[236] vdd gnd cell_6t
Xbit_r237_c106 bl[106] br[106] wl[237] vdd gnd cell_6t
Xbit_r238_c106 bl[106] br[106] wl[238] vdd gnd cell_6t
Xbit_r239_c106 bl[106] br[106] wl[239] vdd gnd cell_6t
Xbit_r240_c106 bl[106] br[106] wl[240] vdd gnd cell_6t
Xbit_r241_c106 bl[106] br[106] wl[241] vdd gnd cell_6t
Xbit_r242_c106 bl[106] br[106] wl[242] vdd gnd cell_6t
Xbit_r243_c106 bl[106] br[106] wl[243] vdd gnd cell_6t
Xbit_r244_c106 bl[106] br[106] wl[244] vdd gnd cell_6t
Xbit_r245_c106 bl[106] br[106] wl[245] vdd gnd cell_6t
Xbit_r246_c106 bl[106] br[106] wl[246] vdd gnd cell_6t
Xbit_r247_c106 bl[106] br[106] wl[247] vdd gnd cell_6t
Xbit_r248_c106 bl[106] br[106] wl[248] vdd gnd cell_6t
Xbit_r249_c106 bl[106] br[106] wl[249] vdd gnd cell_6t
Xbit_r250_c106 bl[106] br[106] wl[250] vdd gnd cell_6t
Xbit_r251_c106 bl[106] br[106] wl[251] vdd gnd cell_6t
Xbit_r252_c106 bl[106] br[106] wl[252] vdd gnd cell_6t
Xbit_r253_c106 bl[106] br[106] wl[253] vdd gnd cell_6t
Xbit_r254_c106 bl[106] br[106] wl[254] vdd gnd cell_6t
Xbit_r255_c106 bl[106] br[106] wl[255] vdd gnd cell_6t
Xbit_r0_c107 bl[107] br[107] wl[0] vdd gnd cell_6t
Xbit_r1_c107 bl[107] br[107] wl[1] vdd gnd cell_6t
Xbit_r2_c107 bl[107] br[107] wl[2] vdd gnd cell_6t
Xbit_r3_c107 bl[107] br[107] wl[3] vdd gnd cell_6t
Xbit_r4_c107 bl[107] br[107] wl[4] vdd gnd cell_6t
Xbit_r5_c107 bl[107] br[107] wl[5] vdd gnd cell_6t
Xbit_r6_c107 bl[107] br[107] wl[6] vdd gnd cell_6t
Xbit_r7_c107 bl[107] br[107] wl[7] vdd gnd cell_6t
Xbit_r8_c107 bl[107] br[107] wl[8] vdd gnd cell_6t
Xbit_r9_c107 bl[107] br[107] wl[9] vdd gnd cell_6t
Xbit_r10_c107 bl[107] br[107] wl[10] vdd gnd cell_6t
Xbit_r11_c107 bl[107] br[107] wl[11] vdd gnd cell_6t
Xbit_r12_c107 bl[107] br[107] wl[12] vdd gnd cell_6t
Xbit_r13_c107 bl[107] br[107] wl[13] vdd gnd cell_6t
Xbit_r14_c107 bl[107] br[107] wl[14] vdd gnd cell_6t
Xbit_r15_c107 bl[107] br[107] wl[15] vdd gnd cell_6t
Xbit_r16_c107 bl[107] br[107] wl[16] vdd gnd cell_6t
Xbit_r17_c107 bl[107] br[107] wl[17] vdd gnd cell_6t
Xbit_r18_c107 bl[107] br[107] wl[18] vdd gnd cell_6t
Xbit_r19_c107 bl[107] br[107] wl[19] vdd gnd cell_6t
Xbit_r20_c107 bl[107] br[107] wl[20] vdd gnd cell_6t
Xbit_r21_c107 bl[107] br[107] wl[21] vdd gnd cell_6t
Xbit_r22_c107 bl[107] br[107] wl[22] vdd gnd cell_6t
Xbit_r23_c107 bl[107] br[107] wl[23] vdd gnd cell_6t
Xbit_r24_c107 bl[107] br[107] wl[24] vdd gnd cell_6t
Xbit_r25_c107 bl[107] br[107] wl[25] vdd gnd cell_6t
Xbit_r26_c107 bl[107] br[107] wl[26] vdd gnd cell_6t
Xbit_r27_c107 bl[107] br[107] wl[27] vdd gnd cell_6t
Xbit_r28_c107 bl[107] br[107] wl[28] vdd gnd cell_6t
Xbit_r29_c107 bl[107] br[107] wl[29] vdd gnd cell_6t
Xbit_r30_c107 bl[107] br[107] wl[30] vdd gnd cell_6t
Xbit_r31_c107 bl[107] br[107] wl[31] vdd gnd cell_6t
Xbit_r32_c107 bl[107] br[107] wl[32] vdd gnd cell_6t
Xbit_r33_c107 bl[107] br[107] wl[33] vdd gnd cell_6t
Xbit_r34_c107 bl[107] br[107] wl[34] vdd gnd cell_6t
Xbit_r35_c107 bl[107] br[107] wl[35] vdd gnd cell_6t
Xbit_r36_c107 bl[107] br[107] wl[36] vdd gnd cell_6t
Xbit_r37_c107 bl[107] br[107] wl[37] vdd gnd cell_6t
Xbit_r38_c107 bl[107] br[107] wl[38] vdd gnd cell_6t
Xbit_r39_c107 bl[107] br[107] wl[39] vdd gnd cell_6t
Xbit_r40_c107 bl[107] br[107] wl[40] vdd gnd cell_6t
Xbit_r41_c107 bl[107] br[107] wl[41] vdd gnd cell_6t
Xbit_r42_c107 bl[107] br[107] wl[42] vdd gnd cell_6t
Xbit_r43_c107 bl[107] br[107] wl[43] vdd gnd cell_6t
Xbit_r44_c107 bl[107] br[107] wl[44] vdd gnd cell_6t
Xbit_r45_c107 bl[107] br[107] wl[45] vdd gnd cell_6t
Xbit_r46_c107 bl[107] br[107] wl[46] vdd gnd cell_6t
Xbit_r47_c107 bl[107] br[107] wl[47] vdd gnd cell_6t
Xbit_r48_c107 bl[107] br[107] wl[48] vdd gnd cell_6t
Xbit_r49_c107 bl[107] br[107] wl[49] vdd gnd cell_6t
Xbit_r50_c107 bl[107] br[107] wl[50] vdd gnd cell_6t
Xbit_r51_c107 bl[107] br[107] wl[51] vdd gnd cell_6t
Xbit_r52_c107 bl[107] br[107] wl[52] vdd gnd cell_6t
Xbit_r53_c107 bl[107] br[107] wl[53] vdd gnd cell_6t
Xbit_r54_c107 bl[107] br[107] wl[54] vdd gnd cell_6t
Xbit_r55_c107 bl[107] br[107] wl[55] vdd gnd cell_6t
Xbit_r56_c107 bl[107] br[107] wl[56] vdd gnd cell_6t
Xbit_r57_c107 bl[107] br[107] wl[57] vdd gnd cell_6t
Xbit_r58_c107 bl[107] br[107] wl[58] vdd gnd cell_6t
Xbit_r59_c107 bl[107] br[107] wl[59] vdd gnd cell_6t
Xbit_r60_c107 bl[107] br[107] wl[60] vdd gnd cell_6t
Xbit_r61_c107 bl[107] br[107] wl[61] vdd gnd cell_6t
Xbit_r62_c107 bl[107] br[107] wl[62] vdd gnd cell_6t
Xbit_r63_c107 bl[107] br[107] wl[63] vdd gnd cell_6t
Xbit_r64_c107 bl[107] br[107] wl[64] vdd gnd cell_6t
Xbit_r65_c107 bl[107] br[107] wl[65] vdd gnd cell_6t
Xbit_r66_c107 bl[107] br[107] wl[66] vdd gnd cell_6t
Xbit_r67_c107 bl[107] br[107] wl[67] vdd gnd cell_6t
Xbit_r68_c107 bl[107] br[107] wl[68] vdd gnd cell_6t
Xbit_r69_c107 bl[107] br[107] wl[69] vdd gnd cell_6t
Xbit_r70_c107 bl[107] br[107] wl[70] vdd gnd cell_6t
Xbit_r71_c107 bl[107] br[107] wl[71] vdd gnd cell_6t
Xbit_r72_c107 bl[107] br[107] wl[72] vdd gnd cell_6t
Xbit_r73_c107 bl[107] br[107] wl[73] vdd gnd cell_6t
Xbit_r74_c107 bl[107] br[107] wl[74] vdd gnd cell_6t
Xbit_r75_c107 bl[107] br[107] wl[75] vdd gnd cell_6t
Xbit_r76_c107 bl[107] br[107] wl[76] vdd gnd cell_6t
Xbit_r77_c107 bl[107] br[107] wl[77] vdd gnd cell_6t
Xbit_r78_c107 bl[107] br[107] wl[78] vdd gnd cell_6t
Xbit_r79_c107 bl[107] br[107] wl[79] vdd gnd cell_6t
Xbit_r80_c107 bl[107] br[107] wl[80] vdd gnd cell_6t
Xbit_r81_c107 bl[107] br[107] wl[81] vdd gnd cell_6t
Xbit_r82_c107 bl[107] br[107] wl[82] vdd gnd cell_6t
Xbit_r83_c107 bl[107] br[107] wl[83] vdd gnd cell_6t
Xbit_r84_c107 bl[107] br[107] wl[84] vdd gnd cell_6t
Xbit_r85_c107 bl[107] br[107] wl[85] vdd gnd cell_6t
Xbit_r86_c107 bl[107] br[107] wl[86] vdd gnd cell_6t
Xbit_r87_c107 bl[107] br[107] wl[87] vdd gnd cell_6t
Xbit_r88_c107 bl[107] br[107] wl[88] vdd gnd cell_6t
Xbit_r89_c107 bl[107] br[107] wl[89] vdd gnd cell_6t
Xbit_r90_c107 bl[107] br[107] wl[90] vdd gnd cell_6t
Xbit_r91_c107 bl[107] br[107] wl[91] vdd gnd cell_6t
Xbit_r92_c107 bl[107] br[107] wl[92] vdd gnd cell_6t
Xbit_r93_c107 bl[107] br[107] wl[93] vdd gnd cell_6t
Xbit_r94_c107 bl[107] br[107] wl[94] vdd gnd cell_6t
Xbit_r95_c107 bl[107] br[107] wl[95] vdd gnd cell_6t
Xbit_r96_c107 bl[107] br[107] wl[96] vdd gnd cell_6t
Xbit_r97_c107 bl[107] br[107] wl[97] vdd gnd cell_6t
Xbit_r98_c107 bl[107] br[107] wl[98] vdd gnd cell_6t
Xbit_r99_c107 bl[107] br[107] wl[99] vdd gnd cell_6t
Xbit_r100_c107 bl[107] br[107] wl[100] vdd gnd cell_6t
Xbit_r101_c107 bl[107] br[107] wl[101] vdd gnd cell_6t
Xbit_r102_c107 bl[107] br[107] wl[102] vdd gnd cell_6t
Xbit_r103_c107 bl[107] br[107] wl[103] vdd gnd cell_6t
Xbit_r104_c107 bl[107] br[107] wl[104] vdd gnd cell_6t
Xbit_r105_c107 bl[107] br[107] wl[105] vdd gnd cell_6t
Xbit_r106_c107 bl[107] br[107] wl[106] vdd gnd cell_6t
Xbit_r107_c107 bl[107] br[107] wl[107] vdd gnd cell_6t
Xbit_r108_c107 bl[107] br[107] wl[108] vdd gnd cell_6t
Xbit_r109_c107 bl[107] br[107] wl[109] vdd gnd cell_6t
Xbit_r110_c107 bl[107] br[107] wl[110] vdd gnd cell_6t
Xbit_r111_c107 bl[107] br[107] wl[111] vdd gnd cell_6t
Xbit_r112_c107 bl[107] br[107] wl[112] vdd gnd cell_6t
Xbit_r113_c107 bl[107] br[107] wl[113] vdd gnd cell_6t
Xbit_r114_c107 bl[107] br[107] wl[114] vdd gnd cell_6t
Xbit_r115_c107 bl[107] br[107] wl[115] vdd gnd cell_6t
Xbit_r116_c107 bl[107] br[107] wl[116] vdd gnd cell_6t
Xbit_r117_c107 bl[107] br[107] wl[117] vdd gnd cell_6t
Xbit_r118_c107 bl[107] br[107] wl[118] vdd gnd cell_6t
Xbit_r119_c107 bl[107] br[107] wl[119] vdd gnd cell_6t
Xbit_r120_c107 bl[107] br[107] wl[120] vdd gnd cell_6t
Xbit_r121_c107 bl[107] br[107] wl[121] vdd gnd cell_6t
Xbit_r122_c107 bl[107] br[107] wl[122] vdd gnd cell_6t
Xbit_r123_c107 bl[107] br[107] wl[123] vdd gnd cell_6t
Xbit_r124_c107 bl[107] br[107] wl[124] vdd gnd cell_6t
Xbit_r125_c107 bl[107] br[107] wl[125] vdd gnd cell_6t
Xbit_r126_c107 bl[107] br[107] wl[126] vdd gnd cell_6t
Xbit_r127_c107 bl[107] br[107] wl[127] vdd gnd cell_6t
Xbit_r128_c107 bl[107] br[107] wl[128] vdd gnd cell_6t
Xbit_r129_c107 bl[107] br[107] wl[129] vdd gnd cell_6t
Xbit_r130_c107 bl[107] br[107] wl[130] vdd gnd cell_6t
Xbit_r131_c107 bl[107] br[107] wl[131] vdd gnd cell_6t
Xbit_r132_c107 bl[107] br[107] wl[132] vdd gnd cell_6t
Xbit_r133_c107 bl[107] br[107] wl[133] vdd gnd cell_6t
Xbit_r134_c107 bl[107] br[107] wl[134] vdd gnd cell_6t
Xbit_r135_c107 bl[107] br[107] wl[135] vdd gnd cell_6t
Xbit_r136_c107 bl[107] br[107] wl[136] vdd gnd cell_6t
Xbit_r137_c107 bl[107] br[107] wl[137] vdd gnd cell_6t
Xbit_r138_c107 bl[107] br[107] wl[138] vdd gnd cell_6t
Xbit_r139_c107 bl[107] br[107] wl[139] vdd gnd cell_6t
Xbit_r140_c107 bl[107] br[107] wl[140] vdd gnd cell_6t
Xbit_r141_c107 bl[107] br[107] wl[141] vdd gnd cell_6t
Xbit_r142_c107 bl[107] br[107] wl[142] vdd gnd cell_6t
Xbit_r143_c107 bl[107] br[107] wl[143] vdd gnd cell_6t
Xbit_r144_c107 bl[107] br[107] wl[144] vdd gnd cell_6t
Xbit_r145_c107 bl[107] br[107] wl[145] vdd gnd cell_6t
Xbit_r146_c107 bl[107] br[107] wl[146] vdd gnd cell_6t
Xbit_r147_c107 bl[107] br[107] wl[147] vdd gnd cell_6t
Xbit_r148_c107 bl[107] br[107] wl[148] vdd gnd cell_6t
Xbit_r149_c107 bl[107] br[107] wl[149] vdd gnd cell_6t
Xbit_r150_c107 bl[107] br[107] wl[150] vdd gnd cell_6t
Xbit_r151_c107 bl[107] br[107] wl[151] vdd gnd cell_6t
Xbit_r152_c107 bl[107] br[107] wl[152] vdd gnd cell_6t
Xbit_r153_c107 bl[107] br[107] wl[153] vdd gnd cell_6t
Xbit_r154_c107 bl[107] br[107] wl[154] vdd gnd cell_6t
Xbit_r155_c107 bl[107] br[107] wl[155] vdd gnd cell_6t
Xbit_r156_c107 bl[107] br[107] wl[156] vdd gnd cell_6t
Xbit_r157_c107 bl[107] br[107] wl[157] vdd gnd cell_6t
Xbit_r158_c107 bl[107] br[107] wl[158] vdd gnd cell_6t
Xbit_r159_c107 bl[107] br[107] wl[159] vdd gnd cell_6t
Xbit_r160_c107 bl[107] br[107] wl[160] vdd gnd cell_6t
Xbit_r161_c107 bl[107] br[107] wl[161] vdd gnd cell_6t
Xbit_r162_c107 bl[107] br[107] wl[162] vdd gnd cell_6t
Xbit_r163_c107 bl[107] br[107] wl[163] vdd gnd cell_6t
Xbit_r164_c107 bl[107] br[107] wl[164] vdd gnd cell_6t
Xbit_r165_c107 bl[107] br[107] wl[165] vdd gnd cell_6t
Xbit_r166_c107 bl[107] br[107] wl[166] vdd gnd cell_6t
Xbit_r167_c107 bl[107] br[107] wl[167] vdd gnd cell_6t
Xbit_r168_c107 bl[107] br[107] wl[168] vdd gnd cell_6t
Xbit_r169_c107 bl[107] br[107] wl[169] vdd gnd cell_6t
Xbit_r170_c107 bl[107] br[107] wl[170] vdd gnd cell_6t
Xbit_r171_c107 bl[107] br[107] wl[171] vdd gnd cell_6t
Xbit_r172_c107 bl[107] br[107] wl[172] vdd gnd cell_6t
Xbit_r173_c107 bl[107] br[107] wl[173] vdd gnd cell_6t
Xbit_r174_c107 bl[107] br[107] wl[174] vdd gnd cell_6t
Xbit_r175_c107 bl[107] br[107] wl[175] vdd gnd cell_6t
Xbit_r176_c107 bl[107] br[107] wl[176] vdd gnd cell_6t
Xbit_r177_c107 bl[107] br[107] wl[177] vdd gnd cell_6t
Xbit_r178_c107 bl[107] br[107] wl[178] vdd gnd cell_6t
Xbit_r179_c107 bl[107] br[107] wl[179] vdd gnd cell_6t
Xbit_r180_c107 bl[107] br[107] wl[180] vdd gnd cell_6t
Xbit_r181_c107 bl[107] br[107] wl[181] vdd gnd cell_6t
Xbit_r182_c107 bl[107] br[107] wl[182] vdd gnd cell_6t
Xbit_r183_c107 bl[107] br[107] wl[183] vdd gnd cell_6t
Xbit_r184_c107 bl[107] br[107] wl[184] vdd gnd cell_6t
Xbit_r185_c107 bl[107] br[107] wl[185] vdd gnd cell_6t
Xbit_r186_c107 bl[107] br[107] wl[186] vdd gnd cell_6t
Xbit_r187_c107 bl[107] br[107] wl[187] vdd gnd cell_6t
Xbit_r188_c107 bl[107] br[107] wl[188] vdd gnd cell_6t
Xbit_r189_c107 bl[107] br[107] wl[189] vdd gnd cell_6t
Xbit_r190_c107 bl[107] br[107] wl[190] vdd gnd cell_6t
Xbit_r191_c107 bl[107] br[107] wl[191] vdd gnd cell_6t
Xbit_r192_c107 bl[107] br[107] wl[192] vdd gnd cell_6t
Xbit_r193_c107 bl[107] br[107] wl[193] vdd gnd cell_6t
Xbit_r194_c107 bl[107] br[107] wl[194] vdd gnd cell_6t
Xbit_r195_c107 bl[107] br[107] wl[195] vdd gnd cell_6t
Xbit_r196_c107 bl[107] br[107] wl[196] vdd gnd cell_6t
Xbit_r197_c107 bl[107] br[107] wl[197] vdd gnd cell_6t
Xbit_r198_c107 bl[107] br[107] wl[198] vdd gnd cell_6t
Xbit_r199_c107 bl[107] br[107] wl[199] vdd gnd cell_6t
Xbit_r200_c107 bl[107] br[107] wl[200] vdd gnd cell_6t
Xbit_r201_c107 bl[107] br[107] wl[201] vdd gnd cell_6t
Xbit_r202_c107 bl[107] br[107] wl[202] vdd gnd cell_6t
Xbit_r203_c107 bl[107] br[107] wl[203] vdd gnd cell_6t
Xbit_r204_c107 bl[107] br[107] wl[204] vdd gnd cell_6t
Xbit_r205_c107 bl[107] br[107] wl[205] vdd gnd cell_6t
Xbit_r206_c107 bl[107] br[107] wl[206] vdd gnd cell_6t
Xbit_r207_c107 bl[107] br[107] wl[207] vdd gnd cell_6t
Xbit_r208_c107 bl[107] br[107] wl[208] vdd gnd cell_6t
Xbit_r209_c107 bl[107] br[107] wl[209] vdd gnd cell_6t
Xbit_r210_c107 bl[107] br[107] wl[210] vdd gnd cell_6t
Xbit_r211_c107 bl[107] br[107] wl[211] vdd gnd cell_6t
Xbit_r212_c107 bl[107] br[107] wl[212] vdd gnd cell_6t
Xbit_r213_c107 bl[107] br[107] wl[213] vdd gnd cell_6t
Xbit_r214_c107 bl[107] br[107] wl[214] vdd gnd cell_6t
Xbit_r215_c107 bl[107] br[107] wl[215] vdd gnd cell_6t
Xbit_r216_c107 bl[107] br[107] wl[216] vdd gnd cell_6t
Xbit_r217_c107 bl[107] br[107] wl[217] vdd gnd cell_6t
Xbit_r218_c107 bl[107] br[107] wl[218] vdd gnd cell_6t
Xbit_r219_c107 bl[107] br[107] wl[219] vdd gnd cell_6t
Xbit_r220_c107 bl[107] br[107] wl[220] vdd gnd cell_6t
Xbit_r221_c107 bl[107] br[107] wl[221] vdd gnd cell_6t
Xbit_r222_c107 bl[107] br[107] wl[222] vdd gnd cell_6t
Xbit_r223_c107 bl[107] br[107] wl[223] vdd gnd cell_6t
Xbit_r224_c107 bl[107] br[107] wl[224] vdd gnd cell_6t
Xbit_r225_c107 bl[107] br[107] wl[225] vdd gnd cell_6t
Xbit_r226_c107 bl[107] br[107] wl[226] vdd gnd cell_6t
Xbit_r227_c107 bl[107] br[107] wl[227] vdd gnd cell_6t
Xbit_r228_c107 bl[107] br[107] wl[228] vdd gnd cell_6t
Xbit_r229_c107 bl[107] br[107] wl[229] vdd gnd cell_6t
Xbit_r230_c107 bl[107] br[107] wl[230] vdd gnd cell_6t
Xbit_r231_c107 bl[107] br[107] wl[231] vdd gnd cell_6t
Xbit_r232_c107 bl[107] br[107] wl[232] vdd gnd cell_6t
Xbit_r233_c107 bl[107] br[107] wl[233] vdd gnd cell_6t
Xbit_r234_c107 bl[107] br[107] wl[234] vdd gnd cell_6t
Xbit_r235_c107 bl[107] br[107] wl[235] vdd gnd cell_6t
Xbit_r236_c107 bl[107] br[107] wl[236] vdd gnd cell_6t
Xbit_r237_c107 bl[107] br[107] wl[237] vdd gnd cell_6t
Xbit_r238_c107 bl[107] br[107] wl[238] vdd gnd cell_6t
Xbit_r239_c107 bl[107] br[107] wl[239] vdd gnd cell_6t
Xbit_r240_c107 bl[107] br[107] wl[240] vdd gnd cell_6t
Xbit_r241_c107 bl[107] br[107] wl[241] vdd gnd cell_6t
Xbit_r242_c107 bl[107] br[107] wl[242] vdd gnd cell_6t
Xbit_r243_c107 bl[107] br[107] wl[243] vdd gnd cell_6t
Xbit_r244_c107 bl[107] br[107] wl[244] vdd gnd cell_6t
Xbit_r245_c107 bl[107] br[107] wl[245] vdd gnd cell_6t
Xbit_r246_c107 bl[107] br[107] wl[246] vdd gnd cell_6t
Xbit_r247_c107 bl[107] br[107] wl[247] vdd gnd cell_6t
Xbit_r248_c107 bl[107] br[107] wl[248] vdd gnd cell_6t
Xbit_r249_c107 bl[107] br[107] wl[249] vdd gnd cell_6t
Xbit_r250_c107 bl[107] br[107] wl[250] vdd gnd cell_6t
Xbit_r251_c107 bl[107] br[107] wl[251] vdd gnd cell_6t
Xbit_r252_c107 bl[107] br[107] wl[252] vdd gnd cell_6t
Xbit_r253_c107 bl[107] br[107] wl[253] vdd gnd cell_6t
Xbit_r254_c107 bl[107] br[107] wl[254] vdd gnd cell_6t
Xbit_r255_c107 bl[107] br[107] wl[255] vdd gnd cell_6t
Xbit_r0_c108 bl[108] br[108] wl[0] vdd gnd cell_6t
Xbit_r1_c108 bl[108] br[108] wl[1] vdd gnd cell_6t
Xbit_r2_c108 bl[108] br[108] wl[2] vdd gnd cell_6t
Xbit_r3_c108 bl[108] br[108] wl[3] vdd gnd cell_6t
Xbit_r4_c108 bl[108] br[108] wl[4] vdd gnd cell_6t
Xbit_r5_c108 bl[108] br[108] wl[5] vdd gnd cell_6t
Xbit_r6_c108 bl[108] br[108] wl[6] vdd gnd cell_6t
Xbit_r7_c108 bl[108] br[108] wl[7] vdd gnd cell_6t
Xbit_r8_c108 bl[108] br[108] wl[8] vdd gnd cell_6t
Xbit_r9_c108 bl[108] br[108] wl[9] vdd gnd cell_6t
Xbit_r10_c108 bl[108] br[108] wl[10] vdd gnd cell_6t
Xbit_r11_c108 bl[108] br[108] wl[11] vdd gnd cell_6t
Xbit_r12_c108 bl[108] br[108] wl[12] vdd gnd cell_6t
Xbit_r13_c108 bl[108] br[108] wl[13] vdd gnd cell_6t
Xbit_r14_c108 bl[108] br[108] wl[14] vdd gnd cell_6t
Xbit_r15_c108 bl[108] br[108] wl[15] vdd gnd cell_6t
Xbit_r16_c108 bl[108] br[108] wl[16] vdd gnd cell_6t
Xbit_r17_c108 bl[108] br[108] wl[17] vdd gnd cell_6t
Xbit_r18_c108 bl[108] br[108] wl[18] vdd gnd cell_6t
Xbit_r19_c108 bl[108] br[108] wl[19] vdd gnd cell_6t
Xbit_r20_c108 bl[108] br[108] wl[20] vdd gnd cell_6t
Xbit_r21_c108 bl[108] br[108] wl[21] vdd gnd cell_6t
Xbit_r22_c108 bl[108] br[108] wl[22] vdd gnd cell_6t
Xbit_r23_c108 bl[108] br[108] wl[23] vdd gnd cell_6t
Xbit_r24_c108 bl[108] br[108] wl[24] vdd gnd cell_6t
Xbit_r25_c108 bl[108] br[108] wl[25] vdd gnd cell_6t
Xbit_r26_c108 bl[108] br[108] wl[26] vdd gnd cell_6t
Xbit_r27_c108 bl[108] br[108] wl[27] vdd gnd cell_6t
Xbit_r28_c108 bl[108] br[108] wl[28] vdd gnd cell_6t
Xbit_r29_c108 bl[108] br[108] wl[29] vdd gnd cell_6t
Xbit_r30_c108 bl[108] br[108] wl[30] vdd gnd cell_6t
Xbit_r31_c108 bl[108] br[108] wl[31] vdd gnd cell_6t
Xbit_r32_c108 bl[108] br[108] wl[32] vdd gnd cell_6t
Xbit_r33_c108 bl[108] br[108] wl[33] vdd gnd cell_6t
Xbit_r34_c108 bl[108] br[108] wl[34] vdd gnd cell_6t
Xbit_r35_c108 bl[108] br[108] wl[35] vdd gnd cell_6t
Xbit_r36_c108 bl[108] br[108] wl[36] vdd gnd cell_6t
Xbit_r37_c108 bl[108] br[108] wl[37] vdd gnd cell_6t
Xbit_r38_c108 bl[108] br[108] wl[38] vdd gnd cell_6t
Xbit_r39_c108 bl[108] br[108] wl[39] vdd gnd cell_6t
Xbit_r40_c108 bl[108] br[108] wl[40] vdd gnd cell_6t
Xbit_r41_c108 bl[108] br[108] wl[41] vdd gnd cell_6t
Xbit_r42_c108 bl[108] br[108] wl[42] vdd gnd cell_6t
Xbit_r43_c108 bl[108] br[108] wl[43] vdd gnd cell_6t
Xbit_r44_c108 bl[108] br[108] wl[44] vdd gnd cell_6t
Xbit_r45_c108 bl[108] br[108] wl[45] vdd gnd cell_6t
Xbit_r46_c108 bl[108] br[108] wl[46] vdd gnd cell_6t
Xbit_r47_c108 bl[108] br[108] wl[47] vdd gnd cell_6t
Xbit_r48_c108 bl[108] br[108] wl[48] vdd gnd cell_6t
Xbit_r49_c108 bl[108] br[108] wl[49] vdd gnd cell_6t
Xbit_r50_c108 bl[108] br[108] wl[50] vdd gnd cell_6t
Xbit_r51_c108 bl[108] br[108] wl[51] vdd gnd cell_6t
Xbit_r52_c108 bl[108] br[108] wl[52] vdd gnd cell_6t
Xbit_r53_c108 bl[108] br[108] wl[53] vdd gnd cell_6t
Xbit_r54_c108 bl[108] br[108] wl[54] vdd gnd cell_6t
Xbit_r55_c108 bl[108] br[108] wl[55] vdd gnd cell_6t
Xbit_r56_c108 bl[108] br[108] wl[56] vdd gnd cell_6t
Xbit_r57_c108 bl[108] br[108] wl[57] vdd gnd cell_6t
Xbit_r58_c108 bl[108] br[108] wl[58] vdd gnd cell_6t
Xbit_r59_c108 bl[108] br[108] wl[59] vdd gnd cell_6t
Xbit_r60_c108 bl[108] br[108] wl[60] vdd gnd cell_6t
Xbit_r61_c108 bl[108] br[108] wl[61] vdd gnd cell_6t
Xbit_r62_c108 bl[108] br[108] wl[62] vdd gnd cell_6t
Xbit_r63_c108 bl[108] br[108] wl[63] vdd gnd cell_6t
Xbit_r64_c108 bl[108] br[108] wl[64] vdd gnd cell_6t
Xbit_r65_c108 bl[108] br[108] wl[65] vdd gnd cell_6t
Xbit_r66_c108 bl[108] br[108] wl[66] vdd gnd cell_6t
Xbit_r67_c108 bl[108] br[108] wl[67] vdd gnd cell_6t
Xbit_r68_c108 bl[108] br[108] wl[68] vdd gnd cell_6t
Xbit_r69_c108 bl[108] br[108] wl[69] vdd gnd cell_6t
Xbit_r70_c108 bl[108] br[108] wl[70] vdd gnd cell_6t
Xbit_r71_c108 bl[108] br[108] wl[71] vdd gnd cell_6t
Xbit_r72_c108 bl[108] br[108] wl[72] vdd gnd cell_6t
Xbit_r73_c108 bl[108] br[108] wl[73] vdd gnd cell_6t
Xbit_r74_c108 bl[108] br[108] wl[74] vdd gnd cell_6t
Xbit_r75_c108 bl[108] br[108] wl[75] vdd gnd cell_6t
Xbit_r76_c108 bl[108] br[108] wl[76] vdd gnd cell_6t
Xbit_r77_c108 bl[108] br[108] wl[77] vdd gnd cell_6t
Xbit_r78_c108 bl[108] br[108] wl[78] vdd gnd cell_6t
Xbit_r79_c108 bl[108] br[108] wl[79] vdd gnd cell_6t
Xbit_r80_c108 bl[108] br[108] wl[80] vdd gnd cell_6t
Xbit_r81_c108 bl[108] br[108] wl[81] vdd gnd cell_6t
Xbit_r82_c108 bl[108] br[108] wl[82] vdd gnd cell_6t
Xbit_r83_c108 bl[108] br[108] wl[83] vdd gnd cell_6t
Xbit_r84_c108 bl[108] br[108] wl[84] vdd gnd cell_6t
Xbit_r85_c108 bl[108] br[108] wl[85] vdd gnd cell_6t
Xbit_r86_c108 bl[108] br[108] wl[86] vdd gnd cell_6t
Xbit_r87_c108 bl[108] br[108] wl[87] vdd gnd cell_6t
Xbit_r88_c108 bl[108] br[108] wl[88] vdd gnd cell_6t
Xbit_r89_c108 bl[108] br[108] wl[89] vdd gnd cell_6t
Xbit_r90_c108 bl[108] br[108] wl[90] vdd gnd cell_6t
Xbit_r91_c108 bl[108] br[108] wl[91] vdd gnd cell_6t
Xbit_r92_c108 bl[108] br[108] wl[92] vdd gnd cell_6t
Xbit_r93_c108 bl[108] br[108] wl[93] vdd gnd cell_6t
Xbit_r94_c108 bl[108] br[108] wl[94] vdd gnd cell_6t
Xbit_r95_c108 bl[108] br[108] wl[95] vdd gnd cell_6t
Xbit_r96_c108 bl[108] br[108] wl[96] vdd gnd cell_6t
Xbit_r97_c108 bl[108] br[108] wl[97] vdd gnd cell_6t
Xbit_r98_c108 bl[108] br[108] wl[98] vdd gnd cell_6t
Xbit_r99_c108 bl[108] br[108] wl[99] vdd gnd cell_6t
Xbit_r100_c108 bl[108] br[108] wl[100] vdd gnd cell_6t
Xbit_r101_c108 bl[108] br[108] wl[101] vdd gnd cell_6t
Xbit_r102_c108 bl[108] br[108] wl[102] vdd gnd cell_6t
Xbit_r103_c108 bl[108] br[108] wl[103] vdd gnd cell_6t
Xbit_r104_c108 bl[108] br[108] wl[104] vdd gnd cell_6t
Xbit_r105_c108 bl[108] br[108] wl[105] vdd gnd cell_6t
Xbit_r106_c108 bl[108] br[108] wl[106] vdd gnd cell_6t
Xbit_r107_c108 bl[108] br[108] wl[107] vdd gnd cell_6t
Xbit_r108_c108 bl[108] br[108] wl[108] vdd gnd cell_6t
Xbit_r109_c108 bl[108] br[108] wl[109] vdd gnd cell_6t
Xbit_r110_c108 bl[108] br[108] wl[110] vdd gnd cell_6t
Xbit_r111_c108 bl[108] br[108] wl[111] vdd gnd cell_6t
Xbit_r112_c108 bl[108] br[108] wl[112] vdd gnd cell_6t
Xbit_r113_c108 bl[108] br[108] wl[113] vdd gnd cell_6t
Xbit_r114_c108 bl[108] br[108] wl[114] vdd gnd cell_6t
Xbit_r115_c108 bl[108] br[108] wl[115] vdd gnd cell_6t
Xbit_r116_c108 bl[108] br[108] wl[116] vdd gnd cell_6t
Xbit_r117_c108 bl[108] br[108] wl[117] vdd gnd cell_6t
Xbit_r118_c108 bl[108] br[108] wl[118] vdd gnd cell_6t
Xbit_r119_c108 bl[108] br[108] wl[119] vdd gnd cell_6t
Xbit_r120_c108 bl[108] br[108] wl[120] vdd gnd cell_6t
Xbit_r121_c108 bl[108] br[108] wl[121] vdd gnd cell_6t
Xbit_r122_c108 bl[108] br[108] wl[122] vdd gnd cell_6t
Xbit_r123_c108 bl[108] br[108] wl[123] vdd gnd cell_6t
Xbit_r124_c108 bl[108] br[108] wl[124] vdd gnd cell_6t
Xbit_r125_c108 bl[108] br[108] wl[125] vdd gnd cell_6t
Xbit_r126_c108 bl[108] br[108] wl[126] vdd gnd cell_6t
Xbit_r127_c108 bl[108] br[108] wl[127] vdd gnd cell_6t
Xbit_r128_c108 bl[108] br[108] wl[128] vdd gnd cell_6t
Xbit_r129_c108 bl[108] br[108] wl[129] vdd gnd cell_6t
Xbit_r130_c108 bl[108] br[108] wl[130] vdd gnd cell_6t
Xbit_r131_c108 bl[108] br[108] wl[131] vdd gnd cell_6t
Xbit_r132_c108 bl[108] br[108] wl[132] vdd gnd cell_6t
Xbit_r133_c108 bl[108] br[108] wl[133] vdd gnd cell_6t
Xbit_r134_c108 bl[108] br[108] wl[134] vdd gnd cell_6t
Xbit_r135_c108 bl[108] br[108] wl[135] vdd gnd cell_6t
Xbit_r136_c108 bl[108] br[108] wl[136] vdd gnd cell_6t
Xbit_r137_c108 bl[108] br[108] wl[137] vdd gnd cell_6t
Xbit_r138_c108 bl[108] br[108] wl[138] vdd gnd cell_6t
Xbit_r139_c108 bl[108] br[108] wl[139] vdd gnd cell_6t
Xbit_r140_c108 bl[108] br[108] wl[140] vdd gnd cell_6t
Xbit_r141_c108 bl[108] br[108] wl[141] vdd gnd cell_6t
Xbit_r142_c108 bl[108] br[108] wl[142] vdd gnd cell_6t
Xbit_r143_c108 bl[108] br[108] wl[143] vdd gnd cell_6t
Xbit_r144_c108 bl[108] br[108] wl[144] vdd gnd cell_6t
Xbit_r145_c108 bl[108] br[108] wl[145] vdd gnd cell_6t
Xbit_r146_c108 bl[108] br[108] wl[146] vdd gnd cell_6t
Xbit_r147_c108 bl[108] br[108] wl[147] vdd gnd cell_6t
Xbit_r148_c108 bl[108] br[108] wl[148] vdd gnd cell_6t
Xbit_r149_c108 bl[108] br[108] wl[149] vdd gnd cell_6t
Xbit_r150_c108 bl[108] br[108] wl[150] vdd gnd cell_6t
Xbit_r151_c108 bl[108] br[108] wl[151] vdd gnd cell_6t
Xbit_r152_c108 bl[108] br[108] wl[152] vdd gnd cell_6t
Xbit_r153_c108 bl[108] br[108] wl[153] vdd gnd cell_6t
Xbit_r154_c108 bl[108] br[108] wl[154] vdd gnd cell_6t
Xbit_r155_c108 bl[108] br[108] wl[155] vdd gnd cell_6t
Xbit_r156_c108 bl[108] br[108] wl[156] vdd gnd cell_6t
Xbit_r157_c108 bl[108] br[108] wl[157] vdd gnd cell_6t
Xbit_r158_c108 bl[108] br[108] wl[158] vdd gnd cell_6t
Xbit_r159_c108 bl[108] br[108] wl[159] vdd gnd cell_6t
Xbit_r160_c108 bl[108] br[108] wl[160] vdd gnd cell_6t
Xbit_r161_c108 bl[108] br[108] wl[161] vdd gnd cell_6t
Xbit_r162_c108 bl[108] br[108] wl[162] vdd gnd cell_6t
Xbit_r163_c108 bl[108] br[108] wl[163] vdd gnd cell_6t
Xbit_r164_c108 bl[108] br[108] wl[164] vdd gnd cell_6t
Xbit_r165_c108 bl[108] br[108] wl[165] vdd gnd cell_6t
Xbit_r166_c108 bl[108] br[108] wl[166] vdd gnd cell_6t
Xbit_r167_c108 bl[108] br[108] wl[167] vdd gnd cell_6t
Xbit_r168_c108 bl[108] br[108] wl[168] vdd gnd cell_6t
Xbit_r169_c108 bl[108] br[108] wl[169] vdd gnd cell_6t
Xbit_r170_c108 bl[108] br[108] wl[170] vdd gnd cell_6t
Xbit_r171_c108 bl[108] br[108] wl[171] vdd gnd cell_6t
Xbit_r172_c108 bl[108] br[108] wl[172] vdd gnd cell_6t
Xbit_r173_c108 bl[108] br[108] wl[173] vdd gnd cell_6t
Xbit_r174_c108 bl[108] br[108] wl[174] vdd gnd cell_6t
Xbit_r175_c108 bl[108] br[108] wl[175] vdd gnd cell_6t
Xbit_r176_c108 bl[108] br[108] wl[176] vdd gnd cell_6t
Xbit_r177_c108 bl[108] br[108] wl[177] vdd gnd cell_6t
Xbit_r178_c108 bl[108] br[108] wl[178] vdd gnd cell_6t
Xbit_r179_c108 bl[108] br[108] wl[179] vdd gnd cell_6t
Xbit_r180_c108 bl[108] br[108] wl[180] vdd gnd cell_6t
Xbit_r181_c108 bl[108] br[108] wl[181] vdd gnd cell_6t
Xbit_r182_c108 bl[108] br[108] wl[182] vdd gnd cell_6t
Xbit_r183_c108 bl[108] br[108] wl[183] vdd gnd cell_6t
Xbit_r184_c108 bl[108] br[108] wl[184] vdd gnd cell_6t
Xbit_r185_c108 bl[108] br[108] wl[185] vdd gnd cell_6t
Xbit_r186_c108 bl[108] br[108] wl[186] vdd gnd cell_6t
Xbit_r187_c108 bl[108] br[108] wl[187] vdd gnd cell_6t
Xbit_r188_c108 bl[108] br[108] wl[188] vdd gnd cell_6t
Xbit_r189_c108 bl[108] br[108] wl[189] vdd gnd cell_6t
Xbit_r190_c108 bl[108] br[108] wl[190] vdd gnd cell_6t
Xbit_r191_c108 bl[108] br[108] wl[191] vdd gnd cell_6t
Xbit_r192_c108 bl[108] br[108] wl[192] vdd gnd cell_6t
Xbit_r193_c108 bl[108] br[108] wl[193] vdd gnd cell_6t
Xbit_r194_c108 bl[108] br[108] wl[194] vdd gnd cell_6t
Xbit_r195_c108 bl[108] br[108] wl[195] vdd gnd cell_6t
Xbit_r196_c108 bl[108] br[108] wl[196] vdd gnd cell_6t
Xbit_r197_c108 bl[108] br[108] wl[197] vdd gnd cell_6t
Xbit_r198_c108 bl[108] br[108] wl[198] vdd gnd cell_6t
Xbit_r199_c108 bl[108] br[108] wl[199] vdd gnd cell_6t
Xbit_r200_c108 bl[108] br[108] wl[200] vdd gnd cell_6t
Xbit_r201_c108 bl[108] br[108] wl[201] vdd gnd cell_6t
Xbit_r202_c108 bl[108] br[108] wl[202] vdd gnd cell_6t
Xbit_r203_c108 bl[108] br[108] wl[203] vdd gnd cell_6t
Xbit_r204_c108 bl[108] br[108] wl[204] vdd gnd cell_6t
Xbit_r205_c108 bl[108] br[108] wl[205] vdd gnd cell_6t
Xbit_r206_c108 bl[108] br[108] wl[206] vdd gnd cell_6t
Xbit_r207_c108 bl[108] br[108] wl[207] vdd gnd cell_6t
Xbit_r208_c108 bl[108] br[108] wl[208] vdd gnd cell_6t
Xbit_r209_c108 bl[108] br[108] wl[209] vdd gnd cell_6t
Xbit_r210_c108 bl[108] br[108] wl[210] vdd gnd cell_6t
Xbit_r211_c108 bl[108] br[108] wl[211] vdd gnd cell_6t
Xbit_r212_c108 bl[108] br[108] wl[212] vdd gnd cell_6t
Xbit_r213_c108 bl[108] br[108] wl[213] vdd gnd cell_6t
Xbit_r214_c108 bl[108] br[108] wl[214] vdd gnd cell_6t
Xbit_r215_c108 bl[108] br[108] wl[215] vdd gnd cell_6t
Xbit_r216_c108 bl[108] br[108] wl[216] vdd gnd cell_6t
Xbit_r217_c108 bl[108] br[108] wl[217] vdd gnd cell_6t
Xbit_r218_c108 bl[108] br[108] wl[218] vdd gnd cell_6t
Xbit_r219_c108 bl[108] br[108] wl[219] vdd gnd cell_6t
Xbit_r220_c108 bl[108] br[108] wl[220] vdd gnd cell_6t
Xbit_r221_c108 bl[108] br[108] wl[221] vdd gnd cell_6t
Xbit_r222_c108 bl[108] br[108] wl[222] vdd gnd cell_6t
Xbit_r223_c108 bl[108] br[108] wl[223] vdd gnd cell_6t
Xbit_r224_c108 bl[108] br[108] wl[224] vdd gnd cell_6t
Xbit_r225_c108 bl[108] br[108] wl[225] vdd gnd cell_6t
Xbit_r226_c108 bl[108] br[108] wl[226] vdd gnd cell_6t
Xbit_r227_c108 bl[108] br[108] wl[227] vdd gnd cell_6t
Xbit_r228_c108 bl[108] br[108] wl[228] vdd gnd cell_6t
Xbit_r229_c108 bl[108] br[108] wl[229] vdd gnd cell_6t
Xbit_r230_c108 bl[108] br[108] wl[230] vdd gnd cell_6t
Xbit_r231_c108 bl[108] br[108] wl[231] vdd gnd cell_6t
Xbit_r232_c108 bl[108] br[108] wl[232] vdd gnd cell_6t
Xbit_r233_c108 bl[108] br[108] wl[233] vdd gnd cell_6t
Xbit_r234_c108 bl[108] br[108] wl[234] vdd gnd cell_6t
Xbit_r235_c108 bl[108] br[108] wl[235] vdd gnd cell_6t
Xbit_r236_c108 bl[108] br[108] wl[236] vdd gnd cell_6t
Xbit_r237_c108 bl[108] br[108] wl[237] vdd gnd cell_6t
Xbit_r238_c108 bl[108] br[108] wl[238] vdd gnd cell_6t
Xbit_r239_c108 bl[108] br[108] wl[239] vdd gnd cell_6t
Xbit_r240_c108 bl[108] br[108] wl[240] vdd gnd cell_6t
Xbit_r241_c108 bl[108] br[108] wl[241] vdd gnd cell_6t
Xbit_r242_c108 bl[108] br[108] wl[242] vdd gnd cell_6t
Xbit_r243_c108 bl[108] br[108] wl[243] vdd gnd cell_6t
Xbit_r244_c108 bl[108] br[108] wl[244] vdd gnd cell_6t
Xbit_r245_c108 bl[108] br[108] wl[245] vdd gnd cell_6t
Xbit_r246_c108 bl[108] br[108] wl[246] vdd gnd cell_6t
Xbit_r247_c108 bl[108] br[108] wl[247] vdd gnd cell_6t
Xbit_r248_c108 bl[108] br[108] wl[248] vdd gnd cell_6t
Xbit_r249_c108 bl[108] br[108] wl[249] vdd gnd cell_6t
Xbit_r250_c108 bl[108] br[108] wl[250] vdd gnd cell_6t
Xbit_r251_c108 bl[108] br[108] wl[251] vdd gnd cell_6t
Xbit_r252_c108 bl[108] br[108] wl[252] vdd gnd cell_6t
Xbit_r253_c108 bl[108] br[108] wl[253] vdd gnd cell_6t
Xbit_r254_c108 bl[108] br[108] wl[254] vdd gnd cell_6t
Xbit_r255_c108 bl[108] br[108] wl[255] vdd gnd cell_6t
Xbit_r0_c109 bl[109] br[109] wl[0] vdd gnd cell_6t
Xbit_r1_c109 bl[109] br[109] wl[1] vdd gnd cell_6t
Xbit_r2_c109 bl[109] br[109] wl[2] vdd gnd cell_6t
Xbit_r3_c109 bl[109] br[109] wl[3] vdd gnd cell_6t
Xbit_r4_c109 bl[109] br[109] wl[4] vdd gnd cell_6t
Xbit_r5_c109 bl[109] br[109] wl[5] vdd gnd cell_6t
Xbit_r6_c109 bl[109] br[109] wl[6] vdd gnd cell_6t
Xbit_r7_c109 bl[109] br[109] wl[7] vdd gnd cell_6t
Xbit_r8_c109 bl[109] br[109] wl[8] vdd gnd cell_6t
Xbit_r9_c109 bl[109] br[109] wl[9] vdd gnd cell_6t
Xbit_r10_c109 bl[109] br[109] wl[10] vdd gnd cell_6t
Xbit_r11_c109 bl[109] br[109] wl[11] vdd gnd cell_6t
Xbit_r12_c109 bl[109] br[109] wl[12] vdd gnd cell_6t
Xbit_r13_c109 bl[109] br[109] wl[13] vdd gnd cell_6t
Xbit_r14_c109 bl[109] br[109] wl[14] vdd gnd cell_6t
Xbit_r15_c109 bl[109] br[109] wl[15] vdd gnd cell_6t
Xbit_r16_c109 bl[109] br[109] wl[16] vdd gnd cell_6t
Xbit_r17_c109 bl[109] br[109] wl[17] vdd gnd cell_6t
Xbit_r18_c109 bl[109] br[109] wl[18] vdd gnd cell_6t
Xbit_r19_c109 bl[109] br[109] wl[19] vdd gnd cell_6t
Xbit_r20_c109 bl[109] br[109] wl[20] vdd gnd cell_6t
Xbit_r21_c109 bl[109] br[109] wl[21] vdd gnd cell_6t
Xbit_r22_c109 bl[109] br[109] wl[22] vdd gnd cell_6t
Xbit_r23_c109 bl[109] br[109] wl[23] vdd gnd cell_6t
Xbit_r24_c109 bl[109] br[109] wl[24] vdd gnd cell_6t
Xbit_r25_c109 bl[109] br[109] wl[25] vdd gnd cell_6t
Xbit_r26_c109 bl[109] br[109] wl[26] vdd gnd cell_6t
Xbit_r27_c109 bl[109] br[109] wl[27] vdd gnd cell_6t
Xbit_r28_c109 bl[109] br[109] wl[28] vdd gnd cell_6t
Xbit_r29_c109 bl[109] br[109] wl[29] vdd gnd cell_6t
Xbit_r30_c109 bl[109] br[109] wl[30] vdd gnd cell_6t
Xbit_r31_c109 bl[109] br[109] wl[31] vdd gnd cell_6t
Xbit_r32_c109 bl[109] br[109] wl[32] vdd gnd cell_6t
Xbit_r33_c109 bl[109] br[109] wl[33] vdd gnd cell_6t
Xbit_r34_c109 bl[109] br[109] wl[34] vdd gnd cell_6t
Xbit_r35_c109 bl[109] br[109] wl[35] vdd gnd cell_6t
Xbit_r36_c109 bl[109] br[109] wl[36] vdd gnd cell_6t
Xbit_r37_c109 bl[109] br[109] wl[37] vdd gnd cell_6t
Xbit_r38_c109 bl[109] br[109] wl[38] vdd gnd cell_6t
Xbit_r39_c109 bl[109] br[109] wl[39] vdd gnd cell_6t
Xbit_r40_c109 bl[109] br[109] wl[40] vdd gnd cell_6t
Xbit_r41_c109 bl[109] br[109] wl[41] vdd gnd cell_6t
Xbit_r42_c109 bl[109] br[109] wl[42] vdd gnd cell_6t
Xbit_r43_c109 bl[109] br[109] wl[43] vdd gnd cell_6t
Xbit_r44_c109 bl[109] br[109] wl[44] vdd gnd cell_6t
Xbit_r45_c109 bl[109] br[109] wl[45] vdd gnd cell_6t
Xbit_r46_c109 bl[109] br[109] wl[46] vdd gnd cell_6t
Xbit_r47_c109 bl[109] br[109] wl[47] vdd gnd cell_6t
Xbit_r48_c109 bl[109] br[109] wl[48] vdd gnd cell_6t
Xbit_r49_c109 bl[109] br[109] wl[49] vdd gnd cell_6t
Xbit_r50_c109 bl[109] br[109] wl[50] vdd gnd cell_6t
Xbit_r51_c109 bl[109] br[109] wl[51] vdd gnd cell_6t
Xbit_r52_c109 bl[109] br[109] wl[52] vdd gnd cell_6t
Xbit_r53_c109 bl[109] br[109] wl[53] vdd gnd cell_6t
Xbit_r54_c109 bl[109] br[109] wl[54] vdd gnd cell_6t
Xbit_r55_c109 bl[109] br[109] wl[55] vdd gnd cell_6t
Xbit_r56_c109 bl[109] br[109] wl[56] vdd gnd cell_6t
Xbit_r57_c109 bl[109] br[109] wl[57] vdd gnd cell_6t
Xbit_r58_c109 bl[109] br[109] wl[58] vdd gnd cell_6t
Xbit_r59_c109 bl[109] br[109] wl[59] vdd gnd cell_6t
Xbit_r60_c109 bl[109] br[109] wl[60] vdd gnd cell_6t
Xbit_r61_c109 bl[109] br[109] wl[61] vdd gnd cell_6t
Xbit_r62_c109 bl[109] br[109] wl[62] vdd gnd cell_6t
Xbit_r63_c109 bl[109] br[109] wl[63] vdd gnd cell_6t
Xbit_r64_c109 bl[109] br[109] wl[64] vdd gnd cell_6t
Xbit_r65_c109 bl[109] br[109] wl[65] vdd gnd cell_6t
Xbit_r66_c109 bl[109] br[109] wl[66] vdd gnd cell_6t
Xbit_r67_c109 bl[109] br[109] wl[67] vdd gnd cell_6t
Xbit_r68_c109 bl[109] br[109] wl[68] vdd gnd cell_6t
Xbit_r69_c109 bl[109] br[109] wl[69] vdd gnd cell_6t
Xbit_r70_c109 bl[109] br[109] wl[70] vdd gnd cell_6t
Xbit_r71_c109 bl[109] br[109] wl[71] vdd gnd cell_6t
Xbit_r72_c109 bl[109] br[109] wl[72] vdd gnd cell_6t
Xbit_r73_c109 bl[109] br[109] wl[73] vdd gnd cell_6t
Xbit_r74_c109 bl[109] br[109] wl[74] vdd gnd cell_6t
Xbit_r75_c109 bl[109] br[109] wl[75] vdd gnd cell_6t
Xbit_r76_c109 bl[109] br[109] wl[76] vdd gnd cell_6t
Xbit_r77_c109 bl[109] br[109] wl[77] vdd gnd cell_6t
Xbit_r78_c109 bl[109] br[109] wl[78] vdd gnd cell_6t
Xbit_r79_c109 bl[109] br[109] wl[79] vdd gnd cell_6t
Xbit_r80_c109 bl[109] br[109] wl[80] vdd gnd cell_6t
Xbit_r81_c109 bl[109] br[109] wl[81] vdd gnd cell_6t
Xbit_r82_c109 bl[109] br[109] wl[82] vdd gnd cell_6t
Xbit_r83_c109 bl[109] br[109] wl[83] vdd gnd cell_6t
Xbit_r84_c109 bl[109] br[109] wl[84] vdd gnd cell_6t
Xbit_r85_c109 bl[109] br[109] wl[85] vdd gnd cell_6t
Xbit_r86_c109 bl[109] br[109] wl[86] vdd gnd cell_6t
Xbit_r87_c109 bl[109] br[109] wl[87] vdd gnd cell_6t
Xbit_r88_c109 bl[109] br[109] wl[88] vdd gnd cell_6t
Xbit_r89_c109 bl[109] br[109] wl[89] vdd gnd cell_6t
Xbit_r90_c109 bl[109] br[109] wl[90] vdd gnd cell_6t
Xbit_r91_c109 bl[109] br[109] wl[91] vdd gnd cell_6t
Xbit_r92_c109 bl[109] br[109] wl[92] vdd gnd cell_6t
Xbit_r93_c109 bl[109] br[109] wl[93] vdd gnd cell_6t
Xbit_r94_c109 bl[109] br[109] wl[94] vdd gnd cell_6t
Xbit_r95_c109 bl[109] br[109] wl[95] vdd gnd cell_6t
Xbit_r96_c109 bl[109] br[109] wl[96] vdd gnd cell_6t
Xbit_r97_c109 bl[109] br[109] wl[97] vdd gnd cell_6t
Xbit_r98_c109 bl[109] br[109] wl[98] vdd gnd cell_6t
Xbit_r99_c109 bl[109] br[109] wl[99] vdd gnd cell_6t
Xbit_r100_c109 bl[109] br[109] wl[100] vdd gnd cell_6t
Xbit_r101_c109 bl[109] br[109] wl[101] vdd gnd cell_6t
Xbit_r102_c109 bl[109] br[109] wl[102] vdd gnd cell_6t
Xbit_r103_c109 bl[109] br[109] wl[103] vdd gnd cell_6t
Xbit_r104_c109 bl[109] br[109] wl[104] vdd gnd cell_6t
Xbit_r105_c109 bl[109] br[109] wl[105] vdd gnd cell_6t
Xbit_r106_c109 bl[109] br[109] wl[106] vdd gnd cell_6t
Xbit_r107_c109 bl[109] br[109] wl[107] vdd gnd cell_6t
Xbit_r108_c109 bl[109] br[109] wl[108] vdd gnd cell_6t
Xbit_r109_c109 bl[109] br[109] wl[109] vdd gnd cell_6t
Xbit_r110_c109 bl[109] br[109] wl[110] vdd gnd cell_6t
Xbit_r111_c109 bl[109] br[109] wl[111] vdd gnd cell_6t
Xbit_r112_c109 bl[109] br[109] wl[112] vdd gnd cell_6t
Xbit_r113_c109 bl[109] br[109] wl[113] vdd gnd cell_6t
Xbit_r114_c109 bl[109] br[109] wl[114] vdd gnd cell_6t
Xbit_r115_c109 bl[109] br[109] wl[115] vdd gnd cell_6t
Xbit_r116_c109 bl[109] br[109] wl[116] vdd gnd cell_6t
Xbit_r117_c109 bl[109] br[109] wl[117] vdd gnd cell_6t
Xbit_r118_c109 bl[109] br[109] wl[118] vdd gnd cell_6t
Xbit_r119_c109 bl[109] br[109] wl[119] vdd gnd cell_6t
Xbit_r120_c109 bl[109] br[109] wl[120] vdd gnd cell_6t
Xbit_r121_c109 bl[109] br[109] wl[121] vdd gnd cell_6t
Xbit_r122_c109 bl[109] br[109] wl[122] vdd gnd cell_6t
Xbit_r123_c109 bl[109] br[109] wl[123] vdd gnd cell_6t
Xbit_r124_c109 bl[109] br[109] wl[124] vdd gnd cell_6t
Xbit_r125_c109 bl[109] br[109] wl[125] vdd gnd cell_6t
Xbit_r126_c109 bl[109] br[109] wl[126] vdd gnd cell_6t
Xbit_r127_c109 bl[109] br[109] wl[127] vdd gnd cell_6t
Xbit_r128_c109 bl[109] br[109] wl[128] vdd gnd cell_6t
Xbit_r129_c109 bl[109] br[109] wl[129] vdd gnd cell_6t
Xbit_r130_c109 bl[109] br[109] wl[130] vdd gnd cell_6t
Xbit_r131_c109 bl[109] br[109] wl[131] vdd gnd cell_6t
Xbit_r132_c109 bl[109] br[109] wl[132] vdd gnd cell_6t
Xbit_r133_c109 bl[109] br[109] wl[133] vdd gnd cell_6t
Xbit_r134_c109 bl[109] br[109] wl[134] vdd gnd cell_6t
Xbit_r135_c109 bl[109] br[109] wl[135] vdd gnd cell_6t
Xbit_r136_c109 bl[109] br[109] wl[136] vdd gnd cell_6t
Xbit_r137_c109 bl[109] br[109] wl[137] vdd gnd cell_6t
Xbit_r138_c109 bl[109] br[109] wl[138] vdd gnd cell_6t
Xbit_r139_c109 bl[109] br[109] wl[139] vdd gnd cell_6t
Xbit_r140_c109 bl[109] br[109] wl[140] vdd gnd cell_6t
Xbit_r141_c109 bl[109] br[109] wl[141] vdd gnd cell_6t
Xbit_r142_c109 bl[109] br[109] wl[142] vdd gnd cell_6t
Xbit_r143_c109 bl[109] br[109] wl[143] vdd gnd cell_6t
Xbit_r144_c109 bl[109] br[109] wl[144] vdd gnd cell_6t
Xbit_r145_c109 bl[109] br[109] wl[145] vdd gnd cell_6t
Xbit_r146_c109 bl[109] br[109] wl[146] vdd gnd cell_6t
Xbit_r147_c109 bl[109] br[109] wl[147] vdd gnd cell_6t
Xbit_r148_c109 bl[109] br[109] wl[148] vdd gnd cell_6t
Xbit_r149_c109 bl[109] br[109] wl[149] vdd gnd cell_6t
Xbit_r150_c109 bl[109] br[109] wl[150] vdd gnd cell_6t
Xbit_r151_c109 bl[109] br[109] wl[151] vdd gnd cell_6t
Xbit_r152_c109 bl[109] br[109] wl[152] vdd gnd cell_6t
Xbit_r153_c109 bl[109] br[109] wl[153] vdd gnd cell_6t
Xbit_r154_c109 bl[109] br[109] wl[154] vdd gnd cell_6t
Xbit_r155_c109 bl[109] br[109] wl[155] vdd gnd cell_6t
Xbit_r156_c109 bl[109] br[109] wl[156] vdd gnd cell_6t
Xbit_r157_c109 bl[109] br[109] wl[157] vdd gnd cell_6t
Xbit_r158_c109 bl[109] br[109] wl[158] vdd gnd cell_6t
Xbit_r159_c109 bl[109] br[109] wl[159] vdd gnd cell_6t
Xbit_r160_c109 bl[109] br[109] wl[160] vdd gnd cell_6t
Xbit_r161_c109 bl[109] br[109] wl[161] vdd gnd cell_6t
Xbit_r162_c109 bl[109] br[109] wl[162] vdd gnd cell_6t
Xbit_r163_c109 bl[109] br[109] wl[163] vdd gnd cell_6t
Xbit_r164_c109 bl[109] br[109] wl[164] vdd gnd cell_6t
Xbit_r165_c109 bl[109] br[109] wl[165] vdd gnd cell_6t
Xbit_r166_c109 bl[109] br[109] wl[166] vdd gnd cell_6t
Xbit_r167_c109 bl[109] br[109] wl[167] vdd gnd cell_6t
Xbit_r168_c109 bl[109] br[109] wl[168] vdd gnd cell_6t
Xbit_r169_c109 bl[109] br[109] wl[169] vdd gnd cell_6t
Xbit_r170_c109 bl[109] br[109] wl[170] vdd gnd cell_6t
Xbit_r171_c109 bl[109] br[109] wl[171] vdd gnd cell_6t
Xbit_r172_c109 bl[109] br[109] wl[172] vdd gnd cell_6t
Xbit_r173_c109 bl[109] br[109] wl[173] vdd gnd cell_6t
Xbit_r174_c109 bl[109] br[109] wl[174] vdd gnd cell_6t
Xbit_r175_c109 bl[109] br[109] wl[175] vdd gnd cell_6t
Xbit_r176_c109 bl[109] br[109] wl[176] vdd gnd cell_6t
Xbit_r177_c109 bl[109] br[109] wl[177] vdd gnd cell_6t
Xbit_r178_c109 bl[109] br[109] wl[178] vdd gnd cell_6t
Xbit_r179_c109 bl[109] br[109] wl[179] vdd gnd cell_6t
Xbit_r180_c109 bl[109] br[109] wl[180] vdd gnd cell_6t
Xbit_r181_c109 bl[109] br[109] wl[181] vdd gnd cell_6t
Xbit_r182_c109 bl[109] br[109] wl[182] vdd gnd cell_6t
Xbit_r183_c109 bl[109] br[109] wl[183] vdd gnd cell_6t
Xbit_r184_c109 bl[109] br[109] wl[184] vdd gnd cell_6t
Xbit_r185_c109 bl[109] br[109] wl[185] vdd gnd cell_6t
Xbit_r186_c109 bl[109] br[109] wl[186] vdd gnd cell_6t
Xbit_r187_c109 bl[109] br[109] wl[187] vdd gnd cell_6t
Xbit_r188_c109 bl[109] br[109] wl[188] vdd gnd cell_6t
Xbit_r189_c109 bl[109] br[109] wl[189] vdd gnd cell_6t
Xbit_r190_c109 bl[109] br[109] wl[190] vdd gnd cell_6t
Xbit_r191_c109 bl[109] br[109] wl[191] vdd gnd cell_6t
Xbit_r192_c109 bl[109] br[109] wl[192] vdd gnd cell_6t
Xbit_r193_c109 bl[109] br[109] wl[193] vdd gnd cell_6t
Xbit_r194_c109 bl[109] br[109] wl[194] vdd gnd cell_6t
Xbit_r195_c109 bl[109] br[109] wl[195] vdd gnd cell_6t
Xbit_r196_c109 bl[109] br[109] wl[196] vdd gnd cell_6t
Xbit_r197_c109 bl[109] br[109] wl[197] vdd gnd cell_6t
Xbit_r198_c109 bl[109] br[109] wl[198] vdd gnd cell_6t
Xbit_r199_c109 bl[109] br[109] wl[199] vdd gnd cell_6t
Xbit_r200_c109 bl[109] br[109] wl[200] vdd gnd cell_6t
Xbit_r201_c109 bl[109] br[109] wl[201] vdd gnd cell_6t
Xbit_r202_c109 bl[109] br[109] wl[202] vdd gnd cell_6t
Xbit_r203_c109 bl[109] br[109] wl[203] vdd gnd cell_6t
Xbit_r204_c109 bl[109] br[109] wl[204] vdd gnd cell_6t
Xbit_r205_c109 bl[109] br[109] wl[205] vdd gnd cell_6t
Xbit_r206_c109 bl[109] br[109] wl[206] vdd gnd cell_6t
Xbit_r207_c109 bl[109] br[109] wl[207] vdd gnd cell_6t
Xbit_r208_c109 bl[109] br[109] wl[208] vdd gnd cell_6t
Xbit_r209_c109 bl[109] br[109] wl[209] vdd gnd cell_6t
Xbit_r210_c109 bl[109] br[109] wl[210] vdd gnd cell_6t
Xbit_r211_c109 bl[109] br[109] wl[211] vdd gnd cell_6t
Xbit_r212_c109 bl[109] br[109] wl[212] vdd gnd cell_6t
Xbit_r213_c109 bl[109] br[109] wl[213] vdd gnd cell_6t
Xbit_r214_c109 bl[109] br[109] wl[214] vdd gnd cell_6t
Xbit_r215_c109 bl[109] br[109] wl[215] vdd gnd cell_6t
Xbit_r216_c109 bl[109] br[109] wl[216] vdd gnd cell_6t
Xbit_r217_c109 bl[109] br[109] wl[217] vdd gnd cell_6t
Xbit_r218_c109 bl[109] br[109] wl[218] vdd gnd cell_6t
Xbit_r219_c109 bl[109] br[109] wl[219] vdd gnd cell_6t
Xbit_r220_c109 bl[109] br[109] wl[220] vdd gnd cell_6t
Xbit_r221_c109 bl[109] br[109] wl[221] vdd gnd cell_6t
Xbit_r222_c109 bl[109] br[109] wl[222] vdd gnd cell_6t
Xbit_r223_c109 bl[109] br[109] wl[223] vdd gnd cell_6t
Xbit_r224_c109 bl[109] br[109] wl[224] vdd gnd cell_6t
Xbit_r225_c109 bl[109] br[109] wl[225] vdd gnd cell_6t
Xbit_r226_c109 bl[109] br[109] wl[226] vdd gnd cell_6t
Xbit_r227_c109 bl[109] br[109] wl[227] vdd gnd cell_6t
Xbit_r228_c109 bl[109] br[109] wl[228] vdd gnd cell_6t
Xbit_r229_c109 bl[109] br[109] wl[229] vdd gnd cell_6t
Xbit_r230_c109 bl[109] br[109] wl[230] vdd gnd cell_6t
Xbit_r231_c109 bl[109] br[109] wl[231] vdd gnd cell_6t
Xbit_r232_c109 bl[109] br[109] wl[232] vdd gnd cell_6t
Xbit_r233_c109 bl[109] br[109] wl[233] vdd gnd cell_6t
Xbit_r234_c109 bl[109] br[109] wl[234] vdd gnd cell_6t
Xbit_r235_c109 bl[109] br[109] wl[235] vdd gnd cell_6t
Xbit_r236_c109 bl[109] br[109] wl[236] vdd gnd cell_6t
Xbit_r237_c109 bl[109] br[109] wl[237] vdd gnd cell_6t
Xbit_r238_c109 bl[109] br[109] wl[238] vdd gnd cell_6t
Xbit_r239_c109 bl[109] br[109] wl[239] vdd gnd cell_6t
Xbit_r240_c109 bl[109] br[109] wl[240] vdd gnd cell_6t
Xbit_r241_c109 bl[109] br[109] wl[241] vdd gnd cell_6t
Xbit_r242_c109 bl[109] br[109] wl[242] vdd gnd cell_6t
Xbit_r243_c109 bl[109] br[109] wl[243] vdd gnd cell_6t
Xbit_r244_c109 bl[109] br[109] wl[244] vdd gnd cell_6t
Xbit_r245_c109 bl[109] br[109] wl[245] vdd gnd cell_6t
Xbit_r246_c109 bl[109] br[109] wl[246] vdd gnd cell_6t
Xbit_r247_c109 bl[109] br[109] wl[247] vdd gnd cell_6t
Xbit_r248_c109 bl[109] br[109] wl[248] vdd gnd cell_6t
Xbit_r249_c109 bl[109] br[109] wl[249] vdd gnd cell_6t
Xbit_r250_c109 bl[109] br[109] wl[250] vdd gnd cell_6t
Xbit_r251_c109 bl[109] br[109] wl[251] vdd gnd cell_6t
Xbit_r252_c109 bl[109] br[109] wl[252] vdd gnd cell_6t
Xbit_r253_c109 bl[109] br[109] wl[253] vdd gnd cell_6t
Xbit_r254_c109 bl[109] br[109] wl[254] vdd gnd cell_6t
Xbit_r255_c109 bl[109] br[109] wl[255] vdd gnd cell_6t
Xbit_r0_c110 bl[110] br[110] wl[0] vdd gnd cell_6t
Xbit_r1_c110 bl[110] br[110] wl[1] vdd gnd cell_6t
Xbit_r2_c110 bl[110] br[110] wl[2] vdd gnd cell_6t
Xbit_r3_c110 bl[110] br[110] wl[3] vdd gnd cell_6t
Xbit_r4_c110 bl[110] br[110] wl[4] vdd gnd cell_6t
Xbit_r5_c110 bl[110] br[110] wl[5] vdd gnd cell_6t
Xbit_r6_c110 bl[110] br[110] wl[6] vdd gnd cell_6t
Xbit_r7_c110 bl[110] br[110] wl[7] vdd gnd cell_6t
Xbit_r8_c110 bl[110] br[110] wl[8] vdd gnd cell_6t
Xbit_r9_c110 bl[110] br[110] wl[9] vdd gnd cell_6t
Xbit_r10_c110 bl[110] br[110] wl[10] vdd gnd cell_6t
Xbit_r11_c110 bl[110] br[110] wl[11] vdd gnd cell_6t
Xbit_r12_c110 bl[110] br[110] wl[12] vdd gnd cell_6t
Xbit_r13_c110 bl[110] br[110] wl[13] vdd gnd cell_6t
Xbit_r14_c110 bl[110] br[110] wl[14] vdd gnd cell_6t
Xbit_r15_c110 bl[110] br[110] wl[15] vdd gnd cell_6t
Xbit_r16_c110 bl[110] br[110] wl[16] vdd gnd cell_6t
Xbit_r17_c110 bl[110] br[110] wl[17] vdd gnd cell_6t
Xbit_r18_c110 bl[110] br[110] wl[18] vdd gnd cell_6t
Xbit_r19_c110 bl[110] br[110] wl[19] vdd gnd cell_6t
Xbit_r20_c110 bl[110] br[110] wl[20] vdd gnd cell_6t
Xbit_r21_c110 bl[110] br[110] wl[21] vdd gnd cell_6t
Xbit_r22_c110 bl[110] br[110] wl[22] vdd gnd cell_6t
Xbit_r23_c110 bl[110] br[110] wl[23] vdd gnd cell_6t
Xbit_r24_c110 bl[110] br[110] wl[24] vdd gnd cell_6t
Xbit_r25_c110 bl[110] br[110] wl[25] vdd gnd cell_6t
Xbit_r26_c110 bl[110] br[110] wl[26] vdd gnd cell_6t
Xbit_r27_c110 bl[110] br[110] wl[27] vdd gnd cell_6t
Xbit_r28_c110 bl[110] br[110] wl[28] vdd gnd cell_6t
Xbit_r29_c110 bl[110] br[110] wl[29] vdd gnd cell_6t
Xbit_r30_c110 bl[110] br[110] wl[30] vdd gnd cell_6t
Xbit_r31_c110 bl[110] br[110] wl[31] vdd gnd cell_6t
Xbit_r32_c110 bl[110] br[110] wl[32] vdd gnd cell_6t
Xbit_r33_c110 bl[110] br[110] wl[33] vdd gnd cell_6t
Xbit_r34_c110 bl[110] br[110] wl[34] vdd gnd cell_6t
Xbit_r35_c110 bl[110] br[110] wl[35] vdd gnd cell_6t
Xbit_r36_c110 bl[110] br[110] wl[36] vdd gnd cell_6t
Xbit_r37_c110 bl[110] br[110] wl[37] vdd gnd cell_6t
Xbit_r38_c110 bl[110] br[110] wl[38] vdd gnd cell_6t
Xbit_r39_c110 bl[110] br[110] wl[39] vdd gnd cell_6t
Xbit_r40_c110 bl[110] br[110] wl[40] vdd gnd cell_6t
Xbit_r41_c110 bl[110] br[110] wl[41] vdd gnd cell_6t
Xbit_r42_c110 bl[110] br[110] wl[42] vdd gnd cell_6t
Xbit_r43_c110 bl[110] br[110] wl[43] vdd gnd cell_6t
Xbit_r44_c110 bl[110] br[110] wl[44] vdd gnd cell_6t
Xbit_r45_c110 bl[110] br[110] wl[45] vdd gnd cell_6t
Xbit_r46_c110 bl[110] br[110] wl[46] vdd gnd cell_6t
Xbit_r47_c110 bl[110] br[110] wl[47] vdd gnd cell_6t
Xbit_r48_c110 bl[110] br[110] wl[48] vdd gnd cell_6t
Xbit_r49_c110 bl[110] br[110] wl[49] vdd gnd cell_6t
Xbit_r50_c110 bl[110] br[110] wl[50] vdd gnd cell_6t
Xbit_r51_c110 bl[110] br[110] wl[51] vdd gnd cell_6t
Xbit_r52_c110 bl[110] br[110] wl[52] vdd gnd cell_6t
Xbit_r53_c110 bl[110] br[110] wl[53] vdd gnd cell_6t
Xbit_r54_c110 bl[110] br[110] wl[54] vdd gnd cell_6t
Xbit_r55_c110 bl[110] br[110] wl[55] vdd gnd cell_6t
Xbit_r56_c110 bl[110] br[110] wl[56] vdd gnd cell_6t
Xbit_r57_c110 bl[110] br[110] wl[57] vdd gnd cell_6t
Xbit_r58_c110 bl[110] br[110] wl[58] vdd gnd cell_6t
Xbit_r59_c110 bl[110] br[110] wl[59] vdd gnd cell_6t
Xbit_r60_c110 bl[110] br[110] wl[60] vdd gnd cell_6t
Xbit_r61_c110 bl[110] br[110] wl[61] vdd gnd cell_6t
Xbit_r62_c110 bl[110] br[110] wl[62] vdd gnd cell_6t
Xbit_r63_c110 bl[110] br[110] wl[63] vdd gnd cell_6t
Xbit_r64_c110 bl[110] br[110] wl[64] vdd gnd cell_6t
Xbit_r65_c110 bl[110] br[110] wl[65] vdd gnd cell_6t
Xbit_r66_c110 bl[110] br[110] wl[66] vdd gnd cell_6t
Xbit_r67_c110 bl[110] br[110] wl[67] vdd gnd cell_6t
Xbit_r68_c110 bl[110] br[110] wl[68] vdd gnd cell_6t
Xbit_r69_c110 bl[110] br[110] wl[69] vdd gnd cell_6t
Xbit_r70_c110 bl[110] br[110] wl[70] vdd gnd cell_6t
Xbit_r71_c110 bl[110] br[110] wl[71] vdd gnd cell_6t
Xbit_r72_c110 bl[110] br[110] wl[72] vdd gnd cell_6t
Xbit_r73_c110 bl[110] br[110] wl[73] vdd gnd cell_6t
Xbit_r74_c110 bl[110] br[110] wl[74] vdd gnd cell_6t
Xbit_r75_c110 bl[110] br[110] wl[75] vdd gnd cell_6t
Xbit_r76_c110 bl[110] br[110] wl[76] vdd gnd cell_6t
Xbit_r77_c110 bl[110] br[110] wl[77] vdd gnd cell_6t
Xbit_r78_c110 bl[110] br[110] wl[78] vdd gnd cell_6t
Xbit_r79_c110 bl[110] br[110] wl[79] vdd gnd cell_6t
Xbit_r80_c110 bl[110] br[110] wl[80] vdd gnd cell_6t
Xbit_r81_c110 bl[110] br[110] wl[81] vdd gnd cell_6t
Xbit_r82_c110 bl[110] br[110] wl[82] vdd gnd cell_6t
Xbit_r83_c110 bl[110] br[110] wl[83] vdd gnd cell_6t
Xbit_r84_c110 bl[110] br[110] wl[84] vdd gnd cell_6t
Xbit_r85_c110 bl[110] br[110] wl[85] vdd gnd cell_6t
Xbit_r86_c110 bl[110] br[110] wl[86] vdd gnd cell_6t
Xbit_r87_c110 bl[110] br[110] wl[87] vdd gnd cell_6t
Xbit_r88_c110 bl[110] br[110] wl[88] vdd gnd cell_6t
Xbit_r89_c110 bl[110] br[110] wl[89] vdd gnd cell_6t
Xbit_r90_c110 bl[110] br[110] wl[90] vdd gnd cell_6t
Xbit_r91_c110 bl[110] br[110] wl[91] vdd gnd cell_6t
Xbit_r92_c110 bl[110] br[110] wl[92] vdd gnd cell_6t
Xbit_r93_c110 bl[110] br[110] wl[93] vdd gnd cell_6t
Xbit_r94_c110 bl[110] br[110] wl[94] vdd gnd cell_6t
Xbit_r95_c110 bl[110] br[110] wl[95] vdd gnd cell_6t
Xbit_r96_c110 bl[110] br[110] wl[96] vdd gnd cell_6t
Xbit_r97_c110 bl[110] br[110] wl[97] vdd gnd cell_6t
Xbit_r98_c110 bl[110] br[110] wl[98] vdd gnd cell_6t
Xbit_r99_c110 bl[110] br[110] wl[99] vdd gnd cell_6t
Xbit_r100_c110 bl[110] br[110] wl[100] vdd gnd cell_6t
Xbit_r101_c110 bl[110] br[110] wl[101] vdd gnd cell_6t
Xbit_r102_c110 bl[110] br[110] wl[102] vdd gnd cell_6t
Xbit_r103_c110 bl[110] br[110] wl[103] vdd gnd cell_6t
Xbit_r104_c110 bl[110] br[110] wl[104] vdd gnd cell_6t
Xbit_r105_c110 bl[110] br[110] wl[105] vdd gnd cell_6t
Xbit_r106_c110 bl[110] br[110] wl[106] vdd gnd cell_6t
Xbit_r107_c110 bl[110] br[110] wl[107] vdd gnd cell_6t
Xbit_r108_c110 bl[110] br[110] wl[108] vdd gnd cell_6t
Xbit_r109_c110 bl[110] br[110] wl[109] vdd gnd cell_6t
Xbit_r110_c110 bl[110] br[110] wl[110] vdd gnd cell_6t
Xbit_r111_c110 bl[110] br[110] wl[111] vdd gnd cell_6t
Xbit_r112_c110 bl[110] br[110] wl[112] vdd gnd cell_6t
Xbit_r113_c110 bl[110] br[110] wl[113] vdd gnd cell_6t
Xbit_r114_c110 bl[110] br[110] wl[114] vdd gnd cell_6t
Xbit_r115_c110 bl[110] br[110] wl[115] vdd gnd cell_6t
Xbit_r116_c110 bl[110] br[110] wl[116] vdd gnd cell_6t
Xbit_r117_c110 bl[110] br[110] wl[117] vdd gnd cell_6t
Xbit_r118_c110 bl[110] br[110] wl[118] vdd gnd cell_6t
Xbit_r119_c110 bl[110] br[110] wl[119] vdd gnd cell_6t
Xbit_r120_c110 bl[110] br[110] wl[120] vdd gnd cell_6t
Xbit_r121_c110 bl[110] br[110] wl[121] vdd gnd cell_6t
Xbit_r122_c110 bl[110] br[110] wl[122] vdd gnd cell_6t
Xbit_r123_c110 bl[110] br[110] wl[123] vdd gnd cell_6t
Xbit_r124_c110 bl[110] br[110] wl[124] vdd gnd cell_6t
Xbit_r125_c110 bl[110] br[110] wl[125] vdd gnd cell_6t
Xbit_r126_c110 bl[110] br[110] wl[126] vdd gnd cell_6t
Xbit_r127_c110 bl[110] br[110] wl[127] vdd gnd cell_6t
Xbit_r128_c110 bl[110] br[110] wl[128] vdd gnd cell_6t
Xbit_r129_c110 bl[110] br[110] wl[129] vdd gnd cell_6t
Xbit_r130_c110 bl[110] br[110] wl[130] vdd gnd cell_6t
Xbit_r131_c110 bl[110] br[110] wl[131] vdd gnd cell_6t
Xbit_r132_c110 bl[110] br[110] wl[132] vdd gnd cell_6t
Xbit_r133_c110 bl[110] br[110] wl[133] vdd gnd cell_6t
Xbit_r134_c110 bl[110] br[110] wl[134] vdd gnd cell_6t
Xbit_r135_c110 bl[110] br[110] wl[135] vdd gnd cell_6t
Xbit_r136_c110 bl[110] br[110] wl[136] vdd gnd cell_6t
Xbit_r137_c110 bl[110] br[110] wl[137] vdd gnd cell_6t
Xbit_r138_c110 bl[110] br[110] wl[138] vdd gnd cell_6t
Xbit_r139_c110 bl[110] br[110] wl[139] vdd gnd cell_6t
Xbit_r140_c110 bl[110] br[110] wl[140] vdd gnd cell_6t
Xbit_r141_c110 bl[110] br[110] wl[141] vdd gnd cell_6t
Xbit_r142_c110 bl[110] br[110] wl[142] vdd gnd cell_6t
Xbit_r143_c110 bl[110] br[110] wl[143] vdd gnd cell_6t
Xbit_r144_c110 bl[110] br[110] wl[144] vdd gnd cell_6t
Xbit_r145_c110 bl[110] br[110] wl[145] vdd gnd cell_6t
Xbit_r146_c110 bl[110] br[110] wl[146] vdd gnd cell_6t
Xbit_r147_c110 bl[110] br[110] wl[147] vdd gnd cell_6t
Xbit_r148_c110 bl[110] br[110] wl[148] vdd gnd cell_6t
Xbit_r149_c110 bl[110] br[110] wl[149] vdd gnd cell_6t
Xbit_r150_c110 bl[110] br[110] wl[150] vdd gnd cell_6t
Xbit_r151_c110 bl[110] br[110] wl[151] vdd gnd cell_6t
Xbit_r152_c110 bl[110] br[110] wl[152] vdd gnd cell_6t
Xbit_r153_c110 bl[110] br[110] wl[153] vdd gnd cell_6t
Xbit_r154_c110 bl[110] br[110] wl[154] vdd gnd cell_6t
Xbit_r155_c110 bl[110] br[110] wl[155] vdd gnd cell_6t
Xbit_r156_c110 bl[110] br[110] wl[156] vdd gnd cell_6t
Xbit_r157_c110 bl[110] br[110] wl[157] vdd gnd cell_6t
Xbit_r158_c110 bl[110] br[110] wl[158] vdd gnd cell_6t
Xbit_r159_c110 bl[110] br[110] wl[159] vdd gnd cell_6t
Xbit_r160_c110 bl[110] br[110] wl[160] vdd gnd cell_6t
Xbit_r161_c110 bl[110] br[110] wl[161] vdd gnd cell_6t
Xbit_r162_c110 bl[110] br[110] wl[162] vdd gnd cell_6t
Xbit_r163_c110 bl[110] br[110] wl[163] vdd gnd cell_6t
Xbit_r164_c110 bl[110] br[110] wl[164] vdd gnd cell_6t
Xbit_r165_c110 bl[110] br[110] wl[165] vdd gnd cell_6t
Xbit_r166_c110 bl[110] br[110] wl[166] vdd gnd cell_6t
Xbit_r167_c110 bl[110] br[110] wl[167] vdd gnd cell_6t
Xbit_r168_c110 bl[110] br[110] wl[168] vdd gnd cell_6t
Xbit_r169_c110 bl[110] br[110] wl[169] vdd gnd cell_6t
Xbit_r170_c110 bl[110] br[110] wl[170] vdd gnd cell_6t
Xbit_r171_c110 bl[110] br[110] wl[171] vdd gnd cell_6t
Xbit_r172_c110 bl[110] br[110] wl[172] vdd gnd cell_6t
Xbit_r173_c110 bl[110] br[110] wl[173] vdd gnd cell_6t
Xbit_r174_c110 bl[110] br[110] wl[174] vdd gnd cell_6t
Xbit_r175_c110 bl[110] br[110] wl[175] vdd gnd cell_6t
Xbit_r176_c110 bl[110] br[110] wl[176] vdd gnd cell_6t
Xbit_r177_c110 bl[110] br[110] wl[177] vdd gnd cell_6t
Xbit_r178_c110 bl[110] br[110] wl[178] vdd gnd cell_6t
Xbit_r179_c110 bl[110] br[110] wl[179] vdd gnd cell_6t
Xbit_r180_c110 bl[110] br[110] wl[180] vdd gnd cell_6t
Xbit_r181_c110 bl[110] br[110] wl[181] vdd gnd cell_6t
Xbit_r182_c110 bl[110] br[110] wl[182] vdd gnd cell_6t
Xbit_r183_c110 bl[110] br[110] wl[183] vdd gnd cell_6t
Xbit_r184_c110 bl[110] br[110] wl[184] vdd gnd cell_6t
Xbit_r185_c110 bl[110] br[110] wl[185] vdd gnd cell_6t
Xbit_r186_c110 bl[110] br[110] wl[186] vdd gnd cell_6t
Xbit_r187_c110 bl[110] br[110] wl[187] vdd gnd cell_6t
Xbit_r188_c110 bl[110] br[110] wl[188] vdd gnd cell_6t
Xbit_r189_c110 bl[110] br[110] wl[189] vdd gnd cell_6t
Xbit_r190_c110 bl[110] br[110] wl[190] vdd gnd cell_6t
Xbit_r191_c110 bl[110] br[110] wl[191] vdd gnd cell_6t
Xbit_r192_c110 bl[110] br[110] wl[192] vdd gnd cell_6t
Xbit_r193_c110 bl[110] br[110] wl[193] vdd gnd cell_6t
Xbit_r194_c110 bl[110] br[110] wl[194] vdd gnd cell_6t
Xbit_r195_c110 bl[110] br[110] wl[195] vdd gnd cell_6t
Xbit_r196_c110 bl[110] br[110] wl[196] vdd gnd cell_6t
Xbit_r197_c110 bl[110] br[110] wl[197] vdd gnd cell_6t
Xbit_r198_c110 bl[110] br[110] wl[198] vdd gnd cell_6t
Xbit_r199_c110 bl[110] br[110] wl[199] vdd gnd cell_6t
Xbit_r200_c110 bl[110] br[110] wl[200] vdd gnd cell_6t
Xbit_r201_c110 bl[110] br[110] wl[201] vdd gnd cell_6t
Xbit_r202_c110 bl[110] br[110] wl[202] vdd gnd cell_6t
Xbit_r203_c110 bl[110] br[110] wl[203] vdd gnd cell_6t
Xbit_r204_c110 bl[110] br[110] wl[204] vdd gnd cell_6t
Xbit_r205_c110 bl[110] br[110] wl[205] vdd gnd cell_6t
Xbit_r206_c110 bl[110] br[110] wl[206] vdd gnd cell_6t
Xbit_r207_c110 bl[110] br[110] wl[207] vdd gnd cell_6t
Xbit_r208_c110 bl[110] br[110] wl[208] vdd gnd cell_6t
Xbit_r209_c110 bl[110] br[110] wl[209] vdd gnd cell_6t
Xbit_r210_c110 bl[110] br[110] wl[210] vdd gnd cell_6t
Xbit_r211_c110 bl[110] br[110] wl[211] vdd gnd cell_6t
Xbit_r212_c110 bl[110] br[110] wl[212] vdd gnd cell_6t
Xbit_r213_c110 bl[110] br[110] wl[213] vdd gnd cell_6t
Xbit_r214_c110 bl[110] br[110] wl[214] vdd gnd cell_6t
Xbit_r215_c110 bl[110] br[110] wl[215] vdd gnd cell_6t
Xbit_r216_c110 bl[110] br[110] wl[216] vdd gnd cell_6t
Xbit_r217_c110 bl[110] br[110] wl[217] vdd gnd cell_6t
Xbit_r218_c110 bl[110] br[110] wl[218] vdd gnd cell_6t
Xbit_r219_c110 bl[110] br[110] wl[219] vdd gnd cell_6t
Xbit_r220_c110 bl[110] br[110] wl[220] vdd gnd cell_6t
Xbit_r221_c110 bl[110] br[110] wl[221] vdd gnd cell_6t
Xbit_r222_c110 bl[110] br[110] wl[222] vdd gnd cell_6t
Xbit_r223_c110 bl[110] br[110] wl[223] vdd gnd cell_6t
Xbit_r224_c110 bl[110] br[110] wl[224] vdd gnd cell_6t
Xbit_r225_c110 bl[110] br[110] wl[225] vdd gnd cell_6t
Xbit_r226_c110 bl[110] br[110] wl[226] vdd gnd cell_6t
Xbit_r227_c110 bl[110] br[110] wl[227] vdd gnd cell_6t
Xbit_r228_c110 bl[110] br[110] wl[228] vdd gnd cell_6t
Xbit_r229_c110 bl[110] br[110] wl[229] vdd gnd cell_6t
Xbit_r230_c110 bl[110] br[110] wl[230] vdd gnd cell_6t
Xbit_r231_c110 bl[110] br[110] wl[231] vdd gnd cell_6t
Xbit_r232_c110 bl[110] br[110] wl[232] vdd gnd cell_6t
Xbit_r233_c110 bl[110] br[110] wl[233] vdd gnd cell_6t
Xbit_r234_c110 bl[110] br[110] wl[234] vdd gnd cell_6t
Xbit_r235_c110 bl[110] br[110] wl[235] vdd gnd cell_6t
Xbit_r236_c110 bl[110] br[110] wl[236] vdd gnd cell_6t
Xbit_r237_c110 bl[110] br[110] wl[237] vdd gnd cell_6t
Xbit_r238_c110 bl[110] br[110] wl[238] vdd gnd cell_6t
Xbit_r239_c110 bl[110] br[110] wl[239] vdd gnd cell_6t
Xbit_r240_c110 bl[110] br[110] wl[240] vdd gnd cell_6t
Xbit_r241_c110 bl[110] br[110] wl[241] vdd gnd cell_6t
Xbit_r242_c110 bl[110] br[110] wl[242] vdd gnd cell_6t
Xbit_r243_c110 bl[110] br[110] wl[243] vdd gnd cell_6t
Xbit_r244_c110 bl[110] br[110] wl[244] vdd gnd cell_6t
Xbit_r245_c110 bl[110] br[110] wl[245] vdd gnd cell_6t
Xbit_r246_c110 bl[110] br[110] wl[246] vdd gnd cell_6t
Xbit_r247_c110 bl[110] br[110] wl[247] vdd gnd cell_6t
Xbit_r248_c110 bl[110] br[110] wl[248] vdd gnd cell_6t
Xbit_r249_c110 bl[110] br[110] wl[249] vdd gnd cell_6t
Xbit_r250_c110 bl[110] br[110] wl[250] vdd gnd cell_6t
Xbit_r251_c110 bl[110] br[110] wl[251] vdd gnd cell_6t
Xbit_r252_c110 bl[110] br[110] wl[252] vdd gnd cell_6t
Xbit_r253_c110 bl[110] br[110] wl[253] vdd gnd cell_6t
Xbit_r254_c110 bl[110] br[110] wl[254] vdd gnd cell_6t
Xbit_r255_c110 bl[110] br[110] wl[255] vdd gnd cell_6t
Xbit_r0_c111 bl[111] br[111] wl[0] vdd gnd cell_6t
Xbit_r1_c111 bl[111] br[111] wl[1] vdd gnd cell_6t
Xbit_r2_c111 bl[111] br[111] wl[2] vdd gnd cell_6t
Xbit_r3_c111 bl[111] br[111] wl[3] vdd gnd cell_6t
Xbit_r4_c111 bl[111] br[111] wl[4] vdd gnd cell_6t
Xbit_r5_c111 bl[111] br[111] wl[5] vdd gnd cell_6t
Xbit_r6_c111 bl[111] br[111] wl[6] vdd gnd cell_6t
Xbit_r7_c111 bl[111] br[111] wl[7] vdd gnd cell_6t
Xbit_r8_c111 bl[111] br[111] wl[8] vdd gnd cell_6t
Xbit_r9_c111 bl[111] br[111] wl[9] vdd gnd cell_6t
Xbit_r10_c111 bl[111] br[111] wl[10] vdd gnd cell_6t
Xbit_r11_c111 bl[111] br[111] wl[11] vdd gnd cell_6t
Xbit_r12_c111 bl[111] br[111] wl[12] vdd gnd cell_6t
Xbit_r13_c111 bl[111] br[111] wl[13] vdd gnd cell_6t
Xbit_r14_c111 bl[111] br[111] wl[14] vdd gnd cell_6t
Xbit_r15_c111 bl[111] br[111] wl[15] vdd gnd cell_6t
Xbit_r16_c111 bl[111] br[111] wl[16] vdd gnd cell_6t
Xbit_r17_c111 bl[111] br[111] wl[17] vdd gnd cell_6t
Xbit_r18_c111 bl[111] br[111] wl[18] vdd gnd cell_6t
Xbit_r19_c111 bl[111] br[111] wl[19] vdd gnd cell_6t
Xbit_r20_c111 bl[111] br[111] wl[20] vdd gnd cell_6t
Xbit_r21_c111 bl[111] br[111] wl[21] vdd gnd cell_6t
Xbit_r22_c111 bl[111] br[111] wl[22] vdd gnd cell_6t
Xbit_r23_c111 bl[111] br[111] wl[23] vdd gnd cell_6t
Xbit_r24_c111 bl[111] br[111] wl[24] vdd gnd cell_6t
Xbit_r25_c111 bl[111] br[111] wl[25] vdd gnd cell_6t
Xbit_r26_c111 bl[111] br[111] wl[26] vdd gnd cell_6t
Xbit_r27_c111 bl[111] br[111] wl[27] vdd gnd cell_6t
Xbit_r28_c111 bl[111] br[111] wl[28] vdd gnd cell_6t
Xbit_r29_c111 bl[111] br[111] wl[29] vdd gnd cell_6t
Xbit_r30_c111 bl[111] br[111] wl[30] vdd gnd cell_6t
Xbit_r31_c111 bl[111] br[111] wl[31] vdd gnd cell_6t
Xbit_r32_c111 bl[111] br[111] wl[32] vdd gnd cell_6t
Xbit_r33_c111 bl[111] br[111] wl[33] vdd gnd cell_6t
Xbit_r34_c111 bl[111] br[111] wl[34] vdd gnd cell_6t
Xbit_r35_c111 bl[111] br[111] wl[35] vdd gnd cell_6t
Xbit_r36_c111 bl[111] br[111] wl[36] vdd gnd cell_6t
Xbit_r37_c111 bl[111] br[111] wl[37] vdd gnd cell_6t
Xbit_r38_c111 bl[111] br[111] wl[38] vdd gnd cell_6t
Xbit_r39_c111 bl[111] br[111] wl[39] vdd gnd cell_6t
Xbit_r40_c111 bl[111] br[111] wl[40] vdd gnd cell_6t
Xbit_r41_c111 bl[111] br[111] wl[41] vdd gnd cell_6t
Xbit_r42_c111 bl[111] br[111] wl[42] vdd gnd cell_6t
Xbit_r43_c111 bl[111] br[111] wl[43] vdd gnd cell_6t
Xbit_r44_c111 bl[111] br[111] wl[44] vdd gnd cell_6t
Xbit_r45_c111 bl[111] br[111] wl[45] vdd gnd cell_6t
Xbit_r46_c111 bl[111] br[111] wl[46] vdd gnd cell_6t
Xbit_r47_c111 bl[111] br[111] wl[47] vdd gnd cell_6t
Xbit_r48_c111 bl[111] br[111] wl[48] vdd gnd cell_6t
Xbit_r49_c111 bl[111] br[111] wl[49] vdd gnd cell_6t
Xbit_r50_c111 bl[111] br[111] wl[50] vdd gnd cell_6t
Xbit_r51_c111 bl[111] br[111] wl[51] vdd gnd cell_6t
Xbit_r52_c111 bl[111] br[111] wl[52] vdd gnd cell_6t
Xbit_r53_c111 bl[111] br[111] wl[53] vdd gnd cell_6t
Xbit_r54_c111 bl[111] br[111] wl[54] vdd gnd cell_6t
Xbit_r55_c111 bl[111] br[111] wl[55] vdd gnd cell_6t
Xbit_r56_c111 bl[111] br[111] wl[56] vdd gnd cell_6t
Xbit_r57_c111 bl[111] br[111] wl[57] vdd gnd cell_6t
Xbit_r58_c111 bl[111] br[111] wl[58] vdd gnd cell_6t
Xbit_r59_c111 bl[111] br[111] wl[59] vdd gnd cell_6t
Xbit_r60_c111 bl[111] br[111] wl[60] vdd gnd cell_6t
Xbit_r61_c111 bl[111] br[111] wl[61] vdd gnd cell_6t
Xbit_r62_c111 bl[111] br[111] wl[62] vdd gnd cell_6t
Xbit_r63_c111 bl[111] br[111] wl[63] vdd gnd cell_6t
Xbit_r64_c111 bl[111] br[111] wl[64] vdd gnd cell_6t
Xbit_r65_c111 bl[111] br[111] wl[65] vdd gnd cell_6t
Xbit_r66_c111 bl[111] br[111] wl[66] vdd gnd cell_6t
Xbit_r67_c111 bl[111] br[111] wl[67] vdd gnd cell_6t
Xbit_r68_c111 bl[111] br[111] wl[68] vdd gnd cell_6t
Xbit_r69_c111 bl[111] br[111] wl[69] vdd gnd cell_6t
Xbit_r70_c111 bl[111] br[111] wl[70] vdd gnd cell_6t
Xbit_r71_c111 bl[111] br[111] wl[71] vdd gnd cell_6t
Xbit_r72_c111 bl[111] br[111] wl[72] vdd gnd cell_6t
Xbit_r73_c111 bl[111] br[111] wl[73] vdd gnd cell_6t
Xbit_r74_c111 bl[111] br[111] wl[74] vdd gnd cell_6t
Xbit_r75_c111 bl[111] br[111] wl[75] vdd gnd cell_6t
Xbit_r76_c111 bl[111] br[111] wl[76] vdd gnd cell_6t
Xbit_r77_c111 bl[111] br[111] wl[77] vdd gnd cell_6t
Xbit_r78_c111 bl[111] br[111] wl[78] vdd gnd cell_6t
Xbit_r79_c111 bl[111] br[111] wl[79] vdd gnd cell_6t
Xbit_r80_c111 bl[111] br[111] wl[80] vdd gnd cell_6t
Xbit_r81_c111 bl[111] br[111] wl[81] vdd gnd cell_6t
Xbit_r82_c111 bl[111] br[111] wl[82] vdd gnd cell_6t
Xbit_r83_c111 bl[111] br[111] wl[83] vdd gnd cell_6t
Xbit_r84_c111 bl[111] br[111] wl[84] vdd gnd cell_6t
Xbit_r85_c111 bl[111] br[111] wl[85] vdd gnd cell_6t
Xbit_r86_c111 bl[111] br[111] wl[86] vdd gnd cell_6t
Xbit_r87_c111 bl[111] br[111] wl[87] vdd gnd cell_6t
Xbit_r88_c111 bl[111] br[111] wl[88] vdd gnd cell_6t
Xbit_r89_c111 bl[111] br[111] wl[89] vdd gnd cell_6t
Xbit_r90_c111 bl[111] br[111] wl[90] vdd gnd cell_6t
Xbit_r91_c111 bl[111] br[111] wl[91] vdd gnd cell_6t
Xbit_r92_c111 bl[111] br[111] wl[92] vdd gnd cell_6t
Xbit_r93_c111 bl[111] br[111] wl[93] vdd gnd cell_6t
Xbit_r94_c111 bl[111] br[111] wl[94] vdd gnd cell_6t
Xbit_r95_c111 bl[111] br[111] wl[95] vdd gnd cell_6t
Xbit_r96_c111 bl[111] br[111] wl[96] vdd gnd cell_6t
Xbit_r97_c111 bl[111] br[111] wl[97] vdd gnd cell_6t
Xbit_r98_c111 bl[111] br[111] wl[98] vdd gnd cell_6t
Xbit_r99_c111 bl[111] br[111] wl[99] vdd gnd cell_6t
Xbit_r100_c111 bl[111] br[111] wl[100] vdd gnd cell_6t
Xbit_r101_c111 bl[111] br[111] wl[101] vdd gnd cell_6t
Xbit_r102_c111 bl[111] br[111] wl[102] vdd gnd cell_6t
Xbit_r103_c111 bl[111] br[111] wl[103] vdd gnd cell_6t
Xbit_r104_c111 bl[111] br[111] wl[104] vdd gnd cell_6t
Xbit_r105_c111 bl[111] br[111] wl[105] vdd gnd cell_6t
Xbit_r106_c111 bl[111] br[111] wl[106] vdd gnd cell_6t
Xbit_r107_c111 bl[111] br[111] wl[107] vdd gnd cell_6t
Xbit_r108_c111 bl[111] br[111] wl[108] vdd gnd cell_6t
Xbit_r109_c111 bl[111] br[111] wl[109] vdd gnd cell_6t
Xbit_r110_c111 bl[111] br[111] wl[110] vdd gnd cell_6t
Xbit_r111_c111 bl[111] br[111] wl[111] vdd gnd cell_6t
Xbit_r112_c111 bl[111] br[111] wl[112] vdd gnd cell_6t
Xbit_r113_c111 bl[111] br[111] wl[113] vdd gnd cell_6t
Xbit_r114_c111 bl[111] br[111] wl[114] vdd gnd cell_6t
Xbit_r115_c111 bl[111] br[111] wl[115] vdd gnd cell_6t
Xbit_r116_c111 bl[111] br[111] wl[116] vdd gnd cell_6t
Xbit_r117_c111 bl[111] br[111] wl[117] vdd gnd cell_6t
Xbit_r118_c111 bl[111] br[111] wl[118] vdd gnd cell_6t
Xbit_r119_c111 bl[111] br[111] wl[119] vdd gnd cell_6t
Xbit_r120_c111 bl[111] br[111] wl[120] vdd gnd cell_6t
Xbit_r121_c111 bl[111] br[111] wl[121] vdd gnd cell_6t
Xbit_r122_c111 bl[111] br[111] wl[122] vdd gnd cell_6t
Xbit_r123_c111 bl[111] br[111] wl[123] vdd gnd cell_6t
Xbit_r124_c111 bl[111] br[111] wl[124] vdd gnd cell_6t
Xbit_r125_c111 bl[111] br[111] wl[125] vdd gnd cell_6t
Xbit_r126_c111 bl[111] br[111] wl[126] vdd gnd cell_6t
Xbit_r127_c111 bl[111] br[111] wl[127] vdd gnd cell_6t
Xbit_r128_c111 bl[111] br[111] wl[128] vdd gnd cell_6t
Xbit_r129_c111 bl[111] br[111] wl[129] vdd gnd cell_6t
Xbit_r130_c111 bl[111] br[111] wl[130] vdd gnd cell_6t
Xbit_r131_c111 bl[111] br[111] wl[131] vdd gnd cell_6t
Xbit_r132_c111 bl[111] br[111] wl[132] vdd gnd cell_6t
Xbit_r133_c111 bl[111] br[111] wl[133] vdd gnd cell_6t
Xbit_r134_c111 bl[111] br[111] wl[134] vdd gnd cell_6t
Xbit_r135_c111 bl[111] br[111] wl[135] vdd gnd cell_6t
Xbit_r136_c111 bl[111] br[111] wl[136] vdd gnd cell_6t
Xbit_r137_c111 bl[111] br[111] wl[137] vdd gnd cell_6t
Xbit_r138_c111 bl[111] br[111] wl[138] vdd gnd cell_6t
Xbit_r139_c111 bl[111] br[111] wl[139] vdd gnd cell_6t
Xbit_r140_c111 bl[111] br[111] wl[140] vdd gnd cell_6t
Xbit_r141_c111 bl[111] br[111] wl[141] vdd gnd cell_6t
Xbit_r142_c111 bl[111] br[111] wl[142] vdd gnd cell_6t
Xbit_r143_c111 bl[111] br[111] wl[143] vdd gnd cell_6t
Xbit_r144_c111 bl[111] br[111] wl[144] vdd gnd cell_6t
Xbit_r145_c111 bl[111] br[111] wl[145] vdd gnd cell_6t
Xbit_r146_c111 bl[111] br[111] wl[146] vdd gnd cell_6t
Xbit_r147_c111 bl[111] br[111] wl[147] vdd gnd cell_6t
Xbit_r148_c111 bl[111] br[111] wl[148] vdd gnd cell_6t
Xbit_r149_c111 bl[111] br[111] wl[149] vdd gnd cell_6t
Xbit_r150_c111 bl[111] br[111] wl[150] vdd gnd cell_6t
Xbit_r151_c111 bl[111] br[111] wl[151] vdd gnd cell_6t
Xbit_r152_c111 bl[111] br[111] wl[152] vdd gnd cell_6t
Xbit_r153_c111 bl[111] br[111] wl[153] vdd gnd cell_6t
Xbit_r154_c111 bl[111] br[111] wl[154] vdd gnd cell_6t
Xbit_r155_c111 bl[111] br[111] wl[155] vdd gnd cell_6t
Xbit_r156_c111 bl[111] br[111] wl[156] vdd gnd cell_6t
Xbit_r157_c111 bl[111] br[111] wl[157] vdd gnd cell_6t
Xbit_r158_c111 bl[111] br[111] wl[158] vdd gnd cell_6t
Xbit_r159_c111 bl[111] br[111] wl[159] vdd gnd cell_6t
Xbit_r160_c111 bl[111] br[111] wl[160] vdd gnd cell_6t
Xbit_r161_c111 bl[111] br[111] wl[161] vdd gnd cell_6t
Xbit_r162_c111 bl[111] br[111] wl[162] vdd gnd cell_6t
Xbit_r163_c111 bl[111] br[111] wl[163] vdd gnd cell_6t
Xbit_r164_c111 bl[111] br[111] wl[164] vdd gnd cell_6t
Xbit_r165_c111 bl[111] br[111] wl[165] vdd gnd cell_6t
Xbit_r166_c111 bl[111] br[111] wl[166] vdd gnd cell_6t
Xbit_r167_c111 bl[111] br[111] wl[167] vdd gnd cell_6t
Xbit_r168_c111 bl[111] br[111] wl[168] vdd gnd cell_6t
Xbit_r169_c111 bl[111] br[111] wl[169] vdd gnd cell_6t
Xbit_r170_c111 bl[111] br[111] wl[170] vdd gnd cell_6t
Xbit_r171_c111 bl[111] br[111] wl[171] vdd gnd cell_6t
Xbit_r172_c111 bl[111] br[111] wl[172] vdd gnd cell_6t
Xbit_r173_c111 bl[111] br[111] wl[173] vdd gnd cell_6t
Xbit_r174_c111 bl[111] br[111] wl[174] vdd gnd cell_6t
Xbit_r175_c111 bl[111] br[111] wl[175] vdd gnd cell_6t
Xbit_r176_c111 bl[111] br[111] wl[176] vdd gnd cell_6t
Xbit_r177_c111 bl[111] br[111] wl[177] vdd gnd cell_6t
Xbit_r178_c111 bl[111] br[111] wl[178] vdd gnd cell_6t
Xbit_r179_c111 bl[111] br[111] wl[179] vdd gnd cell_6t
Xbit_r180_c111 bl[111] br[111] wl[180] vdd gnd cell_6t
Xbit_r181_c111 bl[111] br[111] wl[181] vdd gnd cell_6t
Xbit_r182_c111 bl[111] br[111] wl[182] vdd gnd cell_6t
Xbit_r183_c111 bl[111] br[111] wl[183] vdd gnd cell_6t
Xbit_r184_c111 bl[111] br[111] wl[184] vdd gnd cell_6t
Xbit_r185_c111 bl[111] br[111] wl[185] vdd gnd cell_6t
Xbit_r186_c111 bl[111] br[111] wl[186] vdd gnd cell_6t
Xbit_r187_c111 bl[111] br[111] wl[187] vdd gnd cell_6t
Xbit_r188_c111 bl[111] br[111] wl[188] vdd gnd cell_6t
Xbit_r189_c111 bl[111] br[111] wl[189] vdd gnd cell_6t
Xbit_r190_c111 bl[111] br[111] wl[190] vdd gnd cell_6t
Xbit_r191_c111 bl[111] br[111] wl[191] vdd gnd cell_6t
Xbit_r192_c111 bl[111] br[111] wl[192] vdd gnd cell_6t
Xbit_r193_c111 bl[111] br[111] wl[193] vdd gnd cell_6t
Xbit_r194_c111 bl[111] br[111] wl[194] vdd gnd cell_6t
Xbit_r195_c111 bl[111] br[111] wl[195] vdd gnd cell_6t
Xbit_r196_c111 bl[111] br[111] wl[196] vdd gnd cell_6t
Xbit_r197_c111 bl[111] br[111] wl[197] vdd gnd cell_6t
Xbit_r198_c111 bl[111] br[111] wl[198] vdd gnd cell_6t
Xbit_r199_c111 bl[111] br[111] wl[199] vdd gnd cell_6t
Xbit_r200_c111 bl[111] br[111] wl[200] vdd gnd cell_6t
Xbit_r201_c111 bl[111] br[111] wl[201] vdd gnd cell_6t
Xbit_r202_c111 bl[111] br[111] wl[202] vdd gnd cell_6t
Xbit_r203_c111 bl[111] br[111] wl[203] vdd gnd cell_6t
Xbit_r204_c111 bl[111] br[111] wl[204] vdd gnd cell_6t
Xbit_r205_c111 bl[111] br[111] wl[205] vdd gnd cell_6t
Xbit_r206_c111 bl[111] br[111] wl[206] vdd gnd cell_6t
Xbit_r207_c111 bl[111] br[111] wl[207] vdd gnd cell_6t
Xbit_r208_c111 bl[111] br[111] wl[208] vdd gnd cell_6t
Xbit_r209_c111 bl[111] br[111] wl[209] vdd gnd cell_6t
Xbit_r210_c111 bl[111] br[111] wl[210] vdd gnd cell_6t
Xbit_r211_c111 bl[111] br[111] wl[211] vdd gnd cell_6t
Xbit_r212_c111 bl[111] br[111] wl[212] vdd gnd cell_6t
Xbit_r213_c111 bl[111] br[111] wl[213] vdd gnd cell_6t
Xbit_r214_c111 bl[111] br[111] wl[214] vdd gnd cell_6t
Xbit_r215_c111 bl[111] br[111] wl[215] vdd gnd cell_6t
Xbit_r216_c111 bl[111] br[111] wl[216] vdd gnd cell_6t
Xbit_r217_c111 bl[111] br[111] wl[217] vdd gnd cell_6t
Xbit_r218_c111 bl[111] br[111] wl[218] vdd gnd cell_6t
Xbit_r219_c111 bl[111] br[111] wl[219] vdd gnd cell_6t
Xbit_r220_c111 bl[111] br[111] wl[220] vdd gnd cell_6t
Xbit_r221_c111 bl[111] br[111] wl[221] vdd gnd cell_6t
Xbit_r222_c111 bl[111] br[111] wl[222] vdd gnd cell_6t
Xbit_r223_c111 bl[111] br[111] wl[223] vdd gnd cell_6t
Xbit_r224_c111 bl[111] br[111] wl[224] vdd gnd cell_6t
Xbit_r225_c111 bl[111] br[111] wl[225] vdd gnd cell_6t
Xbit_r226_c111 bl[111] br[111] wl[226] vdd gnd cell_6t
Xbit_r227_c111 bl[111] br[111] wl[227] vdd gnd cell_6t
Xbit_r228_c111 bl[111] br[111] wl[228] vdd gnd cell_6t
Xbit_r229_c111 bl[111] br[111] wl[229] vdd gnd cell_6t
Xbit_r230_c111 bl[111] br[111] wl[230] vdd gnd cell_6t
Xbit_r231_c111 bl[111] br[111] wl[231] vdd gnd cell_6t
Xbit_r232_c111 bl[111] br[111] wl[232] vdd gnd cell_6t
Xbit_r233_c111 bl[111] br[111] wl[233] vdd gnd cell_6t
Xbit_r234_c111 bl[111] br[111] wl[234] vdd gnd cell_6t
Xbit_r235_c111 bl[111] br[111] wl[235] vdd gnd cell_6t
Xbit_r236_c111 bl[111] br[111] wl[236] vdd gnd cell_6t
Xbit_r237_c111 bl[111] br[111] wl[237] vdd gnd cell_6t
Xbit_r238_c111 bl[111] br[111] wl[238] vdd gnd cell_6t
Xbit_r239_c111 bl[111] br[111] wl[239] vdd gnd cell_6t
Xbit_r240_c111 bl[111] br[111] wl[240] vdd gnd cell_6t
Xbit_r241_c111 bl[111] br[111] wl[241] vdd gnd cell_6t
Xbit_r242_c111 bl[111] br[111] wl[242] vdd gnd cell_6t
Xbit_r243_c111 bl[111] br[111] wl[243] vdd gnd cell_6t
Xbit_r244_c111 bl[111] br[111] wl[244] vdd gnd cell_6t
Xbit_r245_c111 bl[111] br[111] wl[245] vdd gnd cell_6t
Xbit_r246_c111 bl[111] br[111] wl[246] vdd gnd cell_6t
Xbit_r247_c111 bl[111] br[111] wl[247] vdd gnd cell_6t
Xbit_r248_c111 bl[111] br[111] wl[248] vdd gnd cell_6t
Xbit_r249_c111 bl[111] br[111] wl[249] vdd gnd cell_6t
Xbit_r250_c111 bl[111] br[111] wl[250] vdd gnd cell_6t
Xbit_r251_c111 bl[111] br[111] wl[251] vdd gnd cell_6t
Xbit_r252_c111 bl[111] br[111] wl[252] vdd gnd cell_6t
Xbit_r253_c111 bl[111] br[111] wl[253] vdd gnd cell_6t
Xbit_r254_c111 bl[111] br[111] wl[254] vdd gnd cell_6t
Xbit_r255_c111 bl[111] br[111] wl[255] vdd gnd cell_6t
Xbit_r0_c112 bl[112] br[112] wl[0] vdd gnd cell_6t
Xbit_r1_c112 bl[112] br[112] wl[1] vdd gnd cell_6t
Xbit_r2_c112 bl[112] br[112] wl[2] vdd gnd cell_6t
Xbit_r3_c112 bl[112] br[112] wl[3] vdd gnd cell_6t
Xbit_r4_c112 bl[112] br[112] wl[4] vdd gnd cell_6t
Xbit_r5_c112 bl[112] br[112] wl[5] vdd gnd cell_6t
Xbit_r6_c112 bl[112] br[112] wl[6] vdd gnd cell_6t
Xbit_r7_c112 bl[112] br[112] wl[7] vdd gnd cell_6t
Xbit_r8_c112 bl[112] br[112] wl[8] vdd gnd cell_6t
Xbit_r9_c112 bl[112] br[112] wl[9] vdd gnd cell_6t
Xbit_r10_c112 bl[112] br[112] wl[10] vdd gnd cell_6t
Xbit_r11_c112 bl[112] br[112] wl[11] vdd gnd cell_6t
Xbit_r12_c112 bl[112] br[112] wl[12] vdd gnd cell_6t
Xbit_r13_c112 bl[112] br[112] wl[13] vdd gnd cell_6t
Xbit_r14_c112 bl[112] br[112] wl[14] vdd gnd cell_6t
Xbit_r15_c112 bl[112] br[112] wl[15] vdd gnd cell_6t
Xbit_r16_c112 bl[112] br[112] wl[16] vdd gnd cell_6t
Xbit_r17_c112 bl[112] br[112] wl[17] vdd gnd cell_6t
Xbit_r18_c112 bl[112] br[112] wl[18] vdd gnd cell_6t
Xbit_r19_c112 bl[112] br[112] wl[19] vdd gnd cell_6t
Xbit_r20_c112 bl[112] br[112] wl[20] vdd gnd cell_6t
Xbit_r21_c112 bl[112] br[112] wl[21] vdd gnd cell_6t
Xbit_r22_c112 bl[112] br[112] wl[22] vdd gnd cell_6t
Xbit_r23_c112 bl[112] br[112] wl[23] vdd gnd cell_6t
Xbit_r24_c112 bl[112] br[112] wl[24] vdd gnd cell_6t
Xbit_r25_c112 bl[112] br[112] wl[25] vdd gnd cell_6t
Xbit_r26_c112 bl[112] br[112] wl[26] vdd gnd cell_6t
Xbit_r27_c112 bl[112] br[112] wl[27] vdd gnd cell_6t
Xbit_r28_c112 bl[112] br[112] wl[28] vdd gnd cell_6t
Xbit_r29_c112 bl[112] br[112] wl[29] vdd gnd cell_6t
Xbit_r30_c112 bl[112] br[112] wl[30] vdd gnd cell_6t
Xbit_r31_c112 bl[112] br[112] wl[31] vdd gnd cell_6t
Xbit_r32_c112 bl[112] br[112] wl[32] vdd gnd cell_6t
Xbit_r33_c112 bl[112] br[112] wl[33] vdd gnd cell_6t
Xbit_r34_c112 bl[112] br[112] wl[34] vdd gnd cell_6t
Xbit_r35_c112 bl[112] br[112] wl[35] vdd gnd cell_6t
Xbit_r36_c112 bl[112] br[112] wl[36] vdd gnd cell_6t
Xbit_r37_c112 bl[112] br[112] wl[37] vdd gnd cell_6t
Xbit_r38_c112 bl[112] br[112] wl[38] vdd gnd cell_6t
Xbit_r39_c112 bl[112] br[112] wl[39] vdd gnd cell_6t
Xbit_r40_c112 bl[112] br[112] wl[40] vdd gnd cell_6t
Xbit_r41_c112 bl[112] br[112] wl[41] vdd gnd cell_6t
Xbit_r42_c112 bl[112] br[112] wl[42] vdd gnd cell_6t
Xbit_r43_c112 bl[112] br[112] wl[43] vdd gnd cell_6t
Xbit_r44_c112 bl[112] br[112] wl[44] vdd gnd cell_6t
Xbit_r45_c112 bl[112] br[112] wl[45] vdd gnd cell_6t
Xbit_r46_c112 bl[112] br[112] wl[46] vdd gnd cell_6t
Xbit_r47_c112 bl[112] br[112] wl[47] vdd gnd cell_6t
Xbit_r48_c112 bl[112] br[112] wl[48] vdd gnd cell_6t
Xbit_r49_c112 bl[112] br[112] wl[49] vdd gnd cell_6t
Xbit_r50_c112 bl[112] br[112] wl[50] vdd gnd cell_6t
Xbit_r51_c112 bl[112] br[112] wl[51] vdd gnd cell_6t
Xbit_r52_c112 bl[112] br[112] wl[52] vdd gnd cell_6t
Xbit_r53_c112 bl[112] br[112] wl[53] vdd gnd cell_6t
Xbit_r54_c112 bl[112] br[112] wl[54] vdd gnd cell_6t
Xbit_r55_c112 bl[112] br[112] wl[55] vdd gnd cell_6t
Xbit_r56_c112 bl[112] br[112] wl[56] vdd gnd cell_6t
Xbit_r57_c112 bl[112] br[112] wl[57] vdd gnd cell_6t
Xbit_r58_c112 bl[112] br[112] wl[58] vdd gnd cell_6t
Xbit_r59_c112 bl[112] br[112] wl[59] vdd gnd cell_6t
Xbit_r60_c112 bl[112] br[112] wl[60] vdd gnd cell_6t
Xbit_r61_c112 bl[112] br[112] wl[61] vdd gnd cell_6t
Xbit_r62_c112 bl[112] br[112] wl[62] vdd gnd cell_6t
Xbit_r63_c112 bl[112] br[112] wl[63] vdd gnd cell_6t
Xbit_r64_c112 bl[112] br[112] wl[64] vdd gnd cell_6t
Xbit_r65_c112 bl[112] br[112] wl[65] vdd gnd cell_6t
Xbit_r66_c112 bl[112] br[112] wl[66] vdd gnd cell_6t
Xbit_r67_c112 bl[112] br[112] wl[67] vdd gnd cell_6t
Xbit_r68_c112 bl[112] br[112] wl[68] vdd gnd cell_6t
Xbit_r69_c112 bl[112] br[112] wl[69] vdd gnd cell_6t
Xbit_r70_c112 bl[112] br[112] wl[70] vdd gnd cell_6t
Xbit_r71_c112 bl[112] br[112] wl[71] vdd gnd cell_6t
Xbit_r72_c112 bl[112] br[112] wl[72] vdd gnd cell_6t
Xbit_r73_c112 bl[112] br[112] wl[73] vdd gnd cell_6t
Xbit_r74_c112 bl[112] br[112] wl[74] vdd gnd cell_6t
Xbit_r75_c112 bl[112] br[112] wl[75] vdd gnd cell_6t
Xbit_r76_c112 bl[112] br[112] wl[76] vdd gnd cell_6t
Xbit_r77_c112 bl[112] br[112] wl[77] vdd gnd cell_6t
Xbit_r78_c112 bl[112] br[112] wl[78] vdd gnd cell_6t
Xbit_r79_c112 bl[112] br[112] wl[79] vdd gnd cell_6t
Xbit_r80_c112 bl[112] br[112] wl[80] vdd gnd cell_6t
Xbit_r81_c112 bl[112] br[112] wl[81] vdd gnd cell_6t
Xbit_r82_c112 bl[112] br[112] wl[82] vdd gnd cell_6t
Xbit_r83_c112 bl[112] br[112] wl[83] vdd gnd cell_6t
Xbit_r84_c112 bl[112] br[112] wl[84] vdd gnd cell_6t
Xbit_r85_c112 bl[112] br[112] wl[85] vdd gnd cell_6t
Xbit_r86_c112 bl[112] br[112] wl[86] vdd gnd cell_6t
Xbit_r87_c112 bl[112] br[112] wl[87] vdd gnd cell_6t
Xbit_r88_c112 bl[112] br[112] wl[88] vdd gnd cell_6t
Xbit_r89_c112 bl[112] br[112] wl[89] vdd gnd cell_6t
Xbit_r90_c112 bl[112] br[112] wl[90] vdd gnd cell_6t
Xbit_r91_c112 bl[112] br[112] wl[91] vdd gnd cell_6t
Xbit_r92_c112 bl[112] br[112] wl[92] vdd gnd cell_6t
Xbit_r93_c112 bl[112] br[112] wl[93] vdd gnd cell_6t
Xbit_r94_c112 bl[112] br[112] wl[94] vdd gnd cell_6t
Xbit_r95_c112 bl[112] br[112] wl[95] vdd gnd cell_6t
Xbit_r96_c112 bl[112] br[112] wl[96] vdd gnd cell_6t
Xbit_r97_c112 bl[112] br[112] wl[97] vdd gnd cell_6t
Xbit_r98_c112 bl[112] br[112] wl[98] vdd gnd cell_6t
Xbit_r99_c112 bl[112] br[112] wl[99] vdd gnd cell_6t
Xbit_r100_c112 bl[112] br[112] wl[100] vdd gnd cell_6t
Xbit_r101_c112 bl[112] br[112] wl[101] vdd gnd cell_6t
Xbit_r102_c112 bl[112] br[112] wl[102] vdd gnd cell_6t
Xbit_r103_c112 bl[112] br[112] wl[103] vdd gnd cell_6t
Xbit_r104_c112 bl[112] br[112] wl[104] vdd gnd cell_6t
Xbit_r105_c112 bl[112] br[112] wl[105] vdd gnd cell_6t
Xbit_r106_c112 bl[112] br[112] wl[106] vdd gnd cell_6t
Xbit_r107_c112 bl[112] br[112] wl[107] vdd gnd cell_6t
Xbit_r108_c112 bl[112] br[112] wl[108] vdd gnd cell_6t
Xbit_r109_c112 bl[112] br[112] wl[109] vdd gnd cell_6t
Xbit_r110_c112 bl[112] br[112] wl[110] vdd gnd cell_6t
Xbit_r111_c112 bl[112] br[112] wl[111] vdd gnd cell_6t
Xbit_r112_c112 bl[112] br[112] wl[112] vdd gnd cell_6t
Xbit_r113_c112 bl[112] br[112] wl[113] vdd gnd cell_6t
Xbit_r114_c112 bl[112] br[112] wl[114] vdd gnd cell_6t
Xbit_r115_c112 bl[112] br[112] wl[115] vdd gnd cell_6t
Xbit_r116_c112 bl[112] br[112] wl[116] vdd gnd cell_6t
Xbit_r117_c112 bl[112] br[112] wl[117] vdd gnd cell_6t
Xbit_r118_c112 bl[112] br[112] wl[118] vdd gnd cell_6t
Xbit_r119_c112 bl[112] br[112] wl[119] vdd gnd cell_6t
Xbit_r120_c112 bl[112] br[112] wl[120] vdd gnd cell_6t
Xbit_r121_c112 bl[112] br[112] wl[121] vdd gnd cell_6t
Xbit_r122_c112 bl[112] br[112] wl[122] vdd gnd cell_6t
Xbit_r123_c112 bl[112] br[112] wl[123] vdd gnd cell_6t
Xbit_r124_c112 bl[112] br[112] wl[124] vdd gnd cell_6t
Xbit_r125_c112 bl[112] br[112] wl[125] vdd gnd cell_6t
Xbit_r126_c112 bl[112] br[112] wl[126] vdd gnd cell_6t
Xbit_r127_c112 bl[112] br[112] wl[127] vdd gnd cell_6t
Xbit_r128_c112 bl[112] br[112] wl[128] vdd gnd cell_6t
Xbit_r129_c112 bl[112] br[112] wl[129] vdd gnd cell_6t
Xbit_r130_c112 bl[112] br[112] wl[130] vdd gnd cell_6t
Xbit_r131_c112 bl[112] br[112] wl[131] vdd gnd cell_6t
Xbit_r132_c112 bl[112] br[112] wl[132] vdd gnd cell_6t
Xbit_r133_c112 bl[112] br[112] wl[133] vdd gnd cell_6t
Xbit_r134_c112 bl[112] br[112] wl[134] vdd gnd cell_6t
Xbit_r135_c112 bl[112] br[112] wl[135] vdd gnd cell_6t
Xbit_r136_c112 bl[112] br[112] wl[136] vdd gnd cell_6t
Xbit_r137_c112 bl[112] br[112] wl[137] vdd gnd cell_6t
Xbit_r138_c112 bl[112] br[112] wl[138] vdd gnd cell_6t
Xbit_r139_c112 bl[112] br[112] wl[139] vdd gnd cell_6t
Xbit_r140_c112 bl[112] br[112] wl[140] vdd gnd cell_6t
Xbit_r141_c112 bl[112] br[112] wl[141] vdd gnd cell_6t
Xbit_r142_c112 bl[112] br[112] wl[142] vdd gnd cell_6t
Xbit_r143_c112 bl[112] br[112] wl[143] vdd gnd cell_6t
Xbit_r144_c112 bl[112] br[112] wl[144] vdd gnd cell_6t
Xbit_r145_c112 bl[112] br[112] wl[145] vdd gnd cell_6t
Xbit_r146_c112 bl[112] br[112] wl[146] vdd gnd cell_6t
Xbit_r147_c112 bl[112] br[112] wl[147] vdd gnd cell_6t
Xbit_r148_c112 bl[112] br[112] wl[148] vdd gnd cell_6t
Xbit_r149_c112 bl[112] br[112] wl[149] vdd gnd cell_6t
Xbit_r150_c112 bl[112] br[112] wl[150] vdd gnd cell_6t
Xbit_r151_c112 bl[112] br[112] wl[151] vdd gnd cell_6t
Xbit_r152_c112 bl[112] br[112] wl[152] vdd gnd cell_6t
Xbit_r153_c112 bl[112] br[112] wl[153] vdd gnd cell_6t
Xbit_r154_c112 bl[112] br[112] wl[154] vdd gnd cell_6t
Xbit_r155_c112 bl[112] br[112] wl[155] vdd gnd cell_6t
Xbit_r156_c112 bl[112] br[112] wl[156] vdd gnd cell_6t
Xbit_r157_c112 bl[112] br[112] wl[157] vdd gnd cell_6t
Xbit_r158_c112 bl[112] br[112] wl[158] vdd gnd cell_6t
Xbit_r159_c112 bl[112] br[112] wl[159] vdd gnd cell_6t
Xbit_r160_c112 bl[112] br[112] wl[160] vdd gnd cell_6t
Xbit_r161_c112 bl[112] br[112] wl[161] vdd gnd cell_6t
Xbit_r162_c112 bl[112] br[112] wl[162] vdd gnd cell_6t
Xbit_r163_c112 bl[112] br[112] wl[163] vdd gnd cell_6t
Xbit_r164_c112 bl[112] br[112] wl[164] vdd gnd cell_6t
Xbit_r165_c112 bl[112] br[112] wl[165] vdd gnd cell_6t
Xbit_r166_c112 bl[112] br[112] wl[166] vdd gnd cell_6t
Xbit_r167_c112 bl[112] br[112] wl[167] vdd gnd cell_6t
Xbit_r168_c112 bl[112] br[112] wl[168] vdd gnd cell_6t
Xbit_r169_c112 bl[112] br[112] wl[169] vdd gnd cell_6t
Xbit_r170_c112 bl[112] br[112] wl[170] vdd gnd cell_6t
Xbit_r171_c112 bl[112] br[112] wl[171] vdd gnd cell_6t
Xbit_r172_c112 bl[112] br[112] wl[172] vdd gnd cell_6t
Xbit_r173_c112 bl[112] br[112] wl[173] vdd gnd cell_6t
Xbit_r174_c112 bl[112] br[112] wl[174] vdd gnd cell_6t
Xbit_r175_c112 bl[112] br[112] wl[175] vdd gnd cell_6t
Xbit_r176_c112 bl[112] br[112] wl[176] vdd gnd cell_6t
Xbit_r177_c112 bl[112] br[112] wl[177] vdd gnd cell_6t
Xbit_r178_c112 bl[112] br[112] wl[178] vdd gnd cell_6t
Xbit_r179_c112 bl[112] br[112] wl[179] vdd gnd cell_6t
Xbit_r180_c112 bl[112] br[112] wl[180] vdd gnd cell_6t
Xbit_r181_c112 bl[112] br[112] wl[181] vdd gnd cell_6t
Xbit_r182_c112 bl[112] br[112] wl[182] vdd gnd cell_6t
Xbit_r183_c112 bl[112] br[112] wl[183] vdd gnd cell_6t
Xbit_r184_c112 bl[112] br[112] wl[184] vdd gnd cell_6t
Xbit_r185_c112 bl[112] br[112] wl[185] vdd gnd cell_6t
Xbit_r186_c112 bl[112] br[112] wl[186] vdd gnd cell_6t
Xbit_r187_c112 bl[112] br[112] wl[187] vdd gnd cell_6t
Xbit_r188_c112 bl[112] br[112] wl[188] vdd gnd cell_6t
Xbit_r189_c112 bl[112] br[112] wl[189] vdd gnd cell_6t
Xbit_r190_c112 bl[112] br[112] wl[190] vdd gnd cell_6t
Xbit_r191_c112 bl[112] br[112] wl[191] vdd gnd cell_6t
Xbit_r192_c112 bl[112] br[112] wl[192] vdd gnd cell_6t
Xbit_r193_c112 bl[112] br[112] wl[193] vdd gnd cell_6t
Xbit_r194_c112 bl[112] br[112] wl[194] vdd gnd cell_6t
Xbit_r195_c112 bl[112] br[112] wl[195] vdd gnd cell_6t
Xbit_r196_c112 bl[112] br[112] wl[196] vdd gnd cell_6t
Xbit_r197_c112 bl[112] br[112] wl[197] vdd gnd cell_6t
Xbit_r198_c112 bl[112] br[112] wl[198] vdd gnd cell_6t
Xbit_r199_c112 bl[112] br[112] wl[199] vdd gnd cell_6t
Xbit_r200_c112 bl[112] br[112] wl[200] vdd gnd cell_6t
Xbit_r201_c112 bl[112] br[112] wl[201] vdd gnd cell_6t
Xbit_r202_c112 bl[112] br[112] wl[202] vdd gnd cell_6t
Xbit_r203_c112 bl[112] br[112] wl[203] vdd gnd cell_6t
Xbit_r204_c112 bl[112] br[112] wl[204] vdd gnd cell_6t
Xbit_r205_c112 bl[112] br[112] wl[205] vdd gnd cell_6t
Xbit_r206_c112 bl[112] br[112] wl[206] vdd gnd cell_6t
Xbit_r207_c112 bl[112] br[112] wl[207] vdd gnd cell_6t
Xbit_r208_c112 bl[112] br[112] wl[208] vdd gnd cell_6t
Xbit_r209_c112 bl[112] br[112] wl[209] vdd gnd cell_6t
Xbit_r210_c112 bl[112] br[112] wl[210] vdd gnd cell_6t
Xbit_r211_c112 bl[112] br[112] wl[211] vdd gnd cell_6t
Xbit_r212_c112 bl[112] br[112] wl[212] vdd gnd cell_6t
Xbit_r213_c112 bl[112] br[112] wl[213] vdd gnd cell_6t
Xbit_r214_c112 bl[112] br[112] wl[214] vdd gnd cell_6t
Xbit_r215_c112 bl[112] br[112] wl[215] vdd gnd cell_6t
Xbit_r216_c112 bl[112] br[112] wl[216] vdd gnd cell_6t
Xbit_r217_c112 bl[112] br[112] wl[217] vdd gnd cell_6t
Xbit_r218_c112 bl[112] br[112] wl[218] vdd gnd cell_6t
Xbit_r219_c112 bl[112] br[112] wl[219] vdd gnd cell_6t
Xbit_r220_c112 bl[112] br[112] wl[220] vdd gnd cell_6t
Xbit_r221_c112 bl[112] br[112] wl[221] vdd gnd cell_6t
Xbit_r222_c112 bl[112] br[112] wl[222] vdd gnd cell_6t
Xbit_r223_c112 bl[112] br[112] wl[223] vdd gnd cell_6t
Xbit_r224_c112 bl[112] br[112] wl[224] vdd gnd cell_6t
Xbit_r225_c112 bl[112] br[112] wl[225] vdd gnd cell_6t
Xbit_r226_c112 bl[112] br[112] wl[226] vdd gnd cell_6t
Xbit_r227_c112 bl[112] br[112] wl[227] vdd gnd cell_6t
Xbit_r228_c112 bl[112] br[112] wl[228] vdd gnd cell_6t
Xbit_r229_c112 bl[112] br[112] wl[229] vdd gnd cell_6t
Xbit_r230_c112 bl[112] br[112] wl[230] vdd gnd cell_6t
Xbit_r231_c112 bl[112] br[112] wl[231] vdd gnd cell_6t
Xbit_r232_c112 bl[112] br[112] wl[232] vdd gnd cell_6t
Xbit_r233_c112 bl[112] br[112] wl[233] vdd gnd cell_6t
Xbit_r234_c112 bl[112] br[112] wl[234] vdd gnd cell_6t
Xbit_r235_c112 bl[112] br[112] wl[235] vdd gnd cell_6t
Xbit_r236_c112 bl[112] br[112] wl[236] vdd gnd cell_6t
Xbit_r237_c112 bl[112] br[112] wl[237] vdd gnd cell_6t
Xbit_r238_c112 bl[112] br[112] wl[238] vdd gnd cell_6t
Xbit_r239_c112 bl[112] br[112] wl[239] vdd gnd cell_6t
Xbit_r240_c112 bl[112] br[112] wl[240] vdd gnd cell_6t
Xbit_r241_c112 bl[112] br[112] wl[241] vdd gnd cell_6t
Xbit_r242_c112 bl[112] br[112] wl[242] vdd gnd cell_6t
Xbit_r243_c112 bl[112] br[112] wl[243] vdd gnd cell_6t
Xbit_r244_c112 bl[112] br[112] wl[244] vdd gnd cell_6t
Xbit_r245_c112 bl[112] br[112] wl[245] vdd gnd cell_6t
Xbit_r246_c112 bl[112] br[112] wl[246] vdd gnd cell_6t
Xbit_r247_c112 bl[112] br[112] wl[247] vdd gnd cell_6t
Xbit_r248_c112 bl[112] br[112] wl[248] vdd gnd cell_6t
Xbit_r249_c112 bl[112] br[112] wl[249] vdd gnd cell_6t
Xbit_r250_c112 bl[112] br[112] wl[250] vdd gnd cell_6t
Xbit_r251_c112 bl[112] br[112] wl[251] vdd gnd cell_6t
Xbit_r252_c112 bl[112] br[112] wl[252] vdd gnd cell_6t
Xbit_r253_c112 bl[112] br[112] wl[253] vdd gnd cell_6t
Xbit_r254_c112 bl[112] br[112] wl[254] vdd gnd cell_6t
Xbit_r255_c112 bl[112] br[112] wl[255] vdd gnd cell_6t
Xbit_r0_c113 bl[113] br[113] wl[0] vdd gnd cell_6t
Xbit_r1_c113 bl[113] br[113] wl[1] vdd gnd cell_6t
Xbit_r2_c113 bl[113] br[113] wl[2] vdd gnd cell_6t
Xbit_r3_c113 bl[113] br[113] wl[3] vdd gnd cell_6t
Xbit_r4_c113 bl[113] br[113] wl[4] vdd gnd cell_6t
Xbit_r5_c113 bl[113] br[113] wl[5] vdd gnd cell_6t
Xbit_r6_c113 bl[113] br[113] wl[6] vdd gnd cell_6t
Xbit_r7_c113 bl[113] br[113] wl[7] vdd gnd cell_6t
Xbit_r8_c113 bl[113] br[113] wl[8] vdd gnd cell_6t
Xbit_r9_c113 bl[113] br[113] wl[9] vdd gnd cell_6t
Xbit_r10_c113 bl[113] br[113] wl[10] vdd gnd cell_6t
Xbit_r11_c113 bl[113] br[113] wl[11] vdd gnd cell_6t
Xbit_r12_c113 bl[113] br[113] wl[12] vdd gnd cell_6t
Xbit_r13_c113 bl[113] br[113] wl[13] vdd gnd cell_6t
Xbit_r14_c113 bl[113] br[113] wl[14] vdd gnd cell_6t
Xbit_r15_c113 bl[113] br[113] wl[15] vdd gnd cell_6t
Xbit_r16_c113 bl[113] br[113] wl[16] vdd gnd cell_6t
Xbit_r17_c113 bl[113] br[113] wl[17] vdd gnd cell_6t
Xbit_r18_c113 bl[113] br[113] wl[18] vdd gnd cell_6t
Xbit_r19_c113 bl[113] br[113] wl[19] vdd gnd cell_6t
Xbit_r20_c113 bl[113] br[113] wl[20] vdd gnd cell_6t
Xbit_r21_c113 bl[113] br[113] wl[21] vdd gnd cell_6t
Xbit_r22_c113 bl[113] br[113] wl[22] vdd gnd cell_6t
Xbit_r23_c113 bl[113] br[113] wl[23] vdd gnd cell_6t
Xbit_r24_c113 bl[113] br[113] wl[24] vdd gnd cell_6t
Xbit_r25_c113 bl[113] br[113] wl[25] vdd gnd cell_6t
Xbit_r26_c113 bl[113] br[113] wl[26] vdd gnd cell_6t
Xbit_r27_c113 bl[113] br[113] wl[27] vdd gnd cell_6t
Xbit_r28_c113 bl[113] br[113] wl[28] vdd gnd cell_6t
Xbit_r29_c113 bl[113] br[113] wl[29] vdd gnd cell_6t
Xbit_r30_c113 bl[113] br[113] wl[30] vdd gnd cell_6t
Xbit_r31_c113 bl[113] br[113] wl[31] vdd gnd cell_6t
Xbit_r32_c113 bl[113] br[113] wl[32] vdd gnd cell_6t
Xbit_r33_c113 bl[113] br[113] wl[33] vdd gnd cell_6t
Xbit_r34_c113 bl[113] br[113] wl[34] vdd gnd cell_6t
Xbit_r35_c113 bl[113] br[113] wl[35] vdd gnd cell_6t
Xbit_r36_c113 bl[113] br[113] wl[36] vdd gnd cell_6t
Xbit_r37_c113 bl[113] br[113] wl[37] vdd gnd cell_6t
Xbit_r38_c113 bl[113] br[113] wl[38] vdd gnd cell_6t
Xbit_r39_c113 bl[113] br[113] wl[39] vdd gnd cell_6t
Xbit_r40_c113 bl[113] br[113] wl[40] vdd gnd cell_6t
Xbit_r41_c113 bl[113] br[113] wl[41] vdd gnd cell_6t
Xbit_r42_c113 bl[113] br[113] wl[42] vdd gnd cell_6t
Xbit_r43_c113 bl[113] br[113] wl[43] vdd gnd cell_6t
Xbit_r44_c113 bl[113] br[113] wl[44] vdd gnd cell_6t
Xbit_r45_c113 bl[113] br[113] wl[45] vdd gnd cell_6t
Xbit_r46_c113 bl[113] br[113] wl[46] vdd gnd cell_6t
Xbit_r47_c113 bl[113] br[113] wl[47] vdd gnd cell_6t
Xbit_r48_c113 bl[113] br[113] wl[48] vdd gnd cell_6t
Xbit_r49_c113 bl[113] br[113] wl[49] vdd gnd cell_6t
Xbit_r50_c113 bl[113] br[113] wl[50] vdd gnd cell_6t
Xbit_r51_c113 bl[113] br[113] wl[51] vdd gnd cell_6t
Xbit_r52_c113 bl[113] br[113] wl[52] vdd gnd cell_6t
Xbit_r53_c113 bl[113] br[113] wl[53] vdd gnd cell_6t
Xbit_r54_c113 bl[113] br[113] wl[54] vdd gnd cell_6t
Xbit_r55_c113 bl[113] br[113] wl[55] vdd gnd cell_6t
Xbit_r56_c113 bl[113] br[113] wl[56] vdd gnd cell_6t
Xbit_r57_c113 bl[113] br[113] wl[57] vdd gnd cell_6t
Xbit_r58_c113 bl[113] br[113] wl[58] vdd gnd cell_6t
Xbit_r59_c113 bl[113] br[113] wl[59] vdd gnd cell_6t
Xbit_r60_c113 bl[113] br[113] wl[60] vdd gnd cell_6t
Xbit_r61_c113 bl[113] br[113] wl[61] vdd gnd cell_6t
Xbit_r62_c113 bl[113] br[113] wl[62] vdd gnd cell_6t
Xbit_r63_c113 bl[113] br[113] wl[63] vdd gnd cell_6t
Xbit_r64_c113 bl[113] br[113] wl[64] vdd gnd cell_6t
Xbit_r65_c113 bl[113] br[113] wl[65] vdd gnd cell_6t
Xbit_r66_c113 bl[113] br[113] wl[66] vdd gnd cell_6t
Xbit_r67_c113 bl[113] br[113] wl[67] vdd gnd cell_6t
Xbit_r68_c113 bl[113] br[113] wl[68] vdd gnd cell_6t
Xbit_r69_c113 bl[113] br[113] wl[69] vdd gnd cell_6t
Xbit_r70_c113 bl[113] br[113] wl[70] vdd gnd cell_6t
Xbit_r71_c113 bl[113] br[113] wl[71] vdd gnd cell_6t
Xbit_r72_c113 bl[113] br[113] wl[72] vdd gnd cell_6t
Xbit_r73_c113 bl[113] br[113] wl[73] vdd gnd cell_6t
Xbit_r74_c113 bl[113] br[113] wl[74] vdd gnd cell_6t
Xbit_r75_c113 bl[113] br[113] wl[75] vdd gnd cell_6t
Xbit_r76_c113 bl[113] br[113] wl[76] vdd gnd cell_6t
Xbit_r77_c113 bl[113] br[113] wl[77] vdd gnd cell_6t
Xbit_r78_c113 bl[113] br[113] wl[78] vdd gnd cell_6t
Xbit_r79_c113 bl[113] br[113] wl[79] vdd gnd cell_6t
Xbit_r80_c113 bl[113] br[113] wl[80] vdd gnd cell_6t
Xbit_r81_c113 bl[113] br[113] wl[81] vdd gnd cell_6t
Xbit_r82_c113 bl[113] br[113] wl[82] vdd gnd cell_6t
Xbit_r83_c113 bl[113] br[113] wl[83] vdd gnd cell_6t
Xbit_r84_c113 bl[113] br[113] wl[84] vdd gnd cell_6t
Xbit_r85_c113 bl[113] br[113] wl[85] vdd gnd cell_6t
Xbit_r86_c113 bl[113] br[113] wl[86] vdd gnd cell_6t
Xbit_r87_c113 bl[113] br[113] wl[87] vdd gnd cell_6t
Xbit_r88_c113 bl[113] br[113] wl[88] vdd gnd cell_6t
Xbit_r89_c113 bl[113] br[113] wl[89] vdd gnd cell_6t
Xbit_r90_c113 bl[113] br[113] wl[90] vdd gnd cell_6t
Xbit_r91_c113 bl[113] br[113] wl[91] vdd gnd cell_6t
Xbit_r92_c113 bl[113] br[113] wl[92] vdd gnd cell_6t
Xbit_r93_c113 bl[113] br[113] wl[93] vdd gnd cell_6t
Xbit_r94_c113 bl[113] br[113] wl[94] vdd gnd cell_6t
Xbit_r95_c113 bl[113] br[113] wl[95] vdd gnd cell_6t
Xbit_r96_c113 bl[113] br[113] wl[96] vdd gnd cell_6t
Xbit_r97_c113 bl[113] br[113] wl[97] vdd gnd cell_6t
Xbit_r98_c113 bl[113] br[113] wl[98] vdd gnd cell_6t
Xbit_r99_c113 bl[113] br[113] wl[99] vdd gnd cell_6t
Xbit_r100_c113 bl[113] br[113] wl[100] vdd gnd cell_6t
Xbit_r101_c113 bl[113] br[113] wl[101] vdd gnd cell_6t
Xbit_r102_c113 bl[113] br[113] wl[102] vdd gnd cell_6t
Xbit_r103_c113 bl[113] br[113] wl[103] vdd gnd cell_6t
Xbit_r104_c113 bl[113] br[113] wl[104] vdd gnd cell_6t
Xbit_r105_c113 bl[113] br[113] wl[105] vdd gnd cell_6t
Xbit_r106_c113 bl[113] br[113] wl[106] vdd gnd cell_6t
Xbit_r107_c113 bl[113] br[113] wl[107] vdd gnd cell_6t
Xbit_r108_c113 bl[113] br[113] wl[108] vdd gnd cell_6t
Xbit_r109_c113 bl[113] br[113] wl[109] vdd gnd cell_6t
Xbit_r110_c113 bl[113] br[113] wl[110] vdd gnd cell_6t
Xbit_r111_c113 bl[113] br[113] wl[111] vdd gnd cell_6t
Xbit_r112_c113 bl[113] br[113] wl[112] vdd gnd cell_6t
Xbit_r113_c113 bl[113] br[113] wl[113] vdd gnd cell_6t
Xbit_r114_c113 bl[113] br[113] wl[114] vdd gnd cell_6t
Xbit_r115_c113 bl[113] br[113] wl[115] vdd gnd cell_6t
Xbit_r116_c113 bl[113] br[113] wl[116] vdd gnd cell_6t
Xbit_r117_c113 bl[113] br[113] wl[117] vdd gnd cell_6t
Xbit_r118_c113 bl[113] br[113] wl[118] vdd gnd cell_6t
Xbit_r119_c113 bl[113] br[113] wl[119] vdd gnd cell_6t
Xbit_r120_c113 bl[113] br[113] wl[120] vdd gnd cell_6t
Xbit_r121_c113 bl[113] br[113] wl[121] vdd gnd cell_6t
Xbit_r122_c113 bl[113] br[113] wl[122] vdd gnd cell_6t
Xbit_r123_c113 bl[113] br[113] wl[123] vdd gnd cell_6t
Xbit_r124_c113 bl[113] br[113] wl[124] vdd gnd cell_6t
Xbit_r125_c113 bl[113] br[113] wl[125] vdd gnd cell_6t
Xbit_r126_c113 bl[113] br[113] wl[126] vdd gnd cell_6t
Xbit_r127_c113 bl[113] br[113] wl[127] vdd gnd cell_6t
Xbit_r128_c113 bl[113] br[113] wl[128] vdd gnd cell_6t
Xbit_r129_c113 bl[113] br[113] wl[129] vdd gnd cell_6t
Xbit_r130_c113 bl[113] br[113] wl[130] vdd gnd cell_6t
Xbit_r131_c113 bl[113] br[113] wl[131] vdd gnd cell_6t
Xbit_r132_c113 bl[113] br[113] wl[132] vdd gnd cell_6t
Xbit_r133_c113 bl[113] br[113] wl[133] vdd gnd cell_6t
Xbit_r134_c113 bl[113] br[113] wl[134] vdd gnd cell_6t
Xbit_r135_c113 bl[113] br[113] wl[135] vdd gnd cell_6t
Xbit_r136_c113 bl[113] br[113] wl[136] vdd gnd cell_6t
Xbit_r137_c113 bl[113] br[113] wl[137] vdd gnd cell_6t
Xbit_r138_c113 bl[113] br[113] wl[138] vdd gnd cell_6t
Xbit_r139_c113 bl[113] br[113] wl[139] vdd gnd cell_6t
Xbit_r140_c113 bl[113] br[113] wl[140] vdd gnd cell_6t
Xbit_r141_c113 bl[113] br[113] wl[141] vdd gnd cell_6t
Xbit_r142_c113 bl[113] br[113] wl[142] vdd gnd cell_6t
Xbit_r143_c113 bl[113] br[113] wl[143] vdd gnd cell_6t
Xbit_r144_c113 bl[113] br[113] wl[144] vdd gnd cell_6t
Xbit_r145_c113 bl[113] br[113] wl[145] vdd gnd cell_6t
Xbit_r146_c113 bl[113] br[113] wl[146] vdd gnd cell_6t
Xbit_r147_c113 bl[113] br[113] wl[147] vdd gnd cell_6t
Xbit_r148_c113 bl[113] br[113] wl[148] vdd gnd cell_6t
Xbit_r149_c113 bl[113] br[113] wl[149] vdd gnd cell_6t
Xbit_r150_c113 bl[113] br[113] wl[150] vdd gnd cell_6t
Xbit_r151_c113 bl[113] br[113] wl[151] vdd gnd cell_6t
Xbit_r152_c113 bl[113] br[113] wl[152] vdd gnd cell_6t
Xbit_r153_c113 bl[113] br[113] wl[153] vdd gnd cell_6t
Xbit_r154_c113 bl[113] br[113] wl[154] vdd gnd cell_6t
Xbit_r155_c113 bl[113] br[113] wl[155] vdd gnd cell_6t
Xbit_r156_c113 bl[113] br[113] wl[156] vdd gnd cell_6t
Xbit_r157_c113 bl[113] br[113] wl[157] vdd gnd cell_6t
Xbit_r158_c113 bl[113] br[113] wl[158] vdd gnd cell_6t
Xbit_r159_c113 bl[113] br[113] wl[159] vdd gnd cell_6t
Xbit_r160_c113 bl[113] br[113] wl[160] vdd gnd cell_6t
Xbit_r161_c113 bl[113] br[113] wl[161] vdd gnd cell_6t
Xbit_r162_c113 bl[113] br[113] wl[162] vdd gnd cell_6t
Xbit_r163_c113 bl[113] br[113] wl[163] vdd gnd cell_6t
Xbit_r164_c113 bl[113] br[113] wl[164] vdd gnd cell_6t
Xbit_r165_c113 bl[113] br[113] wl[165] vdd gnd cell_6t
Xbit_r166_c113 bl[113] br[113] wl[166] vdd gnd cell_6t
Xbit_r167_c113 bl[113] br[113] wl[167] vdd gnd cell_6t
Xbit_r168_c113 bl[113] br[113] wl[168] vdd gnd cell_6t
Xbit_r169_c113 bl[113] br[113] wl[169] vdd gnd cell_6t
Xbit_r170_c113 bl[113] br[113] wl[170] vdd gnd cell_6t
Xbit_r171_c113 bl[113] br[113] wl[171] vdd gnd cell_6t
Xbit_r172_c113 bl[113] br[113] wl[172] vdd gnd cell_6t
Xbit_r173_c113 bl[113] br[113] wl[173] vdd gnd cell_6t
Xbit_r174_c113 bl[113] br[113] wl[174] vdd gnd cell_6t
Xbit_r175_c113 bl[113] br[113] wl[175] vdd gnd cell_6t
Xbit_r176_c113 bl[113] br[113] wl[176] vdd gnd cell_6t
Xbit_r177_c113 bl[113] br[113] wl[177] vdd gnd cell_6t
Xbit_r178_c113 bl[113] br[113] wl[178] vdd gnd cell_6t
Xbit_r179_c113 bl[113] br[113] wl[179] vdd gnd cell_6t
Xbit_r180_c113 bl[113] br[113] wl[180] vdd gnd cell_6t
Xbit_r181_c113 bl[113] br[113] wl[181] vdd gnd cell_6t
Xbit_r182_c113 bl[113] br[113] wl[182] vdd gnd cell_6t
Xbit_r183_c113 bl[113] br[113] wl[183] vdd gnd cell_6t
Xbit_r184_c113 bl[113] br[113] wl[184] vdd gnd cell_6t
Xbit_r185_c113 bl[113] br[113] wl[185] vdd gnd cell_6t
Xbit_r186_c113 bl[113] br[113] wl[186] vdd gnd cell_6t
Xbit_r187_c113 bl[113] br[113] wl[187] vdd gnd cell_6t
Xbit_r188_c113 bl[113] br[113] wl[188] vdd gnd cell_6t
Xbit_r189_c113 bl[113] br[113] wl[189] vdd gnd cell_6t
Xbit_r190_c113 bl[113] br[113] wl[190] vdd gnd cell_6t
Xbit_r191_c113 bl[113] br[113] wl[191] vdd gnd cell_6t
Xbit_r192_c113 bl[113] br[113] wl[192] vdd gnd cell_6t
Xbit_r193_c113 bl[113] br[113] wl[193] vdd gnd cell_6t
Xbit_r194_c113 bl[113] br[113] wl[194] vdd gnd cell_6t
Xbit_r195_c113 bl[113] br[113] wl[195] vdd gnd cell_6t
Xbit_r196_c113 bl[113] br[113] wl[196] vdd gnd cell_6t
Xbit_r197_c113 bl[113] br[113] wl[197] vdd gnd cell_6t
Xbit_r198_c113 bl[113] br[113] wl[198] vdd gnd cell_6t
Xbit_r199_c113 bl[113] br[113] wl[199] vdd gnd cell_6t
Xbit_r200_c113 bl[113] br[113] wl[200] vdd gnd cell_6t
Xbit_r201_c113 bl[113] br[113] wl[201] vdd gnd cell_6t
Xbit_r202_c113 bl[113] br[113] wl[202] vdd gnd cell_6t
Xbit_r203_c113 bl[113] br[113] wl[203] vdd gnd cell_6t
Xbit_r204_c113 bl[113] br[113] wl[204] vdd gnd cell_6t
Xbit_r205_c113 bl[113] br[113] wl[205] vdd gnd cell_6t
Xbit_r206_c113 bl[113] br[113] wl[206] vdd gnd cell_6t
Xbit_r207_c113 bl[113] br[113] wl[207] vdd gnd cell_6t
Xbit_r208_c113 bl[113] br[113] wl[208] vdd gnd cell_6t
Xbit_r209_c113 bl[113] br[113] wl[209] vdd gnd cell_6t
Xbit_r210_c113 bl[113] br[113] wl[210] vdd gnd cell_6t
Xbit_r211_c113 bl[113] br[113] wl[211] vdd gnd cell_6t
Xbit_r212_c113 bl[113] br[113] wl[212] vdd gnd cell_6t
Xbit_r213_c113 bl[113] br[113] wl[213] vdd gnd cell_6t
Xbit_r214_c113 bl[113] br[113] wl[214] vdd gnd cell_6t
Xbit_r215_c113 bl[113] br[113] wl[215] vdd gnd cell_6t
Xbit_r216_c113 bl[113] br[113] wl[216] vdd gnd cell_6t
Xbit_r217_c113 bl[113] br[113] wl[217] vdd gnd cell_6t
Xbit_r218_c113 bl[113] br[113] wl[218] vdd gnd cell_6t
Xbit_r219_c113 bl[113] br[113] wl[219] vdd gnd cell_6t
Xbit_r220_c113 bl[113] br[113] wl[220] vdd gnd cell_6t
Xbit_r221_c113 bl[113] br[113] wl[221] vdd gnd cell_6t
Xbit_r222_c113 bl[113] br[113] wl[222] vdd gnd cell_6t
Xbit_r223_c113 bl[113] br[113] wl[223] vdd gnd cell_6t
Xbit_r224_c113 bl[113] br[113] wl[224] vdd gnd cell_6t
Xbit_r225_c113 bl[113] br[113] wl[225] vdd gnd cell_6t
Xbit_r226_c113 bl[113] br[113] wl[226] vdd gnd cell_6t
Xbit_r227_c113 bl[113] br[113] wl[227] vdd gnd cell_6t
Xbit_r228_c113 bl[113] br[113] wl[228] vdd gnd cell_6t
Xbit_r229_c113 bl[113] br[113] wl[229] vdd gnd cell_6t
Xbit_r230_c113 bl[113] br[113] wl[230] vdd gnd cell_6t
Xbit_r231_c113 bl[113] br[113] wl[231] vdd gnd cell_6t
Xbit_r232_c113 bl[113] br[113] wl[232] vdd gnd cell_6t
Xbit_r233_c113 bl[113] br[113] wl[233] vdd gnd cell_6t
Xbit_r234_c113 bl[113] br[113] wl[234] vdd gnd cell_6t
Xbit_r235_c113 bl[113] br[113] wl[235] vdd gnd cell_6t
Xbit_r236_c113 bl[113] br[113] wl[236] vdd gnd cell_6t
Xbit_r237_c113 bl[113] br[113] wl[237] vdd gnd cell_6t
Xbit_r238_c113 bl[113] br[113] wl[238] vdd gnd cell_6t
Xbit_r239_c113 bl[113] br[113] wl[239] vdd gnd cell_6t
Xbit_r240_c113 bl[113] br[113] wl[240] vdd gnd cell_6t
Xbit_r241_c113 bl[113] br[113] wl[241] vdd gnd cell_6t
Xbit_r242_c113 bl[113] br[113] wl[242] vdd gnd cell_6t
Xbit_r243_c113 bl[113] br[113] wl[243] vdd gnd cell_6t
Xbit_r244_c113 bl[113] br[113] wl[244] vdd gnd cell_6t
Xbit_r245_c113 bl[113] br[113] wl[245] vdd gnd cell_6t
Xbit_r246_c113 bl[113] br[113] wl[246] vdd gnd cell_6t
Xbit_r247_c113 bl[113] br[113] wl[247] vdd gnd cell_6t
Xbit_r248_c113 bl[113] br[113] wl[248] vdd gnd cell_6t
Xbit_r249_c113 bl[113] br[113] wl[249] vdd gnd cell_6t
Xbit_r250_c113 bl[113] br[113] wl[250] vdd gnd cell_6t
Xbit_r251_c113 bl[113] br[113] wl[251] vdd gnd cell_6t
Xbit_r252_c113 bl[113] br[113] wl[252] vdd gnd cell_6t
Xbit_r253_c113 bl[113] br[113] wl[253] vdd gnd cell_6t
Xbit_r254_c113 bl[113] br[113] wl[254] vdd gnd cell_6t
Xbit_r255_c113 bl[113] br[113] wl[255] vdd gnd cell_6t
Xbit_r0_c114 bl[114] br[114] wl[0] vdd gnd cell_6t
Xbit_r1_c114 bl[114] br[114] wl[1] vdd gnd cell_6t
Xbit_r2_c114 bl[114] br[114] wl[2] vdd gnd cell_6t
Xbit_r3_c114 bl[114] br[114] wl[3] vdd gnd cell_6t
Xbit_r4_c114 bl[114] br[114] wl[4] vdd gnd cell_6t
Xbit_r5_c114 bl[114] br[114] wl[5] vdd gnd cell_6t
Xbit_r6_c114 bl[114] br[114] wl[6] vdd gnd cell_6t
Xbit_r7_c114 bl[114] br[114] wl[7] vdd gnd cell_6t
Xbit_r8_c114 bl[114] br[114] wl[8] vdd gnd cell_6t
Xbit_r9_c114 bl[114] br[114] wl[9] vdd gnd cell_6t
Xbit_r10_c114 bl[114] br[114] wl[10] vdd gnd cell_6t
Xbit_r11_c114 bl[114] br[114] wl[11] vdd gnd cell_6t
Xbit_r12_c114 bl[114] br[114] wl[12] vdd gnd cell_6t
Xbit_r13_c114 bl[114] br[114] wl[13] vdd gnd cell_6t
Xbit_r14_c114 bl[114] br[114] wl[14] vdd gnd cell_6t
Xbit_r15_c114 bl[114] br[114] wl[15] vdd gnd cell_6t
Xbit_r16_c114 bl[114] br[114] wl[16] vdd gnd cell_6t
Xbit_r17_c114 bl[114] br[114] wl[17] vdd gnd cell_6t
Xbit_r18_c114 bl[114] br[114] wl[18] vdd gnd cell_6t
Xbit_r19_c114 bl[114] br[114] wl[19] vdd gnd cell_6t
Xbit_r20_c114 bl[114] br[114] wl[20] vdd gnd cell_6t
Xbit_r21_c114 bl[114] br[114] wl[21] vdd gnd cell_6t
Xbit_r22_c114 bl[114] br[114] wl[22] vdd gnd cell_6t
Xbit_r23_c114 bl[114] br[114] wl[23] vdd gnd cell_6t
Xbit_r24_c114 bl[114] br[114] wl[24] vdd gnd cell_6t
Xbit_r25_c114 bl[114] br[114] wl[25] vdd gnd cell_6t
Xbit_r26_c114 bl[114] br[114] wl[26] vdd gnd cell_6t
Xbit_r27_c114 bl[114] br[114] wl[27] vdd gnd cell_6t
Xbit_r28_c114 bl[114] br[114] wl[28] vdd gnd cell_6t
Xbit_r29_c114 bl[114] br[114] wl[29] vdd gnd cell_6t
Xbit_r30_c114 bl[114] br[114] wl[30] vdd gnd cell_6t
Xbit_r31_c114 bl[114] br[114] wl[31] vdd gnd cell_6t
Xbit_r32_c114 bl[114] br[114] wl[32] vdd gnd cell_6t
Xbit_r33_c114 bl[114] br[114] wl[33] vdd gnd cell_6t
Xbit_r34_c114 bl[114] br[114] wl[34] vdd gnd cell_6t
Xbit_r35_c114 bl[114] br[114] wl[35] vdd gnd cell_6t
Xbit_r36_c114 bl[114] br[114] wl[36] vdd gnd cell_6t
Xbit_r37_c114 bl[114] br[114] wl[37] vdd gnd cell_6t
Xbit_r38_c114 bl[114] br[114] wl[38] vdd gnd cell_6t
Xbit_r39_c114 bl[114] br[114] wl[39] vdd gnd cell_6t
Xbit_r40_c114 bl[114] br[114] wl[40] vdd gnd cell_6t
Xbit_r41_c114 bl[114] br[114] wl[41] vdd gnd cell_6t
Xbit_r42_c114 bl[114] br[114] wl[42] vdd gnd cell_6t
Xbit_r43_c114 bl[114] br[114] wl[43] vdd gnd cell_6t
Xbit_r44_c114 bl[114] br[114] wl[44] vdd gnd cell_6t
Xbit_r45_c114 bl[114] br[114] wl[45] vdd gnd cell_6t
Xbit_r46_c114 bl[114] br[114] wl[46] vdd gnd cell_6t
Xbit_r47_c114 bl[114] br[114] wl[47] vdd gnd cell_6t
Xbit_r48_c114 bl[114] br[114] wl[48] vdd gnd cell_6t
Xbit_r49_c114 bl[114] br[114] wl[49] vdd gnd cell_6t
Xbit_r50_c114 bl[114] br[114] wl[50] vdd gnd cell_6t
Xbit_r51_c114 bl[114] br[114] wl[51] vdd gnd cell_6t
Xbit_r52_c114 bl[114] br[114] wl[52] vdd gnd cell_6t
Xbit_r53_c114 bl[114] br[114] wl[53] vdd gnd cell_6t
Xbit_r54_c114 bl[114] br[114] wl[54] vdd gnd cell_6t
Xbit_r55_c114 bl[114] br[114] wl[55] vdd gnd cell_6t
Xbit_r56_c114 bl[114] br[114] wl[56] vdd gnd cell_6t
Xbit_r57_c114 bl[114] br[114] wl[57] vdd gnd cell_6t
Xbit_r58_c114 bl[114] br[114] wl[58] vdd gnd cell_6t
Xbit_r59_c114 bl[114] br[114] wl[59] vdd gnd cell_6t
Xbit_r60_c114 bl[114] br[114] wl[60] vdd gnd cell_6t
Xbit_r61_c114 bl[114] br[114] wl[61] vdd gnd cell_6t
Xbit_r62_c114 bl[114] br[114] wl[62] vdd gnd cell_6t
Xbit_r63_c114 bl[114] br[114] wl[63] vdd gnd cell_6t
Xbit_r64_c114 bl[114] br[114] wl[64] vdd gnd cell_6t
Xbit_r65_c114 bl[114] br[114] wl[65] vdd gnd cell_6t
Xbit_r66_c114 bl[114] br[114] wl[66] vdd gnd cell_6t
Xbit_r67_c114 bl[114] br[114] wl[67] vdd gnd cell_6t
Xbit_r68_c114 bl[114] br[114] wl[68] vdd gnd cell_6t
Xbit_r69_c114 bl[114] br[114] wl[69] vdd gnd cell_6t
Xbit_r70_c114 bl[114] br[114] wl[70] vdd gnd cell_6t
Xbit_r71_c114 bl[114] br[114] wl[71] vdd gnd cell_6t
Xbit_r72_c114 bl[114] br[114] wl[72] vdd gnd cell_6t
Xbit_r73_c114 bl[114] br[114] wl[73] vdd gnd cell_6t
Xbit_r74_c114 bl[114] br[114] wl[74] vdd gnd cell_6t
Xbit_r75_c114 bl[114] br[114] wl[75] vdd gnd cell_6t
Xbit_r76_c114 bl[114] br[114] wl[76] vdd gnd cell_6t
Xbit_r77_c114 bl[114] br[114] wl[77] vdd gnd cell_6t
Xbit_r78_c114 bl[114] br[114] wl[78] vdd gnd cell_6t
Xbit_r79_c114 bl[114] br[114] wl[79] vdd gnd cell_6t
Xbit_r80_c114 bl[114] br[114] wl[80] vdd gnd cell_6t
Xbit_r81_c114 bl[114] br[114] wl[81] vdd gnd cell_6t
Xbit_r82_c114 bl[114] br[114] wl[82] vdd gnd cell_6t
Xbit_r83_c114 bl[114] br[114] wl[83] vdd gnd cell_6t
Xbit_r84_c114 bl[114] br[114] wl[84] vdd gnd cell_6t
Xbit_r85_c114 bl[114] br[114] wl[85] vdd gnd cell_6t
Xbit_r86_c114 bl[114] br[114] wl[86] vdd gnd cell_6t
Xbit_r87_c114 bl[114] br[114] wl[87] vdd gnd cell_6t
Xbit_r88_c114 bl[114] br[114] wl[88] vdd gnd cell_6t
Xbit_r89_c114 bl[114] br[114] wl[89] vdd gnd cell_6t
Xbit_r90_c114 bl[114] br[114] wl[90] vdd gnd cell_6t
Xbit_r91_c114 bl[114] br[114] wl[91] vdd gnd cell_6t
Xbit_r92_c114 bl[114] br[114] wl[92] vdd gnd cell_6t
Xbit_r93_c114 bl[114] br[114] wl[93] vdd gnd cell_6t
Xbit_r94_c114 bl[114] br[114] wl[94] vdd gnd cell_6t
Xbit_r95_c114 bl[114] br[114] wl[95] vdd gnd cell_6t
Xbit_r96_c114 bl[114] br[114] wl[96] vdd gnd cell_6t
Xbit_r97_c114 bl[114] br[114] wl[97] vdd gnd cell_6t
Xbit_r98_c114 bl[114] br[114] wl[98] vdd gnd cell_6t
Xbit_r99_c114 bl[114] br[114] wl[99] vdd gnd cell_6t
Xbit_r100_c114 bl[114] br[114] wl[100] vdd gnd cell_6t
Xbit_r101_c114 bl[114] br[114] wl[101] vdd gnd cell_6t
Xbit_r102_c114 bl[114] br[114] wl[102] vdd gnd cell_6t
Xbit_r103_c114 bl[114] br[114] wl[103] vdd gnd cell_6t
Xbit_r104_c114 bl[114] br[114] wl[104] vdd gnd cell_6t
Xbit_r105_c114 bl[114] br[114] wl[105] vdd gnd cell_6t
Xbit_r106_c114 bl[114] br[114] wl[106] vdd gnd cell_6t
Xbit_r107_c114 bl[114] br[114] wl[107] vdd gnd cell_6t
Xbit_r108_c114 bl[114] br[114] wl[108] vdd gnd cell_6t
Xbit_r109_c114 bl[114] br[114] wl[109] vdd gnd cell_6t
Xbit_r110_c114 bl[114] br[114] wl[110] vdd gnd cell_6t
Xbit_r111_c114 bl[114] br[114] wl[111] vdd gnd cell_6t
Xbit_r112_c114 bl[114] br[114] wl[112] vdd gnd cell_6t
Xbit_r113_c114 bl[114] br[114] wl[113] vdd gnd cell_6t
Xbit_r114_c114 bl[114] br[114] wl[114] vdd gnd cell_6t
Xbit_r115_c114 bl[114] br[114] wl[115] vdd gnd cell_6t
Xbit_r116_c114 bl[114] br[114] wl[116] vdd gnd cell_6t
Xbit_r117_c114 bl[114] br[114] wl[117] vdd gnd cell_6t
Xbit_r118_c114 bl[114] br[114] wl[118] vdd gnd cell_6t
Xbit_r119_c114 bl[114] br[114] wl[119] vdd gnd cell_6t
Xbit_r120_c114 bl[114] br[114] wl[120] vdd gnd cell_6t
Xbit_r121_c114 bl[114] br[114] wl[121] vdd gnd cell_6t
Xbit_r122_c114 bl[114] br[114] wl[122] vdd gnd cell_6t
Xbit_r123_c114 bl[114] br[114] wl[123] vdd gnd cell_6t
Xbit_r124_c114 bl[114] br[114] wl[124] vdd gnd cell_6t
Xbit_r125_c114 bl[114] br[114] wl[125] vdd gnd cell_6t
Xbit_r126_c114 bl[114] br[114] wl[126] vdd gnd cell_6t
Xbit_r127_c114 bl[114] br[114] wl[127] vdd gnd cell_6t
Xbit_r128_c114 bl[114] br[114] wl[128] vdd gnd cell_6t
Xbit_r129_c114 bl[114] br[114] wl[129] vdd gnd cell_6t
Xbit_r130_c114 bl[114] br[114] wl[130] vdd gnd cell_6t
Xbit_r131_c114 bl[114] br[114] wl[131] vdd gnd cell_6t
Xbit_r132_c114 bl[114] br[114] wl[132] vdd gnd cell_6t
Xbit_r133_c114 bl[114] br[114] wl[133] vdd gnd cell_6t
Xbit_r134_c114 bl[114] br[114] wl[134] vdd gnd cell_6t
Xbit_r135_c114 bl[114] br[114] wl[135] vdd gnd cell_6t
Xbit_r136_c114 bl[114] br[114] wl[136] vdd gnd cell_6t
Xbit_r137_c114 bl[114] br[114] wl[137] vdd gnd cell_6t
Xbit_r138_c114 bl[114] br[114] wl[138] vdd gnd cell_6t
Xbit_r139_c114 bl[114] br[114] wl[139] vdd gnd cell_6t
Xbit_r140_c114 bl[114] br[114] wl[140] vdd gnd cell_6t
Xbit_r141_c114 bl[114] br[114] wl[141] vdd gnd cell_6t
Xbit_r142_c114 bl[114] br[114] wl[142] vdd gnd cell_6t
Xbit_r143_c114 bl[114] br[114] wl[143] vdd gnd cell_6t
Xbit_r144_c114 bl[114] br[114] wl[144] vdd gnd cell_6t
Xbit_r145_c114 bl[114] br[114] wl[145] vdd gnd cell_6t
Xbit_r146_c114 bl[114] br[114] wl[146] vdd gnd cell_6t
Xbit_r147_c114 bl[114] br[114] wl[147] vdd gnd cell_6t
Xbit_r148_c114 bl[114] br[114] wl[148] vdd gnd cell_6t
Xbit_r149_c114 bl[114] br[114] wl[149] vdd gnd cell_6t
Xbit_r150_c114 bl[114] br[114] wl[150] vdd gnd cell_6t
Xbit_r151_c114 bl[114] br[114] wl[151] vdd gnd cell_6t
Xbit_r152_c114 bl[114] br[114] wl[152] vdd gnd cell_6t
Xbit_r153_c114 bl[114] br[114] wl[153] vdd gnd cell_6t
Xbit_r154_c114 bl[114] br[114] wl[154] vdd gnd cell_6t
Xbit_r155_c114 bl[114] br[114] wl[155] vdd gnd cell_6t
Xbit_r156_c114 bl[114] br[114] wl[156] vdd gnd cell_6t
Xbit_r157_c114 bl[114] br[114] wl[157] vdd gnd cell_6t
Xbit_r158_c114 bl[114] br[114] wl[158] vdd gnd cell_6t
Xbit_r159_c114 bl[114] br[114] wl[159] vdd gnd cell_6t
Xbit_r160_c114 bl[114] br[114] wl[160] vdd gnd cell_6t
Xbit_r161_c114 bl[114] br[114] wl[161] vdd gnd cell_6t
Xbit_r162_c114 bl[114] br[114] wl[162] vdd gnd cell_6t
Xbit_r163_c114 bl[114] br[114] wl[163] vdd gnd cell_6t
Xbit_r164_c114 bl[114] br[114] wl[164] vdd gnd cell_6t
Xbit_r165_c114 bl[114] br[114] wl[165] vdd gnd cell_6t
Xbit_r166_c114 bl[114] br[114] wl[166] vdd gnd cell_6t
Xbit_r167_c114 bl[114] br[114] wl[167] vdd gnd cell_6t
Xbit_r168_c114 bl[114] br[114] wl[168] vdd gnd cell_6t
Xbit_r169_c114 bl[114] br[114] wl[169] vdd gnd cell_6t
Xbit_r170_c114 bl[114] br[114] wl[170] vdd gnd cell_6t
Xbit_r171_c114 bl[114] br[114] wl[171] vdd gnd cell_6t
Xbit_r172_c114 bl[114] br[114] wl[172] vdd gnd cell_6t
Xbit_r173_c114 bl[114] br[114] wl[173] vdd gnd cell_6t
Xbit_r174_c114 bl[114] br[114] wl[174] vdd gnd cell_6t
Xbit_r175_c114 bl[114] br[114] wl[175] vdd gnd cell_6t
Xbit_r176_c114 bl[114] br[114] wl[176] vdd gnd cell_6t
Xbit_r177_c114 bl[114] br[114] wl[177] vdd gnd cell_6t
Xbit_r178_c114 bl[114] br[114] wl[178] vdd gnd cell_6t
Xbit_r179_c114 bl[114] br[114] wl[179] vdd gnd cell_6t
Xbit_r180_c114 bl[114] br[114] wl[180] vdd gnd cell_6t
Xbit_r181_c114 bl[114] br[114] wl[181] vdd gnd cell_6t
Xbit_r182_c114 bl[114] br[114] wl[182] vdd gnd cell_6t
Xbit_r183_c114 bl[114] br[114] wl[183] vdd gnd cell_6t
Xbit_r184_c114 bl[114] br[114] wl[184] vdd gnd cell_6t
Xbit_r185_c114 bl[114] br[114] wl[185] vdd gnd cell_6t
Xbit_r186_c114 bl[114] br[114] wl[186] vdd gnd cell_6t
Xbit_r187_c114 bl[114] br[114] wl[187] vdd gnd cell_6t
Xbit_r188_c114 bl[114] br[114] wl[188] vdd gnd cell_6t
Xbit_r189_c114 bl[114] br[114] wl[189] vdd gnd cell_6t
Xbit_r190_c114 bl[114] br[114] wl[190] vdd gnd cell_6t
Xbit_r191_c114 bl[114] br[114] wl[191] vdd gnd cell_6t
Xbit_r192_c114 bl[114] br[114] wl[192] vdd gnd cell_6t
Xbit_r193_c114 bl[114] br[114] wl[193] vdd gnd cell_6t
Xbit_r194_c114 bl[114] br[114] wl[194] vdd gnd cell_6t
Xbit_r195_c114 bl[114] br[114] wl[195] vdd gnd cell_6t
Xbit_r196_c114 bl[114] br[114] wl[196] vdd gnd cell_6t
Xbit_r197_c114 bl[114] br[114] wl[197] vdd gnd cell_6t
Xbit_r198_c114 bl[114] br[114] wl[198] vdd gnd cell_6t
Xbit_r199_c114 bl[114] br[114] wl[199] vdd gnd cell_6t
Xbit_r200_c114 bl[114] br[114] wl[200] vdd gnd cell_6t
Xbit_r201_c114 bl[114] br[114] wl[201] vdd gnd cell_6t
Xbit_r202_c114 bl[114] br[114] wl[202] vdd gnd cell_6t
Xbit_r203_c114 bl[114] br[114] wl[203] vdd gnd cell_6t
Xbit_r204_c114 bl[114] br[114] wl[204] vdd gnd cell_6t
Xbit_r205_c114 bl[114] br[114] wl[205] vdd gnd cell_6t
Xbit_r206_c114 bl[114] br[114] wl[206] vdd gnd cell_6t
Xbit_r207_c114 bl[114] br[114] wl[207] vdd gnd cell_6t
Xbit_r208_c114 bl[114] br[114] wl[208] vdd gnd cell_6t
Xbit_r209_c114 bl[114] br[114] wl[209] vdd gnd cell_6t
Xbit_r210_c114 bl[114] br[114] wl[210] vdd gnd cell_6t
Xbit_r211_c114 bl[114] br[114] wl[211] vdd gnd cell_6t
Xbit_r212_c114 bl[114] br[114] wl[212] vdd gnd cell_6t
Xbit_r213_c114 bl[114] br[114] wl[213] vdd gnd cell_6t
Xbit_r214_c114 bl[114] br[114] wl[214] vdd gnd cell_6t
Xbit_r215_c114 bl[114] br[114] wl[215] vdd gnd cell_6t
Xbit_r216_c114 bl[114] br[114] wl[216] vdd gnd cell_6t
Xbit_r217_c114 bl[114] br[114] wl[217] vdd gnd cell_6t
Xbit_r218_c114 bl[114] br[114] wl[218] vdd gnd cell_6t
Xbit_r219_c114 bl[114] br[114] wl[219] vdd gnd cell_6t
Xbit_r220_c114 bl[114] br[114] wl[220] vdd gnd cell_6t
Xbit_r221_c114 bl[114] br[114] wl[221] vdd gnd cell_6t
Xbit_r222_c114 bl[114] br[114] wl[222] vdd gnd cell_6t
Xbit_r223_c114 bl[114] br[114] wl[223] vdd gnd cell_6t
Xbit_r224_c114 bl[114] br[114] wl[224] vdd gnd cell_6t
Xbit_r225_c114 bl[114] br[114] wl[225] vdd gnd cell_6t
Xbit_r226_c114 bl[114] br[114] wl[226] vdd gnd cell_6t
Xbit_r227_c114 bl[114] br[114] wl[227] vdd gnd cell_6t
Xbit_r228_c114 bl[114] br[114] wl[228] vdd gnd cell_6t
Xbit_r229_c114 bl[114] br[114] wl[229] vdd gnd cell_6t
Xbit_r230_c114 bl[114] br[114] wl[230] vdd gnd cell_6t
Xbit_r231_c114 bl[114] br[114] wl[231] vdd gnd cell_6t
Xbit_r232_c114 bl[114] br[114] wl[232] vdd gnd cell_6t
Xbit_r233_c114 bl[114] br[114] wl[233] vdd gnd cell_6t
Xbit_r234_c114 bl[114] br[114] wl[234] vdd gnd cell_6t
Xbit_r235_c114 bl[114] br[114] wl[235] vdd gnd cell_6t
Xbit_r236_c114 bl[114] br[114] wl[236] vdd gnd cell_6t
Xbit_r237_c114 bl[114] br[114] wl[237] vdd gnd cell_6t
Xbit_r238_c114 bl[114] br[114] wl[238] vdd gnd cell_6t
Xbit_r239_c114 bl[114] br[114] wl[239] vdd gnd cell_6t
Xbit_r240_c114 bl[114] br[114] wl[240] vdd gnd cell_6t
Xbit_r241_c114 bl[114] br[114] wl[241] vdd gnd cell_6t
Xbit_r242_c114 bl[114] br[114] wl[242] vdd gnd cell_6t
Xbit_r243_c114 bl[114] br[114] wl[243] vdd gnd cell_6t
Xbit_r244_c114 bl[114] br[114] wl[244] vdd gnd cell_6t
Xbit_r245_c114 bl[114] br[114] wl[245] vdd gnd cell_6t
Xbit_r246_c114 bl[114] br[114] wl[246] vdd gnd cell_6t
Xbit_r247_c114 bl[114] br[114] wl[247] vdd gnd cell_6t
Xbit_r248_c114 bl[114] br[114] wl[248] vdd gnd cell_6t
Xbit_r249_c114 bl[114] br[114] wl[249] vdd gnd cell_6t
Xbit_r250_c114 bl[114] br[114] wl[250] vdd gnd cell_6t
Xbit_r251_c114 bl[114] br[114] wl[251] vdd gnd cell_6t
Xbit_r252_c114 bl[114] br[114] wl[252] vdd gnd cell_6t
Xbit_r253_c114 bl[114] br[114] wl[253] vdd gnd cell_6t
Xbit_r254_c114 bl[114] br[114] wl[254] vdd gnd cell_6t
Xbit_r255_c114 bl[114] br[114] wl[255] vdd gnd cell_6t
Xbit_r0_c115 bl[115] br[115] wl[0] vdd gnd cell_6t
Xbit_r1_c115 bl[115] br[115] wl[1] vdd gnd cell_6t
Xbit_r2_c115 bl[115] br[115] wl[2] vdd gnd cell_6t
Xbit_r3_c115 bl[115] br[115] wl[3] vdd gnd cell_6t
Xbit_r4_c115 bl[115] br[115] wl[4] vdd gnd cell_6t
Xbit_r5_c115 bl[115] br[115] wl[5] vdd gnd cell_6t
Xbit_r6_c115 bl[115] br[115] wl[6] vdd gnd cell_6t
Xbit_r7_c115 bl[115] br[115] wl[7] vdd gnd cell_6t
Xbit_r8_c115 bl[115] br[115] wl[8] vdd gnd cell_6t
Xbit_r9_c115 bl[115] br[115] wl[9] vdd gnd cell_6t
Xbit_r10_c115 bl[115] br[115] wl[10] vdd gnd cell_6t
Xbit_r11_c115 bl[115] br[115] wl[11] vdd gnd cell_6t
Xbit_r12_c115 bl[115] br[115] wl[12] vdd gnd cell_6t
Xbit_r13_c115 bl[115] br[115] wl[13] vdd gnd cell_6t
Xbit_r14_c115 bl[115] br[115] wl[14] vdd gnd cell_6t
Xbit_r15_c115 bl[115] br[115] wl[15] vdd gnd cell_6t
Xbit_r16_c115 bl[115] br[115] wl[16] vdd gnd cell_6t
Xbit_r17_c115 bl[115] br[115] wl[17] vdd gnd cell_6t
Xbit_r18_c115 bl[115] br[115] wl[18] vdd gnd cell_6t
Xbit_r19_c115 bl[115] br[115] wl[19] vdd gnd cell_6t
Xbit_r20_c115 bl[115] br[115] wl[20] vdd gnd cell_6t
Xbit_r21_c115 bl[115] br[115] wl[21] vdd gnd cell_6t
Xbit_r22_c115 bl[115] br[115] wl[22] vdd gnd cell_6t
Xbit_r23_c115 bl[115] br[115] wl[23] vdd gnd cell_6t
Xbit_r24_c115 bl[115] br[115] wl[24] vdd gnd cell_6t
Xbit_r25_c115 bl[115] br[115] wl[25] vdd gnd cell_6t
Xbit_r26_c115 bl[115] br[115] wl[26] vdd gnd cell_6t
Xbit_r27_c115 bl[115] br[115] wl[27] vdd gnd cell_6t
Xbit_r28_c115 bl[115] br[115] wl[28] vdd gnd cell_6t
Xbit_r29_c115 bl[115] br[115] wl[29] vdd gnd cell_6t
Xbit_r30_c115 bl[115] br[115] wl[30] vdd gnd cell_6t
Xbit_r31_c115 bl[115] br[115] wl[31] vdd gnd cell_6t
Xbit_r32_c115 bl[115] br[115] wl[32] vdd gnd cell_6t
Xbit_r33_c115 bl[115] br[115] wl[33] vdd gnd cell_6t
Xbit_r34_c115 bl[115] br[115] wl[34] vdd gnd cell_6t
Xbit_r35_c115 bl[115] br[115] wl[35] vdd gnd cell_6t
Xbit_r36_c115 bl[115] br[115] wl[36] vdd gnd cell_6t
Xbit_r37_c115 bl[115] br[115] wl[37] vdd gnd cell_6t
Xbit_r38_c115 bl[115] br[115] wl[38] vdd gnd cell_6t
Xbit_r39_c115 bl[115] br[115] wl[39] vdd gnd cell_6t
Xbit_r40_c115 bl[115] br[115] wl[40] vdd gnd cell_6t
Xbit_r41_c115 bl[115] br[115] wl[41] vdd gnd cell_6t
Xbit_r42_c115 bl[115] br[115] wl[42] vdd gnd cell_6t
Xbit_r43_c115 bl[115] br[115] wl[43] vdd gnd cell_6t
Xbit_r44_c115 bl[115] br[115] wl[44] vdd gnd cell_6t
Xbit_r45_c115 bl[115] br[115] wl[45] vdd gnd cell_6t
Xbit_r46_c115 bl[115] br[115] wl[46] vdd gnd cell_6t
Xbit_r47_c115 bl[115] br[115] wl[47] vdd gnd cell_6t
Xbit_r48_c115 bl[115] br[115] wl[48] vdd gnd cell_6t
Xbit_r49_c115 bl[115] br[115] wl[49] vdd gnd cell_6t
Xbit_r50_c115 bl[115] br[115] wl[50] vdd gnd cell_6t
Xbit_r51_c115 bl[115] br[115] wl[51] vdd gnd cell_6t
Xbit_r52_c115 bl[115] br[115] wl[52] vdd gnd cell_6t
Xbit_r53_c115 bl[115] br[115] wl[53] vdd gnd cell_6t
Xbit_r54_c115 bl[115] br[115] wl[54] vdd gnd cell_6t
Xbit_r55_c115 bl[115] br[115] wl[55] vdd gnd cell_6t
Xbit_r56_c115 bl[115] br[115] wl[56] vdd gnd cell_6t
Xbit_r57_c115 bl[115] br[115] wl[57] vdd gnd cell_6t
Xbit_r58_c115 bl[115] br[115] wl[58] vdd gnd cell_6t
Xbit_r59_c115 bl[115] br[115] wl[59] vdd gnd cell_6t
Xbit_r60_c115 bl[115] br[115] wl[60] vdd gnd cell_6t
Xbit_r61_c115 bl[115] br[115] wl[61] vdd gnd cell_6t
Xbit_r62_c115 bl[115] br[115] wl[62] vdd gnd cell_6t
Xbit_r63_c115 bl[115] br[115] wl[63] vdd gnd cell_6t
Xbit_r64_c115 bl[115] br[115] wl[64] vdd gnd cell_6t
Xbit_r65_c115 bl[115] br[115] wl[65] vdd gnd cell_6t
Xbit_r66_c115 bl[115] br[115] wl[66] vdd gnd cell_6t
Xbit_r67_c115 bl[115] br[115] wl[67] vdd gnd cell_6t
Xbit_r68_c115 bl[115] br[115] wl[68] vdd gnd cell_6t
Xbit_r69_c115 bl[115] br[115] wl[69] vdd gnd cell_6t
Xbit_r70_c115 bl[115] br[115] wl[70] vdd gnd cell_6t
Xbit_r71_c115 bl[115] br[115] wl[71] vdd gnd cell_6t
Xbit_r72_c115 bl[115] br[115] wl[72] vdd gnd cell_6t
Xbit_r73_c115 bl[115] br[115] wl[73] vdd gnd cell_6t
Xbit_r74_c115 bl[115] br[115] wl[74] vdd gnd cell_6t
Xbit_r75_c115 bl[115] br[115] wl[75] vdd gnd cell_6t
Xbit_r76_c115 bl[115] br[115] wl[76] vdd gnd cell_6t
Xbit_r77_c115 bl[115] br[115] wl[77] vdd gnd cell_6t
Xbit_r78_c115 bl[115] br[115] wl[78] vdd gnd cell_6t
Xbit_r79_c115 bl[115] br[115] wl[79] vdd gnd cell_6t
Xbit_r80_c115 bl[115] br[115] wl[80] vdd gnd cell_6t
Xbit_r81_c115 bl[115] br[115] wl[81] vdd gnd cell_6t
Xbit_r82_c115 bl[115] br[115] wl[82] vdd gnd cell_6t
Xbit_r83_c115 bl[115] br[115] wl[83] vdd gnd cell_6t
Xbit_r84_c115 bl[115] br[115] wl[84] vdd gnd cell_6t
Xbit_r85_c115 bl[115] br[115] wl[85] vdd gnd cell_6t
Xbit_r86_c115 bl[115] br[115] wl[86] vdd gnd cell_6t
Xbit_r87_c115 bl[115] br[115] wl[87] vdd gnd cell_6t
Xbit_r88_c115 bl[115] br[115] wl[88] vdd gnd cell_6t
Xbit_r89_c115 bl[115] br[115] wl[89] vdd gnd cell_6t
Xbit_r90_c115 bl[115] br[115] wl[90] vdd gnd cell_6t
Xbit_r91_c115 bl[115] br[115] wl[91] vdd gnd cell_6t
Xbit_r92_c115 bl[115] br[115] wl[92] vdd gnd cell_6t
Xbit_r93_c115 bl[115] br[115] wl[93] vdd gnd cell_6t
Xbit_r94_c115 bl[115] br[115] wl[94] vdd gnd cell_6t
Xbit_r95_c115 bl[115] br[115] wl[95] vdd gnd cell_6t
Xbit_r96_c115 bl[115] br[115] wl[96] vdd gnd cell_6t
Xbit_r97_c115 bl[115] br[115] wl[97] vdd gnd cell_6t
Xbit_r98_c115 bl[115] br[115] wl[98] vdd gnd cell_6t
Xbit_r99_c115 bl[115] br[115] wl[99] vdd gnd cell_6t
Xbit_r100_c115 bl[115] br[115] wl[100] vdd gnd cell_6t
Xbit_r101_c115 bl[115] br[115] wl[101] vdd gnd cell_6t
Xbit_r102_c115 bl[115] br[115] wl[102] vdd gnd cell_6t
Xbit_r103_c115 bl[115] br[115] wl[103] vdd gnd cell_6t
Xbit_r104_c115 bl[115] br[115] wl[104] vdd gnd cell_6t
Xbit_r105_c115 bl[115] br[115] wl[105] vdd gnd cell_6t
Xbit_r106_c115 bl[115] br[115] wl[106] vdd gnd cell_6t
Xbit_r107_c115 bl[115] br[115] wl[107] vdd gnd cell_6t
Xbit_r108_c115 bl[115] br[115] wl[108] vdd gnd cell_6t
Xbit_r109_c115 bl[115] br[115] wl[109] vdd gnd cell_6t
Xbit_r110_c115 bl[115] br[115] wl[110] vdd gnd cell_6t
Xbit_r111_c115 bl[115] br[115] wl[111] vdd gnd cell_6t
Xbit_r112_c115 bl[115] br[115] wl[112] vdd gnd cell_6t
Xbit_r113_c115 bl[115] br[115] wl[113] vdd gnd cell_6t
Xbit_r114_c115 bl[115] br[115] wl[114] vdd gnd cell_6t
Xbit_r115_c115 bl[115] br[115] wl[115] vdd gnd cell_6t
Xbit_r116_c115 bl[115] br[115] wl[116] vdd gnd cell_6t
Xbit_r117_c115 bl[115] br[115] wl[117] vdd gnd cell_6t
Xbit_r118_c115 bl[115] br[115] wl[118] vdd gnd cell_6t
Xbit_r119_c115 bl[115] br[115] wl[119] vdd gnd cell_6t
Xbit_r120_c115 bl[115] br[115] wl[120] vdd gnd cell_6t
Xbit_r121_c115 bl[115] br[115] wl[121] vdd gnd cell_6t
Xbit_r122_c115 bl[115] br[115] wl[122] vdd gnd cell_6t
Xbit_r123_c115 bl[115] br[115] wl[123] vdd gnd cell_6t
Xbit_r124_c115 bl[115] br[115] wl[124] vdd gnd cell_6t
Xbit_r125_c115 bl[115] br[115] wl[125] vdd gnd cell_6t
Xbit_r126_c115 bl[115] br[115] wl[126] vdd gnd cell_6t
Xbit_r127_c115 bl[115] br[115] wl[127] vdd gnd cell_6t
Xbit_r128_c115 bl[115] br[115] wl[128] vdd gnd cell_6t
Xbit_r129_c115 bl[115] br[115] wl[129] vdd gnd cell_6t
Xbit_r130_c115 bl[115] br[115] wl[130] vdd gnd cell_6t
Xbit_r131_c115 bl[115] br[115] wl[131] vdd gnd cell_6t
Xbit_r132_c115 bl[115] br[115] wl[132] vdd gnd cell_6t
Xbit_r133_c115 bl[115] br[115] wl[133] vdd gnd cell_6t
Xbit_r134_c115 bl[115] br[115] wl[134] vdd gnd cell_6t
Xbit_r135_c115 bl[115] br[115] wl[135] vdd gnd cell_6t
Xbit_r136_c115 bl[115] br[115] wl[136] vdd gnd cell_6t
Xbit_r137_c115 bl[115] br[115] wl[137] vdd gnd cell_6t
Xbit_r138_c115 bl[115] br[115] wl[138] vdd gnd cell_6t
Xbit_r139_c115 bl[115] br[115] wl[139] vdd gnd cell_6t
Xbit_r140_c115 bl[115] br[115] wl[140] vdd gnd cell_6t
Xbit_r141_c115 bl[115] br[115] wl[141] vdd gnd cell_6t
Xbit_r142_c115 bl[115] br[115] wl[142] vdd gnd cell_6t
Xbit_r143_c115 bl[115] br[115] wl[143] vdd gnd cell_6t
Xbit_r144_c115 bl[115] br[115] wl[144] vdd gnd cell_6t
Xbit_r145_c115 bl[115] br[115] wl[145] vdd gnd cell_6t
Xbit_r146_c115 bl[115] br[115] wl[146] vdd gnd cell_6t
Xbit_r147_c115 bl[115] br[115] wl[147] vdd gnd cell_6t
Xbit_r148_c115 bl[115] br[115] wl[148] vdd gnd cell_6t
Xbit_r149_c115 bl[115] br[115] wl[149] vdd gnd cell_6t
Xbit_r150_c115 bl[115] br[115] wl[150] vdd gnd cell_6t
Xbit_r151_c115 bl[115] br[115] wl[151] vdd gnd cell_6t
Xbit_r152_c115 bl[115] br[115] wl[152] vdd gnd cell_6t
Xbit_r153_c115 bl[115] br[115] wl[153] vdd gnd cell_6t
Xbit_r154_c115 bl[115] br[115] wl[154] vdd gnd cell_6t
Xbit_r155_c115 bl[115] br[115] wl[155] vdd gnd cell_6t
Xbit_r156_c115 bl[115] br[115] wl[156] vdd gnd cell_6t
Xbit_r157_c115 bl[115] br[115] wl[157] vdd gnd cell_6t
Xbit_r158_c115 bl[115] br[115] wl[158] vdd gnd cell_6t
Xbit_r159_c115 bl[115] br[115] wl[159] vdd gnd cell_6t
Xbit_r160_c115 bl[115] br[115] wl[160] vdd gnd cell_6t
Xbit_r161_c115 bl[115] br[115] wl[161] vdd gnd cell_6t
Xbit_r162_c115 bl[115] br[115] wl[162] vdd gnd cell_6t
Xbit_r163_c115 bl[115] br[115] wl[163] vdd gnd cell_6t
Xbit_r164_c115 bl[115] br[115] wl[164] vdd gnd cell_6t
Xbit_r165_c115 bl[115] br[115] wl[165] vdd gnd cell_6t
Xbit_r166_c115 bl[115] br[115] wl[166] vdd gnd cell_6t
Xbit_r167_c115 bl[115] br[115] wl[167] vdd gnd cell_6t
Xbit_r168_c115 bl[115] br[115] wl[168] vdd gnd cell_6t
Xbit_r169_c115 bl[115] br[115] wl[169] vdd gnd cell_6t
Xbit_r170_c115 bl[115] br[115] wl[170] vdd gnd cell_6t
Xbit_r171_c115 bl[115] br[115] wl[171] vdd gnd cell_6t
Xbit_r172_c115 bl[115] br[115] wl[172] vdd gnd cell_6t
Xbit_r173_c115 bl[115] br[115] wl[173] vdd gnd cell_6t
Xbit_r174_c115 bl[115] br[115] wl[174] vdd gnd cell_6t
Xbit_r175_c115 bl[115] br[115] wl[175] vdd gnd cell_6t
Xbit_r176_c115 bl[115] br[115] wl[176] vdd gnd cell_6t
Xbit_r177_c115 bl[115] br[115] wl[177] vdd gnd cell_6t
Xbit_r178_c115 bl[115] br[115] wl[178] vdd gnd cell_6t
Xbit_r179_c115 bl[115] br[115] wl[179] vdd gnd cell_6t
Xbit_r180_c115 bl[115] br[115] wl[180] vdd gnd cell_6t
Xbit_r181_c115 bl[115] br[115] wl[181] vdd gnd cell_6t
Xbit_r182_c115 bl[115] br[115] wl[182] vdd gnd cell_6t
Xbit_r183_c115 bl[115] br[115] wl[183] vdd gnd cell_6t
Xbit_r184_c115 bl[115] br[115] wl[184] vdd gnd cell_6t
Xbit_r185_c115 bl[115] br[115] wl[185] vdd gnd cell_6t
Xbit_r186_c115 bl[115] br[115] wl[186] vdd gnd cell_6t
Xbit_r187_c115 bl[115] br[115] wl[187] vdd gnd cell_6t
Xbit_r188_c115 bl[115] br[115] wl[188] vdd gnd cell_6t
Xbit_r189_c115 bl[115] br[115] wl[189] vdd gnd cell_6t
Xbit_r190_c115 bl[115] br[115] wl[190] vdd gnd cell_6t
Xbit_r191_c115 bl[115] br[115] wl[191] vdd gnd cell_6t
Xbit_r192_c115 bl[115] br[115] wl[192] vdd gnd cell_6t
Xbit_r193_c115 bl[115] br[115] wl[193] vdd gnd cell_6t
Xbit_r194_c115 bl[115] br[115] wl[194] vdd gnd cell_6t
Xbit_r195_c115 bl[115] br[115] wl[195] vdd gnd cell_6t
Xbit_r196_c115 bl[115] br[115] wl[196] vdd gnd cell_6t
Xbit_r197_c115 bl[115] br[115] wl[197] vdd gnd cell_6t
Xbit_r198_c115 bl[115] br[115] wl[198] vdd gnd cell_6t
Xbit_r199_c115 bl[115] br[115] wl[199] vdd gnd cell_6t
Xbit_r200_c115 bl[115] br[115] wl[200] vdd gnd cell_6t
Xbit_r201_c115 bl[115] br[115] wl[201] vdd gnd cell_6t
Xbit_r202_c115 bl[115] br[115] wl[202] vdd gnd cell_6t
Xbit_r203_c115 bl[115] br[115] wl[203] vdd gnd cell_6t
Xbit_r204_c115 bl[115] br[115] wl[204] vdd gnd cell_6t
Xbit_r205_c115 bl[115] br[115] wl[205] vdd gnd cell_6t
Xbit_r206_c115 bl[115] br[115] wl[206] vdd gnd cell_6t
Xbit_r207_c115 bl[115] br[115] wl[207] vdd gnd cell_6t
Xbit_r208_c115 bl[115] br[115] wl[208] vdd gnd cell_6t
Xbit_r209_c115 bl[115] br[115] wl[209] vdd gnd cell_6t
Xbit_r210_c115 bl[115] br[115] wl[210] vdd gnd cell_6t
Xbit_r211_c115 bl[115] br[115] wl[211] vdd gnd cell_6t
Xbit_r212_c115 bl[115] br[115] wl[212] vdd gnd cell_6t
Xbit_r213_c115 bl[115] br[115] wl[213] vdd gnd cell_6t
Xbit_r214_c115 bl[115] br[115] wl[214] vdd gnd cell_6t
Xbit_r215_c115 bl[115] br[115] wl[215] vdd gnd cell_6t
Xbit_r216_c115 bl[115] br[115] wl[216] vdd gnd cell_6t
Xbit_r217_c115 bl[115] br[115] wl[217] vdd gnd cell_6t
Xbit_r218_c115 bl[115] br[115] wl[218] vdd gnd cell_6t
Xbit_r219_c115 bl[115] br[115] wl[219] vdd gnd cell_6t
Xbit_r220_c115 bl[115] br[115] wl[220] vdd gnd cell_6t
Xbit_r221_c115 bl[115] br[115] wl[221] vdd gnd cell_6t
Xbit_r222_c115 bl[115] br[115] wl[222] vdd gnd cell_6t
Xbit_r223_c115 bl[115] br[115] wl[223] vdd gnd cell_6t
Xbit_r224_c115 bl[115] br[115] wl[224] vdd gnd cell_6t
Xbit_r225_c115 bl[115] br[115] wl[225] vdd gnd cell_6t
Xbit_r226_c115 bl[115] br[115] wl[226] vdd gnd cell_6t
Xbit_r227_c115 bl[115] br[115] wl[227] vdd gnd cell_6t
Xbit_r228_c115 bl[115] br[115] wl[228] vdd gnd cell_6t
Xbit_r229_c115 bl[115] br[115] wl[229] vdd gnd cell_6t
Xbit_r230_c115 bl[115] br[115] wl[230] vdd gnd cell_6t
Xbit_r231_c115 bl[115] br[115] wl[231] vdd gnd cell_6t
Xbit_r232_c115 bl[115] br[115] wl[232] vdd gnd cell_6t
Xbit_r233_c115 bl[115] br[115] wl[233] vdd gnd cell_6t
Xbit_r234_c115 bl[115] br[115] wl[234] vdd gnd cell_6t
Xbit_r235_c115 bl[115] br[115] wl[235] vdd gnd cell_6t
Xbit_r236_c115 bl[115] br[115] wl[236] vdd gnd cell_6t
Xbit_r237_c115 bl[115] br[115] wl[237] vdd gnd cell_6t
Xbit_r238_c115 bl[115] br[115] wl[238] vdd gnd cell_6t
Xbit_r239_c115 bl[115] br[115] wl[239] vdd gnd cell_6t
Xbit_r240_c115 bl[115] br[115] wl[240] vdd gnd cell_6t
Xbit_r241_c115 bl[115] br[115] wl[241] vdd gnd cell_6t
Xbit_r242_c115 bl[115] br[115] wl[242] vdd gnd cell_6t
Xbit_r243_c115 bl[115] br[115] wl[243] vdd gnd cell_6t
Xbit_r244_c115 bl[115] br[115] wl[244] vdd gnd cell_6t
Xbit_r245_c115 bl[115] br[115] wl[245] vdd gnd cell_6t
Xbit_r246_c115 bl[115] br[115] wl[246] vdd gnd cell_6t
Xbit_r247_c115 bl[115] br[115] wl[247] vdd gnd cell_6t
Xbit_r248_c115 bl[115] br[115] wl[248] vdd gnd cell_6t
Xbit_r249_c115 bl[115] br[115] wl[249] vdd gnd cell_6t
Xbit_r250_c115 bl[115] br[115] wl[250] vdd gnd cell_6t
Xbit_r251_c115 bl[115] br[115] wl[251] vdd gnd cell_6t
Xbit_r252_c115 bl[115] br[115] wl[252] vdd gnd cell_6t
Xbit_r253_c115 bl[115] br[115] wl[253] vdd gnd cell_6t
Xbit_r254_c115 bl[115] br[115] wl[254] vdd gnd cell_6t
Xbit_r255_c115 bl[115] br[115] wl[255] vdd gnd cell_6t
Xbit_r0_c116 bl[116] br[116] wl[0] vdd gnd cell_6t
Xbit_r1_c116 bl[116] br[116] wl[1] vdd gnd cell_6t
Xbit_r2_c116 bl[116] br[116] wl[2] vdd gnd cell_6t
Xbit_r3_c116 bl[116] br[116] wl[3] vdd gnd cell_6t
Xbit_r4_c116 bl[116] br[116] wl[4] vdd gnd cell_6t
Xbit_r5_c116 bl[116] br[116] wl[5] vdd gnd cell_6t
Xbit_r6_c116 bl[116] br[116] wl[6] vdd gnd cell_6t
Xbit_r7_c116 bl[116] br[116] wl[7] vdd gnd cell_6t
Xbit_r8_c116 bl[116] br[116] wl[8] vdd gnd cell_6t
Xbit_r9_c116 bl[116] br[116] wl[9] vdd gnd cell_6t
Xbit_r10_c116 bl[116] br[116] wl[10] vdd gnd cell_6t
Xbit_r11_c116 bl[116] br[116] wl[11] vdd gnd cell_6t
Xbit_r12_c116 bl[116] br[116] wl[12] vdd gnd cell_6t
Xbit_r13_c116 bl[116] br[116] wl[13] vdd gnd cell_6t
Xbit_r14_c116 bl[116] br[116] wl[14] vdd gnd cell_6t
Xbit_r15_c116 bl[116] br[116] wl[15] vdd gnd cell_6t
Xbit_r16_c116 bl[116] br[116] wl[16] vdd gnd cell_6t
Xbit_r17_c116 bl[116] br[116] wl[17] vdd gnd cell_6t
Xbit_r18_c116 bl[116] br[116] wl[18] vdd gnd cell_6t
Xbit_r19_c116 bl[116] br[116] wl[19] vdd gnd cell_6t
Xbit_r20_c116 bl[116] br[116] wl[20] vdd gnd cell_6t
Xbit_r21_c116 bl[116] br[116] wl[21] vdd gnd cell_6t
Xbit_r22_c116 bl[116] br[116] wl[22] vdd gnd cell_6t
Xbit_r23_c116 bl[116] br[116] wl[23] vdd gnd cell_6t
Xbit_r24_c116 bl[116] br[116] wl[24] vdd gnd cell_6t
Xbit_r25_c116 bl[116] br[116] wl[25] vdd gnd cell_6t
Xbit_r26_c116 bl[116] br[116] wl[26] vdd gnd cell_6t
Xbit_r27_c116 bl[116] br[116] wl[27] vdd gnd cell_6t
Xbit_r28_c116 bl[116] br[116] wl[28] vdd gnd cell_6t
Xbit_r29_c116 bl[116] br[116] wl[29] vdd gnd cell_6t
Xbit_r30_c116 bl[116] br[116] wl[30] vdd gnd cell_6t
Xbit_r31_c116 bl[116] br[116] wl[31] vdd gnd cell_6t
Xbit_r32_c116 bl[116] br[116] wl[32] vdd gnd cell_6t
Xbit_r33_c116 bl[116] br[116] wl[33] vdd gnd cell_6t
Xbit_r34_c116 bl[116] br[116] wl[34] vdd gnd cell_6t
Xbit_r35_c116 bl[116] br[116] wl[35] vdd gnd cell_6t
Xbit_r36_c116 bl[116] br[116] wl[36] vdd gnd cell_6t
Xbit_r37_c116 bl[116] br[116] wl[37] vdd gnd cell_6t
Xbit_r38_c116 bl[116] br[116] wl[38] vdd gnd cell_6t
Xbit_r39_c116 bl[116] br[116] wl[39] vdd gnd cell_6t
Xbit_r40_c116 bl[116] br[116] wl[40] vdd gnd cell_6t
Xbit_r41_c116 bl[116] br[116] wl[41] vdd gnd cell_6t
Xbit_r42_c116 bl[116] br[116] wl[42] vdd gnd cell_6t
Xbit_r43_c116 bl[116] br[116] wl[43] vdd gnd cell_6t
Xbit_r44_c116 bl[116] br[116] wl[44] vdd gnd cell_6t
Xbit_r45_c116 bl[116] br[116] wl[45] vdd gnd cell_6t
Xbit_r46_c116 bl[116] br[116] wl[46] vdd gnd cell_6t
Xbit_r47_c116 bl[116] br[116] wl[47] vdd gnd cell_6t
Xbit_r48_c116 bl[116] br[116] wl[48] vdd gnd cell_6t
Xbit_r49_c116 bl[116] br[116] wl[49] vdd gnd cell_6t
Xbit_r50_c116 bl[116] br[116] wl[50] vdd gnd cell_6t
Xbit_r51_c116 bl[116] br[116] wl[51] vdd gnd cell_6t
Xbit_r52_c116 bl[116] br[116] wl[52] vdd gnd cell_6t
Xbit_r53_c116 bl[116] br[116] wl[53] vdd gnd cell_6t
Xbit_r54_c116 bl[116] br[116] wl[54] vdd gnd cell_6t
Xbit_r55_c116 bl[116] br[116] wl[55] vdd gnd cell_6t
Xbit_r56_c116 bl[116] br[116] wl[56] vdd gnd cell_6t
Xbit_r57_c116 bl[116] br[116] wl[57] vdd gnd cell_6t
Xbit_r58_c116 bl[116] br[116] wl[58] vdd gnd cell_6t
Xbit_r59_c116 bl[116] br[116] wl[59] vdd gnd cell_6t
Xbit_r60_c116 bl[116] br[116] wl[60] vdd gnd cell_6t
Xbit_r61_c116 bl[116] br[116] wl[61] vdd gnd cell_6t
Xbit_r62_c116 bl[116] br[116] wl[62] vdd gnd cell_6t
Xbit_r63_c116 bl[116] br[116] wl[63] vdd gnd cell_6t
Xbit_r64_c116 bl[116] br[116] wl[64] vdd gnd cell_6t
Xbit_r65_c116 bl[116] br[116] wl[65] vdd gnd cell_6t
Xbit_r66_c116 bl[116] br[116] wl[66] vdd gnd cell_6t
Xbit_r67_c116 bl[116] br[116] wl[67] vdd gnd cell_6t
Xbit_r68_c116 bl[116] br[116] wl[68] vdd gnd cell_6t
Xbit_r69_c116 bl[116] br[116] wl[69] vdd gnd cell_6t
Xbit_r70_c116 bl[116] br[116] wl[70] vdd gnd cell_6t
Xbit_r71_c116 bl[116] br[116] wl[71] vdd gnd cell_6t
Xbit_r72_c116 bl[116] br[116] wl[72] vdd gnd cell_6t
Xbit_r73_c116 bl[116] br[116] wl[73] vdd gnd cell_6t
Xbit_r74_c116 bl[116] br[116] wl[74] vdd gnd cell_6t
Xbit_r75_c116 bl[116] br[116] wl[75] vdd gnd cell_6t
Xbit_r76_c116 bl[116] br[116] wl[76] vdd gnd cell_6t
Xbit_r77_c116 bl[116] br[116] wl[77] vdd gnd cell_6t
Xbit_r78_c116 bl[116] br[116] wl[78] vdd gnd cell_6t
Xbit_r79_c116 bl[116] br[116] wl[79] vdd gnd cell_6t
Xbit_r80_c116 bl[116] br[116] wl[80] vdd gnd cell_6t
Xbit_r81_c116 bl[116] br[116] wl[81] vdd gnd cell_6t
Xbit_r82_c116 bl[116] br[116] wl[82] vdd gnd cell_6t
Xbit_r83_c116 bl[116] br[116] wl[83] vdd gnd cell_6t
Xbit_r84_c116 bl[116] br[116] wl[84] vdd gnd cell_6t
Xbit_r85_c116 bl[116] br[116] wl[85] vdd gnd cell_6t
Xbit_r86_c116 bl[116] br[116] wl[86] vdd gnd cell_6t
Xbit_r87_c116 bl[116] br[116] wl[87] vdd gnd cell_6t
Xbit_r88_c116 bl[116] br[116] wl[88] vdd gnd cell_6t
Xbit_r89_c116 bl[116] br[116] wl[89] vdd gnd cell_6t
Xbit_r90_c116 bl[116] br[116] wl[90] vdd gnd cell_6t
Xbit_r91_c116 bl[116] br[116] wl[91] vdd gnd cell_6t
Xbit_r92_c116 bl[116] br[116] wl[92] vdd gnd cell_6t
Xbit_r93_c116 bl[116] br[116] wl[93] vdd gnd cell_6t
Xbit_r94_c116 bl[116] br[116] wl[94] vdd gnd cell_6t
Xbit_r95_c116 bl[116] br[116] wl[95] vdd gnd cell_6t
Xbit_r96_c116 bl[116] br[116] wl[96] vdd gnd cell_6t
Xbit_r97_c116 bl[116] br[116] wl[97] vdd gnd cell_6t
Xbit_r98_c116 bl[116] br[116] wl[98] vdd gnd cell_6t
Xbit_r99_c116 bl[116] br[116] wl[99] vdd gnd cell_6t
Xbit_r100_c116 bl[116] br[116] wl[100] vdd gnd cell_6t
Xbit_r101_c116 bl[116] br[116] wl[101] vdd gnd cell_6t
Xbit_r102_c116 bl[116] br[116] wl[102] vdd gnd cell_6t
Xbit_r103_c116 bl[116] br[116] wl[103] vdd gnd cell_6t
Xbit_r104_c116 bl[116] br[116] wl[104] vdd gnd cell_6t
Xbit_r105_c116 bl[116] br[116] wl[105] vdd gnd cell_6t
Xbit_r106_c116 bl[116] br[116] wl[106] vdd gnd cell_6t
Xbit_r107_c116 bl[116] br[116] wl[107] vdd gnd cell_6t
Xbit_r108_c116 bl[116] br[116] wl[108] vdd gnd cell_6t
Xbit_r109_c116 bl[116] br[116] wl[109] vdd gnd cell_6t
Xbit_r110_c116 bl[116] br[116] wl[110] vdd gnd cell_6t
Xbit_r111_c116 bl[116] br[116] wl[111] vdd gnd cell_6t
Xbit_r112_c116 bl[116] br[116] wl[112] vdd gnd cell_6t
Xbit_r113_c116 bl[116] br[116] wl[113] vdd gnd cell_6t
Xbit_r114_c116 bl[116] br[116] wl[114] vdd gnd cell_6t
Xbit_r115_c116 bl[116] br[116] wl[115] vdd gnd cell_6t
Xbit_r116_c116 bl[116] br[116] wl[116] vdd gnd cell_6t
Xbit_r117_c116 bl[116] br[116] wl[117] vdd gnd cell_6t
Xbit_r118_c116 bl[116] br[116] wl[118] vdd gnd cell_6t
Xbit_r119_c116 bl[116] br[116] wl[119] vdd gnd cell_6t
Xbit_r120_c116 bl[116] br[116] wl[120] vdd gnd cell_6t
Xbit_r121_c116 bl[116] br[116] wl[121] vdd gnd cell_6t
Xbit_r122_c116 bl[116] br[116] wl[122] vdd gnd cell_6t
Xbit_r123_c116 bl[116] br[116] wl[123] vdd gnd cell_6t
Xbit_r124_c116 bl[116] br[116] wl[124] vdd gnd cell_6t
Xbit_r125_c116 bl[116] br[116] wl[125] vdd gnd cell_6t
Xbit_r126_c116 bl[116] br[116] wl[126] vdd gnd cell_6t
Xbit_r127_c116 bl[116] br[116] wl[127] vdd gnd cell_6t
Xbit_r128_c116 bl[116] br[116] wl[128] vdd gnd cell_6t
Xbit_r129_c116 bl[116] br[116] wl[129] vdd gnd cell_6t
Xbit_r130_c116 bl[116] br[116] wl[130] vdd gnd cell_6t
Xbit_r131_c116 bl[116] br[116] wl[131] vdd gnd cell_6t
Xbit_r132_c116 bl[116] br[116] wl[132] vdd gnd cell_6t
Xbit_r133_c116 bl[116] br[116] wl[133] vdd gnd cell_6t
Xbit_r134_c116 bl[116] br[116] wl[134] vdd gnd cell_6t
Xbit_r135_c116 bl[116] br[116] wl[135] vdd gnd cell_6t
Xbit_r136_c116 bl[116] br[116] wl[136] vdd gnd cell_6t
Xbit_r137_c116 bl[116] br[116] wl[137] vdd gnd cell_6t
Xbit_r138_c116 bl[116] br[116] wl[138] vdd gnd cell_6t
Xbit_r139_c116 bl[116] br[116] wl[139] vdd gnd cell_6t
Xbit_r140_c116 bl[116] br[116] wl[140] vdd gnd cell_6t
Xbit_r141_c116 bl[116] br[116] wl[141] vdd gnd cell_6t
Xbit_r142_c116 bl[116] br[116] wl[142] vdd gnd cell_6t
Xbit_r143_c116 bl[116] br[116] wl[143] vdd gnd cell_6t
Xbit_r144_c116 bl[116] br[116] wl[144] vdd gnd cell_6t
Xbit_r145_c116 bl[116] br[116] wl[145] vdd gnd cell_6t
Xbit_r146_c116 bl[116] br[116] wl[146] vdd gnd cell_6t
Xbit_r147_c116 bl[116] br[116] wl[147] vdd gnd cell_6t
Xbit_r148_c116 bl[116] br[116] wl[148] vdd gnd cell_6t
Xbit_r149_c116 bl[116] br[116] wl[149] vdd gnd cell_6t
Xbit_r150_c116 bl[116] br[116] wl[150] vdd gnd cell_6t
Xbit_r151_c116 bl[116] br[116] wl[151] vdd gnd cell_6t
Xbit_r152_c116 bl[116] br[116] wl[152] vdd gnd cell_6t
Xbit_r153_c116 bl[116] br[116] wl[153] vdd gnd cell_6t
Xbit_r154_c116 bl[116] br[116] wl[154] vdd gnd cell_6t
Xbit_r155_c116 bl[116] br[116] wl[155] vdd gnd cell_6t
Xbit_r156_c116 bl[116] br[116] wl[156] vdd gnd cell_6t
Xbit_r157_c116 bl[116] br[116] wl[157] vdd gnd cell_6t
Xbit_r158_c116 bl[116] br[116] wl[158] vdd gnd cell_6t
Xbit_r159_c116 bl[116] br[116] wl[159] vdd gnd cell_6t
Xbit_r160_c116 bl[116] br[116] wl[160] vdd gnd cell_6t
Xbit_r161_c116 bl[116] br[116] wl[161] vdd gnd cell_6t
Xbit_r162_c116 bl[116] br[116] wl[162] vdd gnd cell_6t
Xbit_r163_c116 bl[116] br[116] wl[163] vdd gnd cell_6t
Xbit_r164_c116 bl[116] br[116] wl[164] vdd gnd cell_6t
Xbit_r165_c116 bl[116] br[116] wl[165] vdd gnd cell_6t
Xbit_r166_c116 bl[116] br[116] wl[166] vdd gnd cell_6t
Xbit_r167_c116 bl[116] br[116] wl[167] vdd gnd cell_6t
Xbit_r168_c116 bl[116] br[116] wl[168] vdd gnd cell_6t
Xbit_r169_c116 bl[116] br[116] wl[169] vdd gnd cell_6t
Xbit_r170_c116 bl[116] br[116] wl[170] vdd gnd cell_6t
Xbit_r171_c116 bl[116] br[116] wl[171] vdd gnd cell_6t
Xbit_r172_c116 bl[116] br[116] wl[172] vdd gnd cell_6t
Xbit_r173_c116 bl[116] br[116] wl[173] vdd gnd cell_6t
Xbit_r174_c116 bl[116] br[116] wl[174] vdd gnd cell_6t
Xbit_r175_c116 bl[116] br[116] wl[175] vdd gnd cell_6t
Xbit_r176_c116 bl[116] br[116] wl[176] vdd gnd cell_6t
Xbit_r177_c116 bl[116] br[116] wl[177] vdd gnd cell_6t
Xbit_r178_c116 bl[116] br[116] wl[178] vdd gnd cell_6t
Xbit_r179_c116 bl[116] br[116] wl[179] vdd gnd cell_6t
Xbit_r180_c116 bl[116] br[116] wl[180] vdd gnd cell_6t
Xbit_r181_c116 bl[116] br[116] wl[181] vdd gnd cell_6t
Xbit_r182_c116 bl[116] br[116] wl[182] vdd gnd cell_6t
Xbit_r183_c116 bl[116] br[116] wl[183] vdd gnd cell_6t
Xbit_r184_c116 bl[116] br[116] wl[184] vdd gnd cell_6t
Xbit_r185_c116 bl[116] br[116] wl[185] vdd gnd cell_6t
Xbit_r186_c116 bl[116] br[116] wl[186] vdd gnd cell_6t
Xbit_r187_c116 bl[116] br[116] wl[187] vdd gnd cell_6t
Xbit_r188_c116 bl[116] br[116] wl[188] vdd gnd cell_6t
Xbit_r189_c116 bl[116] br[116] wl[189] vdd gnd cell_6t
Xbit_r190_c116 bl[116] br[116] wl[190] vdd gnd cell_6t
Xbit_r191_c116 bl[116] br[116] wl[191] vdd gnd cell_6t
Xbit_r192_c116 bl[116] br[116] wl[192] vdd gnd cell_6t
Xbit_r193_c116 bl[116] br[116] wl[193] vdd gnd cell_6t
Xbit_r194_c116 bl[116] br[116] wl[194] vdd gnd cell_6t
Xbit_r195_c116 bl[116] br[116] wl[195] vdd gnd cell_6t
Xbit_r196_c116 bl[116] br[116] wl[196] vdd gnd cell_6t
Xbit_r197_c116 bl[116] br[116] wl[197] vdd gnd cell_6t
Xbit_r198_c116 bl[116] br[116] wl[198] vdd gnd cell_6t
Xbit_r199_c116 bl[116] br[116] wl[199] vdd gnd cell_6t
Xbit_r200_c116 bl[116] br[116] wl[200] vdd gnd cell_6t
Xbit_r201_c116 bl[116] br[116] wl[201] vdd gnd cell_6t
Xbit_r202_c116 bl[116] br[116] wl[202] vdd gnd cell_6t
Xbit_r203_c116 bl[116] br[116] wl[203] vdd gnd cell_6t
Xbit_r204_c116 bl[116] br[116] wl[204] vdd gnd cell_6t
Xbit_r205_c116 bl[116] br[116] wl[205] vdd gnd cell_6t
Xbit_r206_c116 bl[116] br[116] wl[206] vdd gnd cell_6t
Xbit_r207_c116 bl[116] br[116] wl[207] vdd gnd cell_6t
Xbit_r208_c116 bl[116] br[116] wl[208] vdd gnd cell_6t
Xbit_r209_c116 bl[116] br[116] wl[209] vdd gnd cell_6t
Xbit_r210_c116 bl[116] br[116] wl[210] vdd gnd cell_6t
Xbit_r211_c116 bl[116] br[116] wl[211] vdd gnd cell_6t
Xbit_r212_c116 bl[116] br[116] wl[212] vdd gnd cell_6t
Xbit_r213_c116 bl[116] br[116] wl[213] vdd gnd cell_6t
Xbit_r214_c116 bl[116] br[116] wl[214] vdd gnd cell_6t
Xbit_r215_c116 bl[116] br[116] wl[215] vdd gnd cell_6t
Xbit_r216_c116 bl[116] br[116] wl[216] vdd gnd cell_6t
Xbit_r217_c116 bl[116] br[116] wl[217] vdd gnd cell_6t
Xbit_r218_c116 bl[116] br[116] wl[218] vdd gnd cell_6t
Xbit_r219_c116 bl[116] br[116] wl[219] vdd gnd cell_6t
Xbit_r220_c116 bl[116] br[116] wl[220] vdd gnd cell_6t
Xbit_r221_c116 bl[116] br[116] wl[221] vdd gnd cell_6t
Xbit_r222_c116 bl[116] br[116] wl[222] vdd gnd cell_6t
Xbit_r223_c116 bl[116] br[116] wl[223] vdd gnd cell_6t
Xbit_r224_c116 bl[116] br[116] wl[224] vdd gnd cell_6t
Xbit_r225_c116 bl[116] br[116] wl[225] vdd gnd cell_6t
Xbit_r226_c116 bl[116] br[116] wl[226] vdd gnd cell_6t
Xbit_r227_c116 bl[116] br[116] wl[227] vdd gnd cell_6t
Xbit_r228_c116 bl[116] br[116] wl[228] vdd gnd cell_6t
Xbit_r229_c116 bl[116] br[116] wl[229] vdd gnd cell_6t
Xbit_r230_c116 bl[116] br[116] wl[230] vdd gnd cell_6t
Xbit_r231_c116 bl[116] br[116] wl[231] vdd gnd cell_6t
Xbit_r232_c116 bl[116] br[116] wl[232] vdd gnd cell_6t
Xbit_r233_c116 bl[116] br[116] wl[233] vdd gnd cell_6t
Xbit_r234_c116 bl[116] br[116] wl[234] vdd gnd cell_6t
Xbit_r235_c116 bl[116] br[116] wl[235] vdd gnd cell_6t
Xbit_r236_c116 bl[116] br[116] wl[236] vdd gnd cell_6t
Xbit_r237_c116 bl[116] br[116] wl[237] vdd gnd cell_6t
Xbit_r238_c116 bl[116] br[116] wl[238] vdd gnd cell_6t
Xbit_r239_c116 bl[116] br[116] wl[239] vdd gnd cell_6t
Xbit_r240_c116 bl[116] br[116] wl[240] vdd gnd cell_6t
Xbit_r241_c116 bl[116] br[116] wl[241] vdd gnd cell_6t
Xbit_r242_c116 bl[116] br[116] wl[242] vdd gnd cell_6t
Xbit_r243_c116 bl[116] br[116] wl[243] vdd gnd cell_6t
Xbit_r244_c116 bl[116] br[116] wl[244] vdd gnd cell_6t
Xbit_r245_c116 bl[116] br[116] wl[245] vdd gnd cell_6t
Xbit_r246_c116 bl[116] br[116] wl[246] vdd gnd cell_6t
Xbit_r247_c116 bl[116] br[116] wl[247] vdd gnd cell_6t
Xbit_r248_c116 bl[116] br[116] wl[248] vdd gnd cell_6t
Xbit_r249_c116 bl[116] br[116] wl[249] vdd gnd cell_6t
Xbit_r250_c116 bl[116] br[116] wl[250] vdd gnd cell_6t
Xbit_r251_c116 bl[116] br[116] wl[251] vdd gnd cell_6t
Xbit_r252_c116 bl[116] br[116] wl[252] vdd gnd cell_6t
Xbit_r253_c116 bl[116] br[116] wl[253] vdd gnd cell_6t
Xbit_r254_c116 bl[116] br[116] wl[254] vdd gnd cell_6t
Xbit_r255_c116 bl[116] br[116] wl[255] vdd gnd cell_6t
Xbit_r0_c117 bl[117] br[117] wl[0] vdd gnd cell_6t
Xbit_r1_c117 bl[117] br[117] wl[1] vdd gnd cell_6t
Xbit_r2_c117 bl[117] br[117] wl[2] vdd gnd cell_6t
Xbit_r3_c117 bl[117] br[117] wl[3] vdd gnd cell_6t
Xbit_r4_c117 bl[117] br[117] wl[4] vdd gnd cell_6t
Xbit_r5_c117 bl[117] br[117] wl[5] vdd gnd cell_6t
Xbit_r6_c117 bl[117] br[117] wl[6] vdd gnd cell_6t
Xbit_r7_c117 bl[117] br[117] wl[7] vdd gnd cell_6t
Xbit_r8_c117 bl[117] br[117] wl[8] vdd gnd cell_6t
Xbit_r9_c117 bl[117] br[117] wl[9] vdd gnd cell_6t
Xbit_r10_c117 bl[117] br[117] wl[10] vdd gnd cell_6t
Xbit_r11_c117 bl[117] br[117] wl[11] vdd gnd cell_6t
Xbit_r12_c117 bl[117] br[117] wl[12] vdd gnd cell_6t
Xbit_r13_c117 bl[117] br[117] wl[13] vdd gnd cell_6t
Xbit_r14_c117 bl[117] br[117] wl[14] vdd gnd cell_6t
Xbit_r15_c117 bl[117] br[117] wl[15] vdd gnd cell_6t
Xbit_r16_c117 bl[117] br[117] wl[16] vdd gnd cell_6t
Xbit_r17_c117 bl[117] br[117] wl[17] vdd gnd cell_6t
Xbit_r18_c117 bl[117] br[117] wl[18] vdd gnd cell_6t
Xbit_r19_c117 bl[117] br[117] wl[19] vdd gnd cell_6t
Xbit_r20_c117 bl[117] br[117] wl[20] vdd gnd cell_6t
Xbit_r21_c117 bl[117] br[117] wl[21] vdd gnd cell_6t
Xbit_r22_c117 bl[117] br[117] wl[22] vdd gnd cell_6t
Xbit_r23_c117 bl[117] br[117] wl[23] vdd gnd cell_6t
Xbit_r24_c117 bl[117] br[117] wl[24] vdd gnd cell_6t
Xbit_r25_c117 bl[117] br[117] wl[25] vdd gnd cell_6t
Xbit_r26_c117 bl[117] br[117] wl[26] vdd gnd cell_6t
Xbit_r27_c117 bl[117] br[117] wl[27] vdd gnd cell_6t
Xbit_r28_c117 bl[117] br[117] wl[28] vdd gnd cell_6t
Xbit_r29_c117 bl[117] br[117] wl[29] vdd gnd cell_6t
Xbit_r30_c117 bl[117] br[117] wl[30] vdd gnd cell_6t
Xbit_r31_c117 bl[117] br[117] wl[31] vdd gnd cell_6t
Xbit_r32_c117 bl[117] br[117] wl[32] vdd gnd cell_6t
Xbit_r33_c117 bl[117] br[117] wl[33] vdd gnd cell_6t
Xbit_r34_c117 bl[117] br[117] wl[34] vdd gnd cell_6t
Xbit_r35_c117 bl[117] br[117] wl[35] vdd gnd cell_6t
Xbit_r36_c117 bl[117] br[117] wl[36] vdd gnd cell_6t
Xbit_r37_c117 bl[117] br[117] wl[37] vdd gnd cell_6t
Xbit_r38_c117 bl[117] br[117] wl[38] vdd gnd cell_6t
Xbit_r39_c117 bl[117] br[117] wl[39] vdd gnd cell_6t
Xbit_r40_c117 bl[117] br[117] wl[40] vdd gnd cell_6t
Xbit_r41_c117 bl[117] br[117] wl[41] vdd gnd cell_6t
Xbit_r42_c117 bl[117] br[117] wl[42] vdd gnd cell_6t
Xbit_r43_c117 bl[117] br[117] wl[43] vdd gnd cell_6t
Xbit_r44_c117 bl[117] br[117] wl[44] vdd gnd cell_6t
Xbit_r45_c117 bl[117] br[117] wl[45] vdd gnd cell_6t
Xbit_r46_c117 bl[117] br[117] wl[46] vdd gnd cell_6t
Xbit_r47_c117 bl[117] br[117] wl[47] vdd gnd cell_6t
Xbit_r48_c117 bl[117] br[117] wl[48] vdd gnd cell_6t
Xbit_r49_c117 bl[117] br[117] wl[49] vdd gnd cell_6t
Xbit_r50_c117 bl[117] br[117] wl[50] vdd gnd cell_6t
Xbit_r51_c117 bl[117] br[117] wl[51] vdd gnd cell_6t
Xbit_r52_c117 bl[117] br[117] wl[52] vdd gnd cell_6t
Xbit_r53_c117 bl[117] br[117] wl[53] vdd gnd cell_6t
Xbit_r54_c117 bl[117] br[117] wl[54] vdd gnd cell_6t
Xbit_r55_c117 bl[117] br[117] wl[55] vdd gnd cell_6t
Xbit_r56_c117 bl[117] br[117] wl[56] vdd gnd cell_6t
Xbit_r57_c117 bl[117] br[117] wl[57] vdd gnd cell_6t
Xbit_r58_c117 bl[117] br[117] wl[58] vdd gnd cell_6t
Xbit_r59_c117 bl[117] br[117] wl[59] vdd gnd cell_6t
Xbit_r60_c117 bl[117] br[117] wl[60] vdd gnd cell_6t
Xbit_r61_c117 bl[117] br[117] wl[61] vdd gnd cell_6t
Xbit_r62_c117 bl[117] br[117] wl[62] vdd gnd cell_6t
Xbit_r63_c117 bl[117] br[117] wl[63] vdd gnd cell_6t
Xbit_r64_c117 bl[117] br[117] wl[64] vdd gnd cell_6t
Xbit_r65_c117 bl[117] br[117] wl[65] vdd gnd cell_6t
Xbit_r66_c117 bl[117] br[117] wl[66] vdd gnd cell_6t
Xbit_r67_c117 bl[117] br[117] wl[67] vdd gnd cell_6t
Xbit_r68_c117 bl[117] br[117] wl[68] vdd gnd cell_6t
Xbit_r69_c117 bl[117] br[117] wl[69] vdd gnd cell_6t
Xbit_r70_c117 bl[117] br[117] wl[70] vdd gnd cell_6t
Xbit_r71_c117 bl[117] br[117] wl[71] vdd gnd cell_6t
Xbit_r72_c117 bl[117] br[117] wl[72] vdd gnd cell_6t
Xbit_r73_c117 bl[117] br[117] wl[73] vdd gnd cell_6t
Xbit_r74_c117 bl[117] br[117] wl[74] vdd gnd cell_6t
Xbit_r75_c117 bl[117] br[117] wl[75] vdd gnd cell_6t
Xbit_r76_c117 bl[117] br[117] wl[76] vdd gnd cell_6t
Xbit_r77_c117 bl[117] br[117] wl[77] vdd gnd cell_6t
Xbit_r78_c117 bl[117] br[117] wl[78] vdd gnd cell_6t
Xbit_r79_c117 bl[117] br[117] wl[79] vdd gnd cell_6t
Xbit_r80_c117 bl[117] br[117] wl[80] vdd gnd cell_6t
Xbit_r81_c117 bl[117] br[117] wl[81] vdd gnd cell_6t
Xbit_r82_c117 bl[117] br[117] wl[82] vdd gnd cell_6t
Xbit_r83_c117 bl[117] br[117] wl[83] vdd gnd cell_6t
Xbit_r84_c117 bl[117] br[117] wl[84] vdd gnd cell_6t
Xbit_r85_c117 bl[117] br[117] wl[85] vdd gnd cell_6t
Xbit_r86_c117 bl[117] br[117] wl[86] vdd gnd cell_6t
Xbit_r87_c117 bl[117] br[117] wl[87] vdd gnd cell_6t
Xbit_r88_c117 bl[117] br[117] wl[88] vdd gnd cell_6t
Xbit_r89_c117 bl[117] br[117] wl[89] vdd gnd cell_6t
Xbit_r90_c117 bl[117] br[117] wl[90] vdd gnd cell_6t
Xbit_r91_c117 bl[117] br[117] wl[91] vdd gnd cell_6t
Xbit_r92_c117 bl[117] br[117] wl[92] vdd gnd cell_6t
Xbit_r93_c117 bl[117] br[117] wl[93] vdd gnd cell_6t
Xbit_r94_c117 bl[117] br[117] wl[94] vdd gnd cell_6t
Xbit_r95_c117 bl[117] br[117] wl[95] vdd gnd cell_6t
Xbit_r96_c117 bl[117] br[117] wl[96] vdd gnd cell_6t
Xbit_r97_c117 bl[117] br[117] wl[97] vdd gnd cell_6t
Xbit_r98_c117 bl[117] br[117] wl[98] vdd gnd cell_6t
Xbit_r99_c117 bl[117] br[117] wl[99] vdd gnd cell_6t
Xbit_r100_c117 bl[117] br[117] wl[100] vdd gnd cell_6t
Xbit_r101_c117 bl[117] br[117] wl[101] vdd gnd cell_6t
Xbit_r102_c117 bl[117] br[117] wl[102] vdd gnd cell_6t
Xbit_r103_c117 bl[117] br[117] wl[103] vdd gnd cell_6t
Xbit_r104_c117 bl[117] br[117] wl[104] vdd gnd cell_6t
Xbit_r105_c117 bl[117] br[117] wl[105] vdd gnd cell_6t
Xbit_r106_c117 bl[117] br[117] wl[106] vdd gnd cell_6t
Xbit_r107_c117 bl[117] br[117] wl[107] vdd gnd cell_6t
Xbit_r108_c117 bl[117] br[117] wl[108] vdd gnd cell_6t
Xbit_r109_c117 bl[117] br[117] wl[109] vdd gnd cell_6t
Xbit_r110_c117 bl[117] br[117] wl[110] vdd gnd cell_6t
Xbit_r111_c117 bl[117] br[117] wl[111] vdd gnd cell_6t
Xbit_r112_c117 bl[117] br[117] wl[112] vdd gnd cell_6t
Xbit_r113_c117 bl[117] br[117] wl[113] vdd gnd cell_6t
Xbit_r114_c117 bl[117] br[117] wl[114] vdd gnd cell_6t
Xbit_r115_c117 bl[117] br[117] wl[115] vdd gnd cell_6t
Xbit_r116_c117 bl[117] br[117] wl[116] vdd gnd cell_6t
Xbit_r117_c117 bl[117] br[117] wl[117] vdd gnd cell_6t
Xbit_r118_c117 bl[117] br[117] wl[118] vdd gnd cell_6t
Xbit_r119_c117 bl[117] br[117] wl[119] vdd gnd cell_6t
Xbit_r120_c117 bl[117] br[117] wl[120] vdd gnd cell_6t
Xbit_r121_c117 bl[117] br[117] wl[121] vdd gnd cell_6t
Xbit_r122_c117 bl[117] br[117] wl[122] vdd gnd cell_6t
Xbit_r123_c117 bl[117] br[117] wl[123] vdd gnd cell_6t
Xbit_r124_c117 bl[117] br[117] wl[124] vdd gnd cell_6t
Xbit_r125_c117 bl[117] br[117] wl[125] vdd gnd cell_6t
Xbit_r126_c117 bl[117] br[117] wl[126] vdd gnd cell_6t
Xbit_r127_c117 bl[117] br[117] wl[127] vdd gnd cell_6t
Xbit_r128_c117 bl[117] br[117] wl[128] vdd gnd cell_6t
Xbit_r129_c117 bl[117] br[117] wl[129] vdd gnd cell_6t
Xbit_r130_c117 bl[117] br[117] wl[130] vdd gnd cell_6t
Xbit_r131_c117 bl[117] br[117] wl[131] vdd gnd cell_6t
Xbit_r132_c117 bl[117] br[117] wl[132] vdd gnd cell_6t
Xbit_r133_c117 bl[117] br[117] wl[133] vdd gnd cell_6t
Xbit_r134_c117 bl[117] br[117] wl[134] vdd gnd cell_6t
Xbit_r135_c117 bl[117] br[117] wl[135] vdd gnd cell_6t
Xbit_r136_c117 bl[117] br[117] wl[136] vdd gnd cell_6t
Xbit_r137_c117 bl[117] br[117] wl[137] vdd gnd cell_6t
Xbit_r138_c117 bl[117] br[117] wl[138] vdd gnd cell_6t
Xbit_r139_c117 bl[117] br[117] wl[139] vdd gnd cell_6t
Xbit_r140_c117 bl[117] br[117] wl[140] vdd gnd cell_6t
Xbit_r141_c117 bl[117] br[117] wl[141] vdd gnd cell_6t
Xbit_r142_c117 bl[117] br[117] wl[142] vdd gnd cell_6t
Xbit_r143_c117 bl[117] br[117] wl[143] vdd gnd cell_6t
Xbit_r144_c117 bl[117] br[117] wl[144] vdd gnd cell_6t
Xbit_r145_c117 bl[117] br[117] wl[145] vdd gnd cell_6t
Xbit_r146_c117 bl[117] br[117] wl[146] vdd gnd cell_6t
Xbit_r147_c117 bl[117] br[117] wl[147] vdd gnd cell_6t
Xbit_r148_c117 bl[117] br[117] wl[148] vdd gnd cell_6t
Xbit_r149_c117 bl[117] br[117] wl[149] vdd gnd cell_6t
Xbit_r150_c117 bl[117] br[117] wl[150] vdd gnd cell_6t
Xbit_r151_c117 bl[117] br[117] wl[151] vdd gnd cell_6t
Xbit_r152_c117 bl[117] br[117] wl[152] vdd gnd cell_6t
Xbit_r153_c117 bl[117] br[117] wl[153] vdd gnd cell_6t
Xbit_r154_c117 bl[117] br[117] wl[154] vdd gnd cell_6t
Xbit_r155_c117 bl[117] br[117] wl[155] vdd gnd cell_6t
Xbit_r156_c117 bl[117] br[117] wl[156] vdd gnd cell_6t
Xbit_r157_c117 bl[117] br[117] wl[157] vdd gnd cell_6t
Xbit_r158_c117 bl[117] br[117] wl[158] vdd gnd cell_6t
Xbit_r159_c117 bl[117] br[117] wl[159] vdd gnd cell_6t
Xbit_r160_c117 bl[117] br[117] wl[160] vdd gnd cell_6t
Xbit_r161_c117 bl[117] br[117] wl[161] vdd gnd cell_6t
Xbit_r162_c117 bl[117] br[117] wl[162] vdd gnd cell_6t
Xbit_r163_c117 bl[117] br[117] wl[163] vdd gnd cell_6t
Xbit_r164_c117 bl[117] br[117] wl[164] vdd gnd cell_6t
Xbit_r165_c117 bl[117] br[117] wl[165] vdd gnd cell_6t
Xbit_r166_c117 bl[117] br[117] wl[166] vdd gnd cell_6t
Xbit_r167_c117 bl[117] br[117] wl[167] vdd gnd cell_6t
Xbit_r168_c117 bl[117] br[117] wl[168] vdd gnd cell_6t
Xbit_r169_c117 bl[117] br[117] wl[169] vdd gnd cell_6t
Xbit_r170_c117 bl[117] br[117] wl[170] vdd gnd cell_6t
Xbit_r171_c117 bl[117] br[117] wl[171] vdd gnd cell_6t
Xbit_r172_c117 bl[117] br[117] wl[172] vdd gnd cell_6t
Xbit_r173_c117 bl[117] br[117] wl[173] vdd gnd cell_6t
Xbit_r174_c117 bl[117] br[117] wl[174] vdd gnd cell_6t
Xbit_r175_c117 bl[117] br[117] wl[175] vdd gnd cell_6t
Xbit_r176_c117 bl[117] br[117] wl[176] vdd gnd cell_6t
Xbit_r177_c117 bl[117] br[117] wl[177] vdd gnd cell_6t
Xbit_r178_c117 bl[117] br[117] wl[178] vdd gnd cell_6t
Xbit_r179_c117 bl[117] br[117] wl[179] vdd gnd cell_6t
Xbit_r180_c117 bl[117] br[117] wl[180] vdd gnd cell_6t
Xbit_r181_c117 bl[117] br[117] wl[181] vdd gnd cell_6t
Xbit_r182_c117 bl[117] br[117] wl[182] vdd gnd cell_6t
Xbit_r183_c117 bl[117] br[117] wl[183] vdd gnd cell_6t
Xbit_r184_c117 bl[117] br[117] wl[184] vdd gnd cell_6t
Xbit_r185_c117 bl[117] br[117] wl[185] vdd gnd cell_6t
Xbit_r186_c117 bl[117] br[117] wl[186] vdd gnd cell_6t
Xbit_r187_c117 bl[117] br[117] wl[187] vdd gnd cell_6t
Xbit_r188_c117 bl[117] br[117] wl[188] vdd gnd cell_6t
Xbit_r189_c117 bl[117] br[117] wl[189] vdd gnd cell_6t
Xbit_r190_c117 bl[117] br[117] wl[190] vdd gnd cell_6t
Xbit_r191_c117 bl[117] br[117] wl[191] vdd gnd cell_6t
Xbit_r192_c117 bl[117] br[117] wl[192] vdd gnd cell_6t
Xbit_r193_c117 bl[117] br[117] wl[193] vdd gnd cell_6t
Xbit_r194_c117 bl[117] br[117] wl[194] vdd gnd cell_6t
Xbit_r195_c117 bl[117] br[117] wl[195] vdd gnd cell_6t
Xbit_r196_c117 bl[117] br[117] wl[196] vdd gnd cell_6t
Xbit_r197_c117 bl[117] br[117] wl[197] vdd gnd cell_6t
Xbit_r198_c117 bl[117] br[117] wl[198] vdd gnd cell_6t
Xbit_r199_c117 bl[117] br[117] wl[199] vdd gnd cell_6t
Xbit_r200_c117 bl[117] br[117] wl[200] vdd gnd cell_6t
Xbit_r201_c117 bl[117] br[117] wl[201] vdd gnd cell_6t
Xbit_r202_c117 bl[117] br[117] wl[202] vdd gnd cell_6t
Xbit_r203_c117 bl[117] br[117] wl[203] vdd gnd cell_6t
Xbit_r204_c117 bl[117] br[117] wl[204] vdd gnd cell_6t
Xbit_r205_c117 bl[117] br[117] wl[205] vdd gnd cell_6t
Xbit_r206_c117 bl[117] br[117] wl[206] vdd gnd cell_6t
Xbit_r207_c117 bl[117] br[117] wl[207] vdd gnd cell_6t
Xbit_r208_c117 bl[117] br[117] wl[208] vdd gnd cell_6t
Xbit_r209_c117 bl[117] br[117] wl[209] vdd gnd cell_6t
Xbit_r210_c117 bl[117] br[117] wl[210] vdd gnd cell_6t
Xbit_r211_c117 bl[117] br[117] wl[211] vdd gnd cell_6t
Xbit_r212_c117 bl[117] br[117] wl[212] vdd gnd cell_6t
Xbit_r213_c117 bl[117] br[117] wl[213] vdd gnd cell_6t
Xbit_r214_c117 bl[117] br[117] wl[214] vdd gnd cell_6t
Xbit_r215_c117 bl[117] br[117] wl[215] vdd gnd cell_6t
Xbit_r216_c117 bl[117] br[117] wl[216] vdd gnd cell_6t
Xbit_r217_c117 bl[117] br[117] wl[217] vdd gnd cell_6t
Xbit_r218_c117 bl[117] br[117] wl[218] vdd gnd cell_6t
Xbit_r219_c117 bl[117] br[117] wl[219] vdd gnd cell_6t
Xbit_r220_c117 bl[117] br[117] wl[220] vdd gnd cell_6t
Xbit_r221_c117 bl[117] br[117] wl[221] vdd gnd cell_6t
Xbit_r222_c117 bl[117] br[117] wl[222] vdd gnd cell_6t
Xbit_r223_c117 bl[117] br[117] wl[223] vdd gnd cell_6t
Xbit_r224_c117 bl[117] br[117] wl[224] vdd gnd cell_6t
Xbit_r225_c117 bl[117] br[117] wl[225] vdd gnd cell_6t
Xbit_r226_c117 bl[117] br[117] wl[226] vdd gnd cell_6t
Xbit_r227_c117 bl[117] br[117] wl[227] vdd gnd cell_6t
Xbit_r228_c117 bl[117] br[117] wl[228] vdd gnd cell_6t
Xbit_r229_c117 bl[117] br[117] wl[229] vdd gnd cell_6t
Xbit_r230_c117 bl[117] br[117] wl[230] vdd gnd cell_6t
Xbit_r231_c117 bl[117] br[117] wl[231] vdd gnd cell_6t
Xbit_r232_c117 bl[117] br[117] wl[232] vdd gnd cell_6t
Xbit_r233_c117 bl[117] br[117] wl[233] vdd gnd cell_6t
Xbit_r234_c117 bl[117] br[117] wl[234] vdd gnd cell_6t
Xbit_r235_c117 bl[117] br[117] wl[235] vdd gnd cell_6t
Xbit_r236_c117 bl[117] br[117] wl[236] vdd gnd cell_6t
Xbit_r237_c117 bl[117] br[117] wl[237] vdd gnd cell_6t
Xbit_r238_c117 bl[117] br[117] wl[238] vdd gnd cell_6t
Xbit_r239_c117 bl[117] br[117] wl[239] vdd gnd cell_6t
Xbit_r240_c117 bl[117] br[117] wl[240] vdd gnd cell_6t
Xbit_r241_c117 bl[117] br[117] wl[241] vdd gnd cell_6t
Xbit_r242_c117 bl[117] br[117] wl[242] vdd gnd cell_6t
Xbit_r243_c117 bl[117] br[117] wl[243] vdd gnd cell_6t
Xbit_r244_c117 bl[117] br[117] wl[244] vdd gnd cell_6t
Xbit_r245_c117 bl[117] br[117] wl[245] vdd gnd cell_6t
Xbit_r246_c117 bl[117] br[117] wl[246] vdd gnd cell_6t
Xbit_r247_c117 bl[117] br[117] wl[247] vdd gnd cell_6t
Xbit_r248_c117 bl[117] br[117] wl[248] vdd gnd cell_6t
Xbit_r249_c117 bl[117] br[117] wl[249] vdd gnd cell_6t
Xbit_r250_c117 bl[117] br[117] wl[250] vdd gnd cell_6t
Xbit_r251_c117 bl[117] br[117] wl[251] vdd gnd cell_6t
Xbit_r252_c117 bl[117] br[117] wl[252] vdd gnd cell_6t
Xbit_r253_c117 bl[117] br[117] wl[253] vdd gnd cell_6t
Xbit_r254_c117 bl[117] br[117] wl[254] vdd gnd cell_6t
Xbit_r255_c117 bl[117] br[117] wl[255] vdd gnd cell_6t
Xbit_r0_c118 bl[118] br[118] wl[0] vdd gnd cell_6t
Xbit_r1_c118 bl[118] br[118] wl[1] vdd gnd cell_6t
Xbit_r2_c118 bl[118] br[118] wl[2] vdd gnd cell_6t
Xbit_r3_c118 bl[118] br[118] wl[3] vdd gnd cell_6t
Xbit_r4_c118 bl[118] br[118] wl[4] vdd gnd cell_6t
Xbit_r5_c118 bl[118] br[118] wl[5] vdd gnd cell_6t
Xbit_r6_c118 bl[118] br[118] wl[6] vdd gnd cell_6t
Xbit_r7_c118 bl[118] br[118] wl[7] vdd gnd cell_6t
Xbit_r8_c118 bl[118] br[118] wl[8] vdd gnd cell_6t
Xbit_r9_c118 bl[118] br[118] wl[9] vdd gnd cell_6t
Xbit_r10_c118 bl[118] br[118] wl[10] vdd gnd cell_6t
Xbit_r11_c118 bl[118] br[118] wl[11] vdd gnd cell_6t
Xbit_r12_c118 bl[118] br[118] wl[12] vdd gnd cell_6t
Xbit_r13_c118 bl[118] br[118] wl[13] vdd gnd cell_6t
Xbit_r14_c118 bl[118] br[118] wl[14] vdd gnd cell_6t
Xbit_r15_c118 bl[118] br[118] wl[15] vdd gnd cell_6t
Xbit_r16_c118 bl[118] br[118] wl[16] vdd gnd cell_6t
Xbit_r17_c118 bl[118] br[118] wl[17] vdd gnd cell_6t
Xbit_r18_c118 bl[118] br[118] wl[18] vdd gnd cell_6t
Xbit_r19_c118 bl[118] br[118] wl[19] vdd gnd cell_6t
Xbit_r20_c118 bl[118] br[118] wl[20] vdd gnd cell_6t
Xbit_r21_c118 bl[118] br[118] wl[21] vdd gnd cell_6t
Xbit_r22_c118 bl[118] br[118] wl[22] vdd gnd cell_6t
Xbit_r23_c118 bl[118] br[118] wl[23] vdd gnd cell_6t
Xbit_r24_c118 bl[118] br[118] wl[24] vdd gnd cell_6t
Xbit_r25_c118 bl[118] br[118] wl[25] vdd gnd cell_6t
Xbit_r26_c118 bl[118] br[118] wl[26] vdd gnd cell_6t
Xbit_r27_c118 bl[118] br[118] wl[27] vdd gnd cell_6t
Xbit_r28_c118 bl[118] br[118] wl[28] vdd gnd cell_6t
Xbit_r29_c118 bl[118] br[118] wl[29] vdd gnd cell_6t
Xbit_r30_c118 bl[118] br[118] wl[30] vdd gnd cell_6t
Xbit_r31_c118 bl[118] br[118] wl[31] vdd gnd cell_6t
Xbit_r32_c118 bl[118] br[118] wl[32] vdd gnd cell_6t
Xbit_r33_c118 bl[118] br[118] wl[33] vdd gnd cell_6t
Xbit_r34_c118 bl[118] br[118] wl[34] vdd gnd cell_6t
Xbit_r35_c118 bl[118] br[118] wl[35] vdd gnd cell_6t
Xbit_r36_c118 bl[118] br[118] wl[36] vdd gnd cell_6t
Xbit_r37_c118 bl[118] br[118] wl[37] vdd gnd cell_6t
Xbit_r38_c118 bl[118] br[118] wl[38] vdd gnd cell_6t
Xbit_r39_c118 bl[118] br[118] wl[39] vdd gnd cell_6t
Xbit_r40_c118 bl[118] br[118] wl[40] vdd gnd cell_6t
Xbit_r41_c118 bl[118] br[118] wl[41] vdd gnd cell_6t
Xbit_r42_c118 bl[118] br[118] wl[42] vdd gnd cell_6t
Xbit_r43_c118 bl[118] br[118] wl[43] vdd gnd cell_6t
Xbit_r44_c118 bl[118] br[118] wl[44] vdd gnd cell_6t
Xbit_r45_c118 bl[118] br[118] wl[45] vdd gnd cell_6t
Xbit_r46_c118 bl[118] br[118] wl[46] vdd gnd cell_6t
Xbit_r47_c118 bl[118] br[118] wl[47] vdd gnd cell_6t
Xbit_r48_c118 bl[118] br[118] wl[48] vdd gnd cell_6t
Xbit_r49_c118 bl[118] br[118] wl[49] vdd gnd cell_6t
Xbit_r50_c118 bl[118] br[118] wl[50] vdd gnd cell_6t
Xbit_r51_c118 bl[118] br[118] wl[51] vdd gnd cell_6t
Xbit_r52_c118 bl[118] br[118] wl[52] vdd gnd cell_6t
Xbit_r53_c118 bl[118] br[118] wl[53] vdd gnd cell_6t
Xbit_r54_c118 bl[118] br[118] wl[54] vdd gnd cell_6t
Xbit_r55_c118 bl[118] br[118] wl[55] vdd gnd cell_6t
Xbit_r56_c118 bl[118] br[118] wl[56] vdd gnd cell_6t
Xbit_r57_c118 bl[118] br[118] wl[57] vdd gnd cell_6t
Xbit_r58_c118 bl[118] br[118] wl[58] vdd gnd cell_6t
Xbit_r59_c118 bl[118] br[118] wl[59] vdd gnd cell_6t
Xbit_r60_c118 bl[118] br[118] wl[60] vdd gnd cell_6t
Xbit_r61_c118 bl[118] br[118] wl[61] vdd gnd cell_6t
Xbit_r62_c118 bl[118] br[118] wl[62] vdd gnd cell_6t
Xbit_r63_c118 bl[118] br[118] wl[63] vdd gnd cell_6t
Xbit_r64_c118 bl[118] br[118] wl[64] vdd gnd cell_6t
Xbit_r65_c118 bl[118] br[118] wl[65] vdd gnd cell_6t
Xbit_r66_c118 bl[118] br[118] wl[66] vdd gnd cell_6t
Xbit_r67_c118 bl[118] br[118] wl[67] vdd gnd cell_6t
Xbit_r68_c118 bl[118] br[118] wl[68] vdd gnd cell_6t
Xbit_r69_c118 bl[118] br[118] wl[69] vdd gnd cell_6t
Xbit_r70_c118 bl[118] br[118] wl[70] vdd gnd cell_6t
Xbit_r71_c118 bl[118] br[118] wl[71] vdd gnd cell_6t
Xbit_r72_c118 bl[118] br[118] wl[72] vdd gnd cell_6t
Xbit_r73_c118 bl[118] br[118] wl[73] vdd gnd cell_6t
Xbit_r74_c118 bl[118] br[118] wl[74] vdd gnd cell_6t
Xbit_r75_c118 bl[118] br[118] wl[75] vdd gnd cell_6t
Xbit_r76_c118 bl[118] br[118] wl[76] vdd gnd cell_6t
Xbit_r77_c118 bl[118] br[118] wl[77] vdd gnd cell_6t
Xbit_r78_c118 bl[118] br[118] wl[78] vdd gnd cell_6t
Xbit_r79_c118 bl[118] br[118] wl[79] vdd gnd cell_6t
Xbit_r80_c118 bl[118] br[118] wl[80] vdd gnd cell_6t
Xbit_r81_c118 bl[118] br[118] wl[81] vdd gnd cell_6t
Xbit_r82_c118 bl[118] br[118] wl[82] vdd gnd cell_6t
Xbit_r83_c118 bl[118] br[118] wl[83] vdd gnd cell_6t
Xbit_r84_c118 bl[118] br[118] wl[84] vdd gnd cell_6t
Xbit_r85_c118 bl[118] br[118] wl[85] vdd gnd cell_6t
Xbit_r86_c118 bl[118] br[118] wl[86] vdd gnd cell_6t
Xbit_r87_c118 bl[118] br[118] wl[87] vdd gnd cell_6t
Xbit_r88_c118 bl[118] br[118] wl[88] vdd gnd cell_6t
Xbit_r89_c118 bl[118] br[118] wl[89] vdd gnd cell_6t
Xbit_r90_c118 bl[118] br[118] wl[90] vdd gnd cell_6t
Xbit_r91_c118 bl[118] br[118] wl[91] vdd gnd cell_6t
Xbit_r92_c118 bl[118] br[118] wl[92] vdd gnd cell_6t
Xbit_r93_c118 bl[118] br[118] wl[93] vdd gnd cell_6t
Xbit_r94_c118 bl[118] br[118] wl[94] vdd gnd cell_6t
Xbit_r95_c118 bl[118] br[118] wl[95] vdd gnd cell_6t
Xbit_r96_c118 bl[118] br[118] wl[96] vdd gnd cell_6t
Xbit_r97_c118 bl[118] br[118] wl[97] vdd gnd cell_6t
Xbit_r98_c118 bl[118] br[118] wl[98] vdd gnd cell_6t
Xbit_r99_c118 bl[118] br[118] wl[99] vdd gnd cell_6t
Xbit_r100_c118 bl[118] br[118] wl[100] vdd gnd cell_6t
Xbit_r101_c118 bl[118] br[118] wl[101] vdd gnd cell_6t
Xbit_r102_c118 bl[118] br[118] wl[102] vdd gnd cell_6t
Xbit_r103_c118 bl[118] br[118] wl[103] vdd gnd cell_6t
Xbit_r104_c118 bl[118] br[118] wl[104] vdd gnd cell_6t
Xbit_r105_c118 bl[118] br[118] wl[105] vdd gnd cell_6t
Xbit_r106_c118 bl[118] br[118] wl[106] vdd gnd cell_6t
Xbit_r107_c118 bl[118] br[118] wl[107] vdd gnd cell_6t
Xbit_r108_c118 bl[118] br[118] wl[108] vdd gnd cell_6t
Xbit_r109_c118 bl[118] br[118] wl[109] vdd gnd cell_6t
Xbit_r110_c118 bl[118] br[118] wl[110] vdd gnd cell_6t
Xbit_r111_c118 bl[118] br[118] wl[111] vdd gnd cell_6t
Xbit_r112_c118 bl[118] br[118] wl[112] vdd gnd cell_6t
Xbit_r113_c118 bl[118] br[118] wl[113] vdd gnd cell_6t
Xbit_r114_c118 bl[118] br[118] wl[114] vdd gnd cell_6t
Xbit_r115_c118 bl[118] br[118] wl[115] vdd gnd cell_6t
Xbit_r116_c118 bl[118] br[118] wl[116] vdd gnd cell_6t
Xbit_r117_c118 bl[118] br[118] wl[117] vdd gnd cell_6t
Xbit_r118_c118 bl[118] br[118] wl[118] vdd gnd cell_6t
Xbit_r119_c118 bl[118] br[118] wl[119] vdd gnd cell_6t
Xbit_r120_c118 bl[118] br[118] wl[120] vdd gnd cell_6t
Xbit_r121_c118 bl[118] br[118] wl[121] vdd gnd cell_6t
Xbit_r122_c118 bl[118] br[118] wl[122] vdd gnd cell_6t
Xbit_r123_c118 bl[118] br[118] wl[123] vdd gnd cell_6t
Xbit_r124_c118 bl[118] br[118] wl[124] vdd gnd cell_6t
Xbit_r125_c118 bl[118] br[118] wl[125] vdd gnd cell_6t
Xbit_r126_c118 bl[118] br[118] wl[126] vdd gnd cell_6t
Xbit_r127_c118 bl[118] br[118] wl[127] vdd gnd cell_6t
Xbit_r128_c118 bl[118] br[118] wl[128] vdd gnd cell_6t
Xbit_r129_c118 bl[118] br[118] wl[129] vdd gnd cell_6t
Xbit_r130_c118 bl[118] br[118] wl[130] vdd gnd cell_6t
Xbit_r131_c118 bl[118] br[118] wl[131] vdd gnd cell_6t
Xbit_r132_c118 bl[118] br[118] wl[132] vdd gnd cell_6t
Xbit_r133_c118 bl[118] br[118] wl[133] vdd gnd cell_6t
Xbit_r134_c118 bl[118] br[118] wl[134] vdd gnd cell_6t
Xbit_r135_c118 bl[118] br[118] wl[135] vdd gnd cell_6t
Xbit_r136_c118 bl[118] br[118] wl[136] vdd gnd cell_6t
Xbit_r137_c118 bl[118] br[118] wl[137] vdd gnd cell_6t
Xbit_r138_c118 bl[118] br[118] wl[138] vdd gnd cell_6t
Xbit_r139_c118 bl[118] br[118] wl[139] vdd gnd cell_6t
Xbit_r140_c118 bl[118] br[118] wl[140] vdd gnd cell_6t
Xbit_r141_c118 bl[118] br[118] wl[141] vdd gnd cell_6t
Xbit_r142_c118 bl[118] br[118] wl[142] vdd gnd cell_6t
Xbit_r143_c118 bl[118] br[118] wl[143] vdd gnd cell_6t
Xbit_r144_c118 bl[118] br[118] wl[144] vdd gnd cell_6t
Xbit_r145_c118 bl[118] br[118] wl[145] vdd gnd cell_6t
Xbit_r146_c118 bl[118] br[118] wl[146] vdd gnd cell_6t
Xbit_r147_c118 bl[118] br[118] wl[147] vdd gnd cell_6t
Xbit_r148_c118 bl[118] br[118] wl[148] vdd gnd cell_6t
Xbit_r149_c118 bl[118] br[118] wl[149] vdd gnd cell_6t
Xbit_r150_c118 bl[118] br[118] wl[150] vdd gnd cell_6t
Xbit_r151_c118 bl[118] br[118] wl[151] vdd gnd cell_6t
Xbit_r152_c118 bl[118] br[118] wl[152] vdd gnd cell_6t
Xbit_r153_c118 bl[118] br[118] wl[153] vdd gnd cell_6t
Xbit_r154_c118 bl[118] br[118] wl[154] vdd gnd cell_6t
Xbit_r155_c118 bl[118] br[118] wl[155] vdd gnd cell_6t
Xbit_r156_c118 bl[118] br[118] wl[156] vdd gnd cell_6t
Xbit_r157_c118 bl[118] br[118] wl[157] vdd gnd cell_6t
Xbit_r158_c118 bl[118] br[118] wl[158] vdd gnd cell_6t
Xbit_r159_c118 bl[118] br[118] wl[159] vdd gnd cell_6t
Xbit_r160_c118 bl[118] br[118] wl[160] vdd gnd cell_6t
Xbit_r161_c118 bl[118] br[118] wl[161] vdd gnd cell_6t
Xbit_r162_c118 bl[118] br[118] wl[162] vdd gnd cell_6t
Xbit_r163_c118 bl[118] br[118] wl[163] vdd gnd cell_6t
Xbit_r164_c118 bl[118] br[118] wl[164] vdd gnd cell_6t
Xbit_r165_c118 bl[118] br[118] wl[165] vdd gnd cell_6t
Xbit_r166_c118 bl[118] br[118] wl[166] vdd gnd cell_6t
Xbit_r167_c118 bl[118] br[118] wl[167] vdd gnd cell_6t
Xbit_r168_c118 bl[118] br[118] wl[168] vdd gnd cell_6t
Xbit_r169_c118 bl[118] br[118] wl[169] vdd gnd cell_6t
Xbit_r170_c118 bl[118] br[118] wl[170] vdd gnd cell_6t
Xbit_r171_c118 bl[118] br[118] wl[171] vdd gnd cell_6t
Xbit_r172_c118 bl[118] br[118] wl[172] vdd gnd cell_6t
Xbit_r173_c118 bl[118] br[118] wl[173] vdd gnd cell_6t
Xbit_r174_c118 bl[118] br[118] wl[174] vdd gnd cell_6t
Xbit_r175_c118 bl[118] br[118] wl[175] vdd gnd cell_6t
Xbit_r176_c118 bl[118] br[118] wl[176] vdd gnd cell_6t
Xbit_r177_c118 bl[118] br[118] wl[177] vdd gnd cell_6t
Xbit_r178_c118 bl[118] br[118] wl[178] vdd gnd cell_6t
Xbit_r179_c118 bl[118] br[118] wl[179] vdd gnd cell_6t
Xbit_r180_c118 bl[118] br[118] wl[180] vdd gnd cell_6t
Xbit_r181_c118 bl[118] br[118] wl[181] vdd gnd cell_6t
Xbit_r182_c118 bl[118] br[118] wl[182] vdd gnd cell_6t
Xbit_r183_c118 bl[118] br[118] wl[183] vdd gnd cell_6t
Xbit_r184_c118 bl[118] br[118] wl[184] vdd gnd cell_6t
Xbit_r185_c118 bl[118] br[118] wl[185] vdd gnd cell_6t
Xbit_r186_c118 bl[118] br[118] wl[186] vdd gnd cell_6t
Xbit_r187_c118 bl[118] br[118] wl[187] vdd gnd cell_6t
Xbit_r188_c118 bl[118] br[118] wl[188] vdd gnd cell_6t
Xbit_r189_c118 bl[118] br[118] wl[189] vdd gnd cell_6t
Xbit_r190_c118 bl[118] br[118] wl[190] vdd gnd cell_6t
Xbit_r191_c118 bl[118] br[118] wl[191] vdd gnd cell_6t
Xbit_r192_c118 bl[118] br[118] wl[192] vdd gnd cell_6t
Xbit_r193_c118 bl[118] br[118] wl[193] vdd gnd cell_6t
Xbit_r194_c118 bl[118] br[118] wl[194] vdd gnd cell_6t
Xbit_r195_c118 bl[118] br[118] wl[195] vdd gnd cell_6t
Xbit_r196_c118 bl[118] br[118] wl[196] vdd gnd cell_6t
Xbit_r197_c118 bl[118] br[118] wl[197] vdd gnd cell_6t
Xbit_r198_c118 bl[118] br[118] wl[198] vdd gnd cell_6t
Xbit_r199_c118 bl[118] br[118] wl[199] vdd gnd cell_6t
Xbit_r200_c118 bl[118] br[118] wl[200] vdd gnd cell_6t
Xbit_r201_c118 bl[118] br[118] wl[201] vdd gnd cell_6t
Xbit_r202_c118 bl[118] br[118] wl[202] vdd gnd cell_6t
Xbit_r203_c118 bl[118] br[118] wl[203] vdd gnd cell_6t
Xbit_r204_c118 bl[118] br[118] wl[204] vdd gnd cell_6t
Xbit_r205_c118 bl[118] br[118] wl[205] vdd gnd cell_6t
Xbit_r206_c118 bl[118] br[118] wl[206] vdd gnd cell_6t
Xbit_r207_c118 bl[118] br[118] wl[207] vdd gnd cell_6t
Xbit_r208_c118 bl[118] br[118] wl[208] vdd gnd cell_6t
Xbit_r209_c118 bl[118] br[118] wl[209] vdd gnd cell_6t
Xbit_r210_c118 bl[118] br[118] wl[210] vdd gnd cell_6t
Xbit_r211_c118 bl[118] br[118] wl[211] vdd gnd cell_6t
Xbit_r212_c118 bl[118] br[118] wl[212] vdd gnd cell_6t
Xbit_r213_c118 bl[118] br[118] wl[213] vdd gnd cell_6t
Xbit_r214_c118 bl[118] br[118] wl[214] vdd gnd cell_6t
Xbit_r215_c118 bl[118] br[118] wl[215] vdd gnd cell_6t
Xbit_r216_c118 bl[118] br[118] wl[216] vdd gnd cell_6t
Xbit_r217_c118 bl[118] br[118] wl[217] vdd gnd cell_6t
Xbit_r218_c118 bl[118] br[118] wl[218] vdd gnd cell_6t
Xbit_r219_c118 bl[118] br[118] wl[219] vdd gnd cell_6t
Xbit_r220_c118 bl[118] br[118] wl[220] vdd gnd cell_6t
Xbit_r221_c118 bl[118] br[118] wl[221] vdd gnd cell_6t
Xbit_r222_c118 bl[118] br[118] wl[222] vdd gnd cell_6t
Xbit_r223_c118 bl[118] br[118] wl[223] vdd gnd cell_6t
Xbit_r224_c118 bl[118] br[118] wl[224] vdd gnd cell_6t
Xbit_r225_c118 bl[118] br[118] wl[225] vdd gnd cell_6t
Xbit_r226_c118 bl[118] br[118] wl[226] vdd gnd cell_6t
Xbit_r227_c118 bl[118] br[118] wl[227] vdd gnd cell_6t
Xbit_r228_c118 bl[118] br[118] wl[228] vdd gnd cell_6t
Xbit_r229_c118 bl[118] br[118] wl[229] vdd gnd cell_6t
Xbit_r230_c118 bl[118] br[118] wl[230] vdd gnd cell_6t
Xbit_r231_c118 bl[118] br[118] wl[231] vdd gnd cell_6t
Xbit_r232_c118 bl[118] br[118] wl[232] vdd gnd cell_6t
Xbit_r233_c118 bl[118] br[118] wl[233] vdd gnd cell_6t
Xbit_r234_c118 bl[118] br[118] wl[234] vdd gnd cell_6t
Xbit_r235_c118 bl[118] br[118] wl[235] vdd gnd cell_6t
Xbit_r236_c118 bl[118] br[118] wl[236] vdd gnd cell_6t
Xbit_r237_c118 bl[118] br[118] wl[237] vdd gnd cell_6t
Xbit_r238_c118 bl[118] br[118] wl[238] vdd gnd cell_6t
Xbit_r239_c118 bl[118] br[118] wl[239] vdd gnd cell_6t
Xbit_r240_c118 bl[118] br[118] wl[240] vdd gnd cell_6t
Xbit_r241_c118 bl[118] br[118] wl[241] vdd gnd cell_6t
Xbit_r242_c118 bl[118] br[118] wl[242] vdd gnd cell_6t
Xbit_r243_c118 bl[118] br[118] wl[243] vdd gnd cell_6t
Xbit_r244_c118 bl[118] br[118] wl[244] vdd gnd cell_6t
Xbit_r245_c118 bl[118] br[118] wl[245] vdd gnd cell_6t
Xbit_r246_c118 bl[118] br[118] wl[246] vdd gnd cell_6t
Xbit_r247_c118 bl[118] br[118] wl[247] vdd gnd cell_6t
Xbit_r248_c118 bl[118] br[118] wl[248] vdd gnd cell_6t
Xbit_r249_c118 bl[118] br[118] wl[249] vdd gnd cell_6t
Xbit_r250_c118 bl[118] br[118] wl[250] vdd gnd cell_6t
Xbit_r251_c118 bl[118] br[118] wl[251] vdd gnd cell_6t
Xbit_r252_c118 bl[118] br[118] wl[252] vdd gnd cell_6t
Xbit_r253_c118 bl[118] br[118] wl[253] vdd gnd cell_6t
Xbit_r254_c118 bl[118] br[118] wl[254] vdd gnd cell_6t
Xbit_r255_c118 bl[118] br[118] wl[255] vdd gnd cell_6t
Xbit_r0_c119 bl[119] br[119] wl[0] vdd gnd cell_6t
Xbit_r1_c119 bl[119] br[119] wl[1] vdd gnd cell_6t
Xbit_r2_c119 bl[119] br[119] wl[2] vdd gnd cell_6t
Xbit_r3_c119 bl[119] br[119] wl[3] vdd gnd cell_6t
Xbit_r4_c119 bl[119] br[119] wl[4] vdd gnd cell_6t
Xbit_r5_c119 bl[119] br[119] wl[5] vdd gnd cell_6t
Xbit_r6_c119 bl[119] br[119] wl[6] vdd gnd cell_6t
Xbit_r7_c119 bl[119] br[119] wl[7] vdd gnd cell_6t
Xbit_r8_c119 bl[119] br[119] wl[8] vdd gnd cell_6t
Xbit_r9_c119 bl[119] br[119] wl[9] vdd gnd cell_6t
Xbit_r10_c119 bl[119] br[119] wl[10] vdd gnd cell_6t
Xbit_r11_c119 bl[119] br[119] wl[11] vdd gnd cell_6t
Xbit_r12_c119 bl[119] br[119] wl[12] vdd gnd cell_6t
Xbit_r13_c119 bl[119] br[119] wl[13] vdd gnd cell_6t
Xbit_r14_c119 bl[119] br[119] wl[14] vdd gnd cell_6t
Xbit_r15_c119 bl[119] br[119] wl[15] vdd gnd cell_6t
Xbit_r16_c119 bl[119] br[119] wl[16] vdd gnd cell_6t
Xbit_r17_c119 bl[119] br[119] wl[17] vdd gnd cell_6t
Xbit_r18_c119 bl[119] br[119] wl[18] vdd gnd cell_6t
Xbit_r19_c119 bl[119] br[119] wl[19] vdd gnd cell_6t
Xbit_r20_c119 bl[119] br[119] wl[20] vdd gnd cell_6t
Xbit_r21_c119 bl[119] br[119] wl[21] vdd gnd cell_6t
Xbit_r22_c119 bl[119] br[119] wl[22] vdd gnd cell_6t
Xbit_r23_c119 bl[119] br[119] wl[23] vdd gnd cell_6t
Xbit_r24_c119 bl[119] br[119] wl[24] vdd gnd cell_6t
Xbit_r25_c119 bl[119] br[119] wl[25] vdd gnd cell_6t
Xbit_r26_c119 bl[119] br[119] wl[26] vdd gnd cell_6t
Xbit_r27_c119 bl[119] br[119] wl[27] vdd gnd cell_6t
Xbit_r28_c119 bl[119] br[119] wl[28] vdd gnd cell_6t
Xbit_r29_c119 bl[119] br[119] wl[29] vdd gnd cell_6t
Xbit_r30_c119 bl[119] br[119] wl[30] vdd gnd cell_6t
Xbit_r31_c119 bl[119] br[119] wl[31] vdd gnd cell_6t
Xbit_r32_c119 bl[119] br[119] wl[32] vdd gnd cell_6t
Xbit_r33_c119 bl[119] br[119] wl[33] vdd gnd cell_6t
Xbit_r34_c119 bl[119] br[119] wl[34] vdd gnd cell_6t
Xbit_r35_c119 bl[119] br[119] wl[35] vdd gnd cell_6t
Xbit_r36_c119 bl[119] br[119] wl[36] vdd gnd cell_6t
Xbit_r37_c119 bl[119] br[119] wl[37] vdd gnd cell_6t
Xbit_r38_c119 bl[119] br[119] wl[38] vdd gnd cell_6t
Xbit_r39_c119 bl[119] br[119] wl[39] vdd gnd cell_6t
Xbit_r40_c119 bl[119] br[119] wl[40] vdd gnd cell_6t
Xbit_r41_c119 bl[119] br[119] wl[41] vdd gnd cell_6t
Xbit_r42_c119 bl[119] br[119] wl[42] vdd gnd cell_6t
Xbit_r43_c119 bl[119] br[119] wl[43] vdd gnd cell_6t
Xbit_r44_c119 bl[119] br[119] wl[44] vdd gnd cell_6t
Xbit_r45_c119 bl[119] br[119] wl[45] vdd gnd cell_6t
Xbit_r46_c119 bl[119] br[119] wl[46] vdd gnd cell_6t
Xbit_r47_c119 bl[119] br[119] wl[47] vdd gnd cell_6t
Xbit_r48_c119 bl[119] br[119] wl[48] vdd gnd cell_6t
Xbit_r49_c119 bl[119] br[119] wl[49] vdd gnd cell_6t
Xbit_r50_c119 bl[119] br[119] wl[50] vdd gnd cell_6t
Xbit_r51_c119 bl[119] br[119] wl[51] vdd gnd cell_6t
Xbit_r52_c119 bl[119] br[119] wl[52] vdd gnd cell_6t
Xbit_r53_c119 bl[119] br[119] wl[53] vdd gnd cell_6t
Xbit_r54_c119 bl[119] br[119] wl[54] vdd gnd cell_6t
Xbit_r55_c119 bl[119] br[119] wl[55] vdd gnd cell_6t
Xbit_r56_c119 bl[119] br[119] wl[56] vdd gnd cell_6t
Xbit_r57_c119 bl[119] br[119] wl[57] vdd gnd cell_6t
Xbit_r58_c119 bl[119] br[119] wl[58] vdd gnd cell_6t
Xbit_r59_c119 bl[119] br[119] wl[59] vdd gnd cell_6t
Xbit_r60_c119 bl[119] br[119] wl[60] vdd gnd cell_6t
Xbit_r61_c119 bl[119] br[119] wl[61] vdd gnd cell_6t
Xbit_r62_c119 bl[119] br[119] wl[62] vdd gnd cell_6t
Xbit_r63_c119 bl[119] br[119] wl[63] vdd gnd cell_6t
Xbit_r64_c119 bl[119] br[119] wl[64] vdd gnd cell_6t
Xbit_r65_c119 bl[119] br[119] wl[65] vdd gnd cell_6t
Xbit_r66_c119 bl[119] br[119] wl[66] vdd gnd cell_6t
Xbit_r67_c119 bl[119] br[119] wl[67] vdd gnd cell_6t
Xbit_r68_c119 bl[119] br[119] wl[68] vdd gnd cell_6t
Xbit_r69_c119 bl[119] br[119] wl[69] vdd gnd cell_6t
Xbit_r70_c119 bl[119] br[119] wl[70] vdd gnd cell_6t
Xbit_r71_c119 bl[119] br[119] wl[71] vdd gnd cell_6t
Xbit_r72_c119 bl[119] br[119] wl[72] vdd gnd cell_6t
Xbit_r73_c119 bl[119] br[119] wl[73] vdd gnd cell_6t
Xbit_r74_c119 bl[119] br[119] wl[74] vdd gnd cell_6t
Xbit_r75_c119 bl[119] br[119] wl[75] vdd gnd cell_6t
Xbit_r76_c119 bl[119] br[119] wl[76] vdd gnd cell_6t
Xbit_r77_c119 bl[119] br[119] wl[77] vdd gnd cell_6t
Xbit_r78_c119 bl[119] br[119] wl[78] vdd gnd cell_6t
Xbit_r79_c119 bl[119] br[119] wl[79] vdd gnd cell_6t
Xbit_r80_c119 bl[119] br[119] wl[80] vdd gnd cell_6t
Xbit_r81_c119 bl[119] br[119] wl[81] vdd gnd cell_6t
Xbit_r82_c119 bl[119] br[119] wl[82] vdd gnd cell_6t
Xbit_r83_c119 bl[119] br[119] wl[83] vdd gnd cell_6t
Xbit_r84_c119 bl[119] br[119] wl[84] vdd gnd cell_6t
Xbit_r85_c119 bl[119] br[119] wl[85] vdd gnd cell_6t
Xbit_r86_c119 bl[119] br[119] wl[86] vdd gnd cell_6t
Xbit_r87_c119 bl[119] br[119] wl[87] vdd gnd cell_6t
Xbit_r88_c119 bl[119] br[119] wl[88] vdd gnd cell_6t
Xbit_r89_c119 bl[119] br[119] wl[89] vdd gnd cell_6t
Xbit_r90_c119 bl[119] br[119] wl[90] vdd gnd cell_6t
Xbit_r91_c119 bl[119] br[119] wl[91] vdd gnd cell_6t
Xbit_r92_c119 bl[119] br[119] wl[92] vdd gnd cell_6t
Xbit_r93_c119 bl[119] br[119] wl[93] vdd gnd cell_6t
Xbit_r94_c119 bl[119] br[119] wl[94] vdd gnd cell_6t
Xbit_r95_c119 bl[119] br[119] wl[95] vdd gnd cell_6t
Xbit_r96_c119 bl[119] br[119] wl[96] vdd gnd cell_6t
Xbit_r97_c119 bl[119] br[119] wl[97] vdd gnd cell_6t
Xbit_r98_c119 bl[119] br[119] wl[98] vdd gnd cell_6t
Xbit_r99_c119 bl[119] br[119] wl[99] vdd gnd cell_6t
Xbit_r100_c119 bl[119] br[119] wl[100] vdd gnd cell_6t
Xbit_r101_c119 bl[119] br[119] wl[101] vdd gnd cell_6t
Xbit_r102_c119 bl[119] br[119] wl[102] vdd gnd cell_6t
Xbit_r103_c119 bl[119] br[119] wl[103] vdd gnd cell_6t
Xbit_r104_c119 bl[119] br[119] wl[104] vdd gnd cell_6t
Xbit_r105_c119 bl[119] br[119] wl[105] vdd gnd cell_6t
Xbit_r106_c119 bl[119] br[119] wl[106] vdd gnd cell_6t
Xbit_r107_c119 bl[119] br[119] wl[107] vdd gnd cell_6t
Xbit_r108_c119 bl[119] br[119] wl[108] vdd gnd cell_6t
Xbit_r109_c119 bl[119] br[119] wl[109] vdd gnd cell_6t
Xbit_r110_c119 bl[119] br[119] wl[110] vdd gnd cell_6t
Xbit_r111_c119 bl[119] br[119] wl[111] vdd gnd cell_6t
Xbit_r112_c119 bl[119] br[119] wl[112] vdd gnd cell_6t
Xbit_r113_c119 bl[119] br[119] wl[113] vdd gnd cell_6t
Xbit_r114_c119 bl[119] br[119] wl[114] vdd gnd cell_6t
Xbit_r115_c119 bl[119] br[119] wl[115] vdd gnd cell_6t
Xbit_r116_c119 bl[119] br[119] wl[116] vdd gnd cell_6t
Xbit_r117_c119 bl[119] br[119] wl[117] vdd gnd cell_6t
Xbit_r118_c119 bl[119] br[119] wl[118] vdd gnd cell_6t
Xbit_r119_c119 bl[119] br[119] wl[119] vdd gnd cell_6t
Xbit_r120_c119 bl[119] br[119] wl[120] vdd gnd cell_6t
Xbit_r121_c119 bl[119] br[119] wl[121] vdd gnd cell_6t
Xbit_r122_c119 bl[119] br[119] wl[122] vdd gnd cell_6t
Xbit_r123_c119 bl[119] br[119] wl[123] vdd gnd cell_6t
Xbit_r124_c119 bl[119] br[119] wl[124] vdd gnd cell_6t
Xbit_r125_c119 bl[119] br[119] wl[125] vdd gnd cell_6t
Xbit_r126_c119 bl[119] br[119] wl[126] vdd gnd cell_6t
Xbit_r127_c119 bl[119] br[119] wl[127] vdd gnd cell_6t
Xbit_r128_c119 bl[119] br[119] wl[128] vdd gnd cell_6t
Xbit_r129_c119 bl[119] br[119] wl[129] vdd gnd cell_6t
Xbit_r130_c119 bl[119] br[119] wl[130] vdd gnd cell_6t
Xbit_r131_c119 bl[119] br[119] wl[131] vdd gnd cell_6t
Xbit_r132_c119 bl[119] br[119] wl[132] vdd gnd cell_6t
Xbit_r133_c119 bl[119] br[119] wl[133] vdd gnd cell_6t
Xbit_r134_c119 bl[119] br[119] wl[134] vdd gnd cell_6t
Xbit_r135_c119 bl[119] br[119] wl[135] vdd gnd cell_6t
Xbit_r136_c119 bl[119] br[119] wl[136] vdd gnd cell_6t
Xbit_r137_c119 bl[119] br[119] wl[137] vdd gnd cell_6t
Xbit_r138_c119 bl[119] br[119] wl[138] vdd gnd cell_6t
Xbit_r139_c119 bl[119] br[119] wl[139] vdd gnd cell_6t
Xbit_r140_c119 bl[119] br[119] wl[140] vdd gnd cell_6t
Xbit_r141_c119 bl[119] br[119] wl[141] vdd gnd cell_6t
Xbit_r142_c119 bl[119] br[119] wl[142] vdd gnd cell_6t
Xbit_r143_c119 bl[119] br[119] wl[143] vdd gnd cell_6t
Xbit_r144_c119 bl[119] br[119] wl[144] vdd gnd cell_6t
Xbit_r145_c119 bl[119] br[119] wl[145] vdd gnd cell_6t
Xbit_r146_c119 bl[119] br[119] wl[146] vdd gnd cell_6t
Xbit_r147_c119 bl[119] br[119] wl[147] vdd gnd cell_6t
Xbit_r148_c119 bl[119] br[119] wl[148] vdd gnd cell_6t
Xbit_r149_c119 bl[119] br[119] wl[149] vdd gnd cell_6t
Xbit_r150_c119 bl[119] br[119] wl[150] vdd gnd cell_6t
Xbit_r151_c119 bl[119] br[119] wl[151] vdd gnd cell_6t
Xbit_r152_c119 bl[119] br[119] wl[152] vdd gnd cell_6t
Xbit_r153_c119 bl[119] br[119] wl[153] vdd gnd cell_6t
Xbit_r154_c119 bl[119] br[119] wl[154] vdd gnd cell_6t
Xbit_r155_c119 bl[119] br[119] wl[155] vdd gnd cell_6t
Xbit_r156_c119 bl[119] br[119] wl[156] vdd gnd cell_6t
Xbit_r157_c119 bl[119] br[119] wl[157] vdd gnd cell_6t
Xbit_r158_c119 bl[119] br[119] wl[158] vdd gnd cell_6t
Xbit_r159_c119 bl[119] br[119] wl[159] vdd gnd cell_6t
Xbit_r160_c119 bl[119] br[119] wl[160] vdd gnd cell_6t
Xbit_r161_c119 bl[119] br[119] wl[161] vdd gnd cell_6t
Xbit_r162_c119 bl[119] br[119] wl[162] vdd gnd cell_6t
Xbit_r163_c119 bl[119] br[119] wl[163] vdd gnd cell_6t
Xbit_r164_c119 bl[119] br[119] wl[164] vdd gnd cell_6t
Xbit_r165_c119 bl[119] br[119] wl[165] vdd gnd cell_6t
Xbit_r166_c119 bl[119] br[119] wl[166] vdd gnd cell_6t
Xbit_r167_c119 bl[119] br[119] wl[167] vdd gnd cell_6t
Xbit_r168_c119 bl[119] br[119] wl[168] vdd gnd cell_6t
Xbit_r169_c119 bl[119] br[119] wl[169] vdd gnd cell_6t
Xbit_r170_c119 bl[119] br[119] wl[170] vdd gnd cell_6t
Xbit_r171_c119 bl[119] br[119] wl[171] vdd gnd cell_6t
Xbit_r172_c119 bl[119] br[119] wl[172] vdd gnd cell_6t
Xbit_r173_c119 bl[119] br[119] wl[173] vdd gnd cell_6t
Xbit_r174_c119 bl[119] br[119] wl[174] vdd gnd cell_6t
Xbit_r175_c119 bl[119] br[119] wl[175] vdd gnd cell_6t
Xbit_r176_c119 bl[119] br[119] wl[176] vdd gnd cell_6t
Xbit_r177_c119 bl[119] br[119] wl[177] vdd gnd cell_6t
Xbit_r178_c119 bl[119] br[119] wl[178] vdd gnd cell_6t
Xbit_r179_c119 bl[119] br[119] wl[179] vdd gnd cell_6t
Xbit_r180_c119 bl[119] br[119] wl[180] vdd gnd cell_6t
Xbit_r181_c119 bl[119] br[119] wl[181] vdd gnd cell_6t
Xbit_r182_c119 bl[119] br[119] wl[182] vdd gnd cell_6t
Xbit_r183_c119 bl[119] br[119] wl[183] vdd gnd cell_6t
Xbit_r184_c119 bl[119] br[119] wl[184] vdd gnd cell_6t
Xbit_r185_c119 bl[119] br[119] wl[185] vdd gnd cell_6t
Xbit_r186_c119 bl[119] br[119] wl[186] vdd gnd cell_6t
Xbit_r187_c119 bl[119] br[119] wl[187] vdd gnd cell_6t
Xbit_r188_c119 bl[119] br[119] wl[188] vdd gnd cell_6t
Xbit_r189_c119 bl[119] br[119] wl[189] vdd gnd cell_6t
Xbit_r190_c119 bl[119] br[119] wl[190] vdd gnd cell_6t
Xbit_r191_c119 bl[119] br[119] wl[191] vdd gnd cell_6t
Xbit_r192_c119 bl[119] br[119] wl[192] vdd gnd cell_6t
Xbit_r193_c119 bl[119] br[119] wl[193] vdd gnd cell_6t
Xbit_r194_c119 bl[119] br[119] wl[194] vdd gnd cell_6t
Xbit_r195_c119 bl[119] br[119] wl[195] vdd gnd cell_6t
Xbit_r196_c119 bl[119] br[119] wl[196] vdd gnd cell_6t
Xbit_r197_c119 bl[119] br[119] wl[197] vdd gnd cell_6t
Xbit_r198_c119 bl[119] br[119] wl[198] vdd gnd cell_6t
Xbit_r199_c119 bl[119] br[119] wl[199] vdd gnd cell_6t
Xbit_r200_c119 bl[119] br[119] wl[200] vdd gnd cell_6t
Xbit_r201_c119 bl[119] br[119] wl[201] vdd gnd cell_6t
Xbit_r202_c119 bl[119] br[119] wl[202] vdd gnd cell_6t
Xbit_r203_c119 bl[119] br[119] wl[203] vdd gnd cell_6t
Xbit_r204_c119 bl[119] br[119] wl[204] vdd gnd cell_6t
Xbit_r205_c119 bl[119] br[119] wl[205] vdd gnd cell_6t
Xbit_r206_c119 bl[119] br[119] wl[206] vdd gnd cell_6t
Xbit_r207_c119 bl[119] br[119] wl[207] vdd gnd cell_6t
Xbit_r208_c119 bl[119] br[119] wl[208] vdd gnd cell_6t
Xbit_r209_c119 bl[119] br[119] wl[209] vdd gnd cell_6t
Xbit_r210_c119 bl[119] br[119] wl[210] vdd gnd cell_6t
Xbit_r211_c119 bl[119] br[119] wl[211] vdd gnd cell_6t
Xbit_r212_c119 bl[119] br[119] wl[212] vdd gnd cell_6t
Xbit_r213_c119 bl[119] br[119] wl[213] vdd gnd cell_6t
Xbit_r214_c119 bl[119] br[119] wl[214] vdd gnd cell_6t
Xbit_r215_c119 bl[119] br[119] wl[215] vdd gnd cell_6t
Xbit_r216_c119 bl[119] br[119] wl[216] vdd gnd cell_6t
Xbit_r217_c119 bl[119] br[119] wl[217] vdd gnd cell_6t
Xbit_r218_c119 bl[119] br[119] wl[218] vdd gnd cell_6t
Xbit_r219_c119 bl[119] br[119] wl[219] vdd gnd cell_6t
Xbit_r220_c119 bl[119] br[119] wl[220] vdd gnd cell_6t
Xbit_r221_c119 bl[119] br[119] wl[221] vdd gnd cell_6t
Xbit_r222_c119 bl[119] br[119] wl[222] vdd gnd cell_6t
Xbit_r223_c119 bl[119] br[119] wl[223] vdd gnd cell_6t
Xbit_r224_c119 bl[119] br[119] wl[224] vdd gnd cell_6t
Xbit_r225_c119 bl[119] br[119] wl[225] vdd gnd cell_6t
Xbit_r226_c119 bl[119] br[119] wl[226] vdd gnd cell_6t
Xbit_r227_c119 bl[119] br[119] wl[227] vdd gnd cell_6t
Xbit_r228_c119 bl[119] br[119] wl[228] vdd gnd cell_6t
Xbit_r229_c119 bl[119] br[119] wl[229] vdd gnd cell_6t
Xbit_r230_c119 bl[119] br[119] wl[230] vdd gnd cell_6t
Xbit_r231_c119 bl[119] br[119] wl[231] vdd gnd cell_6t
Xbit_r232_c119 bl[119] br[119] wl[232] vdd gnd cell_6t
Xbit_r233_c119 bl[119] br[119] wl[233] vdd gnd cell_6t
Xbit_r234_c119 bl[119] br[119] wl[234] vdd gnd cell_6t
Xbit_r235_c119 bl[119] br[119] wl[235] vdd gnd cell_6t
Xbit_r236_c119 bl[119] br[119] wl[236] vdd gnd cell_6t
Xbit_r237_c119 bl[119] br[119] wl[237] vdd gnd cell_6t
Xbit_r238_c119 bl[119] br[119] wl[238] vdd gnd cell_6t
Xbit_r239_c119 bl[119] br[119] wl[239] vdd gnd cell_6t
Xbit_r240_c119 bl[119] br[119] wl[240] vdd gnd cell_6t
Xbit_r241_c119 bl[119] br[119] wl[241] vdd gnd cell_6t
Xbit_r242_c119 bl[119] br[119] wl[242] vdd gnd cell_6t
Xbit_r243_c119 bl[119] br[119] wl[243] vdd gnd cell_6t
Xbit_r244_c119 bl[119] br[119] wl[244] vdd gnd cell_6t
Xbit_r245_c119 bl[119] br[119] wl[245] vdd gnd cell_6t
Xbit_r246_c119 bl[119] br[119] wl[246] vdd gnd cell_6t
Xbit_r247_c119 bl[119] br[119] wl[247] vdd gnd cell_6t
Xbit_r248_c119 bl[119] br[119] wl[248] vdd gnd cell_6t
Xbit_r249_c119 bl[119] br[119] wl[249] vdd gnd cell_6t
Xbit_r250_c119 bl[119] br[119] wl[250] vdd gnd cell_6t
Xbit_r251_c119 bl[119] br[119] wl[251] vdd gnd cell_6t
Xbit_r252_c119 bl[119] br[119] wl[252] vdd gnd cell_6t
Xbit_r253_c119 bl[119] br[119] wl[253] vdd gnd cell_6t
Xbit_r254_c119 bl[119] br[119] wl[254] vdd gnd cell_6t
Xbit_r255_c119 bl[119] br[119] wl[255] vdd gnd cell_6t
Xbit_r0_c120 bl[120] br[120] wl[0] vdd gnd cell_6t
Xbit_r1_c120 bl[120] br[120] wl[1] vdd gnd cell_6t
Xbit_r2_c120 bl[120] br[120] wl[2] vdd gnd cell_6t
Xbit_r3_c120 bl[120] br[120] wl[3] vdd gnd cell_6t
Xbit_r4_c120 bl[120] br[120] wl[4] vdd gnd cell_6t
Xbit_r5_c120 bl[120] br[120] wl[5] vdd gnd cell_6t
Xbit_r6_c120 bl[120] br[120] wl[6] vdd gnd cell_6t
Xbit_r7_c120 bl[120] br[120] wl[7] vdd gnd cell_6t
Xbit_r8_c120 bl[120] br[120] wl[8] vdd gnd cell_6t
Xbit_r9_c120 bl[120] br[120] wl[9] vdd gnd cell_6t
Xbit_r10_c120 bl[120] br[120] wl[10] vdd gnd cell_6t
Xbit_r11_c120 bl[120] br[120] wl[11] vdd gnd cell_6t
Xbit_r12_c120 bl[120] br[120] wl[12] vdd gnd cell_6t
Xbit_r13_c120 bl[120] br[120] wl[13] vdd gnd cell_6t
Xbit_r14_c120 bl[120] br[120] wl[14] vdd gnd cell_6t
Xbit_r15_c120 bl[120] br[120] wl[15] vdd gnd cell_6t
Xbit_r16_c120 bl[120] br[120] wl[16] vdd gnd cell_6t
Xbit_r17_c120 bl[120] br[120] wl[17] vdd gnd cell_6t
Xbit_r18_c120 bl[120] br[120] wl[18] vdd gnd cell_6t
Xbit_r19_c120 bl[120] br[120] wl[19] vdd gnd cell_6t
Xbit_r20_c120 bl[120] br[120] wl[20] vdd gnd cell_6t
Xbit_r21_c120 bl[120] br[120] wl[21] vdd gnd cell_6t
Xbit_r22_c120 bl[120] br[120] wl[22] vdd gnd cell_6t
Xbit_r23_c120 bl[120] br[120] wl[23] vdd gnd cell_6t
Xbit_r24_c120 bl[120] br[120] wl[24] vdd gnd cell_6t
Xbit_r25_c120 bl[120] br[120] wl[25] vdd gnd cell_6t
Xbit_r26_c120 bl[120] br[120] wl[26] vdd gnd cell_6t
Xbit_r27_c120 bl[120] br[120] wl[27] vdd gnd cell_6t
Xbit_r28_c120 bl[120] br[120] wl[28] vdd gnd cell_6t
Xbit_r29_c120 bl[120] br[120] wl[29] vdd gnd cell_6t
Xbit_r30_c120 bl[120] br[120] wl[30] vdd gnd cell_6t
Xbit_r31_c120 bl[120] br[120] wl[31] vdd gnd cell_6t
Xbit_r32_c120 bl[120] br[120] wl[32] vdd gnd cell_6t
Xbit_r33_c120 bl[120] br[120] wl[33] vdd gnd cell_6t
Xbit_r34_c120 bl[120] br[120] wl[34] vdd gnd cell_6t
Xbit_r35_c120 bl[120] br[120] wl[35] vdd gnd cell_6t
Xbit_r36_c120 bl[120] br[120] wl[36] vdd gnd cell_6t
Xbit_r37_c120 bl[120] br[120] wl[37] vdd gnd cell_6t
Xbit_r38_c120 bl[120] br[120] wl[38] vdd gnd cell_6t
Xbit_r39_c120 bl[120] br[120] wl[39] vdd gnd cell_6t
Xbit_r40_c120 bl[120] br[120] wl[40] vdd gnd cell_6t
Xbit_r41_c120 bl[120] br[120] wl[41] vdd gnd cell_6t
Xbit_r42_c120 bl[120] br[120] wl[42] vdd gnd cell_6t
Xbit_r43_c120 bl[120] br[120] wl[43] vdd gnd cell_6t
Xbit_r44_c120 bl[120] br[120] wl[44] vdd gnd cell_6t
Xbit_r45_c120 bl[120] br[120] wl[45] vdd gnd cell_6t
Xbit_r46_c120 bl[120] br[120] wl[46] vdd gnd cell_6t
Xbit_r47_c120 bl[120] br[120] wl[47] vdd gnd cell_6t
Xbit_r48_c120 bl[120] br[120] wl[48] vdd gnd cell_6t
Xbit_r49_c120 bl[120] br[120] wl[49] vdd gnd cell_6t
Xbit_r50_c120 bl[120] br[120] wl[50] vdd gnd cell_6t
Xbit_r51_c120 bl[120] br[120] wl[51] vdd gnd cell_6t
Xbit_r52_c120 bl[120] br[120] wl[52] vdd gnd cell_6t
Xbit_r53_c120 bl[120] br[120] wl[53] vdd gnd cell_6t
Xbit_r54_c120 bl[120] br[120] wl[54] vdd gnd cell_6t
Xbit_r55_c120 bl[120] br[120] wl[55] vdd gnd cell_6t
Xbit_r56_c120 bl[120] br[120] wl[56] vdd gnd cell_6t
Xbit_r57_c120 bl[120] br[120] wl[57] vdd gnd cell_6t
Xbit_r58_c120 bl[120] br[120] wl[58] vdd gnd cell_6t
Xbit_r59_c120 bl[120] br[120] wl[59] vdd gnd cell_6t
Xbit_r60_c120 bl[120] br[120] wl[60] vdd gnd cell_6t
Xbit_r61_c120 bl[120] br[120] wl[61] vdd gnd cell_6t
Xbit_r62_c120 bl[120] br[120] wl[62] vdd gnd cell_6t
Xbit_r63_c120 bl[120] br[120] wl[63] vdd gnd cell_6t
Xbit_r64_c120 bl[120] br[120] wl[64] vdd gnd cell_6t
Xbit_r65_c120 bl[120] br[120] wl[65] vdd gnd cell_6t
Xbit_r66_c120 bl[120] br[120] wl[66] vdd gnd cell_6t
Xbit_r67_c120 bl[120] br[120] wl[67] vdd gnd cell_6t
Xbit_r68_c120 bl[120] br[120] wl[68] vdd gnd cell_6t
Xbit_r69_c120 bl[120] br[120] wl[69] vdd gnd cell_6t
Xbit_r70_c120 bl[120] br[120] wl[70] vdd gnd cell_6t
Xbit_r71_c120 bl[120] br[120] wl[71] vdd gnd cell_6t
Xbit_r72_c120 bl[120] br[120] wl[72] vdd gnd cell_6t
Xbit_r73_c120 bl[120] br[120] wl[73] vdd gnd cell_6t
Xbit_r74_c120 bl[120] br[120] wl[74] vdd gnd cell_6t
Xbit_r75_c120 bl[120] br[120] wl[75] vdd gnd cell_6t
Xbit_r76_c120 bl[120] br[120] wl[76] vdd gnd cell_6t
Xbit_r77_c120 bl[120] br[120] wl[77] vdd gnd cell_6t
Xbit_r78_c120 bl[120] br[120] wl[78] vdd gnd cell_6t
Xbit_r79_c120 bl[120] br[120] wl[79] vdd gnd cell_6t
Xbit_r80_c120 bl[120] br[120] wl[80] vdd gnd cell_6t
Xbit_r81_c120 bl[120] br[120] wl[81] vdd gnd cell_6t
Xbit_r82_c120 bl[120] br[120] wl[82] vdd gnd cell_6t
Xbit_r83_c120 bl[120] br[120] wl[83] vdd gnd cell_6t
Xbit_r84_c120 bl[120] br[120] wl[84] vdd gnd cell_6t
Xbit_r85_c120 bl[120] br[120] wl[85] vdd gnd cell_6t
Xbit_r86_c120 bl[120] br[120] wl[86] vdd gnd cell_6t
Xbit_r87_c120 bl[120] br[120] wl[87] vdd gnd cell_6t
Xbit_r88_c120 bl[120] br[120] wl[88] vdd gnd cell_6t
Xbit_r89_c120 bl[120] br[120] wl[89] vdd gnd cell_6t
Xbit_r90_c120 bl[120] br[120] wl[90] vdd gnd cell_6t
Xbit_r91_c120 bl[120] br[120] wl[91] vdd gnd cell_6t
Xbit_r92_c120 bl[120] br[120] wl[92] vdd gnd cell_6t
Xbit_r93_c120 bl[120] br[120] wl[93] vdd gnd cell_6t
Xbit_r94_c120 bl[120] br[120] wl[94] vdd gnd cell_6t
Xbit_r95_c120 bl[120] br[120] wl[95] vdd gnd cell_6t
Xbit_r96_c120 bl[120] br[120] wl[96] vdd gnd cell_6t
Xbit_r97_c120 bl[120] br[120] wl[97] vdd gnd cell_6t
Xbit_r98_c120 bl[120] br[120] wl[98] vdd gnd cell_6t
Xbit_r99_c120 bl[120] br[120] wl[99] vdd gnd cell_6t
Xbit_r100_c120 bl[120] br[120] wl[100] vdd gnd cell_6t
Xbit_r101_c120 bl[120] br[120] wl[101] vdd gnd cell_6t
Xbit_r102_c120 bl[120] br[120] wl[102] vdd gnd cell_6t
Xbit_r103_c120 bl[120] br[120] wl[103] vdd gnd cell_6t
Xbit_r104_c120 bl[120] br[120] wl[104] vdd gnd cell_6t
Xbit_r105_c120 bl[120] br[120] wl[105] vdd gnd cell_6t
Xbit_r106_c120 bl[120] br[120] wl[106] vdd gnd cell_6t
Xbit_r107_c120 bl[120] br[120] wl[107] vdd gnd cell_6t
Xbit_r108_c120 bl[120] br[120] wl[108] vdd gnd cell_6t
Xbit_r109_c120 bl[120] br[120] wl[109] vdd gnd cell_6t
Xbit_r110_c120 bl[120] br[120] wl[110] vdd gnd cell_6t
Xbit_r111_c120 bl[120] br[120] wl[111] vdd gnd cell_6t
Xbit_r112_c120 bl[120] br[120] wl[112] vdd gnd cell_6t
Xbit_r113_c120 bl[120] br[120] wl[113] vdd gnd cell_6t
Xbit_r114_c120 bl[120] br[120] wl[114] vdd gnd cell_6t
Xbit_r115_c120 bl[120] br[120] wl[115] vdd gnd cell_6t
Xbit_r116_c120 bl[120] br[120] wl[116] vdd gnd cell_6t
Xbit_r117_c120 bl[120] br[120] wl[117] vdd gnd cell_6t
Xbit_r118_c120 bl[120] br[120] wl[118] vdd gnd cell_6t
Xbit_r119_c120 bl[120] br[120] wl[119] vdd gnd cell_6t
Xbit_r120_c120 bl[120] br[120] wl[120] vdd gnd cell_6t
Xbit_r121_c120 bl[120] br[120] wl[121] vdd gnd cell_6t
Xbit_r122_c120 bl[120] br[120] wl[122] vdd gnd cell_6t
Xbit_r123_c120 bl[120] br[120] wl[123] vdd gnd cell_6t
Xbit_r124_c120 bl[120] br[120] wl[124] vdd gnd cell_6t
Xbit_r125_c120 bl[120] br[120] wl[125] vdd gnd cell_6t
Xbit_r126_c120 bl[120] br[120] wl[126] vdd gnd cell_6t
Xbit_r127_c120 bl[120] br[120] wl[127] vdd gnd cell_6t
Xbit_r128_c120 bl[120] br[120] wl[128] vdd gnd cell_6t
Xbit_r129_c120 bl[120] br[120] wl[129] vdd gnd cell_6t
Xbit_r130_c120 bl[120] br[120] wl[130] vdd gnd cell_6t
Xbit_r131_c120 bl[120] br[120] wl[131] vdd gnd cell_6t
Xbit_r132_c120 bl[120] br[120] wl[132] vdd gnd cell_6t
Xbit_r133_c120 bl[120] br[120] wl[133] vdd gnd cell_6t
Xbit_r134_c120 bl[120] br[120] wl[134] vdd gnd cell_6t
Xbit_r135_c120 bl[120] br[120] wl[135] vdd gnd cell_6t
Xbit_r136_c120 bl[120] br[120] wl[136] vdd gnd cell_6t
Xbit_r137_c120 bl[120] br[120] wl[137] vdd gnd cell_6t
Xbit_r138_c120 bl[120] br[120] wl[138] vdd gnd cell_6t
Xbit_r139_c120 bl[120] br[120] wl[139] vdd gnd cell_6t
Xbit_r140_c120 bl[120] br[120] wl[140] vdd gnd cell_6t
Xbit_r141_c120 bl[120] br[120] wl[141] vdd gnd cell_6t
Xbit_r142_c120 bl[120] br[120] wl[142] vdd gnd cell_6t
Xbit_r143_c120 bl[120] br[120] wl[143] vdd gnd cell_6t
Xbit_r144_c120 bl[120] br[120] wl[144] vdd gnd cell_6t
Xbit_r145_c120 bl[120] br[120] wl[145] vdd gnd cell_6t
Xbit_r146_c120 bl[120] br[120] wl[146] vdd gnd cell_6t
Xbit_r147_c120 bl[120] br[120] wl[147] vdd gnd cell_6t
Xbit_r148_c120 bl[120] br[120] wl[148] vdd gnd cell_6t
Xbit_r149_c120 bl[120] br[120] wl[149] vdd gnd cell_6t
Xbit_r150_c120 bl[120] br[120] wl[150] vdd gnd cell_6t
Xbit_r151_c120 bl[120] br[120] wl[151] vdd gnd cell_6t
Xbit_r152_c120 bl[120] br[120] wl[152] vdd gnd cell_6t
Xbit_r153_c120 bl[120] br[120] wl[153] vdd gnd cell_6t
Xbit_r154_c120 bl[120] br[120] wl[154] vdd gnd cell_6t
Xbit_r155_c120 bl[120] br[120] wl[155] vdd gnd cell_6t
Xbit_r156_c120 bl[120] br[120] wl[156] vdd gnd cell_6t
Xbit_r157_c120 bl[120] br[120] wl[157] vdd gnd cell_6t
Xbit_r158_c120 bl[120] br[120] wl[158] vdd gnd cell_6t
Xbit_r159_c120 bl[120] br[120] wl[159] vdd gnd cell_6t
Xbit_r160_c120 bl[120] br[120] wl[160] vdd gnd cell_6t
Xbit_r161_c120 bl[120] br[120] wl[161] vdd gnd cell_6t
Xbit_r162_c120 bl[120] br[120] wl[162] vdd gnd cell_6t
Xbit_r163_c120 bl[120] br[120] wl[163] vdd gnd cell_6t
Xbit_r164_c120 bl[120] br[120] wl[164] vdd gnd cell_6t
Xbit_r165_c120 bl[120] br[120] wl[165] vdd gnd cell_6t
Xbit_r166_c120 bl[120] br[120] wl[166] vdd gnd cell_6t
Xbit_r167_c120 bl[120] br[120] wl[167] vdd gnd cell_6t
Xbit_r168_c120 bl[120] br[120] wl[168] vdd gnd cell_6t
Xbit_r169_c120 bl[120] br[120] wl[169] vdd gnd cell_6t
Xbit_r170_c120 bl[120] br[120] wl[170] vdd gnd cell_6t
Xbit_r171_c120 bl[120] br[120] wl[171] vdd gnd cell_6t
Xbit_r172_c120 bl[120] br[120] wl[172] vdd gnd cell_6t
Xbit_r173_c120 bl[120] br[120] wl[173] vdd gnd cell_6t
Xbit_r174_c120 bl[120] br[120] wl[174] vdd gnd cell_6t
Xbit_r175_c120 bl[120] br[120] wl[175] vdd gnd cell_6t
Xbit_r176_c120 bl[120] br[120] wl[176] vdd gnd cell_6t
Xbit_r177_c120 bl[120] br[120] wl[177] vdd gnd cell_6t
Xbit_r178_c120 bl[120] br[120] wl[178] vdd gnd cell_6t
Xbit_r179_c120 bl[120] br[120] wl[179] vdd gnd cell_6t
Xbit_r180_c120 bl[120] br[120] wl[180] vdd gnd cell_6t
Xbit_r181_c120 bl[120] br[120] wl[181] vdd gnd cell_6t
Xbit_r182_c120 bl[120] br[120] wl[182] vdd gnd cell_6t
Xbit_r183_c120 bl[120] br[120] wl[183] vdd gnd cell_6t
Xbit_r184_c120 bl[120] br[120] wl[184] vdd gnd cell_6t
Xbit_r185_c120 bl[120] br[120] wl[185] vdd gnd cell_6t
Xbit_r186_c120 bl[120] br[120] wl[186] vdd gnd cell_6t
Xbit_r187_c120 bl[120] br[120] wl[187] vdd gnd cell_6t
Xbit_r188_c120 bl[120] br[120] wl[188] vdd gnd cell_6t
Xbit_r189_c120 bl[120] br[120] wl[189] vdd gnd cell_6t
Xbit_r190_c120 bl[120] br[120] wl[190] vdd gnd cell_6t
Xbit_r191_c120 bl[120] br[120] wl[191] vdd gnd cell_6t
Xbit_r192_c120 bl[120] br[120] wl[192] vdd gnd cell_6t
Xbit_r193_c120 bl[120] br[120] wl[193] vdd gnd cell_6t
Xbit_r194_c120 bl[120] br[120] wl[194] vdd gnd cell_6t
Xbit_r195_c120 bl[120] br[120] wl[195] vdd gnd cell_6t
Xbit_r196_c120 bl[120] br[120] wl[196] vdd gnd cell_6t
Xbit_r197_c120 bl[120] br[120] wl[197] vdd gnd cell_6t
Xbit_r198_c120 bl[120] br[120] wl[198] vdd gnd cell_6t
Xbit_r199_c120 bl[120] br[120] wl[199] vdd gnd cell_6t
Xbit_r200_c120 bl[120] br[120] wl[200] vdd gnd cell_6t
Xbit_r201_c120 bl[120] br[120] wl[201] vdd gnd cell_6t
Xbit_r202_c120 bl[120] br[120] wl[202] vdd gnd cell_6t
Xbit_r203_c120 bl[120] br[120] wl[203] vdd gnd cell_6t
Xbit_r204_c120 bl[120] br[120] wl[204] vdd gnd cell_6t
Xbit_r205_c120 bl[120] br[120] wl[205] vdd gnd cell_6t
Xbit_r206_c120 bl[120] br[120] wl[206] vdd gnd cell_6t
Xbit_r207_c120 bl[120] br[120] wl[207] vdd gnd cell_6t
Xbit_r208_c120 bl[120] br[120] wl[208] vdd gnd cell_6t
Xbit_r209_c120 bl[120] br[120] wl[209] vdd gnd cell_6t
Xbit_r210_c120 bl[120] br[120] wl[210] vdd gnd cell_6t
Xbit_r211_c120 bl[120] br[120] wl[211] vdd gnd cell_6t
Xbit_r212_c120 bl[120] br[120] wl[212] vdd gnd cell_6t
Xbit_r213_c120 bl[120] br[120] wl[213] vdd gnd cell_6t
Xbit_r214_c120 bl[120] br[120] wl[214] vdd gnd cell_6t
Xbit_r215_c120 bl[120] br[120] wl[215] vdd gnd cell_6t
Xbit_r216_c120 bl[120] br[120] wl[216] vdd gnd cell_6t
Xbit_r217_c120 bl[120] br[120] wl[217] vdd gnd cell_6t
Xbit_r218_c120 bl[120] br[120] wl[218] vdd gnd cell_6t
Xbit_r219_c120 bl[120] br[120] wl[219] vdd gnd cell_6t
Xbit_r220_c120 bl[120] br[120] wl[220] vdd gnd cell_6t
Xbit_r221_c120 bl[120] br[120] wl[221] vdd gnd cell_6t
Xbit_r222_c120 bl[120] br[120] wl[222] vdd gnd cell_6t
Xbit_r223_c120 bl[120] br[120] wl[223] vdd gnd cell_6t
Xbit_r224_c120 bl[120] br[120] wl[224] vdd gnd cell_6t
Xbit_r225_c120 bl[120] br[120] wl[225] vdd gnd cell_6t
Xbit_r226_c120 bl[120] br[120] wl[226] vdd gnd cell_6t
Xbit_r227_c120 bl[120] br[120] wl[227] vdd gnd cell_6t
Xbit_r228_c120 bl[120] br[120] wl[228] vdd gnd cell_6t
Xbit_r229_c120 bl[120] br[120] wl[229] vdd gnd cell_6t
Xbit_r230_c120 bl[120] br[120] wl[230] vdd gnd cell_6t
Xbit_r231_c120 bl[120] br[120] wl[231] vdd gnd cell_6t
Xbit_r232_c120 bl[120] br[120] wl[232] vdd gnd cell_6t
Xbit_r233_c120 bl[120] br[120] wl[233] vdd gnd cell_6t
Xbit_r234_c120 bl[120] br[120] wl[234] vdd gnd cell_6t
Xbit_r235_c120 bl[120] br[120] wl[235] vdd gnd cell_6t
Xbit_r236_c120 bl[120] br[120] wl[236] vdd gnd cell_6t
Xbit_r237_c120 bl[120] br[120] wl[237] vdd gnd cell_6t
Xbit_r238_c120 bl[120] br[120] wl[238] vdd gnd cell_6t
Xbit_r239_c120 bl[120] br[120] wl[239] vdd gnd cell_6t
Xbit_r240_c120 bl[120] br[120] wl[240] vdd gnd cell_6t
Xbit_r241_c120 bl[120] br[120] wl[241] vdd gnd cell_6t
Xbit_r242_c120 bl[120] br[120] wl[242] vdd gnd cell_6t
Xbit_r243_c120 bl[120] br[120] wl[243] vdd gnd cell_6t
Xbit_r244_c120 bl[120] br[120] wl[244] vdd gnd cell_6t
Xbit_r245_c120 bl[120] br[120] wl[245] vdd gnd cell_6t
Xbit_r246_c120 bl[120] br[120] wl[246] vdd gnd cell_6t
Xbit_r247_c120 bl[120] br[120] wl[247] vdd gnd cell_6t
Xbit_r248_c120 bl[120] br[120] wl[248] vdd gnd cell_6t
Xbit_r249_c120 bl[120] br[120] wl[249] vdd gnd cell_6t
Xbit_r250_c120 bl[120] br[120] wl[250] vdd gnd cell_6t
Xbit_r251_c120 bl[120] br[120] wl[251] vdd gnd cell_6t
Xbit_r252_c120 bl[120] br[120] wl[252] vdd gnd cell_6t
Xbit_r253_c120 bl[120] br[120] wl[253] vdd gnd cell_6t
Xbit_r254_c120 bl[120] br[120] wl[254] vdd gnd cell_6t
Xbit_r255_c120 bl[120] br[120] wl[255] vdd gnd cell_6t
Xbit_r0_c121 bl[121] br[121] wl[0] vdd gnd cell_6t
Xbit_r1_c121 bl[121] br[121] wl[1] vdd gnd cell_6t
Xbit_r2_c121 bl[121] br[121] wl[2] vdd gnd cell_6t
Xbit_r3_c121 bl[121] br[121] wl[3] vdd gnd cell_6t
Xbit_r4_c121 bl[121] br[121] wl[4] vdd gnd cell_6t
Xbit_r5_c121 bl[121] br[121] wl[5] vdd gnd cell_6t
Xbit_r6_c121 bl[121] br[121] wl[6] vdd gnd cell_6t
Xbit_r7_c121 bl[121] br[121] wl[7] vdd gnd cell_6t
Xbit_r8_c121 bl[121] br[121] wl[8] vdd gnd cell_6t
Xbit_r9_c121 bl[121] br[121] wl[9] vdd gnd cell_6t
Xbit_r10_c121 bl[121] br[121] wl[10] vdd gnd cell_6t
Xbit_r11_c121 bl[121] br[121] wl[11] vdd gnd cell_6t
Xbit_r12_c121 bl[121] br[121] wl[12] vdd gnd cell_6t
Xbit_r13_c121 bl[121] br[121] wl[13] vdd gnd cell_6t
Xbit_r14_c121 bl[121] br[121] wl[14] vdd gnd cell_6t
Xbit_r15_c121 bl[121] br[121] wl[15] vdd gnd cell_6t
Xbit_r16_c121 bl[121] br[121] wl[16] vdd gnd cell_6t
Xbit_r17_c121 bl[121] br[121] wl[17] vdd gnd cell_6t
Xbit_r18_c121 bl[121] br[121] wl[18] vdd gnd cell_6t
Xbit_r19_c121 bl[121] br[121] wl[19] vdd gnd cell_6t
Xbit_r20_c121 bl[121] br[121] wl[20] vdd gnd cell_6t
Xbit_r21_c121 bl[121] br[121] wl[21] vdd gnd cell_6t
Xbit_r22_c121 bl[121] br[121] wl[22] vdd gnd cell_6t
Xbit_r23_c121 bl[121] br[121] wl[23] vdd gnd cell_6t
Xbit_r24_c121 bl[121] br[121] wl[24] vdd gnd cell_6t
Xbit_r25_c121 bl[121] br[121] wl[25] vdd gnd cell_6t
Xbit_r26_c121 bl[121] br[121] wl[26] vdd gnd cell_6t
Xbit_r27_c121 bl[121] br[121] wl[27] vdd gnd cell_6t
Xbit_r28_c121 bl[121] br[121] wl[28] vdd gnd cell_6t
Xbit_r29_c121 bl[121] br[121] wl[29] vdd gnd cell_6t
Xbit_r30_c121 bl[121] br[121] wl[30] vdd gnd cell_6t
Xbit_r31_c121 bl[121] br[121] wl[31] vdd gnd cell_6t
Xbit_r32_c121 bl[121] br[121] wl[32] vdd gnd cell_6t
Xbit_r33_c121 bl[121] br[121] wl[33] vdd gnd cell_6t
Xbit_r34_c121 bl[121] br[121] wl[34] vdd gnd cell_6t
Xbit_r35_c121 bl[121] br[121] wl[35] vdd gnd cell_6t
Xbit_r36_c121 bl[121] br[121] wl[36] vdd gnd cell_6t
Xbit_r37_c121 bl[121] br[121] wl[37] vdd gnd cell_6t
Xbit_r38_c121 bl[121] br[121] wl[38] vdd gnd cell_6t
Xbit_r39_c121 bl[121] br[121] wl[39] vdd gnd cell_6t
Xbit_r40_c121 bl[121] br[121] wl[40] vdd gnd cell_6t
Xbit_r41_c121 bl[121] br[121] wl[41] vdd gnd cell_6t
Xbit_r42_c121 bl[121] br[121] wl[42] vdd gnd cell_6t
Xbit_r43_c121 bl[121] br[121] wl[43] vdd gnd cell_6t
Xbit_r44_c121 bl[121] br[121] wl[44] vdd gnd cell_6t
Xbit_r45_c121 bl[121] br[121] wl[45] vdd gnd cell_6t
Xbit_r46_c121 bl[121] br[121] wl[46] vdd gnd cell_6t
Xbit_r47_c121 bl[121] br[121] wl[47] vdd gnd cell_6t
Xbit_r48_c121 bl[121] br[121] wl[48] vdd gnd cell_6t
Xbit_r49_c121 bl[121] br[121] wl[49] vdd gnd cell_6t
Xbit_r50_c121 bl[121] br[121] wl[50] vdd gnd cell_6t
Xbit_r51_c121 bl[121] br[121] wl[51] vdd gnd cell_6t
Xbit_r52_c121 bl[121] br[121] wl[52] vdd gnd cell_6t
Xbit_r53_c121 bl[121] br[121] wl[53] vdd gnd cell_6t
Xbit_r54_c121 bl[121] br[121] wl[54] vdd gnd cell_6t
Xbit_r55_c121 bl[121] br[121] wl[55] vdd gnd cell_6t
Xbit_r56_c121 bl[121] br[121] wl[56] vdd gnd cell_6t
Xbit_r57_c121 bl[121] br[121] wl[57] vdd gnd cell_6t
Xbit_r58_c121 bl[121] br[121] wl[58] vdd gnd cell_6t
Xbit_r59_c121 bl[121] br[121] wl[59] vdd gnd cell_6t
Xbit_r60_c121 bl[121] br[121] wl[60] vdd gnd cell_6t
Xbit_r61_c121 bl[121] br[121] wl[61] vdd gnd cell_6t
Xbit_r62_c121 bl[121] br[121] wl[62] vdd gnd cell_6t
Xbit_r63_c121 bl[121] br[121] wl[63] vdd gnd cell_6t
Xbit_r64_c121 bl[121] br[121] wl[64] vdd gnd cell_6t
Xbit_r65_c121 bl[121] br[121] wl[65] vdd gnd cell_6t
Xbit_r66_c121 bl[121] br[121] wl[66] vdd gnd cell_6t
Xbit_r67_c121 bl[121] br[121] wl[67] vdd gnd cell_6t
Xbit_r68_c121 bl[121] br[121] wl[68] vdd gnd cell_6t
Xbit_r69_c121 bl[121] br[121] wl[69] vdd gnd cell_6t
Xbit_r70_c121 bl[121] br[121] wl[70] vdd gnd cell_6t
Xbit_r71_c121 bl[121] br[121] wl[71] vdd gnd cell_6t
Xbit_r72_c121 bl[121] br[121] wl[72] vdd gnd cell_6t
Xbit_r73_c121 bl[121] br[121] wl[73] vdd gnd cell_6t
Xbit_r74_c121 bl[121] br[121] wl[74] vdd gnd cell_6t
Xbit_r75_c121 bl[121] br[121] wl[75] vdd gnd cell_6t
Xbit_r76_c121 bl[121] br[121] wl[76] vdd gnd cell_6t
Xbit_r77_c121 bl[121] br[121] wl[77] vdd gnd cell_6t
Xbit_r78_c121 bl[121] br[121] wl[78] vdd gnd cell_6t
Xbit_r79_c121 bl[121] br[121] wl[79] vdd gnd cell_6t
Xbit_r80_c121 bl[121] br[121] wl[80] vdd gnd cell_6t
Xbit_r81_c121 bl[121] br[121] wl[81] vdd gnd cell_6t
Xbit_r82_c121 bl[121] br[121] wl[82] vdd gnd cell_6t
Xbit_r83_c121 bl[121] br[121] wl[83] vdd gnd cell_6t
Xbit_r84_c121 bl[121] br[121] wl[84] vdd gnd cell_6t
Xbit_r85_c121 bl[121] br[121] wl[85] vdd gnd cell_6t
Xbit_r86_c121 bl[121] br[121] wl[86] vdd gnd cell_6t
Xbit_r87_c121 bl[121] br[121] wl[87] vdd gnd cell_6t
Xbit_r88_c121 bl[121] br[121] wl[88] vdd gnd cell_6t
Xbit_r89_c121 bl[121] br[121] wl[89] vdd gnd cell_6t
Xbit_r90_c121 bl[121] br[121] wl[90] vdd gnd cell_6t
Xbit_r91_c121 bl[121] br[121] wl[91] vdd gnd cell_6t
Xbit_r92_c121 bl[121] br[121] wl[92] vdd gnd cell_6t
Xbit_r93_c121 bl[121] br[121] wl[93] vdd gnd cell_6t
Xbit_r94_c121 bl[121] br[121] wl[94] vdd gnd cell_6t
Xbit_r95_c121 bl[121] br[121] wl[95] vdd gnd cell_6t
Xbit_r96_c121 bl[121] br[121] wl[96] vdd gnd cell_6t
Xbit_r97_c121 bl[121] br[121] wl[97] vdd gnd cell_6t
Xbit_r98_c121 bl[121] br[121] wl[98] vdd gnd cell_6t
Xbit_r99_c121 bl[121] br[121] wl[99] vdd gnd cell_6t
Xbit_r100_c121 bl[121] br[121] wl[100] vdd gnd cell_6t
Xbit_r101_c121 bl[121] br[121] wl[101] vdd gnd cell_6t
Xbit_r102_c121 bl[121] br[121] wl[102] vdd gnd cell_6t
Xbit_r103_c121 bl[121] br[121] wl[103] vdd gnd cell_6t
Xbit_r104_c121 bl[121] br[121] wl[104] vdd gnd cell_6t
Xbit_r105_c121 bl[121] br[121] wl[105] vdd gnd cell_6t
Xbit_r106_c121 bl[121] br[121] wl[106] vdd gnd cell_6t
Xbit_r107_c121 bl[121] br[121] wl[107] vdd gnd cell_6t
Xbit_r108_c121 bl[121] br[121] wl[108] vdd gnd cell_6t
Xbit_r109_c121 bl[121] br[121] wl[109] vdd gnd cell_6t
Xbit_r110_c121 bl[121] br[121] wl[110] vdd gnd cell_6t
Xbit_r111_c121 bl[121] br[121] wl[111] vdd gnd cell_6t
Xbit_r112_c121 bl[121] br[121] wl[112] vdd gnd cell_6t
Xbit_r113_c121 bl[121] br[121] wl[113] vdd gnd cell_6t
Xbit_r114_c121 bl[121] br[121] wl[114] vdd gnd cell_6t
Xbit_r115_c121 bl[121] br[121] wl[115] vdd gnd cell_6t
Xbit_r116_c121 bl[121] br[121] wl[116] vdd gnd cell_6t
Xbit_r117_c121 bl[121] br[121] wl[117] vdd gnd cell_6t
Xbit_r118_c121 bl[121] br[121] wl[118] vdd gnd cell_6t
Xbit_r119_c121 bl[121] br[121] wl[119] vdd gnd cell_6t
Xbit_r120_c121 bl[121] br[121] wl[120] vdd gnd cell_6t
Xbit_r121_c121 bl[121] br[121] wl[121] vdd gnd cell_6t
Xbit_r122_c121 bl[121] br[121] wl[122] vdd gnd cell_6t
Xbit_r123_c121 bl[121] br[121] wl[123] vdd gnd cell_6t
Xbit_r124_c121 bl[121] br[121] wl[124] vdd gnd cell_6t
Xbit_r125_c121 bl[121] br[121] wl[125] vdd gnd cell_6t
Xbit_r126_c121 bl[121] br[121] wl[126] vdd gnd cell_6t
Xbit_r127_c121 bl[121] br[121] wl[127] vdd gnd cell_6t
Xbit_r128_c121 bl[121] br[121] wl[128] vdd gnd cell_6t
Xbit_r129_c121 bl[121] br[121] wl[129] vdd gnd cell_6t
Xbit_r130_c121 bl[121] br[121] wl[130] vdd gnd cell_6t
Xbit_r131_c121 bl[121] br[121] wl[131] vdd gnd cell_6t
Xbit_r132_c121 bl[121] br[121] wl[132] vdd gnd cell_6t
Xbit_r133_c121 bl[121] br[121] wl[133] vdd gnd cell_6t
Xbit_r134_c121 bl[121] br[121] wl[134] vdd gnd cell_6t
Xbit_r135_c121 bl[121] br[121] wl[135] vdd gnd cell_6t
Xbit_r136_c121 bl[121] br[121] wl[136] vdd gnd cell_6t
Xbit_r137_c121 bl[121] br[121] wl[137] vdd gnd cell_6t
Xbit_r138_c121 bl[121] br[121] wl[138] vdd gnd cell_6t
Xbit_r139_c121 bl[121] br[121] wl[139] vdd gnd cell_6t
Xbit_r140_c121 bl[121] br[121] wl[140] vdd gnd cell_6t
Xbit_r141_c121 bl[121] br[121] wl[141] vdd gnd cell_6t
Xbit_r142_c121 bl[121] br[121] wl[142] vdd gnd cell_6t
Xbit_r143_c121 bl[121] br[121] wl[143] vdd gnd cell_6t
Xbit_r144_c121 bl[121] br[121] wl[144] vdd gnd cell_6t
Xbit_r145_c121 bl[121] br[121] wl[145] vdd gnd cell_6t
Xbit_r146_c121 bl[121] br[121] wl[146] vdd gnd cell_6t
Xbit_r147_c121 bl[121] br[121] wl[147] vdd gnd cell_6t
Xbit_r148_c121 bl[121] br[121] wl[148] vdd gnd cell_6t
Xbit_r149_c121 bl[121] br[121] wl[149] vdd gnd cell_6t
Xbit_r150_c121 bl[121] br[121] wl[150] vdd gnd cell_6t
Xbit_r151_c121 bl[121] br[121] wl[151] vdd gnd cell_6t
Xbit_r152_c121 bl[121] br[121] wl[152] vdd gnd cell_6t
Xbit_r153_c121 bl[121] br[121] wl[153] vdd gnd cell_6t
Xbit_r154_c121 bl[121] br[121] wl[154] vdd gnd cell_6t
Xbit_r155_c121 bl[121] br[121] wl[155] vdd gnd cell_6t
Xbit_r156_c121 bl[121] br[121] wl[156] vdd gnd cell_6t
Xbit_r157_c121 bl[121] br[121] wl[157] vdd gnd cell_6t
Xbit_r158_c121 bl[121] br[121] wl[158] vdd gnd cell_6t
Xbit_r159_c121 bl[121] br[121] wl[159] vdd gnd cell_6t
Xbit_r160_c121 bl[121] br[121] wl[160] vdd gnd cell_6t
Xbit_r161_c121 bl[121] br[121] wl[161] vdd gnd cell_6t
Xbit_r162_c121 bl[121] br[121] wl[162] vdd gnd cell_6t
Xbit_r163_c121 bl[121] br[121] wl[163] vdd gnd cell_6t
Xbit_r164_c121 bl[121] br[121] wl[164] vdd gnd cell_6t
Xbit_r165_c121 bl[121] br[121] wl[165] vdd gnd cell_6t
Xbit_r166_c121 bl[121] br[121] wl[166] vdd gnd cell_6t
Xbit_r167_c121 bl[121] br[121] wl[167] vdd gnd cell_6t
Xbit_r168_c121 bl[121] br[121] wl[168] vdd gnd cell_6t
Xbit_r169_c121 bl[121] br[121] wl[169] vdd gnd cell_6t
Xbit_r170_c121 bl[121] br[121] wl[170] vdd gnd cell_6t
Xbit_r171_c121 bl[121] br[121] wl[171] vdd gnd cell_6t
Xbit_r172_c121 bl[121] br[121] wl[172] vdd gnd cell_6t
Xbit_r173_c121 bl[121] br[121] wl[173] vdd gnd cell_6t
Xbit_r174_c121 bl[121] br[121] wl[174] vdd gnd cell_6t
Xbit_r175_c121 bl[121] br[121] wl[175] vdd gnd cell_6t
Xbit_r176_c121 bl[121] br[121] wl[176] vdd gnd cell_6t
Xbit_r177_c121 bl[121] br[121] wl[177] vdd gnd cell_6t
Xbit_r178_c121 bl[121] br[121] wl[178] vdd gnd cell_6t
Xbit_r179_c121 bl[121] br[121] wl[179] vdd gnd cell_6t
Xbit_r180_c121 bl[121] br[121] wl[180] vdd gnd cell_6t
Xbit_r181_c121 bl[121] br[121] wl[181] vdd gnd cell_6t
Xbit_r182_c121 bl[121] br[121] wl[182] vdd gnd cell_6t
Xbit_r183_c121 bl[121] br[121] wl[183] vdd gnd cell_6t
Xbit_r184_c121 bl[121] br[121] wl[184] vdd gnd cell_6t
Xbit_r185_c121 bl[121] br[121] wl[185] vdd gnd cell_6t
Xbit_r186_c121 bl[121] br[121] wl[186] vdd gnd cell_6t
Xbit_r187_c121 bl[121] br[121] wl[187] vdd gnd cell_6t
Xbit_r188_c121 bl[121] br[121] wl[188] vdd gnd cell_6t
Xbit_r189_c121 bl[121] br[121] wl[189] vdd gnd cell_6t
Xbit_r190_c121 bl[121] br[121] wl[190] vdd gnd cell_6t
Xbit_r191_c121 bl[121] br[121] wl[191] vdd gnd cell_6t
Xbit_r192_c121 bl[121] br[121] wl[192] vdd gnd cell_6t
Xbit_r193_c121 bl[121] br[121] wl[193] vdd gnd cell_6t
Xbit_r194_c121 bl[121] br[121] wl[194] vdd gnd cell_6t
Xbit_r195_c121 bl[121] br[121] wl[195] vdd gnd cell_6t
Xbit_r196_c121 bl[121] br[121] wl[196] vdd gnd cell_6t
Xbit_r197_c121 bl[121] br[121] wl[197] vdd gnd cell_6t
Xbit_r198_c121 bl[121] br[121] wl[198] vdd gnd cell_6t
Xbit_r199_c121 bl[121] br[121] wl[199] vdd gnd cell_6t
Xbit_r200_c121 bl[121] br[121] wl[200] vdd gnd cell_6t
Xbit_r201_c121 bl[121] br[121] wl[201] vdd gnd cell_6t
Xbit_r202_c121 bl[121] br[121] wl[202] vdd gnd cell_6t
Xbit_r203_c121 bl[121] br[121] wl[203] vdd gnd cell_6t
Xbit_r204_c121 bl[121] br[121] wl[204] vdd gnd cell_6t
Xbit_r205_c121 bl[121] br[121] wl[205] vdd gnd cell_6t
Xbit_r206_c121 bl[121] br[121] wl[206] vdd gnd cell_6t
Xbit_r207_c121 bl[121] br[121] wl[207] vdd gnd cell_6t
Xbit_r208_c121 bl[121] br[121] wl[208] vdd gnd cell_6t
Xbit_r209_c121 bl[121] br[121] wl[209] vdd gnd cell_6t
Xbit_r210_c121 bl[121] br[121] wl[210] vdd gnd cell_6t
Xbit_r211_c121 bl[121] br[121] wl[211] vdd gnd cell_6t
Xbit_r212_c121 bl[121] br[121] wl[212] vdd gnd cell_6t
Xbit_r213_c121 bl[121] br[121] wl[213] vdd gnd cell_6t
Xbit_r214_c121 bl[121] br[121] wl[214] vdd gnd cell_6t
Xbit_r215_c121 bl[121] br[121] wl[215] vdd gnd cell_6t
Xbit_r216_c121 bl[121] br[121] wl[216] vdd gnd cell_6t
Xbit_r217_c121 bl[121] br[121] wl[217] vdd gnd cell_6t
Xbit_r218_c121 bl[121] br[121] wl[218] vdd gnd cell_6t
Xbit_r219_c121 bl[121] br[121] wl[219] vdd gnd cell_6t
Xbit_r220_c121 bl[121] br[121] wl[220] vdd gnd cell_6t
Xbit_r221_c121 bl[121] br[121] wl[221] vdd gnd cell_6t
Xbit_r222_c121 bl[121] br[121] wl[222] vdd gnd cell_6t
Xbit_r223_c121 bl[121] br[121] wl[223] vdd gnd cell_6t
Xbit_r224_c121 bl[121] br[121] wl[224] vdd gnd cell_6t
Xbit_r225_c121 bl[121] br[121] wl[225] vdd gnd cell_6t
Xbit_r226_c121 bl[121] br[121] wl[226] vdd gnd cell_6t
Xbit_r227_c121 bl[121] br[121] wl[227] vdd gnd cell_6t
Xbit_r228_c121 bl[121] br[121] wl[228] vdd gnd cell_6t
Xbit_r229_c121 bl[121] br[121] wl[229] vdd gnd cell_6t
Xbit_r230_c121 bl[121] br[121] wl[230] vdd gnd cell_6t
Xbit_r231_c121 bl[121] br[121] wl[231] vdd gnd cell_6t
Xbit_r232_c121 bl[121] br[121] wl[232] vdd gnd cell_6t
Xbit_r233_c121 bl[121] br[121] wl[233] vdd gnd cell_6t
Xbit_r234_c121 bl[121] br[121] wl[234] vdd gnd cell_6t
Xbit_r235_c121 bl[121] br[121] wl[235] vdd gnd cell_6t
Xbit_r236_c121 bl[121] br[121] wl[236] vdd gnd cell_6t
Xbit_r237_c121 bl[121] br[121] wl[237] vdd gnd cell_6t
Xbit_r238_c121 bl[121] br[121] wl[238] vdd gnd cell_6t
Xbit_r239_c121 bl[121] br[121] wl[239] vdd gnd cell_6t
Xbit_r240_c121 bl[121] br[121] wl[240] vdd gnd cell_6t
Xbit_r241_c121 bl[121] br[121] wl[241] vdd gnd cell_6t
Xbit_r242_c121 bl[121] br[121] wl[242] vdd gnd cell_6t
Xbit_r243_c121 bl[121] br[121] wl[243] vdd gnd cell_6t
Xbit_r244_c121 bl[121] br[121] wl[244] vdd gnd cell_6t
Xbit_r245_c121 bl[121] br[121] wl[245] vdd gnd cell_6t
Xbit_r246_c121 bl[121] br[121] wl[246] vdd gnd cell_6t
Xbit_r247_c121 bl[121] br[121] wl[247] vdd gnd cell_6t
Xbit_r248_c121 bl[121] br[121] wl[248] vdd gnd cell_6t
Xbit_r249_c121 bl[121] br[121] wl[249] vdd gnd cell_6t
Xbit_r250_c121 bl[121] br[121] wl[250] vdd gnd cell_6t
Xbit_r251_c121 bl[121] br[121] wl[251] vdd gnd cell_6t
Xbit_r252_c121 bl[121] br[121] wl[252] vdd gnd cell_6t
Xbit_r253_c121 bl[121] br[121] wl[253] vdd gnd cell_6t
Xbit_r254_c121 bl[121] br[121] wl[254] vdd gnd cell_6t
Xbit_r255_c121 bl[121] br[121] wl[255] vdd gnd cell_6t
Xbit_r0_c122 bl[122] br[122] wl[0] vdd gnd cell_6t
Xbit_r1_c122 bl[122] br[122] wl[1] vdd gnd cell_6t
Xbit_r2_c122 bl[122] br[122] wl[2] vdd gnd cell_6t
Xbit_r3_c122 bl[122] br[122] wl[3] vdd gnd cell_6t
Xbit_r4_c122 bl[122] br[122] wl[4] vdd gnd cell_6t
Xbit_r5_c122 bl[122] br[122] wl[5] vdd gnd cell_6t
Xbit_r6_c122 bl[122] br[122] wl[6] vdd gnd cell_6t
Xbit_r7_c122 bl[122] br[122] wl[7] vdd gnd cell_6t
Xbit_r8_c122 bl[122] br[122] wl[8] vdd gnd cell_6t
Xbit_r9_c122 bl[122] br[122] wl[9] vdd gnd cell_6t
Xbit_r10_c122 bl[122] br[122] wl[10] vdd gnd cell_6t
Xbit_r11_c122 bl[122] br[122] wl[11] vdd gnd cell_6t
Xbit_r12_c122 bl[122] br[122] wl[12] vdd gnd cell_6t
Xbit_r13_c122 bl[122] br[122] wl[13] vdd gnd cell_6t
Xbit_r14_c122 bl[122] br[122] wl[14] vdd gnd cell_6t
Xbit_r15_c122 bl[122] br[122] wl[15] vdd gnd cell_6t
Xbit_r16_c122 bl[122] br[122] wl[16] vdd gnd cell_6t
Xbit_r17_c122 bl[122] br[122] wl[17] vdd gnd cell_6t
Xbit_r18_c122 bl[122] br[122] wl[18] vdd gnd cell_6t
Xbit_r19_c122 bl[122] br[122] wl[19] vdd gnd cell_6t
Xbit_r20_c122 bl[122] br[122] wl[20] vdd gnd cell_6t
Xbit_r21_c122 bl[122] br[122] wl[21] vdd gnd cell_6t
Xbit_r22_c122 bl[122] br[122] wl[22] vdd gnd cell_6t
Xbit_r23_c122 bl[122] br[122] wl[23] vdd gnd cell_6t
Xbit_r24_c122 bl[122] br[122] wl[24] vdd gnd cell_6t
Xbit_r25_c122 bl[122] br[122] wl[25] vdd gnd cell_6t
Xbit_r26_c122 bl[122] br[122] wl[26] vdd gnd cell_6t
Xbit_r27_c122 bl[122] br[122] wl[27] vdd gnd cell_6t
Xbit_r28_c122 bl[122] br[122] wl[28] vdd gnd cell_6t
Xbit_r29_c122 bl[122] br[122] wl[29] vdd gnd cell_6t
Xbit_r30_c122 bl[122] br[122] wl[30] vdd gnd cell_6t
Xbit_r31_c122 bl[122] br[122] wl[31] vdd gnd cell_6t
Xbit_r32_c122 bl[122] br[122] wl[32] vdd gnd cell_6t
Xbit_r33_c122 bl[122] br[122] wl[33] vdd gnd cell_6t
Xbit_r34_c122 bl[122] br[122] wl[34] vdd gnd cell_6t
Xbit_r35_c122 bl[122] br[122] wl[35] vdd gnd cell_6t
Xbit_r36_c122 bl[122] br[122] wl[36] vdd gnd cell_6t
Xbit_r37_c122 bl[122] br[122] wl[37] vdd gnd cell_6t
Xbit_r38_c122 bl[122] br[122] wl[38] vdd gnd cell_6t
Xbit_r39_c122 bl[122] br[122] wl[39] vdd gnd cell_6t
Xbit_r40_c122 bl[122] br[122] wl[40] vdd gnd cell_6t
Xbit_r41_c122 bl[122] br[122] wl[41] vdd gnd cell_6t
Xbit_r42_c122 bl[122] br[122] wl[42] vdd gnd cell_6t
Xbit_r43_c122 bl[122] br[122] wl[43] vdd gnd cell_6t
Xbit_r44_c122 bl[122] br[122] wl[44] vdd gnd cell_6t
Xbit_r45_c122 bl[122] br[122] wl[45] vdd gnd cell_6t
Xbit_r46_c122 bl[122] br[122] wl[46] vdd gnd cell_6t
Xbit_r47_c122 bl[122] br[122] wl[47] vdd gnd cell_6t
Xbit_r48_c122 bl[122] br[122] wl[48] vdd gnd cell_6t
Xbit_r49_c122 bl[122] br[122] wl[49] vdd gnd cell_6t
Xbit_r50_c122 bl[122] br[122] wl[50] vdd gnd cell_6t
Xbit_r51_c122 bl[122] br[122] wl[51] vdd gnd cell_6t
Xbit_r52_c122 bl[122] br[122] wl[52] vdd gnd cell_6t
Xbit_r53_c122 bl[122] br[122] wl[53] vdd gnd cell_6t
Xbit_r54_c122 bl[122] br[122] wl[54] vdd gnd cell_6t
Xbit_r55_c122 bl[122] br[122] wl[55] vdd gnd cell_6t
Xbit_r56_c122 bl[122] br[122] wl[56] vdd gnd cell_6t
Xbit_r57_c122 bl[122] br[122] wl[57] vdd gnd cell_6t
Xbit_r58_c122 bl[122] br[122] wl[58] vdd gnd cell_6t
Xbit_r59_c122 bl[122] br[122] wl[59] vdd gnd cell_6t
Xbit_r60_c122 bl[122] br[122] wl[60] vdd gnd cell_6t
Xbit_r61_c122 bl[122] br[122] wl[61] vdd gnd cell_6t
Xbit_r62_c122 bl[122] br[122] wl[62] vdd gnd cell_6t
Xbit_r63_c122 bl[122] br[122] wl[63] vdd gnd cell_6t
Xbit_r64_c122 bl[122] br[122] wl[64] vdd gnd cell_6t
Xbit_r65_c122 bl[122] br[122] wl[65] vdd gnd cell_6t
Xbit_r66_c122 bl[122] br[122] wl[66] vdd gnd cell_6t
Xbit_r67_c122 bl[122] br[122] wl[67] vdd gnd cell_6t
Xbit_r68_c122 bl[122] br[122] wl[68] vdd gnd cell_6t
Xbit_r69_c122 bl[122] br[122] wl[69] vdd gnd cell_6t
Xbit_r70_c122 bl[122] br[122] wl[70] vdd gnd cell_6t
Xbit_r71_c122 bl[122] br[122] wl[71] vdd gnd cell_6t
Xbit_r72_c122 bl[122] br[122] wl[72] vdd gnd cell_6t
Xbit_r73_c122 bl[122] br[122] wl[73] vdd gnd cell_6t
Xbit_r74_c122 bl[122] br[122] wl[74] vdd gnd cell_6t
Xbit_r75_c122 bl[122] br[122] wl[75] vdd gnd cell_6t
Xbit_r76_c122 bl[122] br[122] wl[76] vdd gnd cell_6t
Xbit_r77_c122 bl[122] br[122] wl[77] vdd gnd cell_6t
Xbit_r78_c122 bl[122] br[122] wl[78] vdd gnd cell_6t
Xbit_r79_c122 bl[122] br[122] wl[79] vdd gnd cell_6t
Xbit_r80_c122 bl[122] br[122] wl[80] vdd gnd cell_6t
Xbit_r81_c122 bl[122] br[122] wl[81] vdd gnd cell_6t
Xbit_r82_c122 bl[122] br[122] wl[82] vdd gnd cell_6t
Xbit_r83_c122 bl[122] br[122] wl[83] vdd gnd cell_6t
Xbit_r84_c122 bl[122] br[122] wl[84] vdd gnd cell_6t
Xbit_r85_c122 bl[122] br[122] wl[85] vdd gnd cell_6t
Xbit_r86_c122 bl[122] br[122] wl[86] vdd gnd cell_6t
Xbit_r87_c122 bl[122] br[122] wl[87] vdd gnd cell_6t
Xbit_r88_c122 bl[122] br[122] wl[88] vdd gnd cell_6t
Xbit_r89_c122 bl[122] br[122] wl[89] vdd gnd cell_6t
Xbit_r90_c122 bl[122] br[122] wl[90] vdd gnd cell_6t
Xbit_r91_c122 bl[122] br[122] wl[91] vdd gnd cell_6t
Xbit_r92_c122 bl[122] br[122] wl[92] vdd gnd cell_6t
Xbit_r93_c122 bl[122] br[122] wl[93] vdd gnd cell_6t
Xbit_r94_c122 bl[122] br[122] wl[94] vdd gnd cell_6t
Xbit_r95_c122 bl[122] br[122] wl[95] vdd gnd cell_6t
Xbit_r96_c122 bl[122] br[122] wl[96] vdd gnd cell_6t
Xbit_r97_c122 bl[122] br[122] wl[97] vdd gnd cell_6t
Xbit_r98_c122 bl[122] br[122] wl[98] vdd gnd cell_6t
Xbit_r99_c122 bl[122] br[122] wl[99] vdd gnd cell_6t
Xbit_r100_c122 bl[122] br[122] wl[100] vdd gnd cell_6t
Xbit_r101_c122 bl[122] br[122] wl[101] vdd gnd cell_6t
Xbit_r102_c122 bl[122] br[122] wl[102] vdd gnd cell_6t
Xbit_r103_c122 bl[122] br[122] wl[103] vdd gnd cell_6t
Xbit_r104_c122 bl[122] br[122] wl[104] vdd gnd cell_6t
Xbit_r105_c122 bl[122] br[122] wl[105] vdd gnd cell_6t
Xbit_r106_c122 bl[122] br[122] wl[106] vdd gnd cell_6t
Xbit_r107_c122 bl[122] br[122] wl[107] vdd gnd cell_6t
Xbit_r108_c122 bl[122] br[122] wl[108] vdd gnd cell_6t
Xbit_r109_c122 bl[122] br[122] wl[109] vdd gnd cell_6t
Xbit_r110_c122 bl[122] br[122] wl[110] vdd gnd cell_6t
Xbit_r111_c122 bl[122] br[122] wl[111] vdd gnd cell_6t
Xbit_r112_c122 bl[122] br[122] wl[112] vdd gnd cell_6t
Xbit_r113_c122 bl[122] br[122] wl[113] vdd gnd cell_6t
Xbit_r114_c122 bl[122] br[122] wl[114] vdd gnd cell_6t
Xbit_r115_c122 bl[122] br[122] wl[115] vdd gnd cell_6t
Xbit_r116_c122 bl[122] br[122] wl[116] vdd gnd cell_6t
Xbit_r117_c122 bl[122] br[122] wl[117] vdd gnd cell_6t
Xbit_r118_c122 bl[122] br[122] wl[118] vdd gnd cell_6t
Xbit_r119_c122 bl[122] br[122] wl[119] vdd gnd cell_6t
Xbit_r120_c122 bl[122] br[122] wl[120] vdd gnd cell_6t
Xbit_r121_c122 bl[122] br[122] wl[121] vdd gnd cell_6t
Xbit_r122_c122 bl[122] br[122] wl[122] vdd gnd cell_6t
Xbit_r123_c122 bl[122] br[122] wl[123] vdd gnd cell_6t
Xbit_r124_c122 bl[122] br[122] wl[124] vdd gnd cell_6t
Xbit_r125_c122 bl[122] br[122] wl[125] vdd gnd cell_6t
Xbit_r126_c122 bl[122] br[122] wl[126] vdd gnd cell_6t
Xbit_r127_c122 bl[122] br[122] wl[127] vdd gnd cell_6t
Xbit_r128_c122 bl[122] br[122] wl[128] vdd gnd cell_6t
Xbit_r129_c122 bl[122] br[122] wl[129] vdd gnd cell_6t
Xbit_r130_c122 bl[122] br[122] wl[130] vdd gnd cell_6t
Xbit_r131_c122 bl[122] br[122] wl[131] vdd gnd cell_6t
Xbit_r132_c122 bl[122] br[122] wl[132] vdd gnd cell_6t
Xbit_r133_c122 bl[122] br[122] wl[133] vdd gnd cell_6t
Xbit_r134_c122 bl[122] br[122] wl[134] vdd gnd cell_6t
Xbit_r135_c122 bl[122] br[122] wl[135] vdd gnd cell_6t
Xbit_r136_c122 bl[122] br[122] wl[136] vdd gnd cell_6t
Xbit_r137_c122 bl[122] br[122] wl[137] vdd gnd cell_6t
Xbit_r138_c122 bl[122] br[122] wl[138] vdd gnd cell_6t
Xbit_r139_c122 bl[122] br[122] wl[139] vdd gnd cell_6t
Xbit_r140_c122 bl[122] br[122] wl[140] vdd gnd cell_6t
Xbit_r141_c122 bl[122] br[122] wl[141] vdd gnd cell_6t
Xbit_r142_c122 bl[122] br[122] wl[142] vdd gnd cell_6t
Xbit_r143_c122 bl[122] br[122] wl[143] vdd gnd cell_6t
Xbit_r144_c122 bl[122] br[122] wl[144] vdd gnd cell_6t
Xbit_r145_c122 bl[122] br[122] wl[145] vdd gnd cell_6t
Xbit_r146_c122 bl[122] br[122] wl[146] vdd gnd cell_6t
Xbit_r147_c122 bl[122] br[122] wl[147] vdd gnd cell_6t
Xbit_r148_c122 bl[122] br[122] wl[148] vdd gnd cell_6t
Xbit_r149_c122 bl[122] br[122] wl[149] vdd gnd cell_6t
Xbit_r150_c122 bl[122] br[122] wl[150] vdd gnd cell_6t
Xbit_r151_c122 bl[122] br[122] wl[151] vdd gnd cell_6t
Xbit_r152_c122 bl[122] br[122] wl[152] vdd gnd cell_6t
Xbit_r153_c122 bl[122] br[122] wl[153] vdd gnd cell_6t
Xbit_r154_c122 bl[122] br[122] wl[154] vdd gnd cell_6t
Xbit_r155_c122 bl[122] br[122] wl[155] vdd gnd cell_6t
Xbit_r156_c122 bl[122] br[122] wl[156] vdd gnd cell_6t
Xbit_r157_c122 bl[122] br[122] wl[157] vdd gnd cell_6t
Xbit_r158_c122 bl[122] br[122] wl[158] vdd gnd cell_6t
Xbit_r159_c122 bl[122] br[122] wl[159] vdd gnd cell_6t
Xbit_r160_c122 bl[122] br[122] wl[160] vdd gnd cell_6t
Xbit_r161_c122 bl[122] br[122] wl[161] vdd gnd cell_6t
Xbit_r162_c122 bl[122] br[122] wl[162] vdd gnd cell_6t
Xbit_r163_c122 bl[122] br[122] wl[163] vdd gnd cell_6t
Xbit_r164_c122 bl[122] br[122] wl[164] vdd gnd cell_6t
Xbit_r165_c122 bl[122] br[122] wl[165] vdd gnd cell_6t
Xbit_r166_c122 bl[122] br[122] wl[166] vdd gnd cell_6t
Xbit_r167_c122 bl[122] br[122] wl[167] vdd gnd cell_6t
Xbit_r168_c122 bl[122] br[122] wl[168] vdd gnd cell_6t
Xbit_r169_c122 bl[122] br[122] wl[169] vdd gnd cell_6t
Xbit_r170_c122 bl[122] br[122] wl[170] vdd gnd cell_6t
Xbit_r171_c122 bl[122] br[122] wl[171] vdd gnd cell_6t
Xbit_r172_c122 bl[122] br[122] wl[172] vdd gnd cell_6t
Xbit_r173_c122 bl[122] br[122] wl[173] vdd gnd cell_6t
Xbit_r174_c122 bl[122] br[122] wl[174] vdd gnd cell_6t
Xbit_r175_c122 bl[122] br[122] wl[175] vdd gnd cell_6t
Xbit_r176_c122 bl[122] br[122] wl[176] vdd gnd cell_6t
Xbit_r177_c122 bl[122] br[122] wl[177] vdd gnd cell_6t
Xbit_r178_c122 bl[122] br[122] wl[178] vdd gnd cell_6t
Xbit_r179_c122 bl[122] br[122] wl[179] vdd gnd cell_6t
Xbit_r180_c122 bl[122] br[122] wl[180] vdd gnd cell_6t
Xbit_r181_c122 bl[122] br[122] wl[181] vdd gnd cell_6t
Xbit_r182_c122 bl[122] br[122] wl[182] vdd gnd cell_6t
Xbit_r183_c122 bl[122] br[122] wl[183] vdd gnd cell_6t
Xbit_r184_c122 bl[122] br[122] wl[184] vdd gnd cell_6t
Xbit_r185_c122 bl[122] br[122] wl[185] vdd gnd cell_6t
Xbit_r186_c122 bl[122] br[122] wl[186] vdd gnd cell_6t
Xbit_r187_c122 bl[122] br[122] wl[187] vdd gnd cell_6t
Xbit_r188_c122 bl[122] br[122] wl[188] vdd gnd cell_6t
Xbit_r189_c122 bl[122] br[122] wl[189] vdd gnd cell_6t
Xbit_r190_c122 bl[122] br[122] wl[190] vdd gnd cell_6t
Xbit_r191_c122 bl[122] br[122] wl[191] vdd gnd cell_6t
Xbit_r192_c122 bl[122] br[122] wl[192] vdd gnd cell_6t
Xbit_r193_c122 bl[122] br[122] wl[193] vdd gnd cell_6t
Xbit_r194_c122 bl[122] br[122] wl[194] vdd gnd cell_6t
Xbit_r195_c122 bl[122] br[122] wl[195] vdd gnd cell_6t
Xbit_r196_c122 bl[122] br[122] wl[196] vdd gnd cell_6t
Xbit_r197_c122 bl[122] br[122] wl[197] vdd gnd cell_6t
Xbit_r198_c122 bl[122] br[122] wl[198] vdd gnd cell_6t
Xbit_r199_c122 bl[122] br[122] wl[199] vdd gnd cell_6t
Xbit_r200_c122 bl[122] br[122] wl[200] vdd gnd cell_6t
Xbit_r201_c122 bl[122] br[122] wl[201] vdd gnd cell_6t
Xbit_r202_c122 bl[122] br[122] wl[202] vdd gnd cell_6t
Xbit_r203_c122 bl[122] br[122] wl[203] vdd gnd cell_6t
Xbit_r204_c122 bl[122] br[122] wl[204] vdd gnd cell_6t
Xbit_r205_c122 bl[122] br[122] wl[205] vdd gnd cell_6t
Xbit_r206_c122 bl[122] br[122] wl[206] vdd gnd cell_6t
Xbit_r207_c122 bl[122] br[122] wl[207] vdd gnd cell_6t
Xbit_r208_c122 bl[122] br[122] wl[208] vdd gnd cell_6t
Xbit_r209_c122 bl[122] br[122] wl[209] vdd gnd cell_6t
Xbit_r210_c122 bl[122] br[122] wl[210] vdd gnd cell_6t
Xbit_r211_c122 bl[122] br[122] wl[211] vdd gnd cell_6t
Xbit_r212_c122 bl[122] br[122] wl[212] vdd gnd cell_6t
Xbit_r213_c122 bl[122] br[122] wl[213] vdd gnd cell_6t
Xbit_r214_c122 bl[122] br[122] wl[214] vdd gnd cell_6t
Xbit_r215_c122 bl[122] br[122] wl[215] vdd gnd cell_6t
Xbit_r216_c122 bl[122] br[122] wl[216] vdd gnd cell_6t
Xbit_r217_c122 bl[122] br[122] wl[217] vdd gnd cell_6t
Xbit_r218_c122 bl[122] br[122] wl[218] vdd gnd cell_6t
Xbit_r219_c122 bl[122] br[122] wl[219] vdd gnd cell_6t
Xbit_r220_c122 bl[122] br[122] wl[220] vdd gnd cell_6t
Xbit_r221_c122 bl[122] br[122] wl[221] vdd gnd cell_6t
Xbit_r222_c122 bl[122] br[122] wl[222] vdd gnd cell_6t
Xbit_r223_c122 bl[122] br[122] wl[223] vdd gnd cell_6t
Xbit_r224_c122 bl[122] br[122] wl[224] vdd gnd cell_6t
Xbit_r225_c122 bl[122] br[122] wl[225] vdd gnd cell_6t
Xbit_r226_c122 bl[122] br[122] wl[226] vdd gnd cell_6t
Xbit_r227_c122 bl[122] br[122] wl[227] vdd gnd cell_6t
Xbit_r228_c122 bl[122] br[122] wl[228] vdd gnd cell_6t
Xbit_r229_c122 bl[122] br[122] wl[229] vdd gnd cell_6t
Xbit_r230_c122 bl[122] br[122] wl[230] vdd gnd cell_6t
Xbit_r231_c122 bl[122] br[122] wl[231] vdd gnd cell_6t
Xbit_r232_c122 bl[122] br[122] wl[232] vdd gnd cell_6t
Xbit_r233_c122 bl[122] br[122] wl[233] vdd gnd cell_6t
Xbit_r234_c122 bl[122] br[122] wl[234] vdd gnd cell_6t
Xbit_r235_c122 bl[122] br[122] wl[235] vdd gnd cell_6t
Xbit_r236_c122 bl[122] br[122] wl[236] vdd gnd cell_6t
Xbit_r237_c122 bl[122] br[122] wl[237] vdd gnd cell_6t
Xbit_r238_c122 bl[122] br[122] wl[238] vdd gnd cell_6t
Xbit_r239_c122 bl[122] br[122] wl[239] vdd gnd cell_6t
Xbit_r240_c122 bl[122] br[122] wl[240] vdd gnd cell_6t
Xbit_r241_c122 bl[122] br[122] wl[241] vdd gnd cell_6t
Xbit_r242_c122 bl[122] br[122] wl[242] vdd gnd cell_6t
Xbit_r243_c122 bl[122] br[122] wl[243] vdd gnd cell_6t
Xbit_r244_c122 bl[122] br[122] wl[244] vdd gnd cell_6t
Xbit_r245_c122 bl[122] br[122] wl[245] vdd gnd cell_6t
Xbit_r246_c122 bl[122] br[122] wl[246] vdd gnd cell_6t
Xbit_r247_c122 bl[122] br[122] wl[247] vdd gnd cell_6t
Xbit_r248_c122 bl[122] br[122] wl[248] vdd gnd cell_6t
Xbit_r249_c122 bl[122] br[122] wl[249] vdd gnd cell_6t
Xbit_r250_c122 bl[122] br[122] wl[250] vdd gnd cell_6t
Xbit_r251_c122 bl[122] br[122] wl[251] vdd gnd cell_6t
Xbit_r252_c122 bl[122] br[122] wl[252] vdd gnd cell_6t
Xbit_r253_c122 bl[122] br[122] wl[253] vdd gnd cell_6t
Xbit_r254_c122 bl[122] br[122] wl[254] vdd gnd cell_6t
Xbit_r255_c122 bl[122] br[122] wl[255] vdd gnd cell_6t
Xbit_r0_c123 bl[123] br[123] wl[0] vdd gnd cell_6t
Xbit_r1_c123 bl[123] br[123] wl[1] vdd gnd cell_6t
Xbit_r2_c123 bl[123] br[123] wl[2] vdd gnd cell_6t
Xbit_r3_c123 bl[123] br[123] wl[3] vdd gnd cell_6t
Xbit_r4_c123 bl[123] br[123] wl[4] vdd gnd cell_6t
Xbit_r5_c123 bl[123] br[123] wl[5] vdd gnd cell_6t
Xbit_r6_c123 bl[123] br[123] wl[6] vdd gnd cell_6t
Xbit_r7_c123 bl[123] br[123] wl[7] vdd gnd cell_6t
Xbit_r8_c123 bl[123] br[123] wl[8] vdd gnd cell_6t
Xbit_r9_c123 bl[123] br[123] wl[9] vdd gnd cell_6t
Xbit_r10_c123 bl[123] br[123] wl[10] vdd gnd cell_6t
Xbit_r11_c123 bl[123] br[123] wl[11] vdd gnd cell_6t
Xbit_r12_c123 bl[123] br[123] wl[12] vdd gnd cell_6t
Xbit_r13_c123 bl[123] br[123] wl[13] vdd gnd cell_6t
Xbit_r14_c123 bl[123] br[123] wl[14] vdd gnd cell_6t
Xbit_r15_c123 bl[123] br[123] wl[15] vdd gnd cell_6t
Xbit_r16_c123 bl[123] br[123] wl[16] vdd gnd cell_6t
Xbit_r17_c123 bl[123] br[123] wl[17] vdd gnd cell_6t
Xbit_r18_c123 bl[123] br[123] wl[18] vdd gnd cell_6t
Xbit_r19_c123 bl[123] br[123] wl[19] vdd gnd cell_6t
Xbit_r20_c123 bl[123] br[123] wl[20] vdd gnd cell_6t
Xbit_r21_c123 bl[123] br[123] wl[21] vdd gnd cell_6t
Xbit_r22_c123 bl[123] br[123] wl[22] vdd gnd cell_6t
Xbit_r23_c123 bl[123] br[123] wl[23] vdd gnd cell_6t
Xbit_r24_c123 bl[123] br[123] wl[24] vdd gnd cell_6t
Xbit_r25_c123 bl[123] br[123] wl[25] vdd gnd cell_6t
Xbit_r26_c123 bl[123] br[123] wl[26] vdd gnd cell_6t
Xbit_r27_c123 bl[123] br[123] wl[27] vdd gnd cell_6t
Xbit_r28_c123 bl[123] br[123] wl[28] vdd gnd cell_6t
Xbit_r29_c123 bl[123] br[123] wl[29] vdd gnd cell_6t
Xbit_r30_c123 bl[123] br[123] wl[30] vdd gnd cell_6t
Xbit_r31_c123 bl[123] br[123] wl[31] vdd gnd cell_6t
Xbit_r32_c123 bl[123] br[123] wl[32] vdd gnd cell_6t
Xbit_r33_c123 bl[123] br[123] wl[33] vdd gnd cell_6t
Xbit_r34_c123 bl[123] br[123] wl[34] vdd gnd cell_6t
Xbit_r35_c123 bl[123] br[123] wl[35] vdd gnd cell_6t
Xbit_r36_c123 bl[123] br[123] wl[36] vdd gnd cell_6t
Xbit_r37_c123 bl[123] br[123] wl[37] vdd gnd cell_6t
Xbit_r38_c123 bl[123] br[123] wl[38] vdd gnd cell_6t
Xbit_r39_c123 bl[123] br[123] wl[39] vdd gnd cell_6t
Xbit_r40_c123 bl[123] br[123] wl[40] vdd gnd cell_6t
Xbit_r41_c123 bl[123] br[123] wl[41] vdd gnd cell_6t
Xbit_r42_c123 bl[123] br[123] wl[42] vdd gnd cell_6t
Xbit_r43_c123 bl[123] br[123] wl[43] vdd gnd cell_6t
Xbit_r44_c123 bl[123] br[123] wl[44] vdd gnd cell_6t
Xbit_r45_c123 bl[123] br[123] wl[45] vdd gnd cell_6t
Xbit_r46_c123 bl[123] br[123] wl[46] vdd gnd cell_6t
Xbit_r47_c123 bl[123] br[123] wl[47] vdd gnd cell_6t
Xbit_r48_c123 bl[123] br[123] wl[48] vdd gnd cell_6t
Xbit_r49_c123 bl[123] br[123] wl[49] vdd gnd cell_6t
Xbit_r50_c123 bl[123] br[123] wl[50] vdd gnd cell_6t
Xbit_r51_c123 bl[123] br[123] wl[51] vdd gnd cell_6t
Xbit_r52_c123 bl[123] br[123] wl[52] vdd gnd cell_6t
Xbit_r53_c123 bl[123] br[123] wl[53] vdd gnd cell_6t
Xbit_r54_c123 bl[123] br[123] wl[54] vdd gnd cell_6t
Xbit_r55_c123 bl[123] br[123] wl[55] vdd gnd cell_6t
Xbit_r56_c123 bl[123] br[123] wl[56] vdd gnd cell_6t
Xbit_r57_c123 bl[123] br[123] wl[57] vdd gnd cell_6t
Xbit_r58_c123 bl[123] br[123] wl[58] vdd gnd cell_6t
Xbit_r59_c123 bl[123] br[123] wl[59] vdd gnd cell_6t
Xbit_r60_c123 bl[123] br[123] wl[60] vdd gnd cell_6t
Xbit_r61_c123 bl[123] br[123] wl[61] vdd gnd cell_6t
Xbit_r62_c123 bl[123] br[123] wl[62] vdd gnd cell_6t
Xbit_r63_c123 bl[123] br[123] wl[63] vdd gnd cell_6t
Xbit_r64_c123 bl[123] br[123] wl[64] vdd gnd cell_6t
Xbit_r65_c123 bl[123] br[123] wl[65] vdd gnd cell_6t
Xbit_r66_c123 bl[123] br[123] wl[66] vdd gnd cell_6t
Xbit_r67_c123 bl[123] br[123] wl[67] vdd gnd cell_6t
Xbit_r68_c123 bl[123] br[123] wl[68] vdd gnd cell_6t
Xbit_r69_c123 bl[123] br[123] wl[69] vdd gnd cell_6t
Xbit_r70_c123 bl[123] br[123] wl[70] vdd gnd cell_6t
Xbit_r71_c123 bl[123] br[123] wl[71] vdd gnd cell_6t
Xbit_r72_c123 bl[123] br[123] wl[72] vdd gnd cell_6t
Xbit_r73_c123 bl[123] br[123] wl[73] vdd gnd cell_6t
Xbit_r74_c123 bl[123] br[123] wl[74] vdd gnd cell_6t
Xbit_r75_c123 bl[123] br[123] wl[75] vdd gnd cell_6t
Xbit_r76_c123 bl[123] br[123] wl[76] vdd gnd cell_6t
Xbit_r77_c123 bl[123] br[123] wl[77] vdd gnd cell_6t
Xbit_r78_c123 bl[123] br[123] wl[78] vdd gnd cell_6t
Xbit_r79_c123 bl[123] br[123] wl[79] vdd gnd cell_6t
Xbit_r80_c123 bl[123] br[123] wl[80] vdd gnd cell_6t
Xbit_r81_c123 bl[123] br[123] wl[81] vdd gnd cell_6t
Xbit_r82_c123 bl[123] br[123] wl[82] vdd gnd cell_6t
Xbit_r83_c123 bl[123] br[123] wl[83] vdd gnd cell_6t
Xbit_r84_c123 bl[123] br[123] wl[84] vdd gnd cell_6t
Xbit_r85_c123 bl[123] br[123] wl[85] vdd gnd cell_6t
Xbit_r86_c123 bl[123] br[123] wl[86] vdd gnd cell_6t
Xbit_r87_c123 bl[123] br[123] wl[87] vdd gnd cell_6t
Xbit_r88_c123 bl[123] br[123] wl[88] vdd gnd cell_6t
Xbit_r89_c123 bl[123] br[123] wl[89] vdd gnd cell_6t
Xbit_r90_c123 bl[123] br[123] wl[90] vdd gnd cell_6t
Xbit_r91_c123 bl[123] br[123] wl[91] vdd gnd cell_6t
Xbit_r92_c123 bl[123] br[123] wl[92] vdd gnd cell_6t
Xbit_r93_c123 bl[123] br[123] wl[93] vdd gnd cell_6t
Xbit_r94_c123 bl[123] br[123] wl[94] vdd gnd cell_6t
Xbit_r95_c123 bl[123] br[123] wl[95] vdd gnd cell_6t
Xbit_r96_c123 bl[123] br[123] wl[96] vdd gnd cell_6t
Xbit_r97_c123 bl[123] br[123] wl[97] vdd gnd cell_6t
Xbit_r98_c123 bl[123] br[123] wl[98] vdd gnd cell_6t
Xbit_r99_c123 bl[123] br[123] wl[99] vdd gnd cell_6t
Xbit_r100_c123 bl[123] br[123] wl[100] vdd gnd cell_6t
Xbit_r101_c123 bl[123] br[123] wl[101] vdd gnd cell_6t
Xbit_r102_c123 bl[123] br[123] wl[102] vdd gnd cell_6t
Xbit_r103_c123 bl[123] br[123] wl[103] vdd gnd cell_6t
Xbit_r104_c123 bl[123] br[123] wl[104] vdd gnd cell_6t
Xbit_r105_c123 bl[123] br[123] wl[105] vdd gnd cell_6t
Xbit_r106_c123 bl[123] br[123] wl[106] vdd gnd cell_6t
Xbit_r107_c123 bl[123] br[123] wl[107] vdd gnd cell_6t
Xbit_r108_c123 bl[123] br[123] wl[108] vdd gnd cell_6t
Xbit_r109_c123 bl[123] br[123] wl[109] vdd gnd cell_6t
Xbit_r110_c123 bl[123] br[123] wl[110] vdd gnd cell_6t
Xbit_r111_c123 bl[123] br[123] wl[111] vdd gnd cell_6t
Xbit_r112_c123 bl[123] br[123] wl[112] vdd gnd cell_6t
Xbit_r113_c123 bl[123] br[123] wl[113] vdd gnd cell_6t
Xbit_r114_c123 bl[123] br[123] wl[114] vdd gnd cell_6t
Xbit_r115_c123 bl[123] br[123] wl[115] vdd gnd cell_6t
Xbit_r116_c123 bl[123] br[123] wl[116] vdd gnd cell_6t
Xbit_r117_c123 bl[123] br[123] wl[117] vdd gnd cell_6t
Xbit_r118_c123 bl[123] br[123] wl[118] vdd gnd cell_6t
Xbit_r119_c123 bl[123] br[123] wl[119] vdd gnd cell_6t
Xbit_r120_c123 bl[123] br[123] wl[120] vdd gnd cell_6t
Xbit_r121_c123 bl[123] br[123] wl[121] vdd gnd cell_6t
Xbit_r122_c123 bl[123] br[123] wl[122] vdd gnd cell_6t
Xbit_r123_c123 bl[123] br[123] wl[123] vdd gnd cell_6t
Xbit_r124_c123 bl[123] br[123] wl[124] vdd gnd cell_6t
Xbit_r125_c123 bl[123] br[123] wl[125] vdd gnd cell_6t
Xbit_r126_c123 bl[123] br[123] wl[126] vdd gnd cell_6t
Xbit_r127_c123 bl[123] br[123] wl[127] vdd gnd cell_6t
Xbit_r128_c123 bl[123] br[123] wl[128] vdd gnd cell_6t
Xbit_r129_c123 bl[123] br[123] wl[129] vdd gnd cell_6t
Xbit_r130_c123 bl[123] br[123] wl[130] vdd gnd cell_6t
Xbit_r131_c123 bl[123] br[123] wl[131] vdd gnd cell_6t
Xbit_r132_c123 bl[123] br[123] wl[132] vdd gnd cell_6t
Xbit_r133_c123 bl[123] br[123] wl[133] vdd gnd cell_6t
Xbit_r134_c123 bl[123] br[123] wl[134] vdd gnd cell_6t
Xbit_r135_c123 bl[123] br[123] wl[135] vdd gnd cell_6t
Xbit_r136_c123 bl[123] br[123] wl[136] vdd gnd cell_6t
Xbit_r137_c123 bl[123] br[123] wl[137] vdd gnd cell_6t
Xbit_r138_c123 bl[123] br[123] wl[138] vdd gnd cell_6t
Xbit_r139_c123 bl[123] br[123] wl[139] vdd gnd cell_6t
Xbit_r140_c123 bl[123] br[123] wl[140] vdd gnd cell_6t
Xbit_r141_c123 bl[123] br[123] wl[141] vdd gnd cell_6t
Xbit_r142_c123 bl[123] br[123] wl[142] vdd gnd cell_6t
Xbit_r143_c123 bl[123] br[123] wl[143] vdd gnd cell_6t
Xbit_r144_c123 bl[123] br[123] wl[144] vdd gnd cell_6t
Xbit_r145_c123 bl[123] br[123] wl[145] vdd gnd cell_6t
Xbit_r146_c123 bl[123] br[123] wl[146] vdd gnd cell_6t
Xbit_r147_c123 bl[123] br[123] wl[147] vdd gnd cell_6t
Xbit_r148_c123 bl[123] br[123] wl[148] vdd gnd cell_6t
Xbit_r149_c123 bl[123] br[123] wl[149] vdd gnd cell_6t
Xbit_r150_c123 bl[123] br[123] wl[150] vdd gnd cell_6t
Xbit_r151_c123 bl[123] br[123] wl[151] vdd gnd cell_6t
Xbit_r152_c123 bl[123] br[123] wl[152] vdd gnd cell_6t
Xbit_r153_c123 bl[123] br[123] wl[153] vdd gnd cell_6t
Xbit_r154_c123 bl[123] br[123] wl[154] vdd gnd cell_6t
Xbit_r155_c123 bl[123] br[123] wl[155] vdd gnd cell_6t
Xbit_r156_c123 bl[123] br[123] wl[156] vdd gnd cell_6t
Xbit_r157_c123 bl[123] br[123] wl[157] vdd gnd cell_6t
Xbit_r158_c123 bl[123] br[123] wl[158] vdd gnd cell_6t
Xbit_r159_c123 bl[123] br[123] wl[159] vdd gnd cell_6t
Xbit_r160_c123 bl[123] br[123] wl[160] vdd gnd cell_6t
Xbit_r161_c123 bl[123] br[123] wl[161] vdd gnd cell_6t
Xbit_r162_c123 bl[123] br[123] wl[162] vdd gnd cell_6t
Xbit_r163_c123 bl[123] br[123] wl[163] vdd gnd cell_6t
Xbit_r164_c123 bl[123] br[123] wl[164] vdd gnd cell_6t
Xbit_r165_c123 bl[123] br[123] wl[165] vdd gnd cell_6t
Xbit_r166_c123 bl[123] br[123] wl[166] vdd gnd cell_6t
Xbit_r167_c123 bl[123] br[123] wl[167] vdd gnd cell_6t
Xbit_r168_c123 bl[123] br[123] wl[168] vdd gnd cell_6t
Xbit_r169_c123 bl[123] br[123] wl[169] vdd gnd cell_6t
Xbit_r170_c123 bl[123] br[123] wl[170] vdd gnd cell_6t
Xbit_r171_c123 bl[123] br[123] wl[171] vdd gnd cell_6t
Xbit_r172_c123 bl[123] br[123] wl[172] vdd gnd cell_6t
Xbit_r173_c123 bl[123] br[123] wl[173] vdd gnd cell_6t
Xbit_r174_c123 bl[123] br[123] wl[174] vdd gnd cell_6t
Xbit_r175_c123 bl[123] br[123] wl[175] vdd gnd cell_6t
Xbit_r176_c123 bl[123] br[123] wl[176] vdd gnd cell_6t
Xbit_r177_c123 bl[123] br[123] wl[177] vdd gnd cell_6t
Xbit_r178_c123 bl[123] br[123] wl[178] vdd gnd cell_6t
Xbit_r179_c123 bl[123] br[123] wl[179] vdd gnd cell_6t
Xbit_r180_c123 bl[123] br[123] wl[180] vdd gnd cell_6t
Xbit_r181_c123 bl[123] br[123] wl[181] vdd gnd cell_6t
Xbit_r182_c123 bl[123] br[123] wl[182] vdd gnd cell_6t
Xbit_r183_c123 bl[123] br[123] wl[183] vdd gnd cell_6t
Xbit_r184_c123 bl[123] br[123] wl[184] vdd gnd cell_6t
Xbit_r185_c123 bl[123] br[123] wl[185] vdd gnd cell_6t
Xbit_r186_c123 bl[123] br[123] wl[186] vdd gnd cell_6t
Xbit_r187_c123 bl[123] br[123] wl[187] vdd gnd cell_6t
Xbit_r188_c123 bl[123] br[123] wl[188] vdd gnd cell_6t
Xbit_r189_c123 bl[123] br[123] wl[189] vdd gnd cell_6t
Xbit_r190_c123 bl[123] br[123] wl[190] vdd gnd cell_6t
Xbit_r191_c123 bl[123] br[123] wl[191] vdd gnd cell_6t
Xbit_r192_c123 bl[123] br[123] wl[192] vdd gnd cell_6t
Xbit_r193_c123 bl[123] br[123] wl[193] vdd gnd cell_6t
Xbit_r194_c123 bl[123] br[123] wl[194] vdd gnd cell_6t
Xbit_r195_c123 bl[123] br[123] wl[195] vdd gnd cell_6t
Xbit_r196_c123 bl[123] br[123] wl[196] vdd gnd cell_6t
Xbit_r197_c123 bl[123] br[123] wl[197] vdd gnd cell_6t
Xbit_r198_c123 bl[123] br[123] wl[198] vdd gnd cell_6t
Xbit_r199_c123 bl[123] br[123] wl[199] vdd gnd cell_6t
Xbit_r200_c123 bl[123] br[123] wl[200] vdd gnd cell_6t
Xbit_r201_c123 bl[123] br[123] wl[201] vdd gnd cell_6t
Xbit_r202_c123 bl[123] br[123] wl[202] vdd gnd cell_6t
Xbit_r203_c123 bl[123] br[123] wl[203] vdd gnd cell_6t
Xbit_r204_c123 bl[123] br[123] wl[204] vdd gnd cell_6t
Xbit_r205_c123 bl[123] br[123] wl[205] vdd gnd cell_6t
Xbit_r206_c123 bl[123] br[123] wl[206] vdd gnd cell_6t
Xbit_r207_c123 bl[123] br[123] wl[207] vdd gnd cell_6t
Xbit_r208_c123 bl[123] br[123] wl[208] vdd gnd cell_6t
Xbit_r209_c123 bl[123] br[123] wl[209] vdd gnd cell_6t
Xbit_r210_c123 bl[123] br[123] wl[210] vdd gnd cell_6t
Xbit_r211_c123 bl[123] br[123] wl[211] vdd gnd cell_6t
Xbit_r212_c123 bl[123] br[123] wl[212] vdd gnd cell_6t
Xbit_r213_c123 bl[123] br[123] wl[213] vdd gnd cell_6t
Xbit_r214_c123 bl[123] br[123] wl[214] vdd gnd cell_6t
Xbit_r215_c123 bl[123] br[123] wl[215] vdd gnd cell_6t
Xbit_r216_c123 bl[123] br[123] wl[216] vdd gnd cell_6t
Xbit_r217_c123 bl[123] br[123] wl[217] vdd gnd cell_6t
Xbit_r218_c123 bl[123] br[123] wl[218] vdd gnd cell_6t
Xbit_r219_c123 bl[123] br[123] wl[219] vdd gnd cell_6t
Xbit_r220_c123 bl[123] br[123] wl[220] vdd gnd cell_6t
Xbit_r221_c123 bl[123] br[123] wl[221] vdd gnd cell_6t
Xbit_r222_c123 bl[123] br[123] wl[222] vdd gnd cell_6t
Xbit_r223_c123 bl[123] br[123] wl[223] vdd gnd cell_6t
Xbit_r224_c123 bl[123] br[123] wl[224] vdd gnd cell_6t
Xbit_r225_c123 bl[123] br[123] wl[225] vdd gnd cell_6t
Xbit_r226_c123 bl[123] br[123] wl[226] vdd gnd cell_6t
Xbit_r227_c123 bl[123] br[123] wl[227] vdd gnd cell_6t
Xbit_r228_c123 bl[123] br[123] wl[228] vdd gnd cell_6t
Xbit_r229_c123 bl[123] br[123] wl[229] vdd gnd cell_6t
Xbit_r230_c123 bl[123] br[123] wl[230] vdd gnd cell_6t
Xbit_r231_c123 bl[123] br[123] wl[231] vdd gnd cell_6t
Xbit_r232_c123 bl[123] br[123] wl[232] vdd gnd cell_6t
Xbit_r233_c123 bl[123] br[123] wl[233] vdd gnd cell_6t
Xbit_r234_c123 bl[123] br[123] wl[234] vdd gnd cell_6t
Xbit_r235_c123 bl[123] br[123] wl[235] vdd gnd cell_6t
Xbit_r236_c123 bl[123] br[123] wl[236] vdd gnd cell_6t
Xbit_r237_c123 bl[123] br[123] wl[237] vdd gnd cell_6t
Xbit_r238_c123 bl[123] br[123] wl[238] vdd gnd cell_6t
Xbit_r239_c123 bl[123] br[123] wl[239] vdd gnd cell_6t
Xbit_r240_c123 bl[123] br[123] wl[240] vdd gnd cell_6t
Xbit_r241_c123 bl[123] br[123] wl[241] vdd gnd cell_6t
Xbit_r242_c123 bl[123] br[123] wl[242] vdd gnd cell_6t
Xbit_r243_c123 bl[123] br[123] wl[243] vdd gnd cell_6t
Xbit_r244_c123 bl[123] br[123] wl[244] vdd gnd cell_6t
Xbit_r245_c123 bl[123] br[123] wl[245] vdd gnd cell_6t
Xbit_r246_c123 bl[123] br[123] wl[246] vdd gnd cell_6t
Xbit_r247_c123 bl[123] br[123] wl[247] vdd gnd cell_6t
Xbit_r248_c123 bl[123] br[123] wl[248] vdd gnd cell_6t
Xbit_r249_c123 bl[123] br[123] wl[249] vdd gnd cell_6t
Xbit_r250_c123 bl[123] br[123] wl[250] vdd gnd cell_6t
Xbit_r251_c123 bl[123] br[123] wl[251] vdd gnd cell_6t
Xbit_r252_c123 bl[123] br[123] wl[252] vdd gnd cell_6t
Xbit_r253_c123 bl[123] br[123] wl[253] vdd gnd cell_6t
Xbit_r254_c123 bl[123] br[123] wl[254] vdd gnd cell_6t
Xbit_r255_c123 bl[123] br[123] wl[255] vdd gnd cell_6t
Xbit_r0_c124 bl[124] br[124] wl[0] vdd gnd cell_6t
Xbit_r1_c124 bl[124] br[124] wl[1] vdd gnd cell_6t
Xbit_r2_c124 bl[124] br[124] wl[2] vdd gnd cell_6t
Xbit_r3_c124 bl[124] br[124] wl[3] vdd gnd cell_6t
Xbit_r4_c124 bl[124] br[124] wl[4] vdd gnd cell_6t
Xbit_r5_c124 bl[124] br[124] wl[5] vdd gnd cell_6t
Xbit_r6_c124 bl[124] br[124] wl[6] vdd gnd cell_6t
Xbit_r7_c124 bl[124] br[124] wl[7] vdd gnd cell_6t
Xbit_r8_c124 bl[124] br[124] wl[8] vdd gnd cell_6t
Xbit_r9_c124 bl[124] br[124] wl[9] vdd gnd cell_6t
Xbit_r10_c124 bl[124] br[124] wl[10] vdd gnd cell_6t
Xbit_r11_c124 bl[124] br[124] wl[11] vdd gnd cell_6t
Xbit_r12_c124 bl[124] br[124] wl[12] vdd gnd cell_6t
Xbit_r13_c124 bl[124] br[124] wl[13] vdd gnd cell_6t
Xbit_r14_c124 bl[124] br[124] wl[14] vdd gnd cell_6t
Xbit_r15_c124 bl[124] br[124] wl[15] vdd gnd cell_6t
Xbit_r16_c124 bl[124] br[124] wl[16] vdd gnd cell_6t
Xbit_r17_c124 bl[124] br[124] wl[17] vdd gnd cell_6t
Xbit_r18_c124 bl[124] br[124] wl[18] vdd gnd cell_6t
Xbit_r19_c124 bl[124] br[124] wl[19] vdd gnd cell_6t
Xbit_r20_c124 bl[124] br[124] wl[20] vdd gnd cell_6t
Xbit_r21_c124 bl[124] br[124] wl[21] vdd gnd cell_6t
Xbit_r22_c124 bl[124] br[124] wl[22] vdd gnd cell_6t
Xbit_r23_c124 bl[124] br[124] wl[23] vdd gnd cell_6t
Xbit_r24_c124 bl[124] br[124] wl[24] vdd gnd cell_6t
Xbit_r25_c124 bl[124] br[124] wl[25] vdd gnd cell_6t
Xbit_r26_c124 bl[124] br[124] wl[26] vdd gnd cell_6t
Xbit_r27_c124 bl[124] br[124] wl[27] vdd gnd cell_6t
Xbit_r28_c124 bl[124] br[124] wl[28] vdd gnd cell_6t
Xbit_r29_c124 bl[124] br[124] wl[29] vdd gnd cell_6t
Xbit_r30_c124 bl[124] br[124] wl[30] vdd gnd cell_6t
Xbit_r31_c124 bl[124] br[124] wl[31] vdd gnd cell_6t
Xbit_r32_c124 bl[124] br[124] wl[32] vdd gnd cell_6t
Xbit_r33_c124 bl[124] br[124] wl[33] vdd gnd cell_6t
Xbit_r34_c124 bl[124] br[124] wl[34] vdd gnd cell_6t
Xbit_r35_c124 bl[124] br[124] wl[35] vdd gnd cell_6t
Xbit_r36_c124 bl[124] br[124] wl[36] vdd gnd cell_6t
Xbit_r37_c124 bl[124] br[124] wl[37] vdd gnd cell_6t
Xbit_r38_c124 bl[124] br[124] wl[38] vdd gnd cell_6t
Xbit_r39_c124 bl[124] br[124] wl[39] vdd gnd cell_6t
Xbit_r40_c124 bl[124] br[124] wl[40] vdd gnd cell_6t
Xbit_r41_c124 bl[124] br[124] wl[41] vdd gnd cell_6t
Xbit_r42_c124 bl[124] br[124] wl[42] vdd gnd cell_6t
Xbit_r43_c124 bl[124] br[124] wl[43] vdd gnd cell_6t
Xbit_r44_c124 bl[124] br[124] wl[44] vdd gnd cell_6t
Xbit_r45_c124 bl[124] br[124] wl[45] vdd gnd cell_6t
Xbit_r46_c124 bl[124] br[124] wl[46] vdd gnd cell_6t
Xbit_r47_c124 bl[124] br[124] wl[47] vdd gnd cell_6t
Xbit_r48_c124 bl[124] br[124] wl[48] vdd gnd cell_6t
Xbit_r49_c124 bl[124] br[124] wl[49] vdd gnd cell_6t
Xbit_r50_c124 bl[124] br[124] wl[50] vdd gnd cell_6t
Xbit_r51_c124 bl[124] br[124] wl[51] vdd gnd cell_6t
Xbit_r52_c124 bl[124] br[124] wl[52] vdd gnd cell_6t
Xbit_r53_c124 bl[124] br[124] wl[53] vdd gnd cell_6t
Xbit_r54_c124 bl[124] br[124] wl[54] vdd gnd cell_6t
Xbit_r55_c124 bl[124] br[124] wl[55] vdd gnd cell_6t
Xbit_r56_c124 bl[124] br[124] wl[56] vdd gnd cell_6t
Xbit_r57_c124 bl[124] br[124] wl[57] vdd gnd cell_6t
Xbit_r58_c124 bl[124] br[124] wl[58] vdd gnd cell_6t
Xbit_r59_c124 bl[124] br[124] wl[59] vdd gnd cell_6t
Xbit_r60_c124 bl[124] br[124] wl[60] vdd gnd cell_6t
Xbit_r61_c124 bl[124] br[124] wl[61] vdd gnd cell_6t
Xbit_r62_c124 bl[124] br[124] wl[62] vdd gnd cell_6t
Xbit_r63_c124 bl[124] br[124] wl[63] vdd gnd cell_6t
Xbit_r64_c124 bl[124] br[124] wl[64] vdd gnd cell_6t
Xbit_r65_c124 bl[124] br[124] wl[65] vdd gnd cell_6t
Xbit_r66_c124 bl[124] br[124] wl[66] vdd gnd cell_6t
Xbit_r67_c124 bl[124] br[124] wl[67] vdd gnd cell_6t
Xbit_r68_c124 bl[124] br[124] wl[68] vdd gnd cell_6t
Xbit_r69_c124 bl[124] br[124] wl[69] vdd gnd cell_6t
Xbit_r70_c124 bl[124] br[124] wl[70] vdd gnd cell_6t
Xbit_r71_c124 bl[124] br[124] wl[71] vdd gnd cell_6t
Xbit_r72_c124 bl[124] br[124] wl[72] vdd gnd cell_6t
Xbit_r73_c124 bl[124] br[124] wl[73] vdd gnd cell_6t
Xbit_r74_c124 bl[124] br[124] wl[74] vdd gnd cell_6t
Xbit_r75_c124 bl[124] br[124] wl[75] vdd gnd cell_6t
Xbit_r76_c124 bl[124] br[124] wl[76] vdd gnd cell_6t
Xbit_r77_c124 bl[124] br[124] wl[77] vdd gnd cell_6t
Xbit_r78_c124 bl[124] br[124] wl[78] vdd gnd cell_6t
Xbit_r79_c124 bl[124] br[124] wl[79] vdd gnd cell_6t
Xbit_r80_c124 bl[124] br[124] wl[80] vdd gnd cell_6t
Xbit_r81_c124 bl[124] br[124] wl[81] vdd gnd cell_6t
Xbit_r82_c124 bl[124] br[124] wl[82] vdd gnd cell_6t
Xbit_r83_c124 bl[124] br[124] wl[83] vdd gnd cell_6t
Xbit_r84_c124 bl[124] br[124] wl[84] vdd gnd cell_6t
Xbit_r85_c124 bl[124] br[124] wl[85] vdd gnd cell_6t
Xbit_r86_c124 bl[124] br[124] wl[86] vdd gnd cell_6t
Xbit_r87_c124 bl[124] br[124] wl[87] vdd gnd cell_6t
Xbit_r88_c124 bl[124] br[124] wl[88] vdd gnd cell_6t
Xbit_r89_c124 bl[124] br[124] wl[89] vdd gnd cell_6t
Xbit_r90_c124 bl[124] br[124] wl[90] vdd gnd cell_6t
Xbit_r91_c124 bl[124] br[124] wl[91] vdd gnd cell_6t
Xbit_r92_c124 bl[124] br[124] wl[92] vdd gnd cell_6t
Xbit_r93_c124 bl[124] br[124] wl[93] vdd gnd cell_6t
Xbit_r94_c124 bl[124] br[124] wl[94] vdd gnd cell_6t
Xbit_r95_c124 bl[124] br[124] wl[95] vdd gnd cell_6t
Xbit_r96_c124 bl[124] br[124] wl[96] vdd gnd cell_6t
Xbit_r97_c124 bl[124] br[124] wl[97] vdd gnd cell_6t
Xbit_r98_c124 bl[124] br[124] wl[98] vdd gnd cell_6t
Xbit_r99_c124 bl[124] br[124] wl[99] vdd gnd cell_6t
Xbit_r100_c124 bl[124] br[124] wl[100] vdd gnd cell_6t
Xbit_r101_c124 bl[124] br[124] wl[101] vdd gnd cell_6t
Xbit_r102_c124 bl[124] br[124] wl[102] vdd gnd cell_6t
Xbit_r103_c124 bl[124] br[124] wl[103] vdd gnd cell_6t
Xbit_r104_c124 bl[124] br[124] wl[104] vdd gnd cell_6t
Xbit_r105_c124 bl[124] br[124] wl[105] vdd gnd cell_6t
Xbit_r106_c124 bl[124] br[124] wl[106] vdd gnd cell_6t
Xbit_r107_c124 bl[124] br[124] wl[107] vdd gnd cell_6t
Xbit_r108_c124 bl[124] br[124] wl[108] vdd gnd cell_6t
Xbit_r109_c124 bl[124] br[124] wl[109] vdd gnd cell_6t
Xbit_r110_c124 bl[124] br[124] wl[110] vdd gnd cell_6t
Xbit_r111_c124 bl[124] br[124] wl[111] vdd gnd cell_6t
Xbit_r112_c124 bl[124] br[124] wl[112] vdd gnd cell_6t
Xbit_r113_c124 bl[124] br[124] wl[113] vdd gnd cell_6t
Xbit_r114_c124 bl[124] br[124] wl[114] vdd gnd cell_6t
Xbit_r115_c124 bl[124] br[124] wl[115] vdd gnd cell_6t
Xbit_r116_c124 bl[124] br[124] wl[116] vdd gnd cell_6t
Xbit_r117_c124 bl[124] br[124] wl[117] vdd gnd cell_6t
Xbit_r118_c124 bl[124] br[124] wl[118] vdd gnd cell_6t
Xbit_r119_c124 bl[124] br[124] wl[119] vdd gnd cell_6t
Xbit_r120_c124 bl[124] br[124] wl[120] vdd gnd cell_6t
Xbit_r121_c124 bl[124] br[124] wl[121] vdd gnd cell_6t
Xbit_r122_c124 bl[124] br[124] wl[122] vdd gnd cell_6t
Xbit_r123_c124 bl[124] br[124] wl[123] vdd gnd cell_6t
Xbit_r124_c124 bl[124] br[124] wl[124] vdd gnd cell_6t
Xbit_r125_c124 bl[124] br[124] wl[125] vdd gnd cell_6t
Xbit_r126_c124 bl[124] br[124] wl[126] vdd gnd cell_6t
Xbit_r127_c124 bl[124] br[124] wl[127] vdd gnd cell_6t
Xbit_r128_c124 bl[124] br[124] wl[128] vdd gnd cell_6t
Xbit_r129_c124 bl[124] br[124] wl[129] vdd gnd cell_6t
Xbit_r130_c124 bl[124] br[124] wl[130] vdd gnd cell_6t
Xbit_r131_c124 bl[124] br[124] wl[131] vdd gnd cell_6t
Xbit_r132_c124 bl[124] br[124] wl[132] vdd gnd cell_6t
Xbit_r133_c124 bl[124] br[124] wl[133] vdd gnd cell_6t
Xbit_r134_c124 bl[124] br[124] wl[134] vdd gnd cell_6t
Xbit_r135_c124 bl[124] br[124] wl[135] vdd gnd cell_6t
Xbit_r136_c124 bl[124] br[124] wl[136] vdd gnd cell_6t
Xbit_r137_c124 bl[124] br[124] wl[137] vdd gnd cell_6t
Xbit_r138_c124 bl[124] br[124] wl[138] vdd gnd cell_6t
Xbit_r139_c124 bl[124] br[124] wl[139] vdd gnd cell_6t
Xbit_r140_c124 bl[124] br[124] wl[140] vdd gnd cell_6t
Xbit_r141_c124 bl[124] br[124] wl[141] vdd gnd cell_6t
Xbit_r142_c124 bl[124] br[124] wl[142] vdd gnd cell_6t
Xbit_r143_c124 bl[124] br[124] wl[143] vdd gnd cell_6t
Xbit_r144_c124 bl[124] br[124] wl[144] vdd gnd cell_6t
Xbit_r145_c124 bl[124] br[124] wl[145] vdd gnd cell_6t
Xbit_r146_c124 bl[124] br[124] wl[146] vdd gnd cell_6t
Xbit_r147_c124 bl[124] br[124] wl[147] vdd gnd cell_6t
Xbit_r148_c124 bl[124] br[124] wl[148] vdd gnd cell_6t
Xbit_r149_c124 bl[124] br[124] wl[149] vdd gnd cell_6t
Xbit_r150_c124 bl[124] br[124] wl[150] vdd gnd cell_6t
Xbit_r151_c124 bl[124] br[124] wl[151] vdd gnd cell_6t
Xbit_r152_c124 bl[124] br[124] wl[152] vdd gnd cell_6t
Xbit_r153_c124 bl[124] br[124] wl[153] vdd gnd cell_6t
Xbit_r154_c124 bl[124] br[124] wl[154] vdd gnd cell_6t
Xbit_r155_c124 bl[124] br[124] wl[155] vdd gnd cell_6t
Xbit_r156_c124 bl[124] br[124] wl[156] vdd gnd cell_6t
Xbit_r157_c124 bl[124] br[124] wl[157] vdd gnd cell_6t
Xbit_r158_c124 bl[124] br[124] wl[158] vdd gnd cell_6t
Xbit_r159_c124 bl[124] br[124] wl[159] vdd gnd cell_6t
Xbit_r160_c124 bl[124] br[124] wl[160] vdd gnd cell_6t
Xbit_r161_c124 bl[124] br[124] wl[161] vdd gnd cell_6t
Xbit_r162_c124 bl[124] br[124] wl[162] vdd gnd cell_6t
Xbit_r163_c124 bl[124] br[124] wl[163] vdd gnd cell_6t
Xbit_r164_c124 bl[124] br[124] wl[164] vdd gnd cell_6t
Xbit_r165_c124 bl[124] br[124] wl[165] vdd gnd cell_6t
Xbit_r166_c124 bl[124] br[124] wl[166] vdd gnd cell_6t
Xbit_r167_c124 bl[124] br[124] wl[167] vdd gnd cell_6t
Xbit_r168_c124 bl[124] br[124] wl[168] vdd gnd cell_6t
Xbit_r169_c124 bl[124] br[124] wl[169] vdd gnd cell_6t
Xbit_r170_c124 bl[124] br[124] wl[170] vdd gnd cell_6t
Xbit_r171_c124 bl[124] br[124] wl[171] vdd gnd cell_6t
Xbit_r172_c124 bl[124] br[124] wl[172] vdd gnd cell_6t
Xbit_r173_c124 bl[124] br[124] wl[173] vdd gnd cell_6t
Xbit_r174_c124 bl[124] br[124] wl[174] vdd gnd cell_6t
Xbit_r175_c124 bl[124] br[124] wl[175] vdd gnd cell_6t
Xbit_r176_c124 bl[124] br[124] wl[176] vdd gnd cell_6t
Xbit_r177_c124 bl[124] br[124] wl[177] vdd gnd cell_6t
Xbit_r178_c124 bl[124] br[124] wl[178] vdd gnd cell_6t
Xbit_r179_c124 bl[124] br[124] wl[179] vdd gnd cell_6t
Xbit_r180_c124 bl[124] br[124] wl[180] vdd gnd cell_6t
Xbit_r181_c124 bl[124] br[124] wl[181] vdd gnd cell_6t
Xbit_r182_c124 bl[124] br[124] wl[182] vdd gnd cell_6t
Xbit_r183_c124 bl[124] br[124] wl[183] vdd gnd cell_6t
Xbit_r184_c124 bl[124] br[124] wl[184] vdd gnd cell_6t
Xbit_r185_c124 bl[124] br[124] wl[185] vdd gnd cell_6t
Xbit_r186_c124 bl[124] br[124] wl[186] vdd gnd cell_6t
Xbit_r187_c124 bl[124] br[124] wl[187] vdd gnd cell_6t
Xbit_r188_c124 bl[124] br[124] wl[188] vdd gnd cell_6t
Xbit_r189_c124 bl[124] br[124] wl[189] vdd gnd cell_6t
Xbit_r190_c124 bl[124] br[124] wl[190] vdd gnd cell_6t
Xbit_r191_c124 bl[124] br[124] wl[191] vdd gnd cell_6t
Xbit_r192_c124 bl[124] br[124] wl[192] vdd gnd cell_6t
Xbit_r193_c124 bl[124] br[124] wl[193] vdd gnd cell_6t
Xbit_r194_c124 bl[124] br[124] wl[194] vdd gnd cell_6t
Xbit_r195_c124 bl[124] br[124] wl[195] vdd gnd cell_6t
Xbit_r196_c124 bl[124] br[124] wl[196] vdd gnd cell_6t
Xbit_r197_c124 bl[124] br[124] wl[197] vdd gnd cell_6t
Xbit_r198_c124 bl[124] br[124] wl[198] vdd gnd cell_6t
Xbit_r199_c124 bl[124] br[124] wl[199] vdd gnd cell_6t
Xbit_r200_c124 bl[124] br[124] wl[200] vdd gnd cell_6t
Xbit_r201_c124 bl[124] br[124] wl[201] vdd gnd cell_6t
Xbit_r202_c124 bl[124] br[124] wl[202] vdd gnd cell_6t
Xbit_r203_c124 bl[124] br[124] wl[203] vdd gnd cell_6t
Xbit_r204_c124 bl[124] br[124] wl[204] vdd gnd cell_6t
Xbit_r205_c124 bl[124] br[124] wl[205] vdd gnd cell_6t
Xbit_r206_c124 bl[124] br[124] wl[206] vdd gnd cell_6t
Xbit_r207_c124 bl[124] br[124] wl[207] vdd gnd cell_6t
Xbit_r208_c124 bl[124] br[124] wl[208] vdd gnd cell_6t
Xbit_r209_c124 bl[124] br[124] wl[209] vdd gnd cell_6t
Xbit_r210_c124 bl[124] br[124] wl[210] vdd gnd cell_6t
Xbit_r211_c124 bl[124] br[124] wl[211] vdd gnd cell_6t
Xbit_r212_c124 bl[124] br[124] wl[212] vdd gnd cell_6t
Xbit_r213_c124 bl[124] br[124] wl[213] vdd gnd cell_6t
Xbit_r214_c124 bl[124] br[124] wl[214] vdd gnd cell_6t
Xbit_r215_c124 bl[124] br[124] wl[215] vdd gnd cell_6t
Xbit_r216_c124 bl[124] br[124] wl[216] vdd gnd cell_6t
Xbit_r217_c124 bl[124] br[124] wl[217] vdd gnd cell_6t
Xbit_r218_c124 bl[124] br[124] wl[218] vdd gnd cell_6t
Xbit_r219_c124 bl[124] br[124] wl[219] vdd gnd cell_6t
Xbit_r220_c124 bl[124] br[124] wl[220] vdd gnd cell_6t
Xbit_r221_c124 bl[124] br[124] wl[221] vdd gnd cell_6t
Xbit_r222_c124 bl[124] br[124] wl[222] vdd gnd cell_6t
Xbit_r223_c124 bl[124] br[124] wl[223] vdd gnd cell_6t
Xbit_r224_c124 bl[124] br[124] wl[224] vdd gnd cell_6t
Xbit_r225_c124 bl[124] br[124] wl[225] vdd gnd cell_6t
Xbit_r226_c124 bl[124] br[124] wl[226] vdd gnd cell_6t
Xbit_r227_c124 bl[124] br[124] wl[227] vdd gnd cell_6t
Xbit_r228_c124 bl[124] br[124] wl[228] vdd gnd cell_6t
Xbit_r229_c124 bl[124] br[124] wl[229] vdd gnd cell_6t
Xbit_r230_c124 bl[124] br[124] wl[230] vdd gnd cell_6t
Xbit_r231_c124 bl[124] br[124] wl[231] vdd gnd cell_6t
Xbit_r232_c124 bl[124] br[124] wl[232] vdd gnd cell_6t
Xbit_r233_c124 bl[124] br[124] wl[233] vdd gnd cell_6t
Xbit_r234_c124 bl[124] br[124] wl[234] vdd gnd cell_6t
Xbit_r235_c124 bl[124] br[124] wl[235] vdd gnd cell_6t
Xbit_r236_c124 bl[124] br[124] wl[236] vdd gnd cell_6t
Xbit_r237_c124 bl[124] br[124] wl[237] vdd gnd cell_6t
Xbit_r238_c124 bl[124] br[124] wl[238] vdd gnd cell_6t
Xbit_r239_c124 bl[124] br[124] wl[239] vdd gnd cell_6t
Xbit_r240_c124 bl[124] br[124] wl[240] vdd gnd cell_6t
Xbit_r241_c124 bl[124] br[124] wl[241] vdd gnd cell_6t
Xbit_r242_c124 bl[124] br[124] wl[242] vdd gnd cell_6t
Xbit_r243_c124 bl[124] br[124] wl[243] vdd gnd cell_6t
Xbit_r244_c124 bl[124] br[124] wl[244] vdd gnd cell_6t
Xbit_r245_c124 bl[124] br[124] wl[245] vdd gnd cell_6t
Xbit_r246_c124 bl[124] br[124] wl[246] vdd gnd cell_6t
Xbit_r247_c124 bl[124] br[124] wl[247] vdd gnd cell_6t
Xbit_r248_c124 bl[124] br[124] wl[248] vdd gnd cell_6t
Xbit_r249_c124 bl[124] br[124] wl[249] vdd gnd cell_6t
Xbit_r250_c124 bl[124] br[124] wl[250] vdd gnd cell_6t
Xbit_r251_c124 bl[124] br[124] wl[251] vdd gnd cell_6t
Xbit_r252_c124 bl[124] br[124] wl[252] vdd gnd cell_6t
Xbit_r253_c124 bl[124] br[124] wl[253] vdd gnd cell_6t
Xbit_r254_c124 bl[124] br[124] wl[254] vdd gnd cell_6t
Xbit_r255_c124 bl[124] br[124] wl[255] vdd gnd cell_6t
Xbit_r0_c125 bl[125] br[125] wl[0] vdd gnd cell_6t
Xbit_r1_c125 bl[125] br[125] wl[1] vdd gnd cell_6t
Xbit_r2_c125 bl[125] br[125] wl[2] vdd gnd cell_6t
Xbit_r3_c125 bl[125] br[125] wl[3] vdd gnd cell_6t
Xbit_r4_c125 bl[125] br[125] wl[4] vdd gnd cell_6t
Xbit_r5_c125 bl[125] br[125] wl[5] vdd gnd cell_6t
Xbit_r6_c125 bl[125] br[125] wl[6] vdd gnd cell_6t
Xbit_r7_c125 bl[125] br[125] wl[7] vdd gnd cell_6t
Xbit_r8_c125 bl[125] br[125] wl[8] vdd gnd cell_6t
Xbit_r9_c125 bl[125] br[125] wl[9] vdd gnd cell_6t
Xbit_r10_c125 bl[125] br[125] wl[10] vdd gnd cell_6t
Xbit_r11_c125 bl[125] br[125] wl[11] vdd gnd cell_6t
Xbit_r12_c125 bl[125] br[125] wl[12] vdd gnd cell_6t
Xbit_r13_c125 bl[125] br[125] wl[13] vdd gnd cell_6t
Xbit_r14_c125 bl[125] br[125] wl[14] vdd gnd cell_6t
Xbit_r15_c125 bl[125] br[125] wl[15] vdd gnd cell_6t
Xbit_r16_c125 bl[125] br[125] wl[16] vdd gnd cell_6t
Xbit_r17_c125 bl[125] br[125] wl[17] vdd gnd cell_6t
Xbit_r18_c125 bl[125] br[125] wl[18] vdd gnd cell_6t
Xbit_r19_c125 bl[125] br[125] wl[19] vdd gnd cell_6t
Xbit_r20_c125 bl[125] br[125] wl[20] vdd gnd cell_6t
Xbit_r21_c125 bl[125] br[125] wl[21] vdd gnd cell_6t
Xbit_r22_c125 bl[125] br[125] wl[22] vdd gnd cell_6t
Xbit_r23_c125 bl[125] br[125] wl[23] vdd gnd cell_6t
Xbit_r24_c125 bl[125] br[125] wl[24] vdd gnd cell_6t
Xbit_r25_c125 bl[125] br[125] wl[25] vdd gnd cell_6t
Xbit_r26_c125 bl[125] br[125] wl[26] vdd gnd cell_6t
Xbit_r27_c125 bl[125] br[125] wl[27] vdd gnd cell_6t
Xbit_r28_c125 bl[125] br[125] wl[28] vdd gnd cell_6t
Xbit_r29_c125 bl[125] br[125] wl[29] vdd gnd cell_6t
Xbit_r30_c125 bl[125] br[125] wl[30] vdd gnd cell_6t
Xbit_r31_c125 bl[125] br[125] wl[31] vdd gnd cell_6t
Xbit_r32_c125 bl[125] br[125] wl[32] vdd gnd cell_6t
Xbit_r33_c125 bl[125] br[125] wl[33] vdd gnd cell_6t
Xbit_r34_c125 bl[125] br[125] wl[34] vdd gnd cell_6t
Xbit_r35_c125 bl[125] br[125] wl[35] vdd gnd cell_6t
Xbit_r36_c125 bl[125] br[125] wl[36] vdd gnd cell_6t
Xbit_r37_c125 bl[125] br[125] wl[37] vdd gnd cell_6t
Xbit_r38_c125 bl[125] br[125] wl[38] vdd gnd cell_6t
Xbit_r39_c125 bl[125] br[125] wl[39] vdd gnd cell_6t
Xbit_r40_c125 bl[125] br[125] wl[40] vdd gnd cell_6t
Xbit_r41_c125 bl[125] br[125] wl[41] vdd gnd cell_6t
Xbit_r42_c125 bl[125] br[125] wl[42] vdd gnd cell_6t
Xbit_r43_c125 bl[125] br[125] wl[43] vdd gnd cell_6t
Xbit_r44_c125 bl[125] br[125] wl[44] vdd gnd cell_6t
Xbit_r45_c125 bl[125] br[125] wl[45] vdd gnd cell_6t
Xbit_r46_c125 bl[125] br[125] wl[46] vdd gnd cell_6t
Xbit_r47_c125 bl[125] br[125] wl[47] vdd gnd cell_6t
Xbit_r48_c125 bl[125] br[125] wl[48] vdd gnd cell_6t
Xbit_r49_c125 bl[125] br[125] wl[49] vdd gnd cell_6t
Xbit_r50_c125 bl[125] br[125] wl[50] vdd gnd cell_6t
Xbit_r51_c125 bl[125] br[125] wl[51] vdd gnd cell_6t
Xbit_r52_c125 bl[125] br[125] wl[52] vdd gnd cell_6t
Xbit_r53_c125 bl[125] br[125] wl[53] vdd gnd cell_6t
Xbit_r54_c125 bl[125] br[125] wl[54] vdd gnd cell_6t
Xbit_r55_c125 bl[125] br[125] wl[55] vdd gnd cell_6t
Xbit_r56_c125 bl[125] br[125] wl[56] vdd gnd cell_6t
Xbit_r57_c125 bl[125] br[125] wl[57] vdd gnd cell_6t
Xbit_r58_c125 bl[125] br[125] wl[58] vdd gnd cell_6t
Xbit_r59_c125 bl[125] br[125] wl[59] vdd gnd cell_6t
Xbit_r60_c125 bl[125] br[125] wl[60] vdd gnd cell_6t
Xbit_r61_c125 bl[125] br[125] wl[61] vdd gnd cell_6t
Xbit_r62_c125 bl[125] br[125] wl[62] vdd gnd cell_6t
Xbit_r63_c125 bl[125] br[125] wl[63] vdd gnd cell_6t
Xbit_r64_c125 bl[125] br[125] wl[64] vdd gnd cell_6t
Xbit_r65_c125 bl[125] br[125] wl[65] vdd gnd cell_6t
Xbit_r66_c125 bl[125] br[125] wl[66] vdd gnd cell_6t
Xbit_r67_c125 bl[125] br[125] wl[67] vdd gnd cell_6t
Xbit_r68_c125 bl[125] br[125] wl[68] vdd gnd cell_6t
Xbit_r69_c125 bl[125] br[125] wl[69] vdd gnd cell_6t
Xbit_r70_c125 bl[125] br[125] wl[70] vdd gnd cell_6t
Xbit_r71_c125 bl[125] br[125] wl[71] vdd gnd cell_6t
Xbit_r72_c125 bl[125] br[125] wl[72] vdd gnd cell_6t
Xbit_r73_c125 bl[125] br[125] wl[73] vdd gnd cell_6t
Xbit_r74_c125 bl[125] br[125] wl[74] vdd gnd cell_6t
Xbit_r75_c125 bl[125] br[125] wl[75] vdd gnd cell_6t
Xbit_r76_c125 bl[125] br[125] wl[76] vdd gnd cell_6t
Xbit_r77_c125 bl[125] br[125] wl[77] vdd gnd cell_6t
Xbit_r78_c125 bl[125] br[125] wl[78] vdd gnd cell_6t
Xbit_r79_c125 bl[125] br[125] wl[79] vdd gnd cell_6t
Xbit_r80_c125 bl[125] br[125] wl[80] vdd gnd cell_6t
Xbit_r81_c125 bl[125] br[125] wl[81] vdd gnd cell_6t
Xbit_r82_c125 bl[125] br[125] wl[82] vdd gnd cell_6t
Xbit_r83_c125 bl[125] br[125] wl[83] vdd gnd cell_6t
Xbit_r84_c125 bl[125] br[125] wl[84] vdd gnd cell_6t
Xbit_r85_c125 bl[125] br[125] wl[85] vdd gnd cell_6t
Xbit_r86_c125 bl[125] br[125] wl[86] vdd gnd cell_6t
Xbit_r87_c125 bl[125] br[125] wl[87] vdd gnd cell_6t
Xbit_r88_c125 bl[125] br[125] wl[88] vdd gnd cell_6t
Xbit_r89_c125 bl[125] br[125] wl[89] vdd gnd cell_6t
Xbit_r90_c125 bl[125] br[125] wl[90] vdd gnd cell_6t
Xbit_r91_c125 bl[125] br[125] wl[91] vdd gnd cell_6t
Xbit_r92_c125 bl[125] br[125] wl[92] vdd gnd cell_6t
Xbit_r93_c125 bl[125] br[125] wl[93] vdd gnd cell_6t
Xbit_r94_c125 bl[125] br[125] wl[94] vdd gnd cell_6t
Xbit_r95_c125 bl[125] br[125] wl[95] vdd gnd cell_6t
Xbit_r96_c125 bl[125] br[125] wl[96] vdd gnd cell_6t
Xbit_r97_c125 bl[125] br[125] wl[97] vdd gnd cell_6t
Xbit_r98_c125 bl[125] br[125] wl[98] vdd gnd cell_6t
Xbit_r99_c125 bl[125] br[125] wl[99] vdd gnd cell_6t
Xbit_r100_c125 bl[125] br[125] wl[100] vdd gnd cell_6t
Xbit_r101_c125 bl[125] br[125] wl[101] vdd gnd cell_6t
Xbit_r102_c125 bl[125] br[125] wl[102] vdd gnd cell_6t
Xbit_r103_c125 bl[125] br[125] wl[103] vdd gnd cell_6t
Xbit_r104_c125 bl[125] br[125] wl[104] vdd gnd cell_6t
Xbit_r105_c125 bl[125] br[125] wl[105] vdd gnd cell_6t
Xbit_r106_c125 bl[125] br[125] wl[106] vdd gnd cell_6t
Xbit_r107_c125 bl[125] br[125] wl[107] vdd gnd cell_6t
Xbit_r108_c125 bl[125] br[125] wl[108] vdd gnd cell_6t
Xbit_r109_c125 bl[125] br[125] wl[109] vdd gnd cell_6t
Xbit_r110_c125 bl[125] br[125] wl[110] vdd gnd cell_6t
Xbit_r111_c125 bl[125] br[125] wl[111] vdd gnd cell_6t
Xbit_r112_c125 bl[125] br[125] wl[112] vdd gnd cell_6t
Xbit_r113_c125 bl[125] br[125] wl[113] vdd gnd cell_6t
Xbit_r114_c125 bl[125] br[125] wl[114] vdd gnd cell_6t
Xbit_r115_c125 bl[125] br[125] wl[115] vdd gnd cell_6t
Xbit_r116_c125 bl[125] br[125] wl[116] vdd gnd cell_6t
Xbit_r117_c125 bl[125] br[125] wl[117] vdd gnd cell_6t
Xbit_r118_c125 bl[125] br[125] wl[118] vdd gnd cell_6t
Xbit_r119_c125 bl[125] br[125] wl[119] vdd gnd cell_6t
Xbit_r120_c125 bl[125] br[125] wl[120] vdd gnd cell_6t
Xbit_r121_c125 bl[125] br[125] wl[121] vdd gnd cell_6t
Xbit_r122_c125 bl[125] br[125] wl[122] vdd gnd cell_6t
Xbit_r123_c125 bl[125] br[125] wl[123] vdd gnd cell_6t
Xbit_r124_c125 bl[125] br[125] wl[124] vdd gnd cell_6t
Xbit_r125_c125 bl[125] br[125] wl[125] vdd gnd cell_6t
Xbit_r126_c125 bl[125] br[125] wl[126] vdd gnd cell_6t
Xbit_r127_c125 bl[125] br[125] wl[127] vdd gnd cell_6t
Xbit_r128_c125 bl[125] br[125] wl[128] vdd gnd cell_6t
Xbit_r129_c125 bl[125] br[125] wl[129] vdd gnd cell_6t
Xbit_r130_c125 bl[125] br[125] wl[130] vdd gnd cell_6t
Xbit_r131_c125 bl[125] br[125] wl[131] vdd gnd cell_6t
Xbit_r132_c125 bl[125] br[125] wl[132] vdd gnd cell_6t
Xbit_r133_c125 bl[125] br[125] wl[133] vdd gnd cell_6t
Xbit_r134_c125 bl[125] br[125] wl[134] vdd gnd cell_6t
Xbit_r135_c125 bl[125] br[125] wl[135] vdd gnd cell_6t
Xbit_r136_c125 bl[125] br[125] wl[136] vdd gnd cell_6t
Xbit_r137_c125 bl[125] br[125] wl[137] vdd gnd cell_6t
Xbit_r138_c125 bl[125] br[125] wl[138] vdd gnd cell_6t
Xbit_r139_c125 bl[125] br[125] wl[139] vdd gnd cell_6t
Xbit_r140_c125 bl[125] br[125] wl[140] vdd gnd cell_6t
Xbit_r141_c125 bl[125] br[125] wl[141] vdd gnd cell_6t
Xbit_r142_c125 bl[125] br[125] wl[142] vdd gnd cell_6t
Xbit_r143_c125 bl[125] br[125] wl[143] vdd gnd cell_6t
Xbit_r144_c125 bl[125] br[125] wl[144] vdd gnd cell_6t
Xbit_r145_c125 bl[125] br[125] wl[145] vdd gnd cell_6t
Xbit_r146_c125 bl[125] br[125] wl[146] vdd gnd cell_6t
Xbit_r147_c125 bl[125] br[125] wl[147] vdd gnd cell_6t
Xbit_r148_c125 bl[125] br[125] wl[148] vdd gnd cell_6t
Xbit_r149_c125 bl[125] br[125] wl[149] vdd gnd cell_6t
Xbit_r150_c125 bl[125] br[125] wl[150] vdd gnd cell_6t
Xbit_r151_c125 bl[125] br[125] wl[151] vdd gnd cell_6t
Xbit_r152_c125 bl[125] br[125] wl[152] vdd gnd cell_6t
Xbit_r153_c125 bl[125] br[125] wl[153] vdd gnd cell_6t
Xbit_r154_c125 bl[125] br[125] wl[154] vdd gnd cell_6t
Xbit_r155_c125 bl[125] br[125] wl[155] vdd gnd cell_6t
Xbit_r156_c125 bl[125] br[125] wl[156] vdd gnd cell_6t
Xbit_r157_c125 bl[125] br[125] wl[157] vdd gnd cell_6t
Xbit_r158_c125 bl[125] br[125] wl[158] vdd gnd cell_6t
Xbit_r159_c125 bl[125] br[125] wl[159] vdd gnd cell_6t
Xbit_r160_c125 bl[125] br[125] wl[160] vdd gnd cell_6t
Xbit_r161_c125 bl[125] br[125] wl[161] vdd gnd cell_6t
Xbit_r162_c125 bl[125] br[125] wl[162] vdd gnd cell_6t
Xbit_r163_c125 bl[125] br[125] wl[163] vdd gnd cell_6t
Xbit_r164_c125 bl[125] br[125] wl[164] vdd gnd cell_6t
Xbit_r165_c125 bl[125] br[125] wl[165] vdd gnd cell_6t
Xbit_r166_c125 bl[125] br[125] wl[166] vdd gnd cell_6t
Xbit_r167_c125 bl[125] br[125] wl[167] vdd gnd cell_6t
Xbit_r168_c125 bl[125] br[125] wl[168] vdd gnd cell_6t
Xbit_r169_c125 bl[125] br[125] wl[169] vdd gnd cell_6t
Xbit_r170_c125 bl[125] br[125] wl[170] vdd gnd cell_6t
Xbit_r171_c125 bl[125] br[125] wl[171] vdd gnd cell_6t
Xbit_r172_c125 bl[125] br[125] wl[172] vdd gnd cell_6t
Xbit_r173_c125 bl[125] br[125] wl[173] vdd gnd cell_6t
Xbit_r174_c125 bl[125] br[125] wl[174] vdd gnd cell_6t
Xbit_r175_c125 bl[125] br[125] wl[175] vdd gnd cell_6t
Xbit_r176_c125 bl[125] br[125] wl[176] vdd gnd cell_6t
Xbit_r177_c125 bl[125] br[125] wl[177] vdd gnd cell_6t
Xbit_r178_c125 bl[125] br[125] wl[178] vdd gnd cell_6t
Xbit_r179_c125 bl[125] br[125] wl[179] vdd gnd cell_6t
Xbit_r180_c125 bl[125] br[125] wl[180] vdd gnd cell_6t
Xbit_r181_c125 bl[125] br[125] wl[181] vdd gnd cell_6t
Xbit_r182_c125 bl[125] br[125] wl[182] vdd gnd cell_6t
Xbit_r183_c125 bl[125] br[125] wl[183] vdd gnd cell_6t
Xbit_r184_c125 bl[125] br[125] wl[184] vdd gnd cell_6t
Xbit_r185_c125 bl[125] br[125] wl[185] vdd gnd cell_6t
Xbit_r186_c125 bl[125] br[125] wl[186] vdd gnd cell_6t
Xbit_r187_c125 bl[125] br[125] wl[187] vdd gnd cell_6t
Xbit_r188_c125 bl[125] br[125] wl[188] vdd gnd cell_6t
Xbit_r189_c125 bl[125] br[125] wl[189] vdd gnd cell_6t
Xbit_r190_c125 bl[125] br[125] wl[190] vdd gnd cell_6t
Xbit_r191_c125 bl[125] br[125] wl[191] vdd gnd cell_6t
Xbit_r192_c125 bl[125] br[125] wl[192] vdd gnd cell_6t
Xbit_r193_c125 bl[125] br[125] wl[193] vdd gnd cell_6t
Xbit_r194_c125 bl[125] br[125] wl[194] vdd gnd cell_6t
Xbit_r195_c125 bl[125] br[125] wl[195] vdd gnd cell_6t
Xbit_r196_c125 bl[125] br[125] wl[196] vdd gnd cell_6t
Xbit_r197_c125 bl[125] br[125] wl[197] vdd gnd cell_6t
Xbit_r198_c125 bl[125] br[125] wl[198] vdd gnd cell_6t
Xbit_r199_c125 bl[125] br[125] wl[199] vdd gnd cell_6t
Xbit_r200_c125 bl[125] br[125] wl[200] vdd gnd cell_6t
Xbit_r201_c125 bl[125] br[125] wl[201] vdd gnd cell_6t
Xbit_r202_c125 bl[125] br[125] wl[202] vdd gnd cell_6t
Xbit_r203_c125 bl[125] br[125] wl[203] vdd gnd cell_6t
Xbit_r204_c125 bl[125] br[125] wl[204] vdd gnd cell_6t
Xbit_r205_c125 bl[125] br[125] wl[205] vdd gnd cell_6t
Xbit_r206_c125 bl[125] br[125] wl[206] vdd gnd cell_6t
Xbit_r207_c125 bl[125] br[125] wl[207] vdd gnd cell_6t
Xbit_r208_c125 bl[125] br[125] wl[208] vdd gnd cell_6t
Xbit_r209_c125 bl[125] br[125] wl[209] vdd gnd cell_6t
Xbit_r210_c125 bl[125] br[125] wl[210] vdd gnd cell_6t
Xbit_r211_c125 bl[125] br[125] wl[211] vdd gnd cell_6t
Xbit_r212_c125 bl[125] br[125] wl[212] vdd gnd cell_6t
Xbit_r213_c125 bl[125] br[125] wl[213] vdd gnd cell_6t
Xbit_r214_c125 bl[125] br[125] wl[214] vdd gnd cell_6t
Xbit_r215_c125 bl[125] br[125] wl[215] vdd gnd cell_6t
Xbit_r216_c125 bl[125] br[125] wl[216] vdd gnd cell_6t
Xbit_r217_c125 bl[125] br[125] wl[217] vdd gnd cell_6t
Xbit_r218_c125 bl[125] br[125] wl[218] vdd gnd cell_6t
Xbit_r219_c125 bl[125] br[125] wl[219] vdd gnd cell_6t
Xbit_r220_c125 bl[125] br[125] wl[220] vdd gnd cell_6t
Xbit_r221_c125 bl[125] br[125] wl[221] vdd gnd cell_6t
Xbit_r222_c125 bl[125] br[125] wl[222] vdd gnd cell_6t
Xbit_r223_c125 bl[125] br[125] wl[223] vdd gnd cell_6t
Xbit_r224_c125 bl[125] br[125] wl[224] vdd gnd cell_6t
Xbit_r225_c125 bl[125] br[125] wl[225] vdd gnd cell_6t
Xbit_r226_c125 bl[125] br[125] wl[226] vdd gnd cell_6t
Xbit_r227_c125 bl[125] br[125] wl[227] vdd gnd cell_6t
Xbit_r228_c125 bl[125] br[125] wl[228] vdd gnd cell_6t
Xbit_r229_c125 bl[125] br[125] wl[229] vdd gnd cell_6t
Xbit_r230_c125 bl[125] br[125] wl[230] vdd gnd cell_6t
Xbit_r231_c125 bl[125] br[125] wl[231] vdd gnd cell_6t
Xbit_r232_c125 bl[125] br[125] wl[232] vdd gnd cell_6t
Xbit_r233_c125 bl[125] br[125] wl[233] vdd gnd cell_6t
Xbit_r234_c125 bl[125] br[125] wl[234] vdd gnd cell_6t
Xbit_r235_c125 bl[125] br[125] wl[235] vdd gnd cell_6t
Xbit_r236_c125 bl[125] br[125] wl[236] vdd gnd cell_6t
Xbit_r237_c125 bl[125] br[125] wl[237] vdd gnd cell_6t
Xbit_r238_c125 bl[125] br[125] wl[238] vdd gnd cell_6t
Xbit_r239_c125 bl[125] br[125] wl[239] vdd gnd cell_6t
Xbit_r240_c125 bl[125] br[125] wl[240] vdd gnd cell_6t
Xbit_r241_c125 bl[125] br[125] wl[241] vdd gnd cell_6t
Xbit_r242_c125 bl[125] br[125] wl[242] vdd gnd cell_6t
Xbit_r243_c125 bl[125] br[125] wl[243] vdd gnd cell_6t
Xbit_r244_c125 bl[125] br[125] wl[244] vdd gnd cell_6t
Xbit_r245_c125 bl[125] br[125] wl[245] vdd gnd cell_6t
Xbit_r246_c125 bl[125] br[125] wl[246] vdd gnd cell_6t
Xbit_r247_c125 bl[125] br[125] wl[247] vdd gnd cell_6t
Xbit_r248_c125 bl[125] br[125] wl[248] vdd gnd cell_6t
Xbit_r249_c125 bl[125] br[125] wl[249] vdd gnd cell_6t
Xbit_r250_c125 bl[125] br[125] wl[250] vdd gnd cell_6t
Xbit_r251_c125 bl[125] br[125] wl[251] vdd gnd cell_6t
Xbit_r252_c125 bl[125] br[125] wl[252] vdd gnd cell_6t
Xbit_r253_c125 bl[125] br[125] wl[253] vdd gnd cell_6t
Xbit_r254_c125 bl[125] br[125] wl[254] vdd gnd cell_6t
Xbit_r255_c125 bl[125] br[125] wl[255] vdd gnd cell_6t
Xbit_r0_c126 bl[126] br[126] wl[0] vdd gnd cell_6t
Xbit_r1_c126 bl[126] br[126] wl[1] vdd gnd cell_6t
Xbit_r2_c126 bl[126] br[126] wl[2] vdd gnd cell_6t
Xbit_r3_c126 bl[126] br[126] wl[3] vdd gnd cell_6t
Xbit_r4_c126 bl[126] br[126] wl[4] vdd gnd cell_6t
Xbit_r5_c126 bl[126] br[126] wl[5] vdd gnd cell_6t
Xbit_r6_c126 bl[126] br[126] wl[6] vdd gnd cell_6t
Xbit_r7_c126 bl[126] br[126] wl[7] vdd gnd cell_6t
Xbit_r8_c126 bl[126] br[126] wl[8] vdd gnd cell_6t
Xbit_r9_c126 bl[126] br[126] wl[9] vdd gnd cell_6t
Xbit_r10_c126 bl[126] br[126] wl[10] vdd gnd cell_6t
Xbit_r11_c126 bl[126] br[126] wl[11] vdd gnd cell_6t
Xbit_r12_c126 bl[126] br[126] wl[12] vdd gnd cell_6t
Xbit_r13_c126 bl[126] br[126] wl[13] vdd gnd cell_6t
Xbit_r14_c126 bl[126] br[126] wl[14] vdd gnd cell_6t
Xbit_r15_c126 bl[126] br[126] wl[15] vdd gnd cell_6t
Xbit_r16_c126 bl[126] br[126] wl[16] vdd gnd cell_6t
Xbit_r17_c126 bl[126] br[126] wl[17] vdd gnd cell_6t
Xbit_r18_c126 bl[126] br[126] wl[18] vdd gnd cell_6t
Xbit_r19_c126 bl[126] br[126] wl[19] vdd gnd cell_6t
Xbit_r20_c126 bl[126] br[126] wl[20] vdd gnd cell_6t
Xbit_r21_c126 bl[126] br[126] wl[21] vdd gnd cell_6t
Xbit_r22_c126 bl[126] br[126] wl[22] vdd gnd cell_6t
Xbit_r23_c126 bl[126] br[126] wl[23] vdd gnd cell_6t
Xbit_r24_c126 bl[126] br[126] wl[24] vdd gnd cell_6t
Xbit_r25_c126 bl[126] br[126] wl[25] vdd gnd cell_6t
Xbit_r26_c126 bl[126] br[126] wl[26] vdd gnd cell_6t
Xbit_r27_c126 bl[126] br[126] wl[27] vdd gnd cell_6t
Xbit_r28_c126 bl[126] br[126] wl[28] vdd gnd cell_6t
Xbit_r29_c126 bl[126] br[126] wl[29] vdd gnd cell_6t
Xbit_r30_c126 bl[126] br[126] wl[30] vdd gnd cell_6t
Xbit_r31_c126 bl[126] br[126] wl[31] vdd gnd cell_6t
Xbit_r32_c126 bl[126] br[126] wl[32] vdd gnd cell_6t
Xbit_r33_c126 bl[126] br[126] wl[33] vdd gnd cell_6t
Xbit_r34_c126 bl[126] br[126] wl[34] vdd gnd cell_6t
Xbit_r35_c126 bl[126] br[126] wl[35] vdd gnd cell_6t
Xbit_r36_c126 bl[126] br[126] wl[36] vdd gnd cell_6t
Xbit_r37_c126 bl[126] br[126] wl[37] vdd gnd cell_6t
Xbit_r38_c126 bl[126] br[126] wl[38] vdd gnd cell_6t
Xbit_r39_c126 bl[126] br[126] wl[39] vdd gnd cell_6t
Xbit_r40_c126 bl[126] br[126] wl[40] vdd gnd cell_6t
Xbit_r41_c126 bl[126] br[126] wl[41] vdd gnd cell_6t
Xbit_r42_c126 bl[126] br[126] wl[42] vdd gnd cell_6t
Xbit_r43_c126 bl[126] br[126] wl[43] vdd gnd cell_6t
Xbit_r44_c126 bl[126] br[126] wl[44] vdd gnd cell_6t
Xbit_r45_c126 bl[126] br[126] wl[45] vdd gnd cell_6t
Xbit_r46_c126 bl[126] br[126] wl[46] vdd gnd cell_6t
Xbit_r47_c126 bl[126] br[126] wl[47] vdd gnd cell_6t
Xbit_r48_c126 bl[126] br[126] wl[48] vdd gnd cell_6t
Xbit_r49_c126 bl[126] br[126] wl[49] vdd gnd cell_6t
Xbit_r50_c126 bl[126] br[126] wl[50] vdd gnd cell_6t
Xbit_r51_c126 bl[126] br[126] wl[51] vdd gnd cell_6t
Xbit_r52_c126 bl[126] br[126] wl[52] vdd gnd cell_6t
Xbit_r53_c126 bl[126] br[126] wl[53] vdd gnd cell_6t
Xbit_r54_c126 bl[126] br[126] wl[54] vdd gnd cell_6t
Xbit_r55_c126 bl[126] br[126] wl[55] vdd gnd cell_6t
Xbit_r56_c126 bl[126] br[126] wl[56] vdd gnd cell_6t
Xbit_r57_c126 bl[126] br[126] wl[57] vdd gnd cell_6t
Xbit_r58_c126 bl[126] br[126] wl[58] vdd gnd cell_6t
Xbit_r59_c126 bl[126] br[126] wl[59] vdd gnd cell_6t
Xbit_r60_c126 bl[126] br[126] wl[60] vdd gnd cell_6t
Xbit_r61_c126 bl[126] br[126] wl[61] vdd gnd cell_6t
Xbit_r62_c126 bl[126] br[126] wl[62] vdd gnd cell_6t
Xbit_r63_c126 bl[126] br[126] wl[63] vdd gnd cell_6t
Xbit_r64_c126 bl[126] br[126] wl[64] vdd gnd cell_6t
Xbit_r65_c126 bl[126] br[126] wl[65] vdd gnd cell_6t
Xbit_r66_c126 bl[126] br[126] wl[66] vdd gnd cell_6t
Xbit_r67_c126 bl[126] br[126] wl[67] vdd gnd cell_6t
Xbit_r68_c126 bl[126] br[126] wl[68] vdd gnd cell_6t
Xbit_r69_c126 bl[126] br[126] wl[69] vdd gnd cell_6t
Xbit_r70_c126 bl[126] br[126] wl[70] vdd gnd cell_6t
Xbit_r71_c126 bl[126] br[126] wl[71] vdd gnd cell_6t
Xbit_r72_c126 bl[126] br[126] wl[72] vdd gnd cell_6t
Xbit_r73_c126 bl[126] br[126] wl[73] vdd gnd cell_6t
Xbit_r74_c126 bl[126] br[126] wl[74] vdd gnd cell_6t
Xbit_r75_c126 bl[126] br[126] wl[75] vdd gnd cell_6t
Xbit_r76_c126 bl[126] br[126] wl[76] vdd gnd cell_6t
Xbit_r77_c126 bl[126] br[126] wl[77] vdd gnd cell_6t
Xbit_r78_c126 bl[126] br[126] wl[78] vdd gnd cell_6t
Xbit_r79_c126 bl[126] br[126] wl[79] vdd gnd cell_6t
Xbit_r80_c126 bl[126] br[126] wl[80] vdd gnd cell_6t
Xbit_r81_c126 bl[126] br[126] wl[81] vdd gnd cell_6t
Xbit_r82_c126 bl[126] br[126] wl[82] vdd gnd cell_6t
Xbit_r83_c126 bl[126] br[126] wl[83] vdd gnd cell_6t
Xbit_r84_c126 bl[126] br[126] wl[84] vdd gnd cell_6t
Xbit_r85_c126 bl[126] br[126] wl[85] vdd gnd cell_6t
Xbit_r86_c126 bl[126] br[126] wl[86] vdd gnd cell_6t
Xbit_r87_c126 bl[126] br[126] wl[87] vdd gnd cell_6t
Xbit_r88_c126 bl[126] br[126] wl[88] vdd gnd cell_6t
Xbit_r89_c126 bl[126] br[126] wl[89] vdd gnd cell_6t
Xbit_r90_c126 bl[126] br[126] wl[90] vdd gnd cell_6t
Xbit_r91_c126 bl[126] br[126] wl[91] vdd gnd cell_6t
Xbit_r92_c126 bl[126] br[126] wl[92] vdd gnd cell_6t
Xbit_r93_c126 bl[126] br[126] wl[93] vdd gnd cell_6t
Xbit_r94_c126 bl[126] br[126] wl[94] vdd gnd cell_6t
Xbit_r95_c126 bl[126] br[126] wl[95] vdd gnd cell_6t
Xbit_r96_c126 bl[126] br[126] wl[96] vdd gnd cell_6t
Xbit_r97_c126 bl[126] br[126] wl[97] vdd gnd cell_6t
Xbit_r98_c126 bl[126] br[126] wl[98] vdd gnd cell_6t
Xbit_r99_c126 bl[126] br[126] wl[99] vdd gnd cell_6t
Xbit_r100_c126 bl[126] br[126] wl[100] vdd gnd cell_6t
Xbit_r101_c126 bl[126] br[126] wl[101] vdd gnd cell_6t
Xbit_r102_c126 bl[126] br[126] wl[102] vdd gnd cell_6t
Xbit_r103_c126 bl[126] br[126] wl[103] vdd gnd cell_6t
Xbit_r104_c126 bl[126] br[126] wl[104] vdd gnd cell_6t
Xbit_r105_c126 bl[126] br[126] wl[105] vdd gnd cell_6t
Xbit_r106_c126 bl[126] br[126] wl[106] vdd gnd cell_6t
Xbit_r107_c126 bl[126] br[126] wl[107] vdd gnd cell_6t
Xbit_r108_c126 bl[126] br[126] wl[108] vdd gnd cell_6t
Xbit_r109_c126 bl[126] br[126] wl[109] vdd gnd cell_6t
Xbit_r110_c126 bl[126] br[126] wl[110] vdd gnd cell_6t
Xbit_r111_c126 bl[126] br[126] wl[111] vdd gnd cell_6t
Xbit_r112_c126 bl[126] br[126] wl[112] vdd gnd cell_6t
Xbit_r113_c126 bl[126] br[126] wl[113] vdd gnd cell_6t
Xbit_r114_c126 bl[126] br[126] wl[114] vdd gnd cell_6t
Xbit_r115_c126 bl[126] br[126] wl[115] vdd gnd cell_6t
Xbit_r116_c126 bl[126] br[126] wl[116] vdd gnd cell_6t
Xbit_r117_c126 bl[126] br[126] wl[117] vdd gnd cell_6t
Xbit_r118_c126 bl[126] br[126] wl[118] vdd gnd cell_6t
Xbit_r119_c126 bl[126] br[126] wl[119] vdd gnd cell_6t
Xbit_r120_c126 bl[126] br[126] wl[120] vdd gnd cell_6t
Xbit_r121_c126 bl[126] br[126] wl[121] vdd gnd cell_6t
Xbit_r122_c126 bl[126] br[126] wl[122] vdd gnd cell_6t
Xbit_r123_c126 bl[126] br[126] wl[123] vdd gnd cell_6t
Xbit_r124_c126 bl[126] br[126] wl[124] vdd gnd cell_6t
Xbit_r125_c126 bl[126] br[126] wl[125] vdd gnd cell_6t
Xbit_r126_c126 bl[126] br[126] wl[126] vdd gnd cell_6t
Xbit_r127_c126 bl[126] br[126] wl[127] vdd gnd cell_6t
Xbit_r128_c126 bl[126] br[126] wl[128] vdd gnd cell_6t
Xbit_r129_c126 bl[126] br[126] wl[129] vdd gnd cell_6t
Xbit_r130_c126 bl[126] br[126] wl[130] vdd gnd cell_6t
Xbit_r131_c126 bl[126] br[126] wl[131] vdd gnd cell_6t
Xbit_r132_c126 bl[126] br[126] wl[132] vdd gnd cell_6t
Xbit_r133_c126 bl[126] br[126] wl[133] vdd gnd cell_6t
Xbit_r134_c126 bl[126] br[126] wl[134] vdd gnd cell_6t
Xbit_r135_c126 bl[126] br[126] wl[135] vdd gnd cell_6t
Xbit_r136_c126 bl[126] br[126] wl[136] vdd gnd cell_6t
Xbit_r137_c126 bl[126] br[126] wl[137] vdd gnd cell_6t
Xbit_r138_c126 bl[126] br[126] wl[138] vdd gnd cell_6t
Xbit_r139_c126 bl[126] br[126] wl[139] vdd gnd cell_6t
Xbit_r140_c126 bl[126] br[126] wl[140] vdd gnd cell_6t
Xbit_r141_c126 bl[126] br[126] wl[141] vdd gnd cell_6t
Xbit_r142_c126 bl[126] br[126] wl[142] vdd gnd cell_6t
Xbit_r143_c126 bl[126] br[126] wl[143] vdd gnd cell_6t
Xbit_r144_c126 bl[126] br[126] wl[144] vdd gnd cell_6t
Xbit_r145_c126 bl[126] br[126] wl[145] vdd gnd cell_6t
Xbit_r146_c126 bl[126] br[126] wl[146] vdd gnd cell_6t
Xbit_r147_c126 bl[126] br[126] wl[147] vdd gnd cell_6t
Xbit_r148_c126 bl[126] br[126] wl[148] vdd gnd cell_6t
Xbit_r149_c126 bl[126] br[126] wl[149] vdd gnd cell_6t
Xbit_r150_c126 bl[126] br[126] wl[150] vdd gnd cell_6t
Xbit_r151_c126 bl[126] br[126] wl[151] vdd gnd cell_6t
Xbit_r152_c126 bl[126] br[126] wl[152] vdd gnd cell_6t
Xbit_r153_c126 bl[126] br[126] wl[153] vdd gnd cell_6t
Xbit_r154_c126 bl[126] br[126] wl[154] vdd gnd cell_6t
Xbit_r155_c126 bl[126] br[126] wl[155] vdd gnd cell_6t
Xbit_r156_c126 bl[126] br[126] wl[156] vdd gnd cell_6t
Xbit_r157_c126 bl[126] br[126] wl[157] vdd gnd cell_6t
Xbit_r158_c126 bl[126] br[126] wl[158] vdd gnd cell_6t
Xbit_r159_c126 bl[126] br[126] wl[159] vdd gnd cell_6t
Xbit_r160_c126 bl[126] br[126] wl[160] vdd gnd cell_6t
Xbit_r161_c126 bl[126] br[126] wl[161] vdd gnd cell_6t
Xbit_r162_c126 bl[126] br[126] wl[162] vdd gnd cell_6t
Xbit_r163_c126 bl[126] br[126] wl[163] vdd gnd cell_6t
Xbit_r164_c126 bl[126] br[126] wl[164] vdd gnd cell_6t
Xbit_r165_c126 bl[126] br[126] wl[165] vdd gnd cell_6t
Xbit_r166_c126 bl[126] br[126] wl[166] vdd gnd cell_6t
Xbit_r167_c126 bl[126] br[126] wl[167] vdd gnd cell_6t
Xbit_r168_c126 bl[126] br[126] wl[168] vdd gnd cell_6t
Xbit_r169_c126 bl[126] br[126] wl[169] vdd gnd cell_6t
Xbit_r170_c126 bl[126] br[126] wl[170] vdd gnd cell_6t
Xbit_r171_c126 bl[126] br[126] wl[171] vdd gnd cell_6t
Xbit_r172_c126 bl[126] br[126] wl[172] vdd gnd cell_6t
Xbit_r173_c126 bl[126] br[126] wl[173] vdd gnd cell_6t
Xbit_r174_c126 bl[126] br[126] wl[174] vdd gnd cell_6t
Xbit_r175_c126 bl[126] br[126] wl[175] vdd gnd cell_6t
Xbit_r176_c126 bl[126] br[126] wl[176] vdd gnd cell_6t
Xbit_r177_c126 bl[126] br[126] wl[177] vdd gnd cell_6t
Xbit_r178_c126 bl[126] br[126] wl[178] vdd gnd cell_6t
Xbit_r179_c126 bl[126] br[126] wl[179] vdd gnd cell_6t
Xbit_r180_c126 bl[126] br[126] wl[180] vdd gnd cell_6t
Xbit_r181_c126 bl[126] br[126] wl[181] vdd gnd cell_6t
Xbit_r182_c126 bl[126] br[126] wl[182] vdd gnd cell_6t
Xbit_r183_c126 bl[126] br[126] wl[183] vdd gnd cell_6t
Xbit_r184_c126 bl[126] br[126] wl[184] vdd gnd cell_6t
Xbit_r185_c126 bl[126] br[126] wl[185] vdd gnd cell_6t
Xbit_r186_c126 bl[126] br[126] wl[186] vdd gnd cell_6t
Xbit_r187_c126 bl[126] br[126] wl[187] vdd gnd cell_6t
Xbit_r188_c126 bl[126] br[126] wl[188] vdd gnd cell_6t
Xbit_r189_c126 bl[126] br[126] wl[189] vdd gnd cell_6t
Xbit_r190_c126 bl[126] br[126] wl[190] vdd gnd cell_6t
Xbit_r191_c126 bl[126] br[126] wl[191] vdd gnd cell_6t
Xbit_r192_c126 bl[126] br[126] wl[192] vdd gnd cell_6t
Xbit_r193_c126 bl[126] br[126] wl[193] vdd gnd cell_6t
Xbit_r194_c126 bl[126] br[126] wl[194] vdd gnd cell_6t
Xbit_r195_c126 bl[126] br[126] wl[195] vdd gnd cell_6t
Xbit_r196_c126 bl[126] br[126] wl[196] vdd gnd cell_6t
Xbit_r197_c126 bl[126] br[126] wl[197] vdd gnd cell_6t
Xbit_r198_c126 bl[126] br[126] wl[198] vdd gnd cell_6t
Xbit_r199_c126 bl[126] br[126] wl[199] vdd gnd cell_6t
Xbit_r200_c126 bl[126] br[126] wl[200] vdd gnd cell_6t
Xbit_r201_c126 bl[126] br[126] wl[201] vdd gnd cell_6t
Xbit_r202_c126 bl[126] br[126] wl[202] vdd gnd cell_6t
Xbit_r203_c126 bl[126] br[126] wl[203] vdd gnd cell_6t
Xbit_r204_c126 bl[126] br[126] wl[204] vdd gnd cell_6t
Xbit_r205_c126 bl[126] br[126] wl[205] vdd gnd cell_6t
Xbit_r206_c126 bl[126] br[126] wl[206] vdd gnd cell_6t
Xbit_r207_c126 bl[126] br[126] wl[207] vdd gnd cell_6t
Xbit_r208_c126 bl[126] br[126] wl[208] vdd gnd cell_6t
Xbit_r209_c126 bl[126] br[126] wl[209] vdd gnd cell_6t
Xbit_r210_c126 bl[126] br[126] wl[210] vdd gnd cell_6t
Xbit_r211_c126 bl[126] br[126] wl[211] vdd gnd cell_6t
Xbit_r212_c126 bl[126] br[126] wl[212] vdd gnd cell_6t
Xbit_r213_c126 bl[126] br[126] wl[213] vdd gnd cell_6t
Xbit_r214_c126 bl[126] br[126] wl[214] vdd gnd cell_6t
Xbit_r215_c126 bl[126] br[126] wl[215] vdd gnd cell_6t
Xbit_r216_c126 bl[126] br[126] wl[216] vdd gnd cell_6t
Xbit_r217_c126 bl[126] br[126] wl[217] vdd gnd cell_6t
Xbit_r218_c126 bl[126] br[126] wl[218] vdd gnd cell_6t
Xbit_r219_c126 bl[126] br[126] wl[219] vdd gnd cell_6t
Xbit_r220_c126 bl[126] br[126] wl[220] vdd gnd cell_6t
Xbit_r221_c126 bl[126] br[126] wl[221] vdd gnd cell_6t
Xbit_r222_c126 bl[126] br[126] wl[222] vdd gnd cell_6t
Xbit_r223_c126 bl[126] br[126] wl[223] vdd gnd cell_6t
Xbit_r224_c126 bl[126] br[126] wl[224] vdd gnd cell_6t
Xbit_r225_c126 bl[126] br[126] wl[225] vdd gnd cell_6t
Xbit_r226_c126 bl[126] br[126] wl[226] vdd gnd cell_6t
Xbit_r227_c126 bl[126] br[126] wl[227] vdd gnd cell_6t
Xbit_r228_c126 bl[126] br[126] wl[228] vdd gnd cell_6t
Xbit_r229_c126 bl[126] br[126] wl[229] vdd gnd cell_6t
Xbit_r230_c126 bl[126] br[126] wl[230] vdd gnd cell_6t
Xbit_r231_c126 bl[126] br[126] wl[231] vdd gnd cell_6t
Xbit_r232_c126 bl[126] br[126] wl[232] vdd gnd cell_6t
Xbit_r233_c126 bl[126] br[126] wl[233] vdd gnd cell_6t
Xbit_r234_c126 bl[126] br[126] wl[234] vdd gnd cell_6t
Xbit_r235_c126 bl[126] br[126] wl[235] vdd gnd cell_6t
Xbit_r236_c126 bl[126] br[126] wl[236] vdd gnd cell_6t
Xbit_r237_c126 bl[126] br[126] wl[237] vdd gnd cell_6t
Xbit_r238_c126 bl[126] br[126] wl[238] vdd gnd cell_6t
Xbit_r239_c126 bl[126] br[126] wl[239] vdd gnd cell_6t
Xbit_r240_c126 bl[126] br[126] wl[240] vdd gnd cell_6t
Xbit_r241_c126 bl[126] br[126] wl[241] vdd gnd cell_6t
Xbit_r242_c126 bl[126] br[126] wl[242] vdd gnd cell_6t
Xbit_r243_c126 bl[126] br[126] wl[243] vdd gnd cell_6t
Xbit_r244_c126 bl[126] br[126] wl[244] vdd gnd cell_6t
Xbit_r245_c126 bl[126] br[126] wl[245] vdd gnd cell_6t
Xbit_r246_c126 bl[126] br[126] wl[246] vdd gnd cell_6t
Xbit_r247_c126 bl[126] br[126] wl[247] vdd gnd cell_6t
Xbit_r248_c126 bl[126] br[126] wl[248] vdd gnd cell_6t
Xbit_r249_c126 bl[126] br[126] wl[249] vdd gnd cell_6t
Xbit_r250_c126 bl[126] br[126] wl[250] vdd gnd cell_6t
Xbit_r251_c126 bl[126] br[126] wl[251] vdd gnd cell_6t
Xbit_r252_c126 bl[126] br[126] wl[252] vdd gnd cell_6t
Xbit_r253_c126 bl[126] br[126] wl[253] vdd gnd cell_6t
Xbit_r254_c126 bl[126] br[126] wl[254] vdd gnd cell_6t
Xbit_r255_c126 bl[126] br[126] wl[255] vdd gnd cell_6t
Xbit_r0_c127 bl[127] br[127] wl[0] vdd gnd cell_6t
Xbit_r1_c127 bl[127] br[127] wl[1] vdd gnd cell_6t
Xbit_r2_c127 bl[127] br[127] wl[2] vdd gnd cell_6t
Xbit_r3_c127 bl[127] br[127] wl[3] vdd gnd cell_6t
Xbit_r4_c127 bl[127] br[127] wl[4] vdd gnd cell_6t
Xbit_r5_c127 bl[127] br[127] wl[5] vdd gnd cell_6t
Xbit_r6_c127 bl[127] br[127] wl[6] vdd gnd cell_6t
Xbit_r7_c127 bl[127] br[127] wl[7] vdd gnd cell_6t
Xbit_r8_c127 bl[127] br[127] wl[8] vdd gnd cell_6t
Xbit_r9_c127 bl[127] br[127] wl[9] vdd gnd cell_6t
Xbit_r10_c127 bl[127] br[127] wl[10] vdd gnd cell_6t
Xbit_r11_c127 bl[127] br[127] wl[11] vdd gnd cell_6t
Xbit_r12_c127 bl[127] br[127] wl[12] vdd gnd cell_6t
Xbit_r13_c127 bl[127] br[127] wl[13] vdd gnd cell_6t
Xbit_r14_c127 bl[127] br[127] wl[14] vdd gnd cell_6t
Xbit_r15_c127 bl[127] br[127] wl[15] vdd gnd cell_6t
Xbit_r16_c127 bl[127] br[127] wl[16] vdd gnd cell_6t
Xbit_r17_c127 bl[127] br[127] wl[17] vdd gnd cell_6t
Xbit_r18_c127 bl[127] br[127] wl[18] vdd gnd cell_6t
Xbit_r19_c127 bl[127] br[127] wl[19] vdd gnd cell_6t
Xbit_r20_c127 bl[127] br[127] wl[20] vdd gnd cell_6t
Xbit_r21_c127 bl[127] br[127] wl[21] vdd gnd cell_6t
Xbit_r22_c127 bl[127] br[127] wl[22] vdd gnd cell_6t
Xbit_r23_c127 bl[127] br[127] wl[23] vdd gnd cell_6t
Xbit_r24_c127 bl[127] br[127] wl[24] vdd gnd cell_6t
Xbit_r25_c127 bl[127] br[127] wl[25] vdd gnd cell_6t
Xbit_r26_c127 bl[127] br[127] wl[26] vdd gnd cell_6t
Xbit_r27_c127 bl[127] br[127] wl[27] vdd gnd cell_6t
Xbit_r28_c127 bl[127] br[127] wl[28] vdd gnd cell_6t
Xbit_r29_c127 bl[127] br[127] wl[29] vdd gnd cell_6t
Xbit_r30_c127 bl[127] br[127] wl[30] vdd gnd cell_6t
Xbit_r31_c127 bl[127] br[127] wl[31] vdd gnd cell_6t
Xbit_r32_c127 bl[127] br[127] wl[32] vdd gnd cell_6t
Xbit_r33_c127 bl[127] br[127] wl[33] vdd gnd cell_6t
Xbit_r34_c127 bl[127] br[127] wl[34] vdd gnd cell_6t
Xbit_r35_c127 bl[127] br[127] wl[35] vdd gnd cell_6t
Xbit_r36_c127 bl[127] br[127] wl[36] vdd gnd cell_6t
Xbit_r37_c127 bl[127] br[127] wl[37] vdd gnd cell_6t
Xbit_r38_c127 bl[127] br[127] wl[38] vdd gnd cell_6t
Xbit_r39_c127 bl[127] br[127] wl[39] vdd gnd cell_6t
Xbit_r40_c127 bl[127] br[127] wl[40] vdd gnd cell_6t
Xbit_r41_c127 bl[127] br[127] wl[41] vdd gnd cell_6t
Xbit_r42_c127 bl[127] br[127] wl[42] vdd gnd cell_6t
Xbit_r43_c127 bl[127] br[127] wl[43] vdd gnd cell_6t
Xbit_r44_c127 bl[127] br[127] wl[44] vdd gnd cell_6t
Xbit_r45_c127 bl[127] br[127] wl[45] vdd gnd cell_6t
Xbit_r46_c127 bl[127] br[127] wl[46] vdd gnd cell_6t
Xbit_r47_c127 bl[127] br[127] wl[47] vdd gnd cell_6t
Xbit_r48_c127 bl[127] br[127] wl[48] vdd gnd cell_6t
Xbit_r49_c127 bl[127] br[127] wl[49] vdd gnd cell_6t
Xbit_r50_c127 bl[127] br[127] wl[50] vdd gnd cell_6t
Xbit_r51_c127 bl[127] br[127] wl[51] vdd gnd cell_6t
Xbit_r52_c127 bl[127] br[127] wl[52] vdd gnd cell_6t
Xbit_r53_c127 bl[127] br[127] wl[53] vdd gnd cell_6t
Xbit_r54_c127 bl[127] br[127] wl[54] vdd gnd cell_6t
Xbit_r55_c127 bl[127] br[127] wl[55] vdd gnd cell_6t
Xbit_r56_c127 bl[127] br[127] wl[56] vdd gnd cell_6t
Xbit_r57_c127 bl[127] br[127] wl[57] vdd gnd cell_6t
Xbit_r58_c127 bl[127] br[127] wl[58] vdd gnd cell_6t
Xbit_r59_c127 bl[127] br[127] wl[59] vdd gnd cell_6t
Xbit_r60_c127 bl[127] br[127] wl[60] vdd gnd cell_6t
Xbit_r61_c127 bl[127] br[127] wl[61] vdd gnd cell_6t
Xbit_r62_c127 bl[127] br[127] wl[62] vdd gnd cell_6t
Xbit_r63_c127 bl[127] br[127] wl[63] vdd gnd cell_6t
Xbit_r64_c127 bl[127] br[127] wl[64] vdd gnd cell_6t
Xbit_r65_c127 bl[127] br[127] wl[65] vdd gnd cell_6t
Xbit_r66_c127 bl[127] br[127] wl[66] vdd gnd cell_6t
Xbit_r67_c127 bl[127] br[127] wl[67] vdd gnd cell_6t
Xbit_r68_c127 bl[127] br[127] wl[68] vdd gnd cell_6t
Xbit_r69_c127 bl[127] br[127] wl[69] vdd gnd cell_6t
Xbit_r70_c127 bl[127] br[127] wl[70] vdd gnd cell_6t
Xbit_r71_c127 bl[127] br[127] wl[71] vdd gnd cell_6t
Xbit_r72_c127 bl[127] br[127] wl[72] vdd gnd cell_6t
Xbit_r73_c127 bl[127] br[127] wl[73] vdd gnd cell_6t
Xbit_r74_c127 bl[127] br[127] wl[74] vdd gnd cell_6t
Xbit_r75_c127 bl[127] br[127] wl[75] vdd gnd cell_6t
Xbit_r76_c127 bl[127] br[127] wl[76] vdd gnd cell_6t
Xbit_r77_c127 bl[127] br[127] wl[77] vdd gnd cell_6t
Xbit_r78_c127 bl[127] br[127] wl[78] vdd gnd cell_6t
Xbit_r79_c127 bl[127] br[127] wl[79] vdd gnd cell_6t
Xbit_r80_c127 bl[127] br[127] wl[80] vdd gnd cell_6t
Xbit_r81_c127 bl[127] br[127] wl[81] vdd gnd cell_6t
Xbit_r82_c127 bl[127] br[127] wl[82] vdd gnd cell_6t
Xbit_r83_c127 bl[127] br[127] wl[83] vdd gnd cell_6t
Xbit_r84_c127 bl[127] br[127] wl[84] vdd gnd cell_6t
Xbit_r85_c127 bl[127] br[127] wl[85] vdd gnd cell_6t
Xbit_r86_c127 bl[127] br[127] wl[86] vdd gnd cell_6t
Xbit_r87_c127 bl[127] br[127] wl[87] vdd gnd cell_6t
Xbit_r88_c127 bl[127] br[127] wl[88] vdd gnd cell_6t
Xbit_r89_c127 bl[127] br[127] wl[89] vdd gnd cell_6t
Xbit_r90_c127 bl[127] br[127] wl[90] vdd gnd cell_6t
Xbit_r91_c127 bl[127] br[127] wl[91] vdd gnd cell_6t
Xbit_r92_c127 bl[127] br[127] wl[92] vdd gnd cell_6t
Xbit_r93_c127 bl[127] br[127] wl[93] vdd gnd cell_6t
Xbit_r94_c127 bl[127] br[127] wl[94] vdd gnd cell_6t
Xbit_r95_c127 bl[127] br[127] wl[95] vdd gnd cell_6t
Xbit_r96_c127 bl[127] br[127] wl[96] vdd gnd cell_6t
Xbit_r97_c127 bl[127] br[127] wl[97] vdd gnd cell_6t
Xbit_r98_c127 bl[127] br[127] wl[98] vdd gnd cell_6t
Xbit_r99_c127 bl[127] br[127] wl[99] vdd gnd cell_6t
Xbit_r100_c127 bl[127] br[127] wl[100] vdd gnd cell_6t
Xbit_r101_c127 bl[127] br[127] wl[101] vdd gnd cell_6t
Xbit_r102_c127 bl[127] br[127] wl[102] vdd gnd cell_6t
Xbit_r103_c127 bl[127] br[127] wl[103] vdd gnd cell_6t
Xbit_r104_c127 bl[127] br[127] wl[104] vdd gnd cell_6t
Xbit_r105_c127 bl[127] br[127] wl[105] vdd gnd cell_6t
Xbit_r106_c127 bl[127] br[127] wl[106] vdd gnd cell_6t
Xbit_r107_c127 bl[127] br[127] wl[107] vdd gnd cell_6t
Xbit_r108_c127 bl[127] br[127] wl[108] vdd gnd cell_6t
Xbit_r109_c127 bl[127] br[127] wl[109] vdd gnd cell_6t
Xbit_r110_c127 bl[127] br[127] wl[110] vdd gnd cell_6t
Xbit_r111_c127 bl[127] br[127] wl[111] vdd gnd cell_6t
Xbit_r112_c127 bl[127] br[127] wl[112] vdd gnd cell_6t
Xbit_r113_c127 bl[127] br[127] wl[113] vdd gnd cell_6t
Xbit_r114_c127 bl[127] br[127] wl[114] vdd gnd cell_6t
Xbit_r115_c127 bl[127] br[127] wl[115] vdd gnd cell_6t
Xbit_r116_c127 bl[127] br[127] wl[116] vdd gnd cell_6t
Xbit_r117_c127 bl[127] br[127] wl[117] vdd gnd cell_6t
Xbit_r118_c127 bl[127] br[127] wl[118] vdd gnd cell_6t
Xbit_r119_c127 bl[127] br[127] wl[119] vdd gnd cell_6t
Xbit_r120_c127 bl[127] br[127] wl[120] vdd gnd cell_6t
Xbit_r121_c127 bl[127] br[127] wl[121] vdd gnd cell_6t
Xbit_r122_c127 bl[127] br[127] wl[122] vdd gnd cell_6t
Xbit_r123_c127 bl[127] br[127] wl[123] vdd gnd cell_6t
Xbit_r124_c127 bl[127] br[127] wl[124] vdd gnd cell_6t
Xbit_r125_c127 bl[127] br[127] wl[125] vdd gnd cell_6t
Xbit_r126_c127 bl[127] br[127] wl[126] vdd gnd cell_6t
Xbit_r127_c127 bl[127] br[127] wl[127] vdd gnd cell_6t
Xbit_r128_c127 bl[127] br[127] wl[128] vdd gnd cell_6t
Xbit_r129_c127 bl[127] br[127] wl[129] vdd gnd cell_6t
Xbit_r130_c127 bl[127] br[127] wl[130] vdd gnd cell_6t
Xbit_r131_c127 bl[127] br[127] wl[131] vdd gnd cell_6t
Xbit_r132_c127 bl[127] br[127] wl[132] vdd gnd cell_6t
Xbit_r133_c127 bl[127] br[127] wl[133] vdd gnd cell_6t
Xbit_r134_c127 bl[127] br[127] wl[134] vdd gnd cell_6t
Xbit_r135_c127 bl[127] br[127] wl[135] vdd gnd cell_6t
Xbit_r136_c127 bl[127] br[127] wl[136] vdd gnd cell_6t
Xbit_r137_c127 bl[127] br[127] wl[137] vdd gnd cell_6t
Xbit_r138_c127 bl[127] br[127] wl[138] vdd gnd cell_6t
Xbit_r139_c127 bl[127] br[127] wl[139] vdd gnd cell_6t
Xbit_r140_c127 bl[127] br[127] wl[140] vdd gnd cell_6t
Xbit_r141_c127 bl[127] br[127] wl[141] vdd gnd cell_6t
Xbit_r142_c127 bl[127] br[127] wl[142] vdd gnd cell_6t
Xbit_r143_c127 bl[127] br[127] wl[143] vdd gnd cell_6t
Xbit_r144_c127 bl[127] br[127] wl[144] vdd gnd cell_6t
Xbit_r145_c127 bl[127] br[127] wl[145] vdd gnd cell_6t
Xbit_r146_c127 bl[127] br[127] wl[146] vdd gnd cell_6t
Xbit_r147_c127 bl[127] br[127] wl[147] vdd gnd cell_6t
Xbit_r148_c127 bl[127] br[127] wl[148] vdd gnd cell_6t
Xbit_r149_c127 bl[127] br[127] wl[149] vdd gnd cell_6t
Xbit_r150_c127 bl[127] br[127] wl[150] vdd gnd cell_6t
Xbit_r151_c127 bl[127] br[127] wl[151] vdd gnd cell_6t
Xbit_r152_c127 bl[127] br[127] wl[152] vdd gnd cell_6t
Xbit_r153_c127 bl[127] br[127] wl[153] vdd gnd cell_6t
Xbit_r154_c127 bl[127] br[127] wl[154] vdd gnd cell_6t
Xbit_r155_c127 bl[127] br[127] wl[155] vdd gnd cell_6t
Xbit_r156_c127 bl[127] br[127] wl[156] vdd gnd cell_6t
Xbit_r157_c127 bl[127] br[127] wl[157] vdd gnd cell_6t
Xbit_r158_c127 bl[127] br[127] wl[158] vdd gnd cell_6t
Xbit_r159_c127 bl[127] br[127] wl[159] vdd gnd cell_6t
Xbit_r160_c127 bl[127] br[127] wl[160] vdd gnd cell_6t
Xbit_r161_c127 bl[127] br[127] wl[161] vdd gnd cell_6t
Xbit_r162_c127 bl[127] br[127] wl[162] vdd gnd cell_6t
Xbit_r163_c127 bl[127] br[127] wl[163] vdd gnd cell_6t
Xbit_r164_c127 bl[127] br[127] wl[164] vdd gnd cell_6t
Xbit_r165_c127 bl[127] br[127] wl[165] vdd gnd cell_6t
Xbit_r166_c127 bl[127] br[127] wl[166] vdd gnd cell_6t
Xbit_r167_c127 bl[127] br[127] wl[167] vdd gnd cell_6t
Xbit_r168_c127 bl[127] br[127] wl[168] vdd gnd cell_6t
Xbit_r169_c127 bl[127] br[127] wl[169] vdd gnd cell_6t
Xbit_r170_c127 bl[127] br[127] wl[170] vdd gnd cell_6t
Xbit_r171_c127 bl[127] br[127] wl[171] vdd gnd cell_6t
Xbit_r172_c127 bl[127] br[127] wl[172] vdd gnd cell_6t
Xbit_r173_c127 bl[127] br[127] wl[173] vdd gnd cell_6t
Xbit_r174_c127 bl[127] br[127] wl[174] vdd gnd cell_6t
Xbit_r175_c127 bl[127] br[127] wl[175] vdd gnd cell_6t
Xbit_r176_c127 bl[127] br[127] wl[176] vdd gnd cell_6t
Xbit_r177_c127 bl[127] br[127] wl[177] vdd gnd cell_6t
Xbit_r178_c127 bl[127] br[127] wl[178] vdd gnd cell_6t
Xbit_r179_c127 bl[127] br[127] wl[179] vdd gnd cell_6t
Xbit_r180_c127 bl[127] br[127] wl[180] vdd gnd cell_6t
Xbit_r181_c127 bl[127] br[127] wl[181] vdd gnd cell_6t
Xbit_r182_c127 bl[127] br[127] wl[182] vdd gnd cell_6t
Xbit_r183_c127 bl[127] br[127] wl[183] vdd gnd cell_6t
Xbit_r184_c127 bl[127] br[127] wl[184] vdd gnd cell_6t
Xbit_r185_c127 bl[127] br[127] wl[185] vdd gnd cell_6t
Xbit_r186_c127 bl[127] br[127] wl[186] vdd gnd cell_6t
Xbit_r187_c127 bl[127] br[127] wl[187] vdd gnd cell_6t
Xbit_r188_c127 bl[127] br[127] wl[188] vdd gnd cell_6t
Xbit_r189_c127 bl[127] br[127] wl[189] vdd gnd cell_6t
Xbit_r190_c127 bl[127] br[127] wl[190] vdd gnd cell_6t
Xbit_r191_c127 bl[127] br[127] wl[191] vdd gnd cell_6t
Xbit_r192_c127 bl[127] br[127] wl[192] vdd gnd cell_6t
Xbit_r193_c127 bl[127] br[127] wl[193] vdd gnd cell_6t
Xbit_r194_c127 bl[127] br[127] wl[194] vdd gnd cell_6t
Xbit_r195_c127 bl[127] br[127] wl[195] vdd gnd cell_6t
Xbit_r196_c127 bl[127] br[127] wl[196] vdd gnd cell_6t
Xbit_r197_c127 bl[127] br[127] wl[197] vdd gnd cell_6t
Xbit_r198_c127 bl[127] br[127] wl[198] vdd gnd cell_6t
Xbit_r199_c127 bl[127] br[127] wl[199] vdd gnd cell_6t
Xbit_r200_c127 bl[127] br[127] wl[200] vdd gnd cell_6t
Xbit_r201_c127 bl[127] br[127] wl[201] vdd gnd cell_6t
Xbit_r202_c127 bl[127] br[127] wl[202] vdd gnd cell_6t
Xbit_r203_c127 bl[127] br[127] wl[203] vdd gnd cell_6t
Xbit_r204_c127 bl[127] br[127] wl[204] vdd gnd cell_6t
Xbit_r205_c127 bl[127] br[127] wl[205] vdd gnd cell_6t
Xbit_r206_c127 bl[127] br[127] wl[206] vdd gnd cell_6t
Xbit_r207_c127 bl[127] br[127] wl[207] vdd gnd cell_6t
Xbit_r208_c127 bl[127] br[127] wl[208] vdd gnd cell_6t
Xbit_r209_c127 bl[127] br[127] wl[209] vdd gnd cell_6t
Xbit_r210_c127 bl[127] br[127] wl[210] vdd gnd cell_6t
Xbit_r211_c127 bl[127] br[127] wl[211] vdd gnd cell_6t
Xbit_r212_c127 bl[127] br[127] wl[212] vdd gnd cell_6t
Xbit_r213_c127 bl[127] br[127] wl[213] vdd gnd cell_6t
Xbit_r214_c127 bl[127] br[127] wl[214] vdd gnd cell_6t
Xbit_r215_c127 bl[127] br[127] wl[215] vdd gnd cell_6t
Xbit_r216_c127 bl[127] br[127] wl[216] vdd gnd cell_6t
Xbit_r217_c127 bl[127] br[127] wl[217] vdd gnd cell_6t
Xbit_r218_c127 bl[127] br[127] wl[218] vdd gnd cell_6t
Xbit_r219_c127 bl[127] br[127] wl[219] vdd gnd cell_6t
Xbit_r220_c127 bl[127] br[127] wl[220] vdd gnd cell_6t
Xbit_r221_c127 bl[127] br[127] wl[221] vdd gnd cell_6t
Xbit_r222_c127 bl[127] br[127] wl[222] vdd gnd cell_6t
Xbit_r223_c127 bl[127] br[127] wl[223] vdd gnd cell_6t
Xbit_r224_c127 bl[127] br[127] wl[224] vdd gnd cell_6t
Xbit_r225_c127 bl[127] br[127] wl[225] vdd gnd cell_6t
Xbit_r226_c127 bl[127] br[127] wl[226] vdd gnd cell_6t
Xbit_r227_c127 bl[127] br[127] wl[227] vdd gnd cell_6t
Xbit_r228_c127 bl[127] br[127] wl[228] vdd gnd cell_6t
Xbit_r229_c127 bl[127] br[127] wl[229] vdd gnd cell_6t
Xbit_r230_c127 bl[127] br[127] wl[230] vdd gnd cell_6t
Xbit_r231_c127 bl[127] br[127] wl[231] vdd gnd cell_6t
Xbit_r232_c127 bl[127] br[127] wl[232] vdd gnd cell_6t
Xbit_r233_c127 bl[127] br[127] wl[233] vdd gnd cell_6t
Xbit_r234_c127 bl[127] br[127] wl[234] vdd gnd cell_6t
Xbit_r235_c127 bl[127] br[127] wl[235] vdd gnd cell_6t
Xbit_r236_c127 bl[127] br[127] wl[236] vdd gnd cell_6t
Xbit_r237_c127 bl[127] br[127] wl[237] vdd gnd cell_6t
Xbit_r238_c127 bl[127] br[127] wl[238] vdd gnd cell_6t
Xbit_r239_c127 bl[127] br[127] wl[239] vdd gnd cell_6t
Xbit_r240_c127 bl[127] br[127] wl[240] vdd gnd cell_6t
Xbit_r241_c127 bl[127] br[127] wl[241] vdd gnd cell_6t
Xbit_r242_c127 bl[127] br[127] wl[242] vdd gnd cell_6t
Xbit_r243_c127 bl[127] br[127] wl[243] vdd gnd cell_6t
Xbit_r244_c127 bl[127] br[127] wl[244] vdd gnd cell_6t
Xbit_r245_c127 bl[127] br[127] wl[245] vdd gnd cell_6t
Xbit_r246_c127 bl[127] br[127] wl[246] vdd gnd cell_6t
Xbit_r247_c127 bl[127] br[127] wl[247] vdd gnd cell_6t
Xbit_r248_c127 bl[127] br[127] wl[248] vdd gnd cell_6t
Xbit_r249_c127 bl[127] br[127] wl[249] vdd gnd cell_6t
Xbit_r250_c127 bl[127] br[127] wl[250] vdd gnd cell_6t
Xbit_r251_c127 bl[127] br[127] wl[251] vdd gnd cell_6t
Xbit_r252_c127 bl[127] br[127] wl[252] vdd gnd cell_6t
Xbit_r253_c127 bl[127] br[127] wl[253] vdd gnd cell_6t
Xbit_r254_c127 bl[127] br[127] wl[254] vdd gnd cell_6t
Xbit_r255_c127 bl[127] br[127] wl[255] vdd gnd cell_6t
.ENDS bitcell_array

* ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p

.SUBCKT precharge bl br en vdd
Mlower_pmos bl en BR vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mupper_pmos1 bl en vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mupper_pmos2 br en vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
.ENDS precharge

.SUBCKT precharge_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] en vdd
Xpre_column_0 bl[0] br[0] en vdd precharge
Xpre_column_1 bl[1] br[1] en vdd precharge
Xpre_column_2 bl[2] br[2] en vdd precharge
Xpre_column_3 bl[3] br[3] en vdd precharge
Xpre_column_4 bl[4] br[4] en vdd precharge
Xpre_column_5 bl[5] br[5] en vdd precharge
Xpre_column_6 bl[6] br[6] en vdd precharge
Xpre_column_7 bl[7] br[7] en vdd precharge
Xpre_column_8 bl[8] br[8] en vdd precharge
Xpre_column_9 bl[9] br[9] en vdd precharge
Xpre_column_10 bl[10] br[10] en vdd precharge
Xpre_column_11 bl[11] br[11] en vdd precharge
Xpre_column_12 bl[12] br[12] en vdd precharge
Xpre_column_13 bl[13] br[13] en vdd precharge
Xpre_column_14 bl[14] br[14] en vdd precharge
Xpre_column_15 bl[15] br[15] en vdd precharge
Xpre_column_16 bl[16] br[16] en vdd precharge
Xpre_column_17 bl[17] br[17] en vdd precharge
Xpre_column_18 bl[18] br[18] en vdd precharge
Xpre_column_19 bl[19] br[19] en vdd precharge
Xpre_column_20 bl[20] br[20] en vdd precharge
Xpre_column_21 bl[21] br[21] en vdd precharge
Xpre_column_22 bl[22] br[22] en vdd precharge
Xpre_column_23 bl[23] br[23] en vdd precharge
Xpre_column_24 bl[24] br[24] en vdd precharge
Xpre_column_25 bl[25] br[25] en vdd precharge
Xpre_column_26 bl[26] br[26] en vdd precharge
Xpre_column_27 bl[27] br[27] en vdd precharge
Xpre_column_28 bl[28] br[28] en vdd precharge
Xpre_column_29 bl[29] br[29] en vdd precharge
Xpre_column_30 bl[30] br[30] en vdd precharge
Xpre_column_31 bl[31] br[31] en vdd precharge
Xpre_column_32 bl[32] br[32] en vdd precharge
Xpre_column_33 bl[33] br[33] en vdd precharge
Xpre_column_34 bl[34] br[34] en vdd precharge
Xpre_column_35 bl[35] br[35] en vdd precharge
Xpre_column_36 bl[36] br[36] en vdd precharge
Xpre_column_37 bl[37] br[37] en vdd precharge
Xpre_column_38 bl[38] br[38] en vdd precharge
Xpre_column_39 bl[39] br[39] en vdd precharge
Xpre_column_40 bl[40] br[40] en vdd precharge
Xpre_column_41 bl[41] br[41] en vdd precharge
Xpre_column_42 bl[42] br[42] en vdd precharge
Xpre_column_43 bl[43] br[43] en vdd precharge
Xpre_column_44 bl[44] br[44] en vdd precharge
Xpre_column_45 bl[45] br[45] en vdd precharge
Xpre_column_46 bl[46] br[46] en vdd precharge
Xpre_column_47 bl[47] br[47] en vdd precharge
Xpre_column_48 bl[48] br[48] en vdd precharge
Xpre_column_49 bl[49] br[49] en vdd precharge
Xpre_column_50 bl[50] br[50] en vdd precharge
Xpre_column_51 bl[51] br[51] en vdd precharge
Xpre_column_52 bl[52] br[52] en vdd precharge
Xpre_column_53 bl[53] br[53] en vdd precharge
Xpre_column_54 bl[54] br[54] en vdd precharge
Xpre_column_55 bl[55] br[55] en vdd precharge
Xpre_column_56 bl[56] br[56] en vdd precharge
Xpre_column_57 bl[57] br[57] en vdd precharge
Xpre_column_58 bl[58] br[58] en vdd precharge
Xpre_column_59 bl[59] br[59] en vdd precharge
Xpre_column_60 bl[60] br[60] en vdd precharge
Xpre_column_61 bl[61] br[61] en vdd precharge
Xpre_column_62 bl[62] br[62] en vdd precharge
Xpre_column_63 bl[63] br[63] en vdd precharge
Xpre_column_64 bl[64] br[64] en vdd precharge
Xpre_column_65 bl[65] br[65] en vdd precharge
Xpre_column_66 bl[66] br[66] en vdd precharge
Xpre_column_67 bl[67] br[67] en vdd precharge
Xpre_column_68 bl[68] br[68] en vdd precharge
Xpre_column_69 bl[69] br[69] en vdd precharge
Xpre_column_70 bl[70] br[70] en vdd precharge
Xpre_column_71 bl[71] br[71] en vdd precharge
Xpre_column_72 bl[72] br[72] en vdd precharge
Xpre_column_73 bl[73] br[73] en vdd precharge
Xpre_column_74 bl[74] br[74] en vdd precharge
Xpre_column_75 bl[75] br[75] en vdd precharge
Xpre_column_76 bl[76] br[76] en vdd precharge
Xpre_column_77 bl[77] br[77] en vdd precharge
Xpre_column_78 bl[78] br[78] en vdd precharge
Xpre_column_79 bl[79] br[79] en vdd precharge
Xpre_column_80 bl[80] br[80] en vdd precharge
Xpre_column_81 bl[81] br[81] en vdd precharge
Xpre_column_82 bl[82] br[82] en vdd precharge
Xpre_column_83 bl[83] br[83] en vdd precharge
Xpre_column_84 bl[84] br[84] en vdd precharge
Xpre_column_85 bl[85] br[85] en vdd precharge
Xpre_column_86 bl[86] br[86] en vdd precharge
Xpre_column_87 bl[87] br[87] en vdd precharge
Xpre_column_88 bl[88] br[88] en vdd precharge
Xpre_column_89 bl[89] br[89] en vdd precharge
Xpre_column_90 bl[90] br[90] en vdd precharge
Xpre_column_91 bl[91] br[91] en vdd precharge
Xpre_column_92 bl[92] br[92] en vdd precharge
Xpre_column_93 bl[93] br[93] en vdd precharge
Xpre_column_94 bl[94] br[94] en vdd precharge
Xpre_column_95 bl[95] br[95] en vdd precharge
Xpre_column_96 bl[96] br[96] en vdd precharge
Xpre_column_97 bl[97] br[97] en vdd precharge
Xpre_column_98 bl[98] br[98] en vdd precharge
Xpre_column_99 bl[99] br[99] en vdd precharge
Xpre_column_100 bl[100] br[100] en vdd precharge
Xpre_column_101 bl[101] br[101] en vdd precharge
Xpre_column_102 bl[102] br[102] en vdd precharge
Xpre_column_103 bl[103] br[103] en vdd precharge
Xpre_column_104 bl[104] br[104] en vdd precharge
Xpre_column_105 bl[105] br[105] en vdd precharge
Xpre_column_106 bl[106] br[106] en vdd precharge
Xpre_column_107 bl[107] br[107] en vdd precharge
Xpre_column_108 bl[108] br[108] en vdd precharge
Xpre_column_109 bl[109] br[109] en vdd precharge
Xpre_column_110 bl[110] br[110] en vdd precharge
Xpre_column_111 bl[111] br[111] en vdd precharge
Xpre_column_112 bl[112] br[112] en vdd precharge
Xpre_column_113 bl[113] br[113] en vdd precharge
Xpre_column_114 bl[114] br[114] en vdd precharge
Xpre_column_115 bl[115] br[115] en vdd precharge
Xpre_column_116 bl[116] br[116] en vdd precharge
Xpre_column_117 bl[117] br[117] en vdd precharge
Xpre_column_118 bl[118] br[118] en vdd precharge
Xpre_column_119 bl[119] br[119] en vdd precharge
Xpre_column_120 bl[120] br[120] en vdd precharge
Xpre_column_121 bl[121] br[121] en vdd precharge
Xpre_column_122 bl[122] br[122] en vdd precharge
Xpre_column_123 bl[123] br[123] en vdd precharge
Xpre_column_124 bl[124] br[124] en vdd precharge
Xpre_column_125 bl[125] br[125] en vdd precharge
Xpre_column_126 bl[126] br[126] en vdd precharge
Xpre_column_127 bl[127] br[127] en vdd precharge
.ENDS precharge_array

* ptx M{0} {1} nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p

.SUBCKT single_level_column_mux_8 bl br bl_out br_out sel gnd
Mmux_tx1 bl sel bl_out gnd nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p
Mmux_tx2 br sel br_out gnd nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p
.ENDS single_level_column_mux_8

.SUBCKT columnmux_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] sel[0] sel[1] sel[2] sel[3] bl_out[0] br_out[0] bl_out[1] br_out[1] bl_out[2] br_out[2] bl_out[3] br_out[3] bl_out[4] br_out[4] bl_out[5] br_out[5] bl_out[6] br_out[6] bl_out[7] br_out[7] bl_out[8] br_out[8] bl_out[9] br_out[9] bl_out[10] br_out[10] bl_out[11] br_out[11] bl_out[12] br_out[12] bl_out[13] br_out[13] bl_out[14] br_out[14] bl_out[15] br_out[15] bl_out[16] br_out[16] bl_out[17] br_out[17] bl_out[18] br_out[18] bl_out[19] br_out[19] bl_out[20] br_out[20] bl_out[21] br_out[21] bl_out[22] br_out[22] bl_out[23] br_out[23] bl_out[24] br_out[24] bl_out[25] br_out[25] bl_out[26] br_out[26] bl_out[27] br_out[27] bl_out[28] br_out[28] bl_out[29] br_out[29] bl_out[30] br_out[30] bl_out[31] br_out[31] gnd
XXMUX0 bl[0] br[0] bl_out[0] br_out[0] sel[0] gnd single_level_column_mux_8
XXMUX1 bl[1] br[1] bl_out[0] br_out[0] sel[1] gnd single_level_column_mux_8
XXMUX2 bl[2] br[2] bl_out[0] br_out[0] sel[2] gnd single_level_column_mux_8
XXMUX3 bl[3] br[3] bl_out[0] br_out[0] sel[3] gnd single_level_column_mux_8
XXMUX4 bl[4] br[4] bl_out[1] br_out[1] sel[0] gnd single_level_column_mux_8
XXMUX5 bl[5] br[5] bl_out[1] br_out[1] sel[1] gnd single_level_column_mux_8
XXMUX6 bl[6] br[6] bl_out[1] br_out[1] sel[2] gnd single_level_column_mux_8
XXMUX7 bl[7] br[7] bl_out[1] br_out[1] sel[3] gnd single_level_column_mux_8
XXMUX8 bl[8] br[8] bl_out[2] br_out[2] sel[0] gnd single_level_column_mux_8
XXMUX9 bl[9] br[9] bl_out[2] br_out[2] sel[1] gnd single_level_column_mux_8
XXMUX10 bl[10] br[10] bl_out[2] br_out[2] sel[2] gnd single_level_column_mux_8
XXMUX11 bl[11] br[11] bl_out[2] br_out[2] sel[3] gnd single_level_column_mux_8
XXMUX12 bl[12] br[12] bl_out[3] br_out[3] sel[0] gnd single_level_column_mux_8
XXMUX13 bl[13] br[13] bl_out[3] br_out[3] sel[1] gnd single_level_column_mux_8
XXMUX14 bl[14] br[14] bl_out[3] br_out[3] sel[2] gnd single_level_column_mux_8
XXMUX15 bl[15] br[15] bl_out[3] br_out[3] sel[3] gnd single_level_column_mux_8
XXMUX16 bl[16] br[16] bl_out[4] br_out[4] sel[0] gnd single_level_column_mux_8
XXMUX17 bl[17] br[17] bl_out[4] br_out[4] sel[1] gnd single_level_column_mux_8
XXMUX18 bl[18] br[18] bl_out[4] br_out[4] sel[2] gnd single_level_column_mux_8
XXMUX19 bl[19] br[19] bl_out[4] br_out[4] sel[3] gnd single_level_column_mux_8
XXMUX20 bl[20] br[20] bl_out[5] br_out[5] sel[0] gnd single_level_column_mux_8
XXMUX21 bl[21] br[21] bl_out[5] br_out[5] sel[1] gnd single_level_column_mux_8
XXMUX22 bl[22] br[22] bl_out[5] br_out[5] sel[2] gnd single_level_column_mux_8
XXMUX23 bl[23] br[23] bl_out[5] br_out[5] sel[3] gnd single_level_column_mux_8
XXMUX24 bl[24] br[24] bl_out[6] br_out[6] sel[0] gnd single_level_column_mux_8
XXMUX25 bl[25] br[25] bl_out[6] br_out[6] sel[1] gnd single_level_column_mux_8
XXMUX26 bl[26] br[26] bl_out[6] br_out[6] sel[2] gnd single_level_column_mux_8
XXMUX27 bl[27] br[27] bl_out[6] br_out[6] sel[3] gnd single_level_column_mux_8
XXMUX28 bl[28] br[28] bl_out[7] br_out[7] sel[0] gnd single_level_column_mux_8
XXMUX29 bl[29] br[29] bl_out[7] br_out[7] sel[1] gnd single_level_column_mux_8
XXMUX30 bl[30] br[30] bl_out[7] br_out[7] sel[2] gnd single_level_column_mux_8
XXMUX31 bl[31] br[31] bl_out[7] br_out[7] sel[3] gnd single_level_column_mux_8
XXMUX32 bl[32] br[32] bl_out[8] br_out[8] sel[0] gnd single_level_column_mux_8
XXMUX33 bl[33] br[33] bl_out[8] br_out[8] sel[1] gnd single_level_column_mux_8
XXMUX34 bl[34] br[34] bl_out[8] br_out[8] sel[2] gnd single_level_column_mux_8
XXMUX35 bl[35] br[35] bl_out[8] br_out[8] sel[3] gnd single_level_column_mux_8
XXMUX36 bl[36] br[36] bl_out[9] br_out[9] sel[0] gnd single_level_column_mux_8
XXMUX37 bl[37] br[37] bl_out[9] br_out[9] sel[1] gnd single_level_column_mux_8
XXMUX38 bl[38] br[38] bl_out[9] br_out[9] sel[2] gnd single_level_column_mux_8
XXMUX39 bl[39] br[39] bl_out[9] br_out[9] sel[3] gnd single_level_column_mux_8
XXMUX40 bl[40] br[40] bl_out[10] br_out[10] sel[0] gnd single_level_column_mux_8
XXMUX41 bl[41] br[41] bl_out[10] br_out[10] sel[1] gnd single_level_column_mux_8
XXMUX42 bl[42] br[42] bl_out[10] br_out[10] sel[2] gnd single_level_column_mux_8
XXMUX43 bl[43] br[43] bl_out[10] br_out[10] sel[3] gnd single_level_column_mux_8
XXMUX44 bl[44] br[44] bl_out[11] br_out[11] sel[0] gnd single_level_column_mux_8
XXMUX45 bl[45] br[45] bl_out[11] br_out[11] sel[1] gnd single_level_column_mux_8
XXMUX46 bl[46] br[46] bl_out[11] br_out[11] sel[2] gnd single_level_column_mux_8
XXMUX47 bl[47] br[47] bl_out[11] br_out[11] sel[3] gnd single_level_column_mux_8
XXMUX48 bl[48] br[48] bl_out[12] br_out[12] sel[0] gnd single_level_column_mux_8
XXMUX49 bl[49] br[49] bl_out[12] br_out[12] sel[1] gnd single_level_column_mux_8
XXMUX50 bl[50] br[50] bl_out[12] br_out[12] sel[2] gnd single_level_column_mux_8
XXMUX51 bl[51] br[51] bl_out[12] br_out[12] sel[3] gnd single_level_column_mux_8
XXMUX52 bl[52] br[52] bl_out[13] br_out[13] sel[0] gnd single_level_column_mux_8
XXMUX53 bl[53] br[53] bl_out[13] br_out[13] sel[1] gnd single_level_column_mux_8
XXMUX54 bl[54] br[54] bl_out[13] br_out[13] sel[2] gnd single_level_column_mux_8
XXMUX55 bl[55] br[55] bl_out[13] br_out[13] sel[3] gnd single_level_column_mux_8
XXMUX56 bl[56] br[56] bl_out[14] br_out[14] sel[0] gnd single_level_column_mux_8
XXMUX57 bl[57] br[57] bl_out[14] br_out[14] sel[1] gnd single_level_column_mux_8
XXMUX58 bl[58] br[58] bl_out[14] br_out[14] sel[2] gnd single_level_column_mux_8
XXMUX59 bl[59] br[59] bl_out[14] br_out[14] sel[3] gnd single_level_column_mux_8
XXMUX60 bl[60] br[60] bl_out[15] br_out[15] sel[0] gnd single_level_column_mux_8
XXMUX61 bl[61] br[61] bl_out[15] br_out[15] sel[1] gnd single_level_column_mux_8
XXMUX62 bl[62] br[62] bl_out[15] br_out[15] sel[2] gnd single_level_column_mux_8
XXMUX63 bl[63] br[63] bl_out[15] br_out[15] sel[3] gnd single_level_column_mux_8
XXMUX64 bl[64] br[64] bl_out[16] br_out[16] sel[0] gnd single_level_column_mux_8
XXMUX65 bl[65] br[65] bl_out[16] br_out[16] sel[1] gnd single_level_column_mux_8
XXMUX66 bl[66] br[66] bl_out[16] br_out[16] sel[2] gnd single_level_column_mux_8
XXMUX67 bl[67] br[67] bl_out[16] br_out[16] sel[3] gnd single_level_column_mux_8
XXMUX68 bl[68] br[68] bl_out[17] br_out[17] sel[0] gnd single_level_column_mux_8
XXMUX69 bl[69] br[69] bl_out[17] br_out[17] sel[1] gnd single_level_column_mux_8
XXMUX70 bl[70] br[70] bl_out[17] br_out[17] sel[2] gnd single_level_column_mux_8
XXMUX71 bl[71] br[71] bl_out[17] br_out[17] sel[3] gnd single_level_column_mux_8
XXMUX72 bl[72] br[72] bl_out[18] br_out[18] sel[0] gnd single_level_column_mux_8
XXMUX73 bl[73] br[73] bl_out[18] br_out[18] sel[1] gnd single_level_column_mux_8
XXMUX74 bl[74] br[74] bl_out[18] br_out[18] sel[2] gnd single_level_column_mux_8
XXMUX75 bl[75] br[75] bl_out[18] br_out[18] sel[3] gnd single_level_column_mux_8
XXMUX76 bl[76] br[76] bl_out[19] br_out[19] sel[0] gnd single_level_column_mux_8
XXMUX77 bl[77] br[77] bl_out[19] br_out[19] sel[1] gnd single_level_column_mux_8
XXMUX78 bl[78] br[78] bl_out[19] br_out[19] sel[2] gnd single_level_column_mux_8
XXMUX79 bl[79] br[79] bl_out[19] br_out[19] sel[3] gnd single_level_column_mux_8
XXMUX80 bl[80] br[80] bl_out[20] br_out[20] sel[0] gnd single_level_column_mux_8
XXMUX81 bl[81] br[81] bl_out[20] br_out[20] sel[1] gnd single_level_column_mux_8
XXMUX82 bl[82] br[82] bl_out[20] br_out[20] sel[2] gnd single_level_column_mux_8
XXMUX83 bl[83] br[83] bl_out[20] br_out[20] sel[3] gnd single_level_column_mux_8
XXMUX84 bl[84] br[84] bl_out[21] br_out[21] sel[0] gnd single_level_column_mux_8
XXMUX85 bl[85] br[85] bl_out[21] br_out[21] sel[1] gnd single_level_column_mux_8
XXMUX86 bl[86] br[86] bl_out[21] br_out[21] sel[2] gnd single_level_column_mux_8
XXMUX87 bl[87] br[87] bl_out[21] br_out[21] sel[3] gnd single_level_column_mux_8
XXMUX88 bl[88] br[88] bl_out[22] br_out[22] sel[0] gnd single_level_column_mux_8
XXMUX89 bl[89] br[89] bl_out[22] br_out[22] sel[1] gnd single_level_column_mux_8
XXMUX90 bl[90] br[90] bl_out[22] br_out[22] sel[2] gnd single_level_column_mux_8
XXMUX91 bl[91] br[91] bl_out[22] br_out[22] sel[3] gnd single_level_column_mux_8
XXMUX92 bl[92] br[92] bl_out[23] br_out[23] sel[0] gnd single_level_column_mux_8
XXMUX93 bl[93] br[93] bl_out[23] br_out[23] sel[1] gnd single_level_column_mux_8
XXMUX94 bl[94] br[94] bl_out[23] br_out[23] sel[2] gnd single_level_column_mux_8
XXMUX95 bl[95] br[95] bl_out[23] br_out[23] sel[3] gnd single_level_column_mux_8
XXMUX96 bl[96] br[96] bl_out[24] br_out[24] sel[0] gnd single_level_column_mux_8
XXMUX97 bl[97] br[97] bl_out[24] br_out[24] sel[1] gnd single_level_column_mux_8
XXMUX98 bl[98] br[98] bl_out[24] br_out[24] sel[2] gnd single_level_column_mux_8
XXMUX99 bl[99] br[99] bl_out[24] br_out[24] sel[3] gnd single_level_column_mux_8
XXMUX100 bl[100] br[100] bl_out[25] br_out[25] sel[0] gnd single_level_column_mux_8
XXMUX101 bl[101] br[101] bl_out[25] br_out[25] sel[1] gnd single_level_column_mux_8
XXMUX102 bl[102] br[102] bl_out[25] br_out[25] sel[2] gnd single_level_column_mux_8
XXMUX103 bl[103] br[103] bl_out[25] br_out[25] sel[3] gnd single_level_column_mux_8
XXMUX104 bl[104] br[104] bl_out[26] br_out[26] sel[0] gnd single_level_column_mux_8
XXMUX105 bl[105] br[105] bl_out[26] br_out[26] sel[1] gnd single_level_column_mux_8
XXMUX106 bl[106] br[106] bl_out[26] br_out[26] sel[2] gnd single_level_column_mux_8
XXMUX107 bl[107] br[107] bl_out[26] br_out[26] sel[3] gnd single_level_column_mux_8
XXMUX108 bl[108] br[108] bl_out[27] br_out[27] sel[0] gnd single_level_column_mux_8
XXMUX109 bl[109] br[109] bl_out[27] br_out[27] sel[1] gnd single_level_column_mux_8
XXMUX110 bl[110] br[110] bl_out[27] br_out[27] sel[2] gnd single_level_column_mux_8
XXMUX111 bl[111] br[111] bl_out[27] br_out[27] sel[3] gnd single_level_column_mux_8
XXMUX112 bl[112] br[112] bl_out[28] br_out[28] sel[0] gnd single_level_column_mux_8
XXMUX113 bl[113] br[113] bl_out[28] br_out[28] sel[1] gnd single_level_column_mux_8
XXMUX114 bl[114] br[114] bl_out[28] br_out[28] sel[2] gnd single_level_column_mux_8
XXMUX115 bl[115] br[115] bl_out[28] br_out[28] sel[3] gnd single_level_column_mux_8
XXMUX116 bl[116] br[116] bl_out[29] br_out[29] sel[0] gnd single_level_column_mux_8
XXMUX117 bl[117] br[117] bl_out[29] br_out[29] sel[1] gnd single_level_column_mux_8
XXMUX118 bl[118] br[118] bl_out[29] br_out[29] sel[2] gnd single_level_column_mux_8
XXMUX119 bl[119] br[119] bl_out[29] br_out[29] sel[3] gnd single_level_column_mux_8
XXMUX120 bl[120] br[120] bl_out[30] br_out[30] sel[0] gnd single_level_column_mux_8
XXMUX121 bl[121] br[121] bl_out[30] br_out[30] sel[1] gnd single_level_column_mux_8
XXMUX122 bl[122] br[122] bl_out[30] br_out[30] sel[2] gnd single_level_column_mux_8
XXMUX123 bl[123] br[123] bl_out[30] br_out[30] sel[3] gnd single_level_column_mux_8
XXMUX124 bl[124] br[124] bl_out[31] br_out[31] sel[0] gnd single_level_column_mux_8
XXMUX125 bl[125] br[125] bl_out[31] br_out[31] sel[1] gnd single_level_column_mux_8
XXMUX126 bl[126] br[126] bl_out[31] br_out[31] sel[2] gnd single_level_column_mux_8
XXMUX127 bl[127] br[127] bl_out[31] br_out[31] sel[3] gnd single_level_column_mux_8
.ENDS columnmux_array

.SUBCKT sense_amp bl br dout en vdd gnd
M_1 dout net_1 vdd vdd pmos_vtg w=540.0n l=50.0n
M_3 net_1 dout vdd vdd pmos_vtg w=540.0n l=50.0n
M_2 dout net_1 net_2 gnd nmos_vtg w=270.0n l=50.0n
M_8 net_1 dout net_2 gnd nmos_vtg w=270.0n l=50.0n
M_5 bl en dout vdd pmos_vtg w=720.0n l=50.0n
M_6 br en net_1 vdd pmos_vtg w=720.0n l=50.0n
M_7 net_2 en gnd gnd nmos_vtg w=270.0n l=50.0n
.ENDS sense_amp


.SUBCKT sense_amp_array data[0] bl[0] br[0] data[1] bl[4] br[4] data[2] bl[8] br[8] data[3] bl[12] br[12] data[4] bl[16] br[16] data[5] bl[20] br[20] data[6] bl[24] br[24] data[7] bl[28] br[28] data[8] bl[32] br[32] data[9] bl[36] br[36] data[10] bl[40] br[40] data[11] bl[44] br[44] data[12] bl[48] br[48] data[13] bl[52] br[52] data[14] bl[56] br[56] data[15] bl[60] br[60] data[16] bl[64] br[64] data[17] bl[68] br[68] data[18] bl[72] br[72] data[19] bl[76] br[76] data[20] bl[80] br[80] data[21] bl[84] br[84] data[22] bl[88] br[88] data[23] bl[92] br[92] data[24] bl[96] br[96] data[25] bl[100] br[100] data[26] bl[104] br[104] data[27] bl[108] br[108] data[28] bl[112] br[112] data[29] bl[116] br[116] data[30] bl[120] br[120] data[31] bl[124] br[124] en vdd gnd
Xsa_d0 bl[0] br[0] data[0] en vdd gnd sense_amp
Xsa_d4 bl[4] br[4] data[1] en vdd gnd sense_amp
Xsa_d8 bl[8] br[8] data[2] en vdd gnd sense_amp
Xsa_d12 bl[12] br[12] data[3] en vdd gnd sense_amp
Xsa_d16 bl[16] br[16] data[4] en vdd gnd sense_amp
Xsa_d20 bl[20] br[20] data[5] en vdd gnd sense_amp
Xsa_d24 bl[24] br[24] data[6] en vdd gnd sense_amp
Xsa_d28 bl[28] br[28] data[7] en vdd gnd sense_amp
Xsa_d32 bl[32] br[32] data[8] en vdd gnd sense_amp
Xsa_d36 bl[36] br[36] data[9] en vdd gnd sense_amp
Xsa_d40 bl[40] br[40] data[10] en vdd gnd sense_amp
Xsa_d44 bl[44] br[44] data[11] en vdd gnd sense_amp
Xsa_d48 bl[48] br[48] data[12] en vdd gnd sense_amp
Xsa_d52 bl[52] br[52] data[13] en vdd gnd sense_amp
Xsa_d56 bl[56] br[56] data[14] en vdd gnd sense_amp
Xsa_d60 bl[60] br[60] data[15] en vdd gnd sense_amp
Xsa_d64 bl[64] br[64] data[16] en vdd gnd sense_amp
Xsa_d68 bl[68] br[68] data[17] en vdd gnd sense_amp
Xsa_d72 bl[72] br[72] data[18] en vdd gnd sense_amp
Xsa_d76 bl[76] br[76] data[19] en vdd gnd sense_amp
Xsa_d80 bl[80] br[80] data[20] en vdd gnd sense_amp
Xsa_d84 bl[84] br[84] data[21] en vdd gnd sense_amp
Xsa_d88 bl[88] br[88] data[22] en vdd gnd sense_amp
Xsa_d92 bl[92] br[92] data[23] en vdd gnd sense_amp
Xsa_d96 bl[96] br[96] data[24] en vdd gnd sense_amp
Xsa_d100 bl[100] br[100] data[25] en vdd gnd sense_amp
Xsa_d104 bl[104] br[104] data[26] en vdd gnd sense_amp
Xsa_d108 bl[108] br[108] data[27] en vdd gnd sense_amp
Xsa_d112 bl[112] br[112] data[28] en vdd gnd sense_amp
Xsa_d116 bl[116] br[116] data[29] en vdd gnd sense_amp
Xsa_d120 bl[120] br[120] data[30] en vdd gnd sense_amp
Xsa_d124 bl[124] br[124] data[31] en vdd gnd sense_amp
.ENDS sense_amp_array

.SUBCKT write_driver din bl br en vdd gnd
*inverters for enable and data input
minP bl_bar din vdd vdd pmos_vtg w=360.000000n l=50.000000n
minN bl_bar din gnd gnd nmos_vtg w=180.000000n l=50.000000n
moutP en_bar en vdd vdd pmos_vtg w=360.000000n l=50.000000n
moutN en_bar en gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BL
mout0P int1 bl_bar vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout0P2 bl en_bar int1 vdd pmos_vtg w=360.000000n l=50.000000n
mout0N bl en int2 gnd nmos_vtg w=180.000000n l=50.000000n
mout0N2 int2 bl_bar gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BR
mout1P int3 din vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout1P2 br en_bar int3 vdd pmos_vtg w=360.000000n l=50.000000n
mout1N br en int4 gnd nmos_vtg w=180.000000n l=50.000000n
mout1N2 int4 din gnd gnd nmos_vtg w=180.000000n l=50.000000n
.ENDS write_driver


.SUBCKT write_driver_array data[0] data[1] data[2] data[3] data[4] data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] data[29] data[30] data[31] bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] en vdd gnd
XXwrite_driver0 data[0] bl[0] br[0] en vdd gnd write_driver
XXwrite_driver4 data[1] bl[1] br[1] en vdd gnd write_driver
XXwrite_driver8 data[2] bl[2] br[2] en vdd gnd write_driver
XXwrite_driver12 data[3] bl[3] br[3] en vdd gnd write_driver
XXwrite_driver16 data[4] bl[4] br[4] en vdd gnd write_driver
XXwrite_driver20 data[5] bl[5] br[5] en vdd gnd write_driver
XXwrite_driver24 data[6] bl[6] br[6] en vdd gnd write_driver
XXwrite_driver28 data[7] bl[7] br[7] en vdd gnd write_driver
XXwrite_driver32 data[8] bl[8] br[8] en vdd gnd write_driver
XXwrite_driver36 data[9] bl[9] br[9] en vdd gnd write_driver
XXwrite_driver40 data[10] bl[10] br[10] en vdd gnd write_driver
XXwrite_driver44 data[11] bl[11] br[11] en vdd gnd write_driver
XXwrite_driver48 data[12] bl[12] br[12] en vdd gnd write_driver
XXwrite_driver52 data[13] bl[13] br[13] en vdd gnd write_driver
XXwrite_driver56 data[14] bl[14] br[14] en vdd gnd write_driver
XXwrite_driver60 data[15] bl[15] br[15] en vdd gnd write_driver
XXwrite_driver64 data[16] bl[16] br[16] en vdd gnd write_driver
XXwrite_driver68 data[17] bl[17] br[17] en vdd gnd write_driver
XXwrite_driver72 data[18] bl[18] br[18] en vdd gnd write_driver
XXwrite_driver76 data[19] bl[19] br[19] en vdd gnd write_driver
XXwrite_driver80 data[20] bl[20] br[20] en vdd gnd write_driver
XXwrite_driver84 data[21] bl[21] br[21] en vdd gnd write_driver
XXwrite_driver88 data[22] bl[22] br[22] en vdd gnd write_driver
XXwrite_driver92 data[23] bl[23] br[23] en vdd gnd write_driver
XXwrite_driver96 data[24] bl[24] br[24] en vdd gnd write_driver
XXwrite_driver100 data[25] bl[25] br[25] en vdd gnd write_driver
XXwrite_driver104 data[26] bl[26] br[26] en vdd gnd write_driver
XXwrite_driver108 data[27] bl[27] br[27] en vdd gnd write_driver
XXwrite_driver112 data[28] bl[28] br[28] en vdd gnd write_driver
XXwrite_driver116 data[29] bl[29] br[29] en vdd gnd write_driver
XXwrite_driver120 data[30] bl[30] br[30] en vdd gnd write_driver
XXwrite_driver124 data[31] bl[31] br[31] en vdd gnd write_driver
.ENDS write_driver_array

.SUBCKT pinv_8 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_8

.SUBCKT pnand2_2 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand2_2

.SUBCKT pnand3_2 A B C Z vdd gnd
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand3_2

.SUBCKT pinv_9 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_9

.SUBCKT pnand2_3 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand2_3

.SUBCKT pre2x4 in[0] in[1] out[0] out[1] out[2] out[3] vdd gnd
XXpre_inv[0] in[0] inbar[0] vdd gnd pinv_9
XXpre_inv[1] in[1] inbar[1] vdd gnd pinv_9
XXpre_nand_inv[0] Z[0] out[0] vdd gnd pinv_9
XXpre_nand_inv[1] Z[1] out[1] vdd gnd pinv_9
XXpre_nand_inv[2] Z[2] out[2] vdd gnd pinv_9
XXpre_nand_inv[3] Z[3] out[3] vdd gnd pinv_9
XXpre2x4_nand[0] inbar[0] inbar[1] Z[0] vdd gnd pnand2_3
XXpre2x4_nand[1] in[0] inbar[1] Z[1] vdd gnd pnand2_3
XXpre2x4_nand[2] inbar[0] in[1] Z[2] vdd gnd pnand2_3
XXpre2x4_nand[3] in[0] in[1] Z[3] vdd gnd pnand2_3
.ENDS pre2x4

.SUBCKT pinv_10 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_10

.SUBCKT pnand3_3 A B C Z vdd gnd
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand3_3

.SUBCKT pre3x8 in[0] in[1] in[2] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] vdd gnd
XXpre_inv[0] in[0] inbar[0] vdd gnd pinv_10
XXpre_inv[1] in[1] inbar[1] vdd gnd pinv_10
XXpre_inv[2] in[2] inbar[2] vdd gnd pinv_10
XXpre_nand_inv[0] Z[0] out[0] vdd gnd pinv_10
XXpre_nand_inv[1] Z[1] out[1] vdd gnd pinv_10
XXpre_nand_inv[2] Z[2] out[2] vdd gnd pinv_10
XXpre_nand_inv[3] Z[3] out[3] vdd gnd pinv_10
XXpre_nand_inv[4] Z[4] out[4] vdd gnd pinv_10
XXpre_nand_inv[5] Z[5] out[5] vdd gnd pinv_10
XXpre_nand_inv[6] Z[6] out[6] vdd gnd pinv_10
XXpre_nand_inv[7] Z[7] out[7] vdd gnd pinv_10
XXpre3x8_nand[0] inbar[0] inbar[1] inbar[2] Z[0] vdd gnd pnand3_3
XXpre3x8_nand[1] in[0] inbar[1] inbar[2] Z[1] vdd gnd pnand3_3
XXpre3x8_nand[2] inbar[0] in[1] inbar[2] Z[2] vdd gnd pnand3_3
XXpre3x8_nand[3] in[0] in[1] inbar[2] Z[3] vdd gnd pnand3_3
XXpre3x8_nand[4] inbar[0] inbar[1] in[2] Z[4] vdd gnd pnand3_3
XXpre3x8_nand[5] in[0] inbar[1] in[2] Z[5] vdd gnd pnand3_3
XXpre3x8_nand[6] inbar[0] in[1] in[2] Z[6] vdd gnd pnand3_3
XXpre3x8_nand[7] in[0] in[1] in[2] Z[7] vdd gnd pnand3_3
.ENDS pre3x8

.SUBCKT hierarchical_decoder_256rows A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] decode[0] decode[1] decode[2] decode[3] decode[4] decode[5] decode[6] decode[7] decode[8] decode[9] decode[10] decode[11] decode[12] decode[13] decode[14] decode[15] decode[16] decode[17] decode[18] decode[19] decode[20] decode[21] decode[22] decode[23] decode[24] decode[25] decode[26] decode[27] decode[28] decode[29] decode[30] decode[31] decode[32] decode[33] decode[34] decode[35] decode[36] decode[37] decode[38] decode[39] decode[40] decode[41] decode[42] decode[43] decode[44] decode[45] decode[46] decode[47] decode[48] decode[49] decode[50] decode[51] decode[52] decode[53] decode[54] decode[55] decode[56] decode[57] decode[58] decode[59] decode[60] decode[61] decode[62] decode[63] decode[64] decode[65] decode[66] decode[67] decode[68] decode[69] decode[70] decode[71] decode[72] decode[73] decode[74] decode[75] decode[76] decode[77] decode[78] decode[79] decode[80] decode[81] decode[82] decode[83] decode[84] decode[85] decode[86] decode[87] decode[88] decode[89] decode[90] decode[91] decode[92] decode[93] decode[94] decode[95] decode[96] decode[97] decode[98] decode[99] decode[100] decode[101] decode[102] decode[103] decode[104] decode[105] decode[106] decode[107] decode[108] decode[109] decode[110] decode[111] decode[112] decode[113] decode[114] decode[115] decode[116] decode[117] decode[118] decode[119] decode[120] decode[121] decode[122] decode[123] decode[124] decode[125] decode[126] decode[127] decode[128] decode[129] decode[130] decode[131] decode[132] decode[133] decode[134] decode[135] decode[136] decode[137] decode[138] decode[139] decode[140] decode[141] decode[142] decode[143] decode[144] decode[145] decode[146] decode[147] decode[148] decode[149] decode[150] decode[151] decode[152] decode[153] decode[154] decode[155] decode[156] decode[157] decode[158] decode[159] decode[160] decode[161] decode[162] decode[163] decode[164] decode[165] decode[166] decode[167] decode[168] decode[169] decode[170] decode[171] decode[172] decode[173] decode[174] decode[175] decode[176] decode[177] decode[178] decode[179] decode[180] decode[181] decode[182] decode[183] decode[184] decode[185] decode[186] decode[187] decode[188] decode[189] decode[190] decode[191] decode[192] decode[193] decode[194] decode[195] decode[196] decode[197] decode[198] decode[199] decode[200] decode[201] decode[202] decode[203] decode[204] decode[205] decode[206] decode[207] decode[208] decode[209] decode[210] decode[211] decode[212] decode[213] decode[214] decode[215] decode[216] decode[217] decode[218] decode[219] decode[220] decode[221] decode[222] decode[223] decode[224] decode[225] decode[226] decode[227] decode[228] decode[229] decode[230] decode[231] decode[232] decode[233] decode[234] decode[235] decode[236] decode[237] decode[238] decode[239] decode[240] decode[241] decode[242] decode[243] decode[244] decode[245] decode[246] decode[247] decode[248] decode[249] decode[250] decode[251] decode[252] decode[253] decode[254] decode[255] vdd gnd
Xpre[0] A[0] A[1] out[0] out[1] out[2] out[3] vdd gnd pre2x4
Xpre3x8[0] A[2] A[3] A[4] out[4] out[5] out[6] out[7] out[8] out[9] out[10] out[11] vdd gnd pre3x8
Xpre3x8[1] A[5] A[6] A[7] out[12] out[13] out[14] out[15] out[16] out[17] out[18] out[19] vdd gnd pre3x8
XDEC_NAND[0] out[0] out[4] out[12] Z[0] vdd gnd pnand3_2
XDEC_NAND[1] out[0] out[4] out[13] Z[1] vdd gnd pnand3_2
XDEC_NAND[2] out[0] out[4] out[14] Z[2] vdd gnd pnand3_2
XDEC_NAND[3] out[0] out[4] out[15] Z[3] vdd gnd pnand3_2
XDEC_NAND[4] out[0] out[4] out[16] Z[4] vdd gnd pnand3_2
XDEC_NAND[5] out[0] out[4] out[17] Z[5] vdd gnd pnand3_2
XDEC_NAND[6] out[0] out[4] out[18] Z[6] vdd gnd pnand3_2
XDEC_NAND[7] out[0] out[4] out[19] Z[7] vdd gnd pnand3_2
XDEC_NAND[8] out[0] out[5] out[12] Z[8] vdd gnd pnand3_2
XDEC_NAND[9] out[0] out[5] out[13] Z[9] vdd gnd pnand3_2
XDEC_NAND[10] out[0] out[5] out[14] Z[10] vdd gnd pnand3_2
XDEC_NAND[11] out[0] out[5] out[15] Z[11] vdd gnd pnand3_2
XDEC_NAND[12] out[0] out[5] out[16] Z[12] vdd gnd pnand3_2
XDEC_NAND[13] out[0] out[5] out[17] Z[13] vdd gnd pnand3_2
XDEC_NAND[14] out[0] out[5] out[18] Z[14] vdd gnd pnand3_2
XDEC_NAND[15] out[0] out[5] out[19] Z[15] vdd gnd pnand3_2
XDEC_NAND[16] out[0] out[6] out[12] Z[16] vdd gnd pnand3_2
XDEC_NAND[17] out[0] out[6] out[13] Z[17] vdd gnd pnand3_2
XDEC_NAND[18] out[0] out[6] out[14] Z[18] vdd gnd pnand3_2
XDEC_NAND[19] out[0] out[6] out[15] Z[19] vdd gnd pnand3_2
XDEC_NAND[20] out[0] out[6] out[16] Z[20] vdd gnd pnand3_2
XDEC_NAND[21] out[0] out[6] out[17] Z[21] vdd gnd pnand3_2
XDEC_NAND[22] out[0] out[6] out[18] Z[22] vdd gnd pnand3_2
XDEC_NAND[23] out[0] out[6] out[19] Z[23] vdd gnd pnand3_2
XDEC_NAND[24] out[0] out[7] out[12] Z[24] vdd gnd pnand3_2
XDEC_NAND[25] out[0] out[7] out[13] Z[25] vdd gnd pnand3_2
XDEC_NAND[26] out[0] out[7] out[14] Z[26] vdd gnd pnand3_2
XDEC_NAND[27] out[0] out[7] out[15] Z[27] vdd gnd pnand3_2
XDEC_NAND[28] out[0] out[7] out[16] Z[28] vdd gnd pnand3_2
XDEC_NAND[29] out[0] out[7] out[17] Z[29] vdd gnd pnand3_2
XDEC_NAND[30] out[0] out[7] out[18] Z[30] vdd gnd pnand3_2
XDEC_NAND[31] out[0] out[7] out[19] Z[31] vdd gnd pnand3_2
XDEC_NAND[32] out[0] out[8] out[12] Z[32] vdd gnd pnand3_2
XDEC_NAND[33] out[0] out[8] out[13] Z[33] vdd gnd pnand3_2
XDEC_NAND[34] out[0] out[8] out[14] Z[34] vdd gnd pnand3_2
XDEC_NAND[35] out[0] out[8] out[15] Z[35] vdd gnd pnand3_2
XDEC_NAND[36] out[0] out[8] out[16] Z[36] vdd gnd pnand3_2
XDEC_NAND[37] out[0] out[8] out[17] Z[37] vdd gnd pnand3_2
XDEC_NAND[38] out[0] out[8] out[18] Z[38] vdd gnd pnand3_2
XDEC_NAND[39] out[0] out[8] out[19] Z[39] vdd gnd pnand3_2
XDEC_NAND[40] out[0] out[9] out[12] Z[40] vdd gnd pnand3_2
XDEC_NAND[41] out[0] out[9] out[13] Z[41] vdd gnd pnand3_2
XDEC_NAND[42] out[0] out[9] out[14] Z[42] vdd gnd pnand3_2
XDEC_NAND[43] out[0] out[9] out[15] Z[43] vdd gnd pnand3_2
XDEC_NAND[44] out[0] out[9] out[16] Z[44] vdd gnd pnand3_2
XDEC_NAND[45] out[0] out[9] out[17] Z[45] vdd gnd pnand3_2
XDEC_NAND[46] out[0] out[9] out[18] Z[46] vdd gnd pnand3_2
XDEC_NAND[47] out[0] out[9] out[19] Z[47] vdd gnd pnand3_2
XDEC_NAND[48] out[0] out[10] out[12] Z[48] vdd gnd pnand3_2
XDEC_NAND[49] out[0] out[10] out[13] Z[49] vdd gnd pnand3_2
XDEC_NAND[50] out[0] out[10] out[14] Z[50] vdd gnd pnand3_2
XDEC_NAND[51] out[0] out[10] out[15] Z[51] vdd gnd pnand3_2
XDEC_NAND[52] out[0] out[10] out[16] Z[52] vdd gnd pnand3_2
XDEC_NAND[53] out[0] out[10] out[17] Z[53] vdd gnd pnand3_2
XDEC_NAND[54] out[0] out[10] out[18] Z[54] vdd gnd pnand3_2
XDEC_NAND[55] out[0] out[10] out[19] Z[55] vdd gnd pnand3_2
XDEC_NAND[56] out[0] out[11] out[12] Z[56] vdd gnd pnand3_2
XDEC_NAND[57] out[0] out[11] out[13] Z[57] vdd gnd pnand3_2
XDEC_NAND[58] out[0] out[11] out[14] Z[58] vdd gnd pnand3_2
XDEC_NAND[59] out[0] out[11] out[15] Z[59] vdd gnd pnand3_2
XDEC_NAND[60] out[0] out[11] out[16] Z[60] vdd gnd pnand3_2
XDEC_NAND[61] out[0] out[11] out[17] Z[61] vdd gnd pnand3_2
XDEC_NAND[62] out[0] out[11] out[18] Z[62] vdd gnd pnand3_2
XDEC_NAND[63] out[0] out[11] out[19] Z[63] vdd gnd pnand3_2
XDEC_NAND[64] out[1] out[4] out[12] Z[64] vdd gnd pnand3_2
XDEC_NAND[65] out[1] out[4] out[13] Z[65] vdd gnd pnand3_2
XDEC_NAND[66] out[1] out[4] out[14] Z[66] vdd gnd pnand3_2
XDEC_NAND[67] out[1] out[4] out[15] Z[67] vdd gnd pnand3_2
XDEC_NAND[68] out[1] out[4] out[16] Z[68] vdd gnd pnand3_2
XDEC_NAND[69] out[1] out[4] out[17] Z[69] vdd gnd pnand3_2
XDEC_NAND[70] out[1] out[4] out[18] Z[70] vdd gnd pnand3_2
XDEC_NAND[71] out[1] out[4] out[19] Z[71] vdd gnd pnand3_2
XDEC_NAND[72] out[1] out[5] out[12] Z[72] vdd gnd pnand3_2
XDEC_NAND[73] out[1] out[5] out[13] Z[73] vdd gnd pnand3_2
XDEC_NAND[74] out[1] out[5] out[14] Z[74] vdd gnd pnand3_2
XDEC_NAND[75] out[1] out[5] out[15] Z[75] vdd gnd pnand3_2
XDEC_NAND[76] out[1] out[5] out[16] Z[76] vdd gnd pnand3_2
XDEC_NAND[77] out[1] out[5] out[17] Z[77] vdd gnd pnand3_2
XDEC_NAND[78] out[1] out[5] out[18] Z[78] vdd gnd pnand3_2
XDEC_NAND[79] out[1] out[5] out[19] Z[79] vdd gnd pnand3_2
XDEC_NAND[80] out[1] out[6] out[12] Z[80] vdd gnd pnand3_2
XDEC_NAND[81] out[1] out[6] out[13] Z[81] vdd gnd pnand3_2
XDEC_NAND[82] out[1] out[6] out[14] Z[82] vdd gnd pnand3_2
XDEC_NAND[83] out[1] out[6] out[15] Z[83] vdd gnd pnand3_2
XDEC_NAND[84] out[1] out[6] out[16] Z[84] vdd gnd pnand3_2
XDEC_NAND[85] out[1] out[6] out[17] Z[85] vdd gnd pnand3_2
XDEC_NAND[86] out[1] out[6] out[18] Z[86] vdd gnd pnand3_2
XDEC_NAND[87] out[1] out[6] out[19] Z[87] vdd gnd pnand3_2
XDEC_NAND[88] out[1] out[7] out[12] Z[88] vdd gnd pnand3_2
XDEC_NAND[89] out[1] out[7] out[13] Z[89] vdd gnd pnand3_2
XDEC_NAND[90] out[1] out[7] out[14] Z[90] vdd gnd pnand3_2
XDEC_NAND[91] out[1] out[7] out[15] Z[91] vdd gnd pnand3_2
XDEC_NAND[92] out[1] out[7] out[16] Z[92] vdd gnd pnand3_2
XDEC_NAND[93] out[1] out[7] out[17] Z[93] vdd gnd pnand3_2
XDEC_NAND[94] out[1] out[7] out[18] Z[94] vdd gnd pnand3_2
XDEC_NAND[95] out[1] out[7] out[19] Z[95] vdd gnd pnand3_2
XDEC_NAND[96] out[1] out[8] out[12] Z[96] vdd gnd pnand3_2
XDEC_NAND[97] out[1] out[8] out[13] Z[97] vdd gnd pnand3_2
XDEC_NAND[98] out[1] out[8] out[14] Z[98] vdd gnd pnand3_2
XDEC_NAND[99] out[1] out[8] out[15] Z[99] vdd gnd pnand3_2
XDEC_NAND[100] out[1] out[8] out[16] Z[100] vdd gnd pnand3_2
XDEC_NAND[101] out[1] out[8] out[17] Z[101] vdd gnd pnand3_2
XDEC_NAND[102] out[1] out[8] out[18] Z[102] vdd gnd pnand3_2
XDEC_NAND[103] out[1] out[8] out[19] Z[103] vdd gnd pnand3_2
XDEC_NAND[104] out[1] out[9] out[12] Z[104] vdd gnd pnand3_2
XDEC_NAND[105] out[1] out[9] out[13] Z[105] vdd gnd pnand3_2
XDEC_NAND[106] out[1] out[9] out[14] Z[106] vdd gnd pnand3_2
XDEC_NAND[107] out[1] out[9] out[15] Z[107] vdd gnd pnand3_2
XDEC_NAND[108] out[1] out[9] out[16] Z[108] vdd gnd pnand3_2
XDEC_NAND[109] out[1] out[9] out[17] Z[109] vdd gnd pnand3_2
XDEC_NAND[110] out[1] out[9] out[18] Z[110] vdd gnd pnand3_2
XDEC_NAND[111] out[1] out[9] out[19] Z[111] vdd gnd pnand3_2
XDEC_NAND[112] out[1] out[10] out[12] Z[112] vdd gnd pnand3_2
XDEC_NAND[113] out[1] out[10] out[13] Z[113] vdd gnd pnand3_2
XDEC_NAND[114] out[1] out[10] out[14] Z[114] vdd gnd pnand3_2
XDEC_NAND[115] out[1] out[10] out[15] Z[115] vdd gnd pnand3_2
XDEC_NAND[116] out[1] out[10] out[16] Z[116] vdd gnd pnand3_2
XDEC_NAND[117] out[1] out[10] out[17] Z[117] vdd gnd pnand3_2
XDEC_NAND[118] out[1] out[10] out[18] Z[118] vdd gnd pnand3_2
XDEC_NAND[119] out[1] out[10] out[19] Z[119] vdd gnd pnand3_2
XDEC_NAND[120] out[1] out[11] out[12] Z[120] vdd gnd pnand3_2
XDEC_NAND[121] out[1] out[11] out[13] Z[121] vdd gnd pnand3_2
XDEC_NAND[122] out[1] out[11] out[14] Z[122] vdd gnd pnand3_2
XDEC_NAND[123] out[1] out[11] out[15] Z[123] vdd gnd pnand3_2
XDEC_NAND[124] out[1] out[11] out[16] Z[124] vdd gnd pnand3_2
XDEC_NAND[125] out[1] out[11] out[17] Z[125] vdd gnd pnand3_2
XDEC_NAND[126] out[1] out[11] out[18] Z[126] vdd gnd pnand3_2
XDEC_NAND[127] out[1] out[11] out[19] Z[127] vdd gnd pnand3_2
XDEC_NAND[128] out[2] out[4] out[12] Z[128] vdd gnd pnand3_2
XDEC_NAND[129] out[2] out[4] out[13] Z[129] vdd gnd pnand3_2
XDEC_NAND[130] out[2] out[4] out[14] Z[130] vdd gnd pnand3_2
XDEC_NAND[131] out[2] out[4] out[15] Z[131] vdd gnd pnand3_2
XDEC_NAND[132] out[2] out[4] out[16] Z[132] vdd gnd pnand3_2
XDEC_NAND[133] out[2] out[4] out[17] Z[133] vdd gnd pnand3_2
XDEC_NAND[134] out[2] out[4] out[18] Z[134] vdd gnd pnand3_2
XDEC_NAND[135] out[2] out[4] out[19] Z[135] vdd gnd pnand3_2
XDEC_NAND[136] out[2] out[5] out[12] Z[136] vdd gnd pnand3_2
XDEC_NAND[137] out[2] out[5] out[13] Z[137] vdd gnd pnand3_2
XDEC_NAND[138] out[2] out[5] out[14] Z[138] vdd gnd pnand3_2
XDEC_NAND[139] out[2] out[5] out[15] Z[139] vdd gnd pnand3_2
XDEC_NAND[140] out[2] out[5] out[16] Z[140] vdd gnd pnand3_2
XDEC_NAND[141] out[2] out[5] out[17] Z[141] vdd gnd pnand3_2
XDEC_NAND[142] out[2] out[5] out[18] Z[142] vdd gnd pnand3_2
XDEC_NAND[143] out[2] out[5] out[19] Z[143] vdd gnd pnand3_2
XDEC_NAND[144] out[2] out[6] out[12] Z[144] vdd gnd pnand3_2
XDEC_NAND[145] out[2] out[6] out[13] Z[145] vdd gnd pnand3_2
XDEC_NAND[146] out[2] out[6] out[14] Z[146] vdd gnd pnand3_2
XDEC_NAND[147] out[2] out[6] out[15] Z[147] vdd gnd pnand3_2
XDEC_NAND[148] out[2] out[6] out[16] Z[148] vdd gnd pnand3_2
XDEC_NAND[149] out[2] out[6] out[17] Z[149] vdd gnd pnand3_2
XDEC_NAND[150] out[2] out[6] out[18] Z[150] vdd gnd pnand3_2
XDEC_NAND[151] out[2] out[6] out[19] Z[151] vdd gnd pnand3_2
XDEC_NAND[152] out[2] out[7] out[12] Z[152] vdd gnd pnand3_2
XDEC_NAND[153] out[2] out[7] out[13] Z[153] vdd gnd pnand3_2
XDEC_NAND[154] out[2] out[7] out[14] Z[154] vdd gnd pnand3_2
XDEC_NAND[155] out[2] out[7] out[15] Z[155] vdd gnd pnand3_2
XDEC_NAND[156] out[2] out[7] out[16] Z[156] vdd gnd pnand3_2
XDEC_NAND[157] out[2] out[7] out[17] Z[157] vdd gnd pnand3_2
XDEC_NAND[158] out[2] out[7] out[18] Z[158] vdd gnd pnand3_2
XDEC_NAND[159] out[2] out[7] out[19] Z[159] vdd gnd pnand3_2
XDEC_NAND[160] out[2] out[8] out[12] Z[160] vdd gnd pnand3_2
XDEC_NAND[161] out[2] out[8] out[13] Z[161] vdd gnd pnand3_2
XDEC_NAND[162] out[2] out[8] out[14] Z[162] vdd gnd pnand3_2
XDEC_NAND[163] out[2] out[8] out[15] Z[163] vdd gnd pnand3_2
XDEC_NAND[164] out[2] out[8] out[16] Z[164] vdd gnd pnand3_2
XDEC_NAND[165] out[2] out[8] out[17] Z[165] vdd gnd pnand3_2
XDEC_NAND[166] out[2] out[8] out[18] Z[166] vdd gnd pnand3_2
XDEC_NAND[167] out[2] out[8] out[19] Z[167] vdd gnd pnand3_2
XDEC_NAND[168] out[2] out[9] out[12] Z[168] vdd gnd pnand3_2
XDEC_NAND[169] out[2] out[9] out[13] Z[169] vdd gnd pnand3_2
XDEC_NAND[170] out[2] out[9] out[14] Z[170] vdd gnd pnand3_2
XDEC_NAND[171] out[2] out[9] out[15] Z[171] vdd gnd pnand3_2
XDEC_NAND[172] out[2] out[9] out[16] Z[172] vdd gnd pnand3_2
XDEC_NAND[173] out[2] out[9] out[17] Z[173] vdd gnd pnand3_2
XDEC_NAND[174] out[2] out[9] out[18] Z[174] vdd gnd pnand3_2
XDEC_NAND[175] out[2] out[9] out[19] Z[175] vdd gnd pnand3_2
XDEC_NAND[176] out[2] out[10] out[12] Z[176] vdd gnd pnand3_2
XDEC_NAND[177] out[2] out[10] out[13] Z[177] vdd gnd pnand3_2
XDEC_NAND[178] out[2] out[10] out[14] Z[178] vdd gnd pnand3_2
XDEC_NAND[179] out[2] out[10] out[15] Z[179] vdd gnd pnand3_2
XDEC_NAND[180] out[2] out[10] out[16] Z[180] vdd gnd pnand3_2
XDEC_NAND[181] out[2] out[10] out[17] Z[181] vdd gnd pnand3_2
XDEC_NAND[182] out[2] out[10] out[18] Z[182] vdd gnd pnand3_2
XDEC_NAND[183] out[2] out[10] out[19] Z[183] vdd gnd pnand3_2
XDEC_NAND[184] out[2] out[11] out[12] Z[184] vdd gnd pnand3_2
XDEC_NAND[185] out[2] out[11] out[13] Z[185] vdd gnd pnand3_2
XDEC_NAND[186] out[2] out[11] out[14] Z[186] vdd gnd pnand3_2
XDEC_NAND[187] out[2] out[11] out[15] Z[187] vdd gnd pnand3_2
XDEC_NAND[188] out[2] out[11] out[16] Z[188] vdd gnd pnand3_2
XDEC_NAND[189] out[2] out[11] out[17] Z[189] vdd gnd pnand3_2
XDEC_NAND[190] out[2] out[11] out[18] Z[190] vdd gnd pnand3_2
XDEC_NAND[191] out[2] out[11] out[19] Z[191] vdd gnd pnand3_2
XDEC_NAND[192] out[3] out[4] out[12] Z[192] vdd gnd pnand3_2
XDEC_NAND[193] out[3] out[4] out[13] Z[193] vdd gnd pnand3_2
XDEC_NAND[194] out[3] out[4] out[14] Z[194] vdd gnd pnand3_2
XDEC_NAND[195] out[3] out[4] out[15] Z[195] vdd gnd pnand3_2
XDEC_NAND[196] out[3] out[4] out[16] Z[196] vdd gnd pnand3_2
XDEC_NAND[197] out[3] out[4] out[17] Z[197] vdd gnd pnand3_2
XDEC_NAND[198] out[3] out[4] out[18] Z[198] vdd gnd pnand3_2
XDEC_NAND[199] out[3] out[4] out[19] Z[199] vdd gnd pnand3_2
XDEC_NAND[200] out[3] out[5] out[12] Z[200] vdd gnd pnand3_2
XDEC_NAND[201] out[3] out[5] out[13] Z[201] vdd gnd pnand3_2
XDEC_NAND[202] out[3] out[5] out[14] Z[202] vdd gnd pnand3_2
XDEC_NAND[203] out[3] out[5] out[15] Z[203] vdd gnd pnand3_2
XDEC_NAND[204] out[3] out[5] out[16] Z[204] vdd gnd pnand3_2
XDEC_NAND[205] out[3] out[5] out[17] Z[205] vdd gnd pnand3_2
XDEC_NAND[206] out[3] out[5] out[18] Z[206] vdd gnd pnand3_2
XDEC_NAND[207] out[3] out[5] out[19] Z[207] vdd gnd pnand3_2
XDEC_NAND[208] out[3] out[6] out[12] Z[208] vdd gnd pnand3_2
XDEC_NAND[209] out[3] out[6] out[13] Z[209] vdd gnd pnand3_2
XDEC_NAND[210] out[3] out[6] out[14] Z[210] vdd gnd pnand3_2
XDEC_NAND[211] out[3] out[6] out[15] Z[211] vdd gnd pnand3_2
XDEC_NAND[212] out[3] out[6] out[16] Z[212] vdd gnd pnand3_2
XDEC_NAND[213] out[3] out[6] out[17] Z[213] vdd gnd pnand3_2
XDEC_NAND[214] out[3] out[6] out[18] Z[214] vdd gnd pnand3_2
XDEC_NAND[215] out[3] out[6] out[19] Z[215] vdd gnd pnand3_2
XDEC_NAND[216] out[3] out[7] out[12] Z[216] vdd gnd pnand3_2
XDEC_NAND[217] out[3] out[7] out[13] Z[217] vdd gnd pnand3_2
XDEC_NAND[218] out[3] out[7] out[14] Z[218] vdd gnd pnand3_2
XDEC_NAND[219] out[3] out[7] out[15] Z[219] vdd gnd pnand3_2
XDEC_NAND[220] out[3] out[7] out[16] Z[220] vdd gnd pnand3_2
XDEC_NAND[221] out[3] out[7] out[17] Z[221] vdd gnd pnand3_2
XDEC_NAND[222] out[3] out[7] out[18] Z[222] vdd gnd pnand3_2
XDEC_NAND[223] out[3] out[7] out[19] Z[223] vdd gnd pnand3_2
XDEC_NAND[224] out[3] out[8] out[12] Z[224] vdd gnd pnand3_2
XDEC_NAND[225] out[3] out[8] out[13] Z[225] vdd gnd pnand3_2
XDEC_NAND[226] out[3] out[8] out[14] Z[226] vdd gnd pnand3_2
XDEC_NAND[227] out[3] out[8] out[15] Z[227] vdd gnd pnand3_2
XDEC_NAND[228] out[3] out[8] out[16] Z[228] vdd gnd pnand3_2
XDEC_NAND[229] out[3] out[8] out[17] Z[229] vdd gnd pnand3_2
XDEC_NAND[230] out[3] out[8] out[18] Z[230] vdd gnd pnand3_2
XDEC_NAND[231] out[3] out[8] out[19] Z[231] vdd gnd pnand3_2
XDEC_NAND[232] out[3] out[9] out[12] Z[232] vdd gnd pnand3_2
XDEC_NAND[233] out[3] out[9] out[13] Z[233] vdd gnd pnand3_2
XDEC_NAND[234] out[3] out[9] out[14] Z[234] vdd gnd pnand3_2
XDEC_NAND[235] out[3] out[9] out[15] Z[235] vdd gnd pnand3_2
XDEC_NAND[236] out[3] out[9] out[16] Z[236] vdd gnd pnand3_2
XDEC_NAND[237] out[3] out[9] out[17] Z[237] vdd gnd pnand3_2
XDEC_NAND[238] out[3] out[9] out[18] Z[238] vdd gnd pnand3_2
XDEC_NAND[239] out[3] out[9] out[19] Z[239] vdd gnd pnand3_2
XDEC_NAND[240] out[3] out[10] out[12] Z[240] vdd gnd pnand3_2
XDEC_NAND[241] out[3] out[10] out[13] Z[241] vdd gnd pnand3_2
XDEC_NAND[242] out[3] out[10] out[14] Z[242] vdd gnd pnand3_2
XDEC_NAND[243] out[3] out[10] out[15] Z[243] vdd gnd pnand3_2
XDEC_NAND[244] out[3] out[10] out[16] Z[244] vdd gnd pnand3_2
XDEC_NAND[245] out[3] out[10] out[17] Z[245] vdd gnd pnand3_2
XDEC_NAND[246] out[3] out[10] out[18] Z[246] vdd gnd pnand3_2
XDEC_NAND[247] out[3] out[10] out[19] Z[247] vdd gnd pnand3_2
XDEC_NAND[248] out[3] out[11] out[12] Z[248] vdd gnd pnand3_2
XDEC_NAND[249] out[3] out[11] out[13] Z[249] vdd gnd pnand3_2
XDEC_NAND[250] out[3] out[11] out[14] Z[250] vdd gnd pnand3_2
XDEC_NAND[251] out[3] out[11] out[15] Z[251] vdd gnd pnand3_2
XDEC_NAND[252] out[3] out[11] out[16] Z[252] vdd gnd pnand3_2
XDEC_NAND[253] out[3] out[11] out[17] Z[253] vdd gnd pnand3_2
XDEC_NAND[254] out[3] out[11] out[18] Z[254] vdd gnd pnand3_2
XDEC_NAND[255] out[3] out[11] out[19] Z[255] vdd gnd pnand3_2
XDEC_INV_[0] Z[0] decode[0] vdd gnd pinv_8
XDEC_INV_[1] Z[1] decode[1] vdd gnd pinv_8
XDEC_INV_[2] Z[2] decode[2] vdd gnd pinv_8
XDEC_INV_[3] Z[3] decode[3] vdd gnd pinv_8
XDEC_INV_[4] Z[4] decode[4] vdd gnd pinv_8
XDEC_INV_[5] Z[5] decode[5] vdd gnd pinv_8
XDEC_INV_[6] Z[6] decode[6] vdd gnd pinv_8
XDEC_INV_[7] Z[7] decode[7] vdd gnd pinv_8
XDEC_INV_[8] Z[8] decode[8] vdd gnd pinv_8
XDEC_INV_[9] Z[9] decode[9] vdd gnd pinv_8
XDEC_INV_[10] Z[10] decode[10] vdd gnd pinv_8
XDEC_INV_[11] Z[11] decode[11] vdd gnd pinv_8
XDEC_INV_[12] Z[12] decode[12] vdd gnd pinv_8
XDEC_INV_[13] Z[13] decode[13] vdd gnd pinv_8
XDEC_INV_[14] Z[14] decode[14] vdd gnd pinv_8
XDEC_INV_[15] Z[15] decode[15] vdd gnd pinv_8
XDEC_INV_[16] Z[16] decode[16] vdd gnd pinv_8
XDEC_INV_[17] Z[17] decode[17] vdd gnd pinv_8
XDEC_INV_[18] Z[18] decode[18] vdd gnd pinv_8
XDEC_INV_[19] Z[19] decode[19] vdd gnd pinv_8
XDEC_INV_[20] Z[20] decode[20] vdd gnd pinv_8
XDEC_INV_[21] Z[21] decode[21] vdd gnd pinv_8
XDEC_INV_[22] Z[22] decode[22] vdd gnd pinv_8
XDEC_INV_[23] Z[23] decode[23] vdd gnd pinv_8
XDEC_INV_[24] Z[24] decode[24] vdd gnd pinv_8
XDEC_INV_[25] Z[25] decode[25] vdd gnd pinv_8
XDEC_INV_[26] Z[26] decode[26] vdd gnd pinv_8
XDEC_INV_[27] Z[27] decode[27] vdd gnd pinv_8
XDEC_INV_[28] Z[28] decode[28] vdd gnd pinv_8
XDEC_INV_[29] Z[29] decode[29] vdd gnd pinv_8
XDEC_INV_[30] Z[30] decode[30] vdd gnd pinv_8
XDEC_INV_[31] Z[31] decode[31] vdd gnd pinv_8
XDEC_INV_[32] Z[32] decode[32] vdd gnd pinv_8
XDEC_INV_[33] Z[33] decode[33] vdd gnd pinv_8
XDEC_INV_[34] Z[34] decode[34] vdd gnd pinv_8
XDEC_INV_[35] Z[35] decode[35] vdd gnd pinv_8
XDEC_INV_[36] Z[36] decode[36] vdd gnd pinv_8
XDEC_INV_[37] Z[37] decode[37] vdd gnd pinv_8
XDEC_INV_[38] Z[38] decode[38] vdd gnd pinv_8
XDEC_INV_[39] Z[39] decode[39] vdd gnd pinv_8
XDEC_INV_[40] Z[40] decode[40] vdd gnd pinv_8
XDEC_INV_[41] Z[41] decode[41] vdd gnd pinv_8
XDEC_INV_[42] Z[42] decode[42] vdd gnd pinv_8
XDEC_INV_[43] Z[43] decode[43] vdd gnd pinv_8
XDEC_INV_[44] Z[44] decode[44] vdd gnd pinv_8
XDEC_INV_[45] Z[45] decode[45] vdd gnd pinv_8
XDEC_INV_[46] Z[46] decode[46] vdd gnd pinv_8
XDEC_INV_[47] Z[47] decode[47] vdd gnd pinv_8
XDEC_INV_[48] Z[48] decode[48] vdd gnd pinv_8
XDEC_INV_[49] Z[49] decode[49] vdd gnd pinv_8
XDEC_INV_[50] Z[50] decode[50] vdd gnd pinv_8
XDEC_INV_[51] Z[51] decode[51] vdd gnd pinv_8
XDEC_INV_[52] Z[52] decode[52] vdd gnd pinv_8
XDEC_INV_[53] Z[53] decode[53] vdd gnd pinv_8
XDEC_INV_[54] Z[54] decode[54] vdd gnd pinv_8
XDEC_INV_[55] Z[55] decode[55] vdd gnd pinv_8
XDEC_INV_[56] Z[56] decode[56] vdd gnd pinv_8
XDEC_INV_[57] Z[57] decode[57] vdd gnd pinv_8
XDEC_INV_[58] Z[58] decode[58] vdd gnd pinv_8
XDEC_INV_[59] Z[59] decode[59] vdd gnd pinv_8
XDEC_INV_[60] Z[60] decode[60] vdd gnd pinv_8
XDEC_INV_[61] Z[61] decode[61] vdd gnd pinv_8
XDEC_INV_[62] Z[62] decode[62] vdd gnd pinv_8
XDEC_INV_[63] Z[63] decode[63] vdd gnd pinv_8
XDEC_INV_[64] Z[64] decode[64] vdd gnd pinv_8
XDEC_INV_[65] Z[65] decode[65] vdd gnd pinv_8
XDEC_INV_[66] Z[66] decode[66] vdd gnd pinv_8
XDEC_INV_[67] Z[67] decode[67] vdd gnd pinv_8
XDEC_INV_[68] Z[68] decode[68] vdd gnd pinv_8
XDEC_INV_[69] Z[69] decode[69] vdd gnd pinv_8
XDEC_INV_[70] Z[70] decode[70] vdd gnd pinv_8
XDEC_INV_[71] Z[71] decode[71] vdd gnd pinv_8
XDEC_INV_[72] Z[72] decode[72] vdd gnd pinv_8
XDEC_INV_[73] Z[73] decode[73] vdd gnd pinv_8
XDEC_INV_[74] Z[74] decode[74] vdd gnd pinv_8
XDEC_INV_[75] Z[75] decode[75] vdd gnd pinv_8
XDEC_INV_[76] Z[76] decode[76] vdd gnd pinv_8
XDEC_INV_[77] Z[77] decode[77] vdd gnd pinv_8
XDEC_INV_[78] Z[78] decode[78] vdd gnd pinv_8
XDEC_INV_[79] Z[79] decode[79] vdd gnd pinv_8
XDEC_INV_[80] Z[80] decode[80] vdd gnd pinv_8
XDEC_INV_[81] Z[81] decode[81] vdd gnd pinv_8
XDEC_INV_[82] Z[82] decode[82] vdd gnd pinv_8
XDEC_INV_[83] Z[83] decode[83] vdd gnd pinv_8
XDEC_INV_[84] Z[84] decode[84] vdd gnd pinv_8
XDEC_INV_[85] Z[85] decode[85] vdd gnd pinv_8
XDEC_INV_[86] Z[86] decode[86] vdd gnd pinv_8
XDEC_INV_[87] Z[87] decode[87] vdd gnd pinv_8
XDEC_INV_[88] Z[88] decode[88] vdd gnd pinv_8
XDEC_INV_[89] Z[89] decode[89] vdd gnd pinv_8
XDEC_INV_[90] Z[90] decode[90] vdd gnd pinv_8
XDEC_INV_[91] Z[91] decode[91] vdd gnd pinv_8
XDEC_INV_[92] Z[92] decode[92] vdd gnd pinv_8
XDEC_INV_[93] Z[93] decode[93] vdd gnd pinv_8
XDEC_INV_[94] Z[94] decode[94] vdd gnd pinv_8
XDEC_INV_[95] Z[95] decode[95] vdd gnd pinv_8
XDEC_INV_[96] Z[96] decode[96] vdd gnd pinv_8
XDEC_INV_[97] Z[97] decode[97] vdd gnd pinv_8
XDEC_INV_[98] Z[98] decode[98] vdd gnd pinv_8
XDEC_INV_[99] Z[99] decode[99] vdd gnd pinv_8
XDEC_INV_[100] Z[100] decode[100] vdd gnd pinv_8
XDEC_INV_[101] Z[101] decode[101] vdd gnd pinv_8
XDEC_INV_[102] Z[102] decode[102] vdd gnd pinv_8
XDEC_INV_[103] Z[103] decode[103] vdd gnd pinv_8
XDEC_INV_[104] Z[104] decode[104] vdd gnd pinv_8
XDEC_INV_[105] Z[105] decode[105] vdd gnd pinv_8
XDEC_INV_[106] Z[106] decode[106] vdd gnd pinv_8
XDEC_INV_[107] Z[107] decode[107] vdd gnd pinv_8
XDEC_INV_[108] Z[108] decode[108] vdd gnd pinv_8
XDEC_INV_[109] Z[109] decode[109] vdd gnd pinv_8
XDEC_INV_[110] Z[110] decode[110] vdd gnd pinv_8
XDEC_INV_[111] Z[111] decode[111] vdd gnd pinv_8
XDEC_INV_[112] Z[112] decode[112] vdd gnd pinv_8
XDEC_INV_[113] Z[113] decode[113] vdd gnd pinv_8
XDEC_INV_[114] Z[114] decode[114] vdd gnd pinv_8
XDEC_INV_[115] Z[115] decode[115] vdd gnd pinv_8
XDEC_INV_[116] Z[116] decode[116] vdd gnd pinv_8
XDEC_INV_[117] Z[117] decode[117] vdd gnd pinv_8
XDEC_INV_[118] Z[118] decode[118] vdd gnd pinv_8
XDEC_INV_[119] Z[119] decode[119] vdd gnd pinv_8
XDEC_INV_[120] Z[120] decode[120] vdd gnd pinv_8
XDEC_INV_[121] Z[121] decode[121] vdd gnd pinv_8
XDEC_INV_[122] Z[122] decode[122] vdd gnd pinv_8
XDEC_INV_[123] Z[123] decode[123] vdd gnd pinv_8
XDEC_INV_[124] Z[124] decode[124] vdd gnd pinv_8
XDEC_INV_[125] Z[125] decode[125] vdd gnd pinv_8
XDEC_INV_[126] Z[126] decode[126] vdd gnd pinv_8
XDEC_INV_[127] Z[127] decode[127] vdd gnd pinv_8
XDEC_INV_[128] Z[128] decode[128] vdd gnd pinv_8
XDEC_INV_[129] Z[129] decode[129] vdd gnd pinv_8
XDEC_INV_[130] Z[130] decode[130] vdd gnd pinv_8
XDEC_INV_[131] Z[131] decode[131] vdd gnd pinv_8
XDEC_INV_[132] Z[132] decode[132] vdd gnd pinv_8
XDEC_INV_[133] Z[133] decode[133] vdd gnd pinv_8
XDEC_INV_[134] Z[134] decode[134] vdd gnd pinv_8
XDEC_INV_[135] Z[135] decode[135] vdd gnd pinv_8
XDEC_INV_[136] Z[136] decode[136] vdd gnd pinv_8
XDEC_INV_[137] Z[137] decode[137] vdd gnd pinv_8
XDEC_INV_[138] Z[138] decode[138] vdd gnd pinv_8
XDEC_INV_[139] Z[139] decode[139] vdd gnd pinv_8
XDEC_INV_[140] Z[140] decode[140] vdd gnd pinv_8
XDEC_INV_[141] Z[141] decode[141] vdd gnd pinv_8
XDEC_INV_[142] Z[142] decode[142] vdd gnd pinv_8
XDEC_INV_[143] Z[143] decode[143] vdd gnd pinv_8
XDEC_INV_[144] Z[144] decode[144] vdd gnd pinv_8
XDEC_INV_[145] Z[145] decode[145] vdd gnd pinv_8
XDEC_INV_[146] Z[146] decode[146] vdd gnd pinv_8
XDEC_INV_[147] Z[147] decode[147] vdd gnd pinv_8
XDEC_INV_[148] Z[148] decode[148] vdd gnd pinv_8
XDEC_INV_[149] Z[149] decode[149] vdd gnd pinv_8
XDEC_INV_[150] Z[150] decode[150] vdd gnd pinv_8
XDEC_INV_[151] Z[151] decode[151] vdd gnd pinv_8
XDEC_INV_[152] Z[152] decode[152] vdd gnd pinv_8
XDEC_INV_[153] Z[153] decode[153] vdd gnd pinv_8
XDEC_INV_[154] Z[154] decode[154] vdd gnd pinv_8
XDEC_INV_[155] Z[155] decode[155] vdd gnd pinv_8
XDEC_INV_[156] Z[156] decode[156] vdd gnd pinv_8
XDEC_INV_[157] Z[157] decode[157] vdd gnd pinv_8
XDEC_INV_[158] Z[158] decode[158] vdd gnd pinv_8
XDEC_INV_[159] Z[159] decode[159] vdd gnd pinv_8
XDEC_INV_[160] Z[160] decode[160] vdd gnd pinv_8
XDEC_INV_[161] Z[161] decode[161] vdd gnd pinv_8
XDEC_INV_[162] Z[162] decode[162] vdd gnd pinv_8
XDEC_INV_[163] Z[163] decode[163] vdd gnd pinv_8
XDEC_INV_[164] Z[164] decode[164] vdd gnd pinv_8
XDEC_INV_[165] Z[165] decode[165] vdd gnd pinv_8
XDEC_INV_[166] Z[166] decode[166] vdd gnd pinv_8
XDEC_INV_[167] Z[167] decode[167] vdd gnd pinv_8
XDEC_INV_[168] Z[168] decode[168] vdd gnd pinv_8
XDEC_INV_[169] Z[169] decode[169] vdd gnd pinv_8
XDEC_INV_[170] Z[170] decode[170] vdd gnd pinv_8
XDEC_INV_[171] Z[171] decode[171] vdd gnd pinv_8
XDEC_INV_[172] Z[172] decode[172] vdd gnd pinv_8
XDEC_INV_[173] Z[173] decode[173] vdd gnd pinv_8
XDEC_INV_[174] Z[174] decode[174] vdd gnd pinv_8
XDEC_INV_[175] Z[175] decode[175] vdd gnd pinv_8
XDEC_INV_[176] Z[176] decode[176] vdd gnd pinv_8
XDEC_INV_[177] Z[177] decode[177] vdd gnd pinv_8
XDEC_INV_[178] Z[178] decode[178] vdd gnd pinv_8
XDEC_INV_[179] Z[179] decode[179] vdd gnd pinv_8
XDEC_INV_[180] Z[180] decode[180] vdd gnd pinv_8
XDEC_INV_[181] Z[181] decode[181] vdd gnd pinv_8
XDEC_INV_[182] Z[182] decode[182] vdd gnd pinv_8
XDEC_INV_[183] Z[183] decode[183] vdd gnd pinv_8
XDEC_INV_[184] Z[184] decode[184] vdd gnd pinv_8
XDEC_INV_[185] Z[185] decode[185] vdd gnd pinv_8
XDEC_INV_[186] Z[186] decode[186] vdd gnd pinv_8
XDEC_INV_[187] Z[187] decode[187] vdd gnd pinv_8
XDEC_INV_[188] Z[188] decode[188] vdd gnd pinv_8
XDEC_INV_[189] Z[189] decode[189] vdd gnd pinv_8
XDEC_INV_[190] Z[190] decode[190] vdd gnd pinv_8
XDEC_INV_[191] Z[191] decode[191] vdd gnd pinv_8
XDEC_INV_[192] Z[192] decode[192] vdd gnd pinv_8
XDEC_INV_[193] Z[193] decode[193] vdd gnd pinv_8
XDEC_INV_[194] Z[194] decode[194] vdd gnd pinv_8
XDEC_INV_[195] Z[195] decode[195] vdd gnd pinv_8
XDEC_INV_[196] Z[196] decode[196] vdd gnd pinv_8
XDEC_INV_[197] Z[197] decode[197] vdd gnd pinv_8
XDEC_INV_[198] Z[198] decode[198] vdd gnd pinv_8
XDEC_INV_[199] Z[199] decode[199] vdd gnd pinv_8
XDEC_INV_[200] Z[200] decode[200] vdd gnd pinv_8
XDEC_INV_[201] Z[201] decode[201] vdd gnd pinv_8
XDEC_INV_[202] Z[202] decode[202] vdd gnd pinv_8
XDEC_INV_[203] Z[203] decode[203] vdd gnd pinv_8
XDEC_INV_[204] Z[204] decode[204] vdd gnd pinv_8
XDEC_INV_[205] Z[205] decode[205] vdd gnd pinv_8
XDEC_INV_[206] Z[206] decode[206] vdd gnd pinv_8
XDEC_INV_[207] Z[207] decode[207] vdd gnd pinv_8
XDEC_INV_[208] Z[208] decode[208] vdd gnd pinv_8
XDEC_INV_[209] Z[209] decode[209] vdd gnd pinv_8
XDEC_INV_[210] Z[210] decode[210] vdd gnd pinv_8
XDEC_INV_[211] Z[211] decode[211] vdd gnd pinv_8
XDEC_INV_[212] Z[212] decode[212] vdd gnd pinv_8
XDEC_INV_[213] Z[213] decode[213] vdd gnd pinv_8
XDEC_INV_[214] Z[214] decode[214] vdd gnd pinv_8
XDEC_INV_[215] Z[215] decode[215] vdd gnd pinv_8
XDEC_INV_[216] Z[216] decode[216] vdd gnd pinv_8
XDEC_INV_[217] Z[217] decode[217] vdd gnd pinv_8
XDEC_INV_[218] Z[218] decode[218] vdd gnd pinv_8
XDEC_INV_[219] Z[219] decode[219] vdd gnd pinv_8
XDEC_INV_[220] Z[220] decode[220] vdd gnd pinv_8
XDEC_INV_[221] Z[221] decode[221] vdd gnd pinv_8
XDEC_INV_[222] Z[222] decode[222] vdd gnd pinv_8
XDEC_INV_[223] Z[223] decode[223] vdd gnd pinv_8
XDEC_INV_[224] Z[224] decode[224] vdd gnd pinv_8
XDEC_INV_[225] Z[225] decode[225] vdd gnd pinv_8
XDEC_INV_[226] Z[226] decode[226] vdd gnd pinv_8
XDEC_INV_[227] Z[227] decode[227] vdd gnd pinv_8
XDEC_INV_[228] Z[228] decode[228] vdd gnd pinv_8
XDEC_INV_[229] Z[229] decode[229] vdd gnd pinv_8
XDEC_INV_[230] Z[230] decode[230] vdd gnd pinv_8
XDEC_INV_[231] Z[231] decode[231] vdd gnd pinv_8
XDEC_INV_[232] Z[232] decode[232] vdd gnd pinv_8
XDEC_INV_[233] Z[233] decode[233] vdd gnd pinv_8
XDEC_INV_[234] Z[234] decode[234] vdd gnd pinv_8
XDEC_INV_[235] Z[235] decode[235] vdd gnd pinv_8
XDEC_INV_[236] Z[236] decode[236] vdd gnd pinv_8
XDEC_INV_[237] Z[237] decode[237] vdd gnd pinv_8
XDEC_INV_[238] Z[238] decode[238] vdd gnd pinv_8
XDEC_INV_[239] Z[239] decode[239] vdd gnd pinv_8
XDEC_INV_[240] Z[240] decode[240] vdd gnd pinv_8
XDEC_INV_[241] Z[241] decode[241] vdd gnd pinv_8
XDEC_INV_[242] Z[242] decode[242] vdd gnd pinv_8
XDEC_INV_[243] Z[243] decode[243] vdd gnd pinv_8
XDEC_INV_[244] Z[244] decode[244] vdd gnd pinv_8
XDEC_INV_[245] Z[245] decode[245] vdd gnd pinv_8
XDEC_INV_[246] Z[246] decode[246] vdd gnd pinv_8
XDEC_INV_[247] Z[247] decode[247] vdd gnd pinv_8
XDEC_INV_[248] Z[248] decode[248] vdd gnd pinv_8
XDEC_INV_[249] Z[249] decode[249] vdd gnd pinv_8
XDEC_INV_[250] Z[250] decode[250] vdd gnd pinv_8
XDEC_INV_[251] Z[251] decode[251] vdd gnd pinv_8
XDEC_INV_[252] Z[252] decode[252] vdd gnd pinv_8
XDEC_INV_[253] Z[253] decode[253] vdd gnd pinv_8
XDEC_INV_[254] Z[254] decode[254] vdd gnd pinv_8
XDEC_INV_[255] Z[255] decode[255] vdd gnd pinv_8
.ENDS hierarchical_decoder_256rows

.SUBCKT msf_address din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] dout[0] dout_bar[0] dout[1] dout_bar[1] dout[2] dout_bar[2] dout[3] dout_bar[3] dout[4] dout_bar[4] dout[5] dout_bar[5] dout[6] dout_bar[6] dout[7] dout_bar[7] dout[8] dout_bar[8] dout[9] dout_bar[9] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
XXdff1 din[1] dout[1] dout_bar[1] clk vdd gnd ms_flop
XXdff2 din[2] dout[2] dout_bar[2] clk vdd gnd ms_flop
XXdff3 din[3] dout[3] dout_bar[3] clk vdd gnd ms_flop
XXdff4 din[4] dout[4] dout_bar[4] clk vdd gnd ms_flop
XXdff5 din[5] dout[5] dout_bar[5] clk vdd gnd ms_flop
XXdff6 din[6] dout[6] dout_bar[6] clk vdd gnd ms_flop
XXdff7 din[7] dout[7] dout_bar[7] clk vdd gnd ms_flop
XXdff8 din[8] dout[8] dout_bar[8] clk vdd gnd ms_flop
XXdff9 din[9] dout[9] dout_bar[9] clk vdd gnd ms_flop
.ENDS msf_address

.SUBCKT msf_data_in din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] dout[0] dout_bar[0] dout[1] dout_bar[1] dout[2] dout_bar[2] dout[3] dout_bar[3] dout[4] dout_bar[4] dout[5] dout_bar[5] dout[6] dout_bar[6] dout[7] dout_bar[7] dout[8] dout_bar[8] dout[9] dout_bar[9] dout[10] dout_bar[10] dout[11] dout_bar[11] dout[12] dout_bar[12] dout[13] dout_bar[13] dout[14] dout_bar[14] dout[15] dout_bar[15] dout[16] dout_bar[16] dout[17] dout_bar[17] dout[18] dout_bar[18] dout[19] dout_bar[19] dout[20] dout_bar[20] dout[21] dout_bar[21] dout[22] dout_bar[22] dout[23] dout_bar[23] dout[24] dout_bar[24] dout[25] dout_bar[25] dout[26] dout_bar[26] dout[27] dout_bar[27] dout[28] dout_bar[28] dout[29] dout_bar[29] dout[30] dout_bar[30] dout[31] dout_bar[31] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
XXdff4 din[1] dout[1] dout_bar[1] clk vdd gnd ms_flop
XXdff8 din[2] dout[2] dout_bar[2] clk vdd gnd ms_flop
XXdff12 din[3] dout[3] dout_bar[3] clk vdd gnd ms_flop
XXdff16 din[4] dout[4] dout_bar[4] clk vdd gnd ms_flop
XXdff20 din[5] dout[5] dout_bar[5] clk vdd gnd ms_flop
XXdff24 din[6] dout[6] dout_bar[6] clk vdd gnd ms_flop
XXdff28 din[7] dout[7] dout_bar[7] clk vdd gnd ms_flop
XXdff32 din[8] dout[8] dout_bar[8] clk vdd gnd ms_flop
XXdff36 din[9] dout[9] dout_bar[9] clk vdd gnd ms_flop
XXdff40 din[10] dout[10] dout_bar[10] clk vdd gnd ms_flop
XXdff44 din[11] dout[11] dout_bar[11] clk vdd gnd ms_flop
XXdff48 din[12] dout[12] dout_bar[12] clk vdd gnd ms_flop
XXdff52 din[13] dout[13] dout_bar[13] clk vdd gnd ms_flop
XXdff56 din[14] dout[14] dout_bar[14] clk vdd gnd ms_flop
XXdff60 din[15] dout[15] dout_bar[15] clk vdd gnd ms_flop
XXdff64 din[16] dout[16] dout_bar[16] clk vdd gnd ms_flop
XXdff68 din[17] dout[17] dout_bar[17] clk vdd gnd ms_flop
XXdff72 din[18] dout[18] dout_bar[18] clk vdd gnd ms_flop
XXdff76 din[19] dout[19] dout_bar[19] clk vdd gnd ms_flop
XXdff80 din[20] dout[20] dout_bar[20] clk vdd gnd ms_flop
XXdff84 din[21] dout[21] dout_bar[21] clk vdd gnd ms_flop
XXdff88 din[22] dout[22] dout_bar[22] clk vdd gnd ms_flop
XXdff92 din[23] dout[23] dout_bar[23] clk vdd gnd ms_flop
XXdff96 din[24] dout[24] dout_bar[24] clk vdd gnd ms_flop
XXdff100 din[25] dout[25] dout_bar[25] clk vdd gnd ms_flop
XXdff104 din[26] dout[26] dout_bar[26] clk vdd gnd ms_flop
XXdff108 din[27] dout[27] dout_bar[27] clk vdd gnd ms_flop
XXdff112 din[28] dout[28] dout_bar[28] clk vdd gnd ms_flop
XXdff116 din[29] dout[29] dout_bar[29] clk vdd gnd ms_flop
XXdff120 din[30] dout[30] dout_bar[30] clk vdd gnd ms_flop
XXdff124 din[31] dout[31] dout_bar[31] clk vdd gnd ms_flop
.ENDS msf_data_in

.SUBCKT tri_gate in out en en_bar vdd gnd
M_1 net_2 in_inv gnd gnd NMOS_VTG W=180.000000n L=50.000000n
M_2 out en net_2 gnd NMOS_VTG W=180.000000n L=50.000000n
M_3 net_3 in_inv vdd vdd PMOS_VTG W=360.000000n L=50.000000n
M_4 out en_bar net_3 vdd PMOS_VTG W=360.000000n L=50.000000n
M_5 in_inv in vdd vdd PMOS_VTG W=180.000000n L=50.000000n
M_6 in_inv in gnd gnd NMOS_VTG W=90.000000n L=50.000000n
.ENDS


.SUBCKT tri_gate_array in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[18] in[19] in[20] in[21] in[22] in[23] in[24] in[25] in[26] in[27] in[28] in[29] in[30] in[31] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] out[10] out[11] out[12] out[13] out[14] out[15] out[16] out[17] out[18] out[19] out[20] out[21] out[22] out[23] out[24] out[25] out[26] out[27] out[28] out[29] out[30] out[31] en en_bar vdd gnd
XXtri_gate0 in[0] out[0] en en_bar vdd gnd tri_gate
XXtri_gate4 in[1] out[1] en en_bar vdd gnd tri_gate
XXtri_gate8 in[2] out[2] en en_bar vdd gnd tri_gate
XXtri_gate12 in[3] out[3] en en_bar vdd gnd tri_gate
XXtri_gate16 in[4] out[4] en en_bar vdd gnd tri_gate
XXtri_gate20 in[5] out[5] en en_bar vdd gnd tri_gate
XXtri_gate24 in[6] out[6] en en_bar vdd gnd tri_gate
XXtri_gate28 in[7] out[7] en en_bar vdd gnd tri_gate
XXtri_gate32 in[8] out[8] en en_bar vdd gnd tri_gate
XXtri_gate36 in[9] out[9] en en_bar vdd gnd tri_gate
XXtri_gate40 in[10] out[10] en en_bar vdd gnd tri_gate
XXtri_gate44 in[11] out[11] en en_bar vdd gnd tri_gate
XXtri_gate48 in[12] out[12] en en_bar vdd gnd tri_gate
XXtri_gate52 in[13] out[13] en en_bar vdd gnd tri_gate
XXtri_gate56 in[14] out[14] en en_bar vdd gnd tri_gate
XXtri_gate60 in[15] out[15] en en_bar vdd gnd tri_gate
XXtri_gate64 in[16] out[16] en en_bar vdd gnd tri_gate
XXtri_gate68 in[17] out[17] en en_bar vdd gnd tri_gate
XXtri_gate72 in[18] out[18] en en_bar vdd gnd tri_gate
XXtri_gate76 in[19] out[19] en en_bar vdd gnd tri_gate
XXtri_gate80 in[20] out[20] en en_bar vdd gnd tri_gate
XXtri_gate84 in[21] out[21] en en_bar vdd gnd tri_gate
XXtri_gate88 in[22] out[22] en en_bar vdd gnd tri_gate
XXtri_gate92 in[23] out[23] en en_bar vdd gnd tri_gate
XXtri_gate96 in[24] out[24] en en_bar vdd gnd tri_gate
XXtri_gate100 in[25] out[25] en en_bar vdd gnd tri_gate
XXtri_gate104 in[26] out[26] en en_bar vdd gnd tri_gate
XXtri_gate108 in[27] out[27] en en_bar vdd gnd tri_gate
XXtri_gate112 in[28] out[28] en en_bar vdd gnd tri_gate
XXtri_gate116 in[29] out[29] en en_bar vdd gnd tri_gate
XXtri_gate120 in[30] out[30] en en_bar vdd gnd tri_gate
XXtri_gate124 in[31] out[31] en en_bar vdd gnd tri_gate
.ENDS tri_gate_array

.SUBCKT pinv_11 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_11

.SUBCKT pinv_12 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_12

.SUBCKT pnand2_4 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand2_4

.SUBCKT wordline_driver in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[18] in[19] in[20] in[21] in[22] in[23] in[24] in[25] in[26] in[27] in[28] in[29] in[30] in[31] in[32] in[33] in[34] in[35] in[36] in[37] in[38] in[39] in[40] in[41] in[42] in[43] in[44] in[45] in[46] in[47] in[48] in[49] in[50] in[51] in[52] in[53] in[54] in[55] in[56] in[57] in[58] in[59] in[60] in[61] in[62] in[63] in[64] in[65] in[66] in[67] in[68] in[69] in[70] in[71] in[72] in[73] in[74] in[75] in[76] in[77] in[78] in[79] in[80] in[81] in[82] in[83] in[84] in[85] in[86] in[87] in[88] in[89] in[90] in[91] in[92] in[93] in[94] in[95] in[96] in[97] in[98] in[99] in[100] in[101] in[102] in[103] in[104] in[105] in[106] in[107] in[108] in[109] in[110] in[111] in[112] in[113] in[114] in[115] in[116] in[117] in[118] in[119] in[120] in[121] in[122] in[123] in[124] in[125] in[126] in[127] in[128] in[129] in[130] in[131] in[132] in[133] in[134] in[135] in[136] in[137] in[138] in[139] in[140] in[141] in[142] in[143] in[144] in[145] in[146] in[147] in[148] in[149] in[150] in[151] in[152] in[153] in[154] in[155] in[156] in[157] in[158] in[159] in[160] in[161] in[162] in[163] in[164] in[165] in[166] in[167] in[168] in[169] in[170] in[171] in[172] in[173] in[174] in[175] in[176] in[177] in[178] in[179] in[180] in[181] in[182] in[183] in[184] in[185] in[186] in[187] in[188] in[189] in[190] in[191] in[192] in[193] in[194] in[195] in[196] in[197] in[198] in[199] in[200] in[201] in[202] in[203] in[204] in[205] in[206] in[207] in[208] in[209] in[210] in[211] in[212] in[213] in[214] in[215] in[216] in[217] in[218] in[219] in[220] in[221] in[222] in[223] in[224] in[225] in[226] in[227] in[228] in[229] in[230] in[231] in[232] in[233] in[234] in[235] in[236] in[237] in[238] in[239] in[240] in[241] in[242] in[243] in[244] in[245] in[246] in[247] in[248] in[249] in[250] in[251] in[252] in[253] in[254] in[255] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] en vdd gnd
Xwl_driver_inv_en0 en en_bar[0] vdd gnd pinv_12
Xwl_driver_nand0 en_bar[0] in[0] net[0] vdd gnd pnand2_4
Xwl_driver_inv0 net[0] wl[0] vdd gnd pinv_11
Xwl_driver_inv_en1 en en_bar[1] vdd gnd pinv_12
Xwl_driver_nand1 en_bar[1] in[1] net[1] vdd gnd pnand2_4
Xwl_driver_inv1 net[1] wl[1] vdd gnd pinv_11
Xwl_driver_inv_en2 en en_bar[2] vdd gnd pinv_12
Xwl_driver_nand2 en_bar[2] in[2] net[2] vdd gnd pnand2_4
Xwl_driver_inv2 net[2] wl[2] vdd gnd pinv_11
Xwl_driver_inv_en3 en en_bar[3] vdd gnd pinv_12
Xwl_driver_nand3 en_bar[3] in[3] net[3] vdd gnd pnand2_4
Xwl_driver_inv3 net[3] wl[3] vdd gnd pinv_11
Xwl_driver_inv_en4 en en_bar[4] vdd gnd pinv_12
Xwl_driver_nand4 en_bar[4] in[4] net[4] vdd gnd pnand2_4
Xwl_driver_inv4 net[4] wl[4] vdd gnd pinv_11
Xwl_driver_inv_en5 en en_bar[5] vdd gnd pinv_12
Xwl_driver_nand5 en_bar[5] in[5] net[5] vdd gnd pnand2_4
Xwl_driver_inv5 net[5] wl[5] vdd gnd pinv_11
Xwl_driver_inv_en6 en en_bar[6] vdd gnd pinv_12
Xwl_driver_nand6 en_bar[6] in[6] net[6] vdd gnd pnand2_4
Xwl_driver_inv6 net[6] wl[6] vdd gnd pinv_11
Xwl_driver_inv_en7 en en_bar[7] vdd gnd pinv_12
Xwl_driver_nand7 en_bar[7] in[7] net[7] vdd gnd pnand2_4
Xwl_driver_inv7 net[7] wl[7] vdd gnd pinv_11
Xwl_driver_inv_en8 en en_bar[8] vdd gnd pinv_12
Xwl_driver_nand8 en_bar[8] in[8] net[8] vdd gnd pnand2_4
Xwl_driver_inv8 net[8] wl[8] vdd gnd pinv_11
Xwl_driver_inv_en9 en en_bar[9] vdd gnd pinv_12
Xwl_driver_nand9 en_bar[9] in[9] net[9] vdd gnd pnand2_4
Xwl_driver_inv9 net[9] wl[9] vdd gnd pinv_11
Xwl_driver_inv_en10 en en_bar[10] vdd gnd pinv_12
Xwl_driver_nand10 en_bar[10] in[10] net[10] vdd gnd pnand2_4
Xwl_driver_inv10 net[10] wl[10] vdd gnd pinv_11
Xwl_driver_inv_en11 en en_bar[11] vdd gnd pinv_12
Xwl_driver_nand11 en_bar[11] in[11] net[11] vdd gnd pnand2_4
Xwl_driver_inv11 net[11] wl[11] vdd gnd pinv_11
Xwl_driver_inv_en12 en en_bar[12] vdd gnd pinv_12
Xwl_driver_nand12 en_bar[12] in[12] net[12] vdd gnd pnand2_4
Xwl_driver_inv12 net[12] wl[12] vdd gnd pinv_11
Xwl_driver_inv_en13 en en_bar[13] vdd gnd pinv_12
Xwl_driver_nand13 en_bar[13] in[13] net[13] vdd gnd pnand2_4
Xwl_driver_inv13 net[13] wl[13] vdd gnd pinv_11
Xwl_driver_inv_en14 en en_bar[14] vdd gnd pinv_12
Xwl_driver_nand14 en_bar[14] in[14] net[14] vdd gnd pnand2_4
Xwl_driver_inv14 net[14] wl[14] vdd gnd pinv_11
Xwl_driver_inv_en15 en en_bar[15] vdd gnd pinv_12
Xwl_driver_nand15 en_bar[15] in[15] net[15] vdd gnd pnand2_4
Xwl_driver_inv15 net[15] wl[15] vdd gnd pinv_11
Xwl_driver_inv_en16 en en_bar[16] vdd gnd pinv_12
Xwl_driver_nand16 en_bar[16] in[16] net[16] vdd gnd pnand2_4
Xwl_driver_inv16 net[16] wl[16] vdd gnd pinv_11
Xwl_driver_inv_en17 en en_bar[17] vdd gnd pinv_12
Xwl_driver_nand17 en_bar[17] in[17] net[17] vdd gnd pnand2_4
Xwl_driver_inv17 net[17] wl[17] vdd gnd pinv_11
Xwl_driver_inv_en18 en en_bar[18] vdd gnd pinv_12
Xwl_driver_nand18 en_bar[18] in[18] net[18] vdd gnd pnand2_4
Xwl_driver_inv18 net[18] wl[18] vdd gnd pinv_11
Xwl_driver_inv_en19 en en_bar[19] vdd gnd pinv_12
Xwl_driver_nand19 en_bar[19] in[19] net[19] vdd gnd pnand2_4
Xwl_driver_inv19 net[19] wl[19] vdd gnd pinv_11
Xwl_driver_inv_en20 en en_bar[20] vdd gnd pinv_12
Xwl_driver_nand20 en_bar[20] in[20] net[20] vdd gnd pnand2_4
Xwl_driver_inv20 net[20] wl[20] vdd gnd pinv_11
Xwl_driver_inv_en21 en en_bar[21] vdd gnd pinv_12
Xwl_driver_nand21 en_bar[21] in[21] net[21] vdd gnd pnand2_4
Xwl_driver_inv21 net[21] wl[21] vdd gnd pinv_11
Xwl_driver_inv_en22 en en_bar[22] vdd gnd pinv_12
Xwl_driver_nand22 en_bar[22] in[22] net[22] vdd gnd pnand2_4
Xwl_driver_inv22 net[22] wl[22] vdd gnd pinv_11
Xwl_driver_inv_en23 en en_bar[23] vdd gnd pinv_12
Xwl_driver_nand23 en_bar[23] in[23] net[23] vdd gnd pnand2_4
Xwl_driver_inv23 net[23] wl[23] vdd gnd pinv_11
Xwl_driver_inv_en24 en en_bar[24] vdd gnd pinv_12
Xwl_driver_nand24 en_bar[24] in[24] net[24] vdd gnd pnand2_4
Xwl_driver_inv24 net[24] wl[24] vdd gnd pinv_11
Xwl_driver_inv_en25 en en_bar[25] vdd gnd pinv_12
Xwl_driver_nand25 en_bar[25] in[25] net[25] vdd gnd pnand2_4
Xwl_driver_inv25 net[25] wl[25] vdd gnd pinv_11
Xwl_driver_inv_en26 en en_bar[26] vdd gnd pinv_12
Xwl_driver_nand26 en_bar[26] in[26] net[26] vdd gnd pnand2_4
Xwl_driver_inv26 net[26] wl[26] vdd gnd pinv_11
Xwl_driver_inv_en27 en en_bar[27] vdd gnd pinv_12
Xwl_driver_nand27 en_bar[27] in[27] net[27] vdd gnd pnand2_4
Xwl_driver_inv27 net[27] wl[27] vdd gnd pinv_11
Xwl_driver_inv_en28 en en_bar[28] vdd gnd pinv_12
Xwl_driver_nand28 en_bar[28] in[28] net[28] vdd gnd pnand2_4
Xwl_driver_inv28 net[28] wl[28] vdd gnd pinv_11
Xwl_driver_inv_en29 en en_bar[29] vdd gnd pinv_12
Xwl_driver_nand29 en_bar[29] in[29] net[29] vdd gnd pnand2_4
Xwl_driver_inv29 net[29] wl[29] vdd gnd pinv_11
Xwl_driver_inv_en30 en en_bar[30] vdd gnd pinv_12
Xwl_driver_nand30 en_bar[30] in[30] net[30] vdd gnd pnand2_4
Xwl_driver_inv30 net[30] wl[30] vdd gnd pinv_11
Xwl_driver_inv_en31 en en_bar[31] vdd gnd pinv_12
Xwl_driver_nand31 en_bar[31] in[31] net[31] vdd gnd pnand2_4
Xwl_driver_inv31 net[31] wl[31] vdd gnd pinv_11
Xwl_driver_inv_en32 en en_bar[32] vdd gnd pinv_12
Xwl_driver_nand32 en_bar[32] in[32] net[32] vdd gnd pnand2_4
Xwl_driver_inv32 net[32] wl[32] vdd gnd pinv_11
Xwl_driver_inv_en33 en en_bar[33] vdd gnd pinv_12
Xwl_driver_nand33 en_bar[33] in[33] net[33] vdd gnd pnand2_4
Xwl_driver_inv33 net[33] wl[33] vdd gnd pinv_11
Xwl_driver_inv_en34 en en_bar[34] vdd gnd pinv_12
Xwl_driver_nand34 en_bar[34] in[34] net[34] vdd gnd pnand2_4
Xwl_driver_inv34 net[34] wl[34] vdd gnd pinv_11
Xwl_driver_inv_en35 en en_bar[35] vdd gnd pinv_12
Xwl_driver_nand35 en_bar[35] in[35] net[35] vdd gnd pnand2_4
Xwl_driver_inv35 net[35] wl[35] vdd gnd pinv_11
Xwl_driver_inv_en36 en en_bar[36] vdd gnd pinv_12
Xwl_driver_nand36 en_bar[36] in[36] net[36] vdd gnd pnand2_4
Xwl_driver_inv36 net[36] wl[36] vdd gnd pinv_11
Xwl_driver_inv_en37 en en_bar[37] vdd gnd pinv_12
Xwl_driver_nand37 en_bar[37] in[37] net[37] vdd gnd pnand2_4
Xwl_driver_inv37 net[37] wl[37] vdd gnd pinv_11
Xwl_driver_inv_en38 en en_bar[38] vdd gnd pinv_12
Xwl_driver_nand38 en_bar[38] in[38] net[38] vdd gnd pnand2_4
Xwl_driver_inv38 net[38] wl[38] vdd gnd pinv_11
Xwl_driver_inv_en39 en en_bar[39] vdd gnd pinv_12
Xwl_driver_nand39 en_bar[39] in[39] net[39] vdd gnd pnand2_4
Xwl_driver_inv39 net[39] wl[39] vdd gnd pinv_11
Xwl_driver_inv_en40 en en_bar[40] vdd gnd pinv_12
Xwl_driver_nand40 en_bar[40] in[40] net[40] vdd gnd pnand2_4
Xwl_driver_inv40 net[40] wl[40] vdd gnd pinv_11
Xwl_driver_inv_en41 en en_bar[41] vdd gnd pinv_12
Xwl_driver_nand41 en_bar[41] in[41] net[41] vdd gnd pnand2_4
Xwl_driver_inv41 net[41] wl[41] vdd gnd pinv_11
Xwl_driver_inv_en42 en en_bar[42] vdd gnd pinv_12
Xwl_driver_nand42 en_bar[42] in[42] net[42] vdd gnd pnand2_4
Xwl_driver_inv42 net[42] wl[42] vdd gnd pinv_11
Xwl_driver_inv_en43 en en_bar[43] vdd gnd pinv_12
Xwl_driver_nand43 en_bar[43] in[43] net[43] vdd gnd pnand2_4
Xwl_driver_inv43 net[43] wl[43] vdd gnd pinv_11
Xwl_driver_inv_en44 en en_bar[44] vdd gnd pinv_12
Xwl_driver_nand44 en_bar[44] in[44] net[44] vdd gnd pnand2_4
Xwl_driver_inv44 net[44] wl[44] vdd gnd pinv_11
Xwl_driver_inv_en45 en en_bar[45] vdd gnd pinv_12
Xwl_driver_nand45 en_bar[45] in[45] net[45] vdd gnd pnand2_4
Xwl_driver_inv45 net[45] wl[45] vdd gnd pinv_11
Xwl_driver_inv_en46 en en_bar[46] vdd gnd pinv_12
Xwl_driver_nand46 en_bar[46] in[46] net[46] vdd gnd pnand2_4
Xwl_driver_inv46 net[46] wl[46] vdd gnd pinv_11
Xwl_driver_inv_en47 en en_bar[47] vdd gnd pinv_12
Xwl_driver_nand47 en_bar[47] in[47] net[47] vdd gnd pnand2_4
Xwl_driver_inv47 net[47] wl[47] vdd gnd pinv_11
Xwl_driver_inv_en48 en en_bar[48] vdd gnd pinv_12
Xwl_driver_nand48 en_bar[48] in[48] net[48] vdd gnd pnand2_4
Xwl_driver_inv48 net[48] wl[48] vdd gnd pinv_11
Xwl_driver_inv_en49 en en_bar[49] vdd gnd pinv_12
Xwl_driver_nand49 en_bar[49] in[49] net[49] vdd gnd pnand2_4
Xwl_driver_inv49 net[49] wl[49] vdd gnd pinv_11
Xwl_driver_inv_en50 en en_bar[50] vdd gnd pinv_12
Xwl_driver_nand50 en_bar[50] in[50] net[50] vdd gnd pnand2_4
Xwl_driver_inv50 net[50] wl[50] vdd gnd pinv_11
Xwl_driver_inv_en51 en en_bar[51] vdd gnd pinv_12
Xwl_driver_nand51 en_bar[51] in[51] net[51] vdd gnd pnand2_4
Xwl_driver_inv51 net[51] wl[51] vdd gnd pinv_11
Xwl_driver_inv_en52 en en_bar[52] vdd gnd pinv_12
Xwl_driver_nand52 en_bar[52] in[52] net[52] vdd gnd pnand2_4
Xwl_driver_inv52 net[52] wl[52] vdd gnd pinv_11
Xwl_driver_inv_en53 en en_bar[53] vdd gnd pinv_12
Xwl_driver_nand53 en_bar[53] in[53] net[53] vdd gnd pnand2_4
Xwl_driver_inv53 net[53] wl[53] vdd gnd pinv_11
Xwl_driver_inv_en54 en en_bar[54] vdd gnd pinv_12
Xwl_driver_nand54 en_bar[54] in[54] net[54] vdd gnd pnand2_4
Xwl_driver_inv54 net[54] wl[54] vdd gnd pinv_11
Xwl_driver_inv_en55 en en_bar[55] vdd gnd pinv_12
Xwl_driver_nand55 en_bar[55] in[55] net[55] vdd gnd pnand2_4
Xwl_driver_inv55 net[55] wl[55] vdd gnd pinv_11
Xwl_driver_inv_en56 en en_bar[56] vdd gnd pinv_12
Xwl_driver_nand56 en_bar[56] in[56] net[56] vdd gnd pnand2_4
Xwl_driver_inv56 net[56] wl[56] vdd gnd pinv_11
Xwl_driver_inv_en57 en en_bar[57] vdd gnd pinv_12
Xwl_driver_nand57 en_bar[57] in[57] net[57] vdd gnd pnand2_4
Xwl_driver_inv57 net[57] wl[57] vdd gnd pinv_11
Xwl_driver_inv_en58 en en_bar[58] vdd gnd pinv_12
Xwl_driver_nand58 en_bar[58] in[58] net[58] vdd gnd pnand2_4
Xwl_driver_inv58 net[58] wl[58] vdd gnd pinv_11
Xwl_driver_inv_en59 en en_bar[59] vdd gnd pinv_12
Xwl_driver_nand59 en_bar[59] in[59] net[59] vdd gnd pnand2_4
Xwl_driver_inv59 net[59] wl[59] vdd gnd pinv_11
Xwl_driver_inv_en60 en en_bar[60] vdd gnd pinv_12
Xwl_driver_nand60 en_bar[60] in[60] net[60] vdd gnd pnand2_4
Xwl_driver_inv60 net[60] wl[60] vdd gnd pinv_11
Xwl_driver_inv_en61 en en_bar[61] vdd gnd pinv_12
Xwl_driver_nand61 en_bar[61] in[61] net[61] vdd gnd pnand2_4
Xwl_driver_inv61 net[61] wl[61] vdd gnd pinv_11
Xwl_driver_inv_en62 en en_bar[62] vdd gnd pinv_12
Xwl_driver_nand62 en_bar[62] in[62] net[62] vdd gnd pnand2_4
Xwl_driver_inv62 net[62] wl[62] vdd gnd pinv_11
Xwl_driver_inv_en63 en en_bar[63] vdd gnd pinv_12
Xwl_driver_nand63 en_bar[63] in[63] net[63] vdd gnd pnand2_4
Xwl_driver_inv63 net[63] wl[63] vdd gnd pinv_11
Xwl_driver_inv_en64 en en_bar[64] vdd gnd pinv_12
Xwl_driver_nand64 en_bar[64] in[64] net[64] vdd gnd pnand2_4
Xwl_driver_inv64 net[64] wl[64] vdd gnd pinv_11
Xwl_driver_inv_en65 en en_bar[65] vdd gnd pinv_12
Xwl_driver_nand65 en_bar[65] in[65] net[65] vdd gnd pnand2_4
Xwl_driver_inv65 net[65] wl[65] vdd gnd pinv_11
Xwl_driver_inv_en66 en en_bar[66] vdd gnd pinv_12
Xwl_driver_nand66 en_bar[66] in[66] net[66] vdd gnd pnand2_4
Xwl_driver_inv66 net[66] wl[66] vdd gnd pinv_11
Xwl_driver_inv_en67 en en_bar[67] vdd gnd pinv_12
Xwl_driver_nand67 en_bar[67] in[67] net[67] vdd gnd pnand2_4
Xwl_driver_inv67 net[67] wl[67] vdd gnd pinv_11
Xwl_driver_inv_en68 en en_bar[68] vdd gnd pinv_12
Xwl_driver_nand68 en_bar[68] in[68] net[68] vdd gnd pnand2_4
Xwl_driver_inv68 net[68] wl[68] vdd gnd pinv_11
Xwl_driver_inv_en69 en en_bar[69] vdd gnd pinv_12
Xwl_driver_nand69 en_bar[69] in[69] net[69] vdd gnd pnand2_4
Xwl_driver_inv69 net[69] wl[69] vdd gnd pinv_11
Xwl_driver_inv_en70 en en_bar[70] vdd gnd pinv_12
Xwl_driver_nand70 en_bar[70] in[70] net[70] vdd gnd pnand2_4
Xwl_driver_inv70 net[70] wl[70] vdd gnd pinv_11
Xwl_driver_inv_en71 en en_bar[71] vdd gnd pinv_12
Xwl_driver_nand71 en_bar[71] in[71] net[71] vdd gnd pnand2_4
Xwl_driver_inv71 net[71] wl[71] vdd gnd pinv_11
Xwl_driver_inv_en72 en en_bar[72] vdd gnd pinv_12
Xwl_driver_nand72 en_bar[72] in[72] net[72] vdd gnd pnand2_4
Xwl_driver_inv72 net[72] wl[72] vdd gnd pinv_11
Xwl_driver_inv_en73 en en_bar[73] vdd gnd pinv_12
Xwl_driver_nand73 en_bar[73] in[73] net[73] vdd gnd pnand2_4
Xwl_driver_inv73 net[73] wl[73] vdd gnd pinv_11
Xwl_driver_inv_en74 en en_bar[74] vdd gnd pinv_12
Xwl_driver_nand74 en_bar[74] in[74] net[74] vdd gnd pnand2_4
Xwl_driver_inv74 net[74] wl[74] vdd gnd pinv_11
Xwl_driver_inv_en75 en en_bar[75] vdd gnd pinv_12
Xwl_driver_nand75 en_bar[75] in[75] net[75] vdd gnd pnand2_4
Xwl_driver_inv75 net[75] wl[75] vdd gnd pinv_11
Xwl_driver_inv_en76 en en_bar[76] vdd gnd pinv_12
Xwl_driver_nand76 en_bar[76] in[76] net[76] vdd gnd pnand2_4
Xwl_driver_inv76 net[76] wl[76] vdd gnd pinv_11
Xwl_driver_inv_en77 en en_bar[77] vdd gnd pinv_12
Xwl_driver_nand77 en_bar[77] in[77] net[77] vdd gnd pnand2_4
Xwl_driver_inv77 net[77] wl[77] vdd gnd pinv_11
Xwl_driver_inv_en78 en en_bar[78] vdd gnd pinv_12
Xwl_driver_nand78 en_bar[78] in[78] net[78] vdd gnd pnand2_4
Xwl_driver_inv78 net[78] wl[78] vdd gnd pinv_11
Xwl_driver_inv_en79 en en_bar[79] vdd gnd pinv_12
Xwl_driver_nand79 en_bar[79] in[79] net[79] vdd gnd pnand2_4
Xwl_driver_inv79 net[79] wl[79] vdd gnd pinv_11
Xwl_driver_inv_en80 en en_bar[80] vdd gnd pinv_12
Xwl_driver_nand80 en_bar[80] in[80] net[80] vdd gnd pnand2_4
Xwl_driver_inv80 net[80] wl[80] vdd gnd pinv_11
Xwl_driver_inv_en81 en en_bar[81] vdd gnd pinv_12
Xwl_driver_nand81 en_bar[81] in[81] net[81] vdd gnd pnand2_4
Xwl_driver_inv81 net[81] wl[81] vdd gnd pinv_11
Xwl_driver_inv_en82 en en_bar[82] vdd gnd pinv_12
Xwl_driver_nand82 en_bar[82] in[82] net[82] vdd gnd pnand2_4
Xwl_driver_inv82 net[82] wl[82] vdd gnd pinv_11
Xwl_driver_inv_en83 en en_bar[83] vdd gnd pinv_12
Xwl_driver_nand83 en_bar[83] in[83] net[83] vdd gnd pnand2_4
Xwl_driver_inv83 net[83] wl[83] vdd gnd pinv_11
Xwl_driver_inv_en84 en en_bar[84] vdd gnd pinv_12
Xwl_driver_nand84 en_bar[84] in[84] net[84] vdd gnd pnand2_4
Xwl_driver_inv84 net[84] wl[84] vdd gnd pinv_11
Xwl_driver_inv_en85 en en_bar[85] vdd gnd pinv_12
Xwl_driver_nand85 en_bar[85] in[85] net[85] vdd gnd pnand2_4
Xwl_driver_inv85 net[85] wl[85] vdd gnd pinv_11
Xwl_driver_inv_en86 en en_bar[86] vdd gnd pinv_12
Xwl_driver_nand86 en_bar[86] in[86] net[86] vdd gnd pnand2_4
Xwl_driver_inv86 net[86] wl[86] vdd gnd pinv_11
Xwl_driver_inv_en87 en en_bar[87] vdd gnd pinv_12
Xwl_driver_nand87 en_bar[87] in[87] net[87] vdd gnd pnand2_4
Xwl_driver_inv87 net[87] wl[87] vdd gnd pinv_11
Xwl_driver_inv_en88 en en_bar[88] vdd gnd pinv_12
Xwl_driver_nand88 en_bar[88] in[88] net[88] vdd gnd pnand2_4
Xwl_driver_inv88 net[88] wl[88] vdd gnd pinv_11
Xwl_driver_inv_en89 en en_bar[89] vdd gnd pinv_12
Xwl_driver_nand89 en_bar[89] in[89] net[89] vdd gnd pnand2_4
Xwl_driver_inv89 net[89] wl[89] vdd gnd pinv_11
Xwl_driver_inv_en90 en en_bar[90] vdd gnd pinv_12
Xwl_driver_nand90 en_bar[90] in[90] net[90] vdd gnd pnand2_4
Xwl_driver_inv90 net[90] wl[90] vdd gnd pinv_11
Xwl_driver_inv_en91 en en_bar[91] vdd gnd pinv_12
Xwl_driver_nand91 en_bar[91] in[91] net[91] vdd gnd pnand2_4
Xwl_driver_inv91 net[91] wl[91] vdd gnd pinv_11
Xwl_driver_inv_en92 en en_bar[92] vdd gnd pinv_12
Xwl_driver_nand92 en_bar[92] in[92] net[92] vdd gnd pnand2_4
Xwl_driver_inv92 net[92] wl[92] vdd gnd pinv_11
Xwl_driver_inv_en93 en en_bar[93] vdd gnd pinv_12
Xwl_driver_nand93 en_bar[93] in[93] net[93] vdd gnd pnand2_4
Xwl_driver_inv93 net[93] wl[93] vdd gnd pinv_11
Xwl_driver_inv_en94 en en_bar[94] vdd gnd pinv_12
Xwl_driver_nand94 en_bar[94] in[94] net[94] vdd gnd pnand2_4
Xwl_driver_inv94 net[94] wl[94] vdd gnd pinv_11
Xwl_driver_inv_en95 en en_bar[95] vdd gnd pinv_12
Xwl_driver_nand95 en_bar[95] in[95] net[95] vdd gnd pnand2_4
Xwl_driver_inv95 net[95] wl[95] vdd gnd pinv_11
Xwl_driver_inv_en96 en en_bar[96] vdd gnd pinv_12
Xwl_driver_nand96 en_bar[96] in[96] net[96] vdd gnd pnand2_4
Xwl_driver_inv96 net[96] wl[96] vdd gnd pinv_11
Xwl_driver_inv_en97 en en_bar[97] vdd gnd pinv_12
Xwl_driver_nand97 en_bar[97] in[97] net[97] vdd gnd pnand2_4
Xwl_driver_inv97 net[97] wl[97] vdd gnd pinv_11
Xwl_driver_inv_en98 en en_bar[98] vdd gnd pinv_12
Xwl_driver_nand98 en_bar[98] in[98] net[98] vdd gnd pnand2_4
Xwl_driver_inv98 net[98] wl[98] vdd gnd pinv_11
Xwl_driver_inv_en99 en en_bar[99] vdd gnd pinv_12
Xwl_driver_nand99 en_bar[99] in[99] net[99] vdd gnd pnand2_4
Xwl_driver_inv99 net[99] wl[99] vdd gnd pinv_11
Xwl_driver_inv_en100 en en_bar[100] vdd gnd pinv_12
Xwl_driver_nand100 en_bar[100] in[100] net[100] vdd gnd pnand2_4
Xwl_driver_inv100 net[100] wl[100] vdd gnd pinv_11
Xwl_driver_inv_en101 en en_bar[101] vdd gnd pinv_12
Xwl_driver_nand101 en_bar[101] in[101] net[101] vdd gnd pnand2_4
Xwl_driver_inv101 net[101] wl[101] vdd gnd pinv_11
Xwl_driver_inv_en102 en en_bar[102] vdd gnd pinv_12
Xwl_driver_nand102 en_bar[102] in[102] net[102] vdd gnd pnand2_4
Xwl_driver_inv102 net[102] wl[102] vdd gnd pinv_11
Xwl_driver_inv_en103 en en_bar[103] vdd gnd pinv_12
Xwl_driver_nand103 en_bar[103] in[103] net[103] vdd gnd pnand2_4
Xwl_driver_inv103 net[103] wl[103] vdd gnd pinv_11
Xwl_driver_inv_en104 en en_bar[104] vdd gnd pinv_12
Xwl_driver_nand104 en_bar[104] in[104] net[104] vdd gnd pnand2_4
Xwl_driver_inv104 net[104] wl[104] vdd gnd pinv_11
Xwl_driver_inv_en105 en en_bar[105] vdd gnd pinv_12
Xwl_driver_nand105 en_bar[105] in[105] net[105] vdd gnd pnand2_4
Xwl_driver_inv105 net[105] wl[105] vdd gnd pinv_11
Xwl_driver_inv_en106 en en_bar[106] vdd gnd pinv_12
Xwl_driver_nand106 en_bar[106] in[106] net[106] vdd gnd pnand2_4
Xwl_driver_inv106 net[106] wl[106] vdd gnd pinv_11
Xwl_driver_inv_en107 en en_bar[107] vdd gnd pinv_12
Xwl_driver_nand107 en_bar[107] in[107] net[107] vdd gnd pnand2_4
Xwl_driver_inv107 net[107] wl[107] vdd gnd pinv_11
Xwl_driver_inv_en108 en en_bar[108] vdd gnd pinv_12
Xwl_driver_nand108 en_bar[108] in[108] net[108] vdd gnd pnand2_4
Xwl_driver_inv108 net[108] wl[108] vdd gnd pinv_11
Xwl_driver_inv_en109 en en_bar[109] vdd gnd pinv_12
Xwl_driver_nand109 en_bar[109] in[109] net[109] vdd gnd pnand2_4
Xwl_driver_inv109 net[109] wl[109] vdd gnd pinv_11
Xwl_driver_inv_en110 en en_bar[110] vdd gnd pinv_12
Xwl_driver_nand110 en_bar[110] in[110] net[110] vdd gnd pnand2_4
Xwl_driver_inv110 net[110] wl[110] vdd gnd pinv_11
Xwl_driver_inv_en111 en en_bar[111] vdd gnd pinv_12
Xwl_driver_nand111 en_bar[111] in[111] net[111] vdd gnd pnand2_4
Xwl_driver_inv111 net[111] wl[111] vdd gnd pinv_11
Xwl_driver_inv_en112 en en_bar[112] vdd gnd pinv_12
Xwl_driver_nand112 en_bar[112] in[112] net[112] vdd gnd pnand2_4
Xwl_driver_inv112 net[112] wl[112] vdd gnd pinv_11
Xwl_driver_inv_en113 en en_bar[113] vdd gnd pinv_12
Xwl_driver_nand113 en_bar[113] in[113] net[113] vdd gnd pnand2_4
Xwl_driver_inv113 net[113] wl[113] vdd gnd pinv_11
Xwl_driver_inv_en114 en en_bar[114] vdd gnd pinv_12
Xwl_driver_nand114 en_bar[114] in[114] net[114] vdd gnd pnand2_4
Xwl_driver_inv114 net[114] wl[114] vdd gnd pinv_11
Xwl_driver_inv_en115 en en_bar[115] vdd gnd pinv_12
Xwl_driver_nand115 en_bar[115] in[115] net[115] vdd gnd pnand2_4
Xwl_driver_inv115 net[115] wl[115] vdd gnd pinv_11
Xwl_driver_inv_en116 en en_bar[116] vdd gnd pinv_12
Xwl_driver_nand116 en_bar[116] in[116] net[116] vdd gnd pnand2_4
Xwl_driver_inv116 net[116] wl[116] vdd gnd pinv_11
Xwl_driver_inv_en117 en en_bar[117] vdd gnd pinv_12
Xwl_driver_nand117 en_bar[117] in[117] net[117] vdd gnd pnand2_4
Xwl_driver_inv117 net[117] wl[117] vdd gnd pinv_11
Xwl_driver_inv_en118 en en_bar[118] vdd gnd pinv_12
Xwl_driver_nand118 en_bar[118] in[118] net[118] vdd gnd pnand2_4
Xwl_driver_inv118 net[118] wl[118] vdd gnd pinv_11
Xwl_driver_inv_en119 en en_bar[119] vdd gnd pinv_12
Xwl_driver_nand119 en_bar[119] in[119] net[119] vdd gnd pnand2_4
Xwl_driver_inv119 net[119] wl[119] vdd gnd pinv_11
Xwl_driver_inv_en120 en en_bar[120] vdd gnd pinv_12
Xwl_driver_nand120 en_bar[120] in[120] net[120] vdd gnd pnand2_4
Xwl_driver_inv120 net[120] wl[120] vdd gnd pinv_11
Xwl_driver_inv_en121 en en_bar[121] vdd gnd pinv_12
Xwl_driver_nand121 en_bar[121] in[121] net[121] vdd gnd pnand2_4
Xwl_driver_inv121 net[121] wl[121] vdd gnd pinv_11
Xwl_driver_inv_en122 en en_bar[122] vdd gnd pinv_12
Xwl_driver_nand122 en_bar[122] in[122] net[122] vdd gnd pnand2_4
Xwl_driver_inv122 net[122] wl[122] vdd gnd pinv_11
Xwl_driver_inv_en123 en en_bar[123] vdd gnd pinv_12
Xwl_driver_nand123 en_bar[123] in[123] net[123] vdd gnd pnand2_4
Xwl_driver_inv123 net[123] wl[123] vdd gnd pinv_11
Xwl_driver_inv_en124 en en_bar[124] vdd gnd pinv_12
Xwl_driver_nand124 en_bar[124] in[124] net[124] vdd gnd pnand2_4
Xwl_driver_inv124 net[124] wl[124] vdd gnd pinv_11
Xwl_driver_inv_en125 en en_bar[125] vdd gnd pinv_12
Xwl_driver_nand125 en_bar[125] in[125] net[125] vdd gnd pnand2_4
Xwl_driver_inv125 net[125] wl[125] vdd gnd pinv_11
Xwl_driver_inv_en126 en en_bar[126] vdd gnd pinv_12
Xwl_driver_nand126 en_bar[126] in[126] net[126] vdd gnd pnand2_4
Xwl_driver_inv126 net[126] wl[126] vdd gnd pinv_11
Xwl_driver_inv_en127 en en_bar[127] vdd gnd pinv_12
Xwl_driver_nand127 en_bar[127] in[127] net[127] vdd gnd pnand2_4
Xwl_driver_inv127 net[127] wl[127] vdd gnd pinv_11
Xwl_driver_inv_en128 en en_bar[128] vdd gnd pinv_12
Xwl_driver_nand128 en_bar[128] in[128] net[128] vdd gnd pnand2_4
Xwl_driver_inv128 net[128] wl[128] vdd gnd pinv_11
Xwl_driver_inv_en129 en en_bar[129] vdd gnd pinv_12
Xwl_driver_nand129 en_bar[129] in[129] net[129] vdd gnd pnand2_4
Xwl_driver_inv129 net[129] wl[129] vdd gnd pinv_11
Xwl_driver_inv_en130 en en_bar[130] vdd gnd pinv_12
Xwl_driver_nand130 en_bar[130] in[130] net[130] vdd gnd pnand2_4
Xwl_driver_inv130 net[130] wl[130] vdd gnd pinv_11
Xwl_driver_inv_en131 en en_bar[131] vdd gnd pinv_12
Xwl_driver_nand131 en_bar[131] in[131] net[131] vdd gnd pnand2_4
Xwl_driver_inv131 net[131] wl[131] vdd gnd pinv_11
Xwl_driver_inv_en132 en en_bar[132] vdd gnd pinv_12
Xwl_driver_nand132 en_bar[132] in[132] net[132] vdd gnd pnand2_4
Xwl_driver_inv132 net[132] wl[132] vdd gnd pinv_11
Xwl_driver_inv_en133 en en_bar[133] vdd gnd pinv_12
Xwl_driver_nand133 en_bar[133] in[133] net[133] vdd gnd pnand2_4
Xwl_driver_inv133 net[133] wl[133] vdd gnd pinv_11
Xwl_driver_inv_en134 en en_bar[134] vdd gnd pinv_12
Xwl_driver_nand134 en_bar[134] in[134] net[134] vdd gnd pnand2_4
Xwl_driver_inv134 net[134] wl[134] vdd gnd pinv_11
Xwl_driver_inv_en135 en en_bar[135] vdd gnd pinv_12
Xwl_driver_nand135 en_bar[135] in[135] net[135] vdd gnd pnand2_4
Xwl_driver_inv135 net[135] wl[135] vdd gnd pinv_11
Xwl_driver_inv_en136 en en_bar[136] vdd gnd pinv_12
Xwl_driver_nand136 en_bar[136] in[136] net[136] vdd gnd pnand2_4
Xwl_driver_inv136 net[136] wl[136] vdd gnd pinv_11
Xwl_driver_inv_en137 en en_bar[137] vdd gnd pinv_12
Xwl_driver_nand137 en_bar[137] in[137] net[137] vdd gnd pnand2_4
Xwl_driver_inv137 net[137] wl[137] vdd gnd pinv_11
Xwl_driver_inv_en138 en en_bar[138] vdd gnd pinv_12
Xwl_driver_nand138 en_bar[138] in[138] net[138] vdd gnd pnand2_4
Xwl_driver_inv138 net[138] wl[138] vdd gnd pinv_11
Xwl_driver_inv_en139 en en_bar[139] vdd gnd pinv_12
Xwl_driver_nand139 en_bar[139] in[139] net[139] vdd gnd pnand2_4
Xwl_driver_inv139 net[139] wl[139] vdd gnd pinv_11
Xwl_driver_inv_en140 en en_bar[140] vdd gnd pinv_12
Xwl_driver_nand140 en_bar[140] in[140] net[140] vdd gnd pnand2_4
Xwl_driver_inv140 net[140] wl[140] vdd gnd pinv_11
Xwl_driver_inv_en141 en en_bar[141] vdd gnd pinv_12
Xwl_driver_nand141 en_bar[141] in[141] net[141] vdd gnd pnand2_4
Xwl_driver_inv141 net[141] wl[141] vdd gnd pinv_11
Xwl_driver_inv_en142 en en_bar[142] vdd gnd pinv_12
Xwl_driver_nand142 en_bar[142] in[142] net[142] vdd gnd pnand2_4
Xwl_driver_inv142 net[142] wl[142] vdd gnd pinv_11
Xwl_driver_inv_en143 en en_bar[143] vdd gnd pinv_12
Xwl_driver_nand143 en_bar[143] in[143] net[143] vdd gnd pnand2_4
Xwl_driver_inv143 net[143] wl[143] vdd gnd pinv_11
Xwl_driver_inv_en144 en en_bar[144] vdd gnd pinv_12
Xwl_driver_nand144 en_bar[144] in[144] net[144] vdd gnd pnand2_4
Xwl_driver_inv144 net[144] wl[144] vdd gnd pinv_11
Xwl_driver_inv_en145 en en_bar[145] vdd gnd pinv_12
Xwl_driver_nand145 en_bar[145] in[145] net[145] vdd gnd pnand2_4
Xwl_driver_inv145 net[145] wl[145] vdd gnd pinv_11
Xwl_driver_inv_en146 en en_bar[146] vdd gnd pinv_12
Xwl_driver_nand146 en_bar[146] in[146] net[146] vdd gnd pnand2_4
Xwl_driver_inv146 net[146] wl[146] vdd gnd pinv_11
Xwl_driver_inv_en147 en en_bar[147] vdd gnd pinv_12
Xwl_driver_nand147 en_bar[147] in[147] net[147] vdd gnd pnand2_4
Xwl_driver_inv147 net[147] wl[147] vdd gnd pinv_11
Xwl_driver_inv_en148 en en_bar[148] vdd gnd pinv_12
Xwl_driver_nand148 en_bar[148] in[148] net[148] vdd gnd pnand2_4
Xwl_driver_inv148 net[148] wl[148] vdd gnd pinv_11
Xwl_driver_inv_en149 en en_bar[149] vdd gnd pinv_12
Xwl_driver_nand149 en_bar[149] in[149] net[149] vdd gnd pnand2_4
Xwl_driver_inv149 net[149] wl[149] vdd gnd pinv_11
Xwl_driver_inv_en150 en en_bar[150] vdd gnd pinv_12
Xwl_driver_nand150 en_bar[150] in[150] net[150] vdd gnd pnand2_4
Xwl_driver_inv150 net[150] wl[150] vdd gnd pinv_11
Xwl_driver_inv_en151 en en_bar[151] vdd gnd pinv_12
Xwl_driver_nand151 en_bar[151] in[151] net[151] vdd gnd pnand2_4
Xwl_driver_inv151 net[151] wl[151] vdd gnd pinv_11
Xwl_driver_inv_en152 en en_bar[152] vdd gnd pinv_12
Xwl_driver_nand152 en_bar[152] in[152] net[152] vdd gnd pnand2_4
Xwl_driver_inv152 net[152] wl[152] vdd gnd pinv_11
Xwl_driver_inv_en153 en en_bar[153] vdd gnd pinv_12
Xwl_driver_nand153 en_bar[153] in[153] net[153] vdd gnd pnand2_4
Xwl_driver_inv153 net[153] wl[153] vdd gnd pinv_11
Xwl_driver_inv_en154 en en_bar[154] vdd gnd pinv_12
Xwl_driver_nand154 en_bar[154] in[154] net[154] vdd gnd pnand2_4
Xwl_driver_inv154 net[154] wl[154] vdd gnd pinv_11
Xwl_driver_inv_en155 en en_bar[155] vdd gnd pinv_12
Xwl_driver_nand155 en_bar[155] in[155] net[155] vdd gnd pnand2_4
Xwl_driver_inv155 net[155] wl[155] vdd gnd pinv_11
Xwl_driver_inv_en156 en en_bar[156] vdd gnd pinv_12
Xwl_driver_nand156 en_bar[156] in[156] net[156] vdd gnd pnand2_4
Xwl_driver_inv156 net[156] wl[156] vdd gnd pinv_11
Xwl_driver_inv_en157 en en_bar[157] vdd gnd pinv_12
Xwl_driver_nand157 en_bar[157] in[157] net[157] vdd gnd pnand2_4
Xwl_driver_inv157 net[157] wl[157] vdd gnd pinv_11
Xwl_driver_inv_en158 en en_bar[158] vdd gnd pinv_12
Xwl_driver_nand158 en_bar[158] in[158] net[158] vdd gnd pnand2_4
Xwl_driver_inv158 net[158] wl[158] vdd gnd pinv_11
Xwl_driver_inv_en159 en en_bar[159] vdd gnd pinv_12
Xwl_driver_nand159 en_bar[159] in[159] net[159] vdd gnd pnand2_4
Xwl_driver_inv159 net[159] wl[159] vdd gnd pinv_11
Xwl_driver_inv_en160 en en_bar[160] vdd gnd pinv_12
Xwl_driver_nand160 en_bar[160] in[160] net[160] vdd gnd pnand2_4
Xwl_driver_inv160 net[160] wl[160] vdd gnd pinv_11
Xwl_driver_inv_en161 en en_bar[161] vdd gnd pinv_12
Xwl_driver_nand161 en_bar[161] in[161] net[161] vdd gnd pnand2_4
Xwl_driver_inv161 net[161] wl[161] vdd gnd pinv_11
Xwl_driver_inv_en162 en en_bar[162] vdd gnd pinv_12
Xwl_driver_nand162 en_bar[162] in[162] net[162] vdd gnd pnand2_4
Xwl_driver_inv162 net[162] wl[162] vdd gnd pinv_11
Xwl_driver_inv_en163 en en_bar[163] vdd gnd pinv_12
Xwl_driver_nand163 en_bar[163] in[163] net[163] vdd gnd pnand2_4
Xwl_driver_inv163 net[163] wl[163] vdd gnd pinv_11
Xwl_driver_inv_en164 en en_bar[164] vdd gnd pinv_12
Xwl_driver_nand164 en_bar[164] in[164] net[164] vdd gnd pnand2_4
Xwl_driver_inv164 net[164] wl[164] vdd gnd pinv_11
Xwl_driver_inv_en165 en en_bar[165] vdd gnd pinv_12
Xwl_driver_nand165 en_bar[165] in[165] net[165] vdd gnd pnand2_4
Xwl_driver_inv165 net[165] wl[165] vdd gnd pinv_11
Xwl_driver_inv_en166 en en_bar[166] vdd gnd pinv_12
Xwl_driver_nand166 en_bar[166] in[166] net[166] vdd gnd pnand2_4
Xwl_driver_inv166 net[166] wl[166] vdd gnd pinv_11
Xwl_driver_inv_en167 en en_bar[167] vdd gnd pinv_12
Xwl_driver_nand167 en_bar[167] in[167] net[167] vdd gnd pnand2_4
Xwl_driver_inv167 net[167] wl[167] vdd gnd pinv_11
Xwl_driver_inv_en168 en en_bar[168] vdd gnd pinv_12
Xwl_driver_nand168 en_bar[168] in[168] net[168] vdd gnd pnand2_4
Xwl_driver_inv168 net[168] wl[168] vdd gnd pinv_11
Xwl_driver_inv_en169 en en_bar[169] vdd gnd pinv_12
Xwl_driver_nand169 en_bar[169] in[169] net[169] vdd gnd pnand2_4
Xwl_driver_inv169 net[169] wl[169] vdd gnd pinv_11
Xwl_driver_inv_en170 en en_bar[170] vdd gnd pinv_12
Xwl_driver_nand170 en_bar[170] in[170] net[170] vdd gnd pnand2_4
Xwl_driver_inv170 net[170] wl[170] vdd gnd pinv_11
Xwl_driver_inv_en171 en en_bar[171] vdd gnd pinv_12
Xwl_driver_nand171 en_bar[171] in[171] net[171] vdd gnd pnand2_4
Xwl_driver_inv171 net[171] wl[171] vdd gnd pinv_11
Xwl_driver_inv_en172 en en_bar[172] vdd gnd pinv_12
Xwl_driver_nand172 en_bar[172] in[172] net[172] vdd gnd pnand2_4
Xwl_driver_inv172 net[172] wl[172] vdd gnd pinv_11
Xwl_driver_inv_en173 en en_bar[173] vdd gnd pinv_12
Xwl_driver_nand173 en_bar[173] in[173] net[173] vdd gnd pnand2_4
Xwl_driver_inv173 net[173] wl[173] vdd gnd pinv_11
Xwl_driver_inv_en174 en en_bar[174] vdd gnd pinv_12
Xwl_driver_nand174 en_bar[174] in[174] net[174] vdd gnd pnand2_4
Xwl_driver_inv174 net[174] wl[174] vdd gnd pinv_11
Xwl_driver_inv_en175 en en_bar[175] vdd gnd pinv_12
Xwl_driver_nand175 en_bar[175] in[175] net[175] vdd gnd pnand2_4
Xwl_driver_inv175 net[175] wl[175] vdd gnd pinv_11
Xwl_driver_inv_en176 en en_bar[176] vdd gnd pinv_12
Xwl_driver_nand176 en_bar[176] in[176] net[176] vdd gnd pnand2_4
Xwl_driver_inv176 net[176] wl[176] vdd gnd pinv_11
Xwl_driver_inv_en177 en en_bar[177] vdd gnd pinv_12
Xwl_driver_nand177 en_bar[177] in[177] net[177] vdd gnd pnand2_4
Xwl_driver_inv177 net[177] wl[177] vdd gnd pinv_11
Xwl_driver_inv_en178 en en_bar[178] vdd gnd pinv_12
Xwl_driver_nand178 en_bar[178] in[178] net[178] vdd gnd pnand2_4
Xwl_driver_inv178 net[178] wl[178] vdd gnd pinv_11
Xwl_driver_inv_en179 en en_bar[179] vdd gnd pinv_12
Xwl_driver_nand179 en_bar[179] in[179] net[179] vdd gnd pnand2_4
Xwl_driver_inv179 net[179] wl[179] vdd gnd pinv_11
Xwl_driver_inv_en180 en en_bar[180] vdd gnd pinv_12
Xwl_driver_nand180 en_bar[180] in[180] net[180] vdd gnd pnand2_4
Xwl_driver_inv180 net[180] wl[180] vdd gnd pinv_11
Xwl_driver_inv_en181 en en_bar[181] vdd gnd pinv_12
Xwl_driver_nand181 en_bar[181] in[181] net[181] vdd gnd pnand2_4
Xwl_driver_inv181 net[181] wl[181] vdd gnd pinv_11
Xwl_driver_inv_en182 en en_bar[182] vdd gnd pinv_12
Xwl_driver_nand182 en_bar[182] in[182] net[182] vdd gnd pnand2_4
Xwl_driver_inv182 net[182] wl[182] vdd gnd pinv_11
Xwl_driver_inv_en183 en en_bar[183] vdd gnd pinv_12
Xwl_driver_nand183 en_bar[183] in[183] net[183] vdd gnd pnand2_4
Xwl_driver_inv183 net[183] wl[183] vdd gnd pinv_11
Xwl_driver_inv_en184 en en_bar[184] vdd gnd pinv_12
Xwl_driver_nand184 en_bar[184] in[184] net[184] vdd gnd pnand2_4
Xwl_driver_inv184 net[184] wl[184] vdd gnd pinv_11
Xwl_driver_inv_en185 en en_bar[185] vdd gnd pinv_12
Xwl_driver_nand185 en_bar[185] in[185] net[185] vdd gnd pnand2_4
Xwl_driver_inv185 net[185] wl[185] vdd gnd pinv_11
Xwl_driver_inv_en186 en en_bar[186] vdd gnd pinv_12
Xwl_driver_nand186 en_bar[186] in[186] net[186] vdd gnd pnand2_4
Xwl_driver_inv186 net[186] wl[186] vdd gnd pinv_11
Xwl_driver_inv_en187 en en_bar[187] vdd gnd pinv_12
Xwl_driver_nand187 en_bar[187] in[187] net[187] vdd gnd pnand2_4
Xwl_driver_inv187 net[187] wl[187] vdd gnd pinv_11
Xwl_driver_inv_en188 en en_bar[188] vdd gnd pinv_12
Xwl_driver_nand188 en_bar[188] in[188] net[188] vdd gnd pnand2_4
Xwl_driver_inv188 net[188] wl[188] vdd gnd pinv_11
Xwl_driver_inv_en189 en en_bar[189] vdd gnd pinv_12
Xwl_driver_nand189 en_bar[189] in[189] net[189] vdd gnd pnand2_4
Xwl_driver_inv189 net[189] wl[189] vdd gnd pinv_11
Xwl_driver_inv_en190 en en_bar[190] vdd gnd pinv_12
Xwl_driver_nand190 en_bar[190] in[190] net[190] vdd gnd pnand2_4
Xwl_driver_inv190 net[190] wl[190] vdd gnd pinv_11
Xwl_driver_inv_en191 en en_bar[191] vdd gnd pinv_12
Xwl_driver_nand191 en_bar[191] in[191] net[191] vdd gnd pnand2_4
Xwl_driver_inv191 net[191] wl[191] vdd gnd pinv_11
Xwl_driver_inv_en192 en en_bar[192] vdd gnd pinv_12
Xwl_driver_nand192 en_bar[192] in[192] net[192] vdd gnd pnand2_4
Xwl_driver_inv192 net[192] wl[192] vdd gnd pinv_11
Xwl_driver_inv_en193 en en_bar[193] vdd gnd pinv_12
Xwl_driver_nand193 en_bar[193] in[193] net[193] vdd gnd pnand2_4
Xwl_driver_inv193 net[193] wl[193] vdd gnd pinv_11
Xwl_driver_inv_en194 en en_bar[194] vdd gnd pinv_12
Xwl_driver_nand194 en_bar[194] in[194] net[194] vdd gnd pnand2_4
Xwl_driver_inv194 net[194] wl[194] vdd gnd pinv_11
Xwl_driver_inv_en195 en en_bar[195] vdd gnd pinv_12
Xwl_driver_nand195 en_bar[195] in[195] net[195] vdd gnd pnand2_4
Xwl_driver_inv195 net[195] wl[195] vdd gnd pinv_11
Xwl_driver_inv_en196 en en_bar[196] vdd gnd pinv_12
Xwl_driver_nand196 en_bar[196] in[196] net[196] vdd gnd pnand2_4
Xwl_driver_inv196 net[196] wl[196] vdd gnd pinv_11
Xwl_driver_inv_en197 en en_bar[197] vdd gnd pinv_12
Xwl_driver_nand197 en_bar[197] in[197] net[197] vdd gnd pnand2_4
Xwl_driver_inv197 net[197] wl[197] vdd gnd pinv_11
Xwl_driver_inv_en198 en en_bar[198] vdd gnd pinv_12
Xwl_driver_nand198 en_bar[198] in[198] net[198] vdd gnd pnand2_4
Xwl_driver_inv198 net[198] wl[198] vdd gnd pinv_11
Xwl_driver_inv_en199 en en_bar[199] vdd gnd pinv_12
Xwl_driver_nand199 en_bar[199] in[199] net[199] vdd gnd pnand2_4
Xwl_driver_inv199 net[199] wl[199] vdd gnd pinv_11
Xwl_driver_inv_en200 en en_bar[200] vdd gnd pinv_12
Xwl_driver_nand200 en_bar[200] in[200] net[200] vdd gnd pnand2_4
Xwl_driver_inv200 net[200] wl[200] vdd gnd pinv_11
Xwl_driver_inv_en201 en en_bar[201] vdd gnd pinv_12
Xwl_driver_nand201 en_bar[201] in[201] net[201] vdd gnd pnand2_4
Xwl_driver_inv201 net[201] wl[201] vdd gnd pinv_11
Xwl_driver_inv_en202 en en_bar[202] vdd gnd pinv_12
Xwl_driver_nand202 en_bar[202] in[202] net[202] vdd gnd pnand2_4
Xwl_driver_inv202 net[202] wl[202] vdd gnd pinv_11
Xwl_driver_inv_en203 en en_bar[203] vdd gnd pinv_12
Xwl_driver_nand203 en_bar[203] in[203] net[203] vdd gnd pnand2_4
Xwl_driver_inv203 net[203] wl[203] vdd gnd pinv_11
Xwl_driver_inv_en204 en en_bar[204] vdd gnd pinv_12
Xwl_driver_nand204 en_bar[204] in[204] net[204] vdd gnd pnand2_4
Xwl_driver_inv204 net[204] wl[204] vdd gnd pinv_11
Xwl_driver_inv_en205 en en_bar[205] vdd gnd pinv_12
Xwl_driver_nand205 en_bar[205] in[205] net[205] vdd gnd pnand2_4
Xwl_driver_inv205 net[205] wl[205] vdd gnd pinv_11
Xwl_driver_inv_en206 en en_bar[206] vdd gnd pinv_12
Xwl_driver_nand206 en_bar[206] in[206] net[206] vdd gnd pnand2_4
Xwl_driver_inv206 net[206] wl[206] vdd gnd pinv_11
Xwl_driver_inv_en207 en en_bar[207] vdd gnd pinv_12
Xwl_driver_nand207 en_bar[207] in[207] net[207] vdd gnd pnand2_4
Xwl_driver_inv207 net[207] wl[207] vdd gnd pinv_11
Xwl_driver_inv_en208 en en_bar[208] vdd gnd pinv_12
Xwl_driver_nand208 en_bar[208] in[208] net[208] vdd gnd pnand2_4
Xwl_driver_inv208 net[208] wl[208] vdd gnd pinv_11
Xwl_driver_inv_en209 en en_bar[209] vdd gnd pinv_12
Xwl_driver_nand209 en_bar[209] in[209] net[209] vdd gnd pnand2_4
Xwl_driver_inv209 net[209] wl[209] vdd gnd pinv_11
Xwl_driver_inv_en210 en en_bar[210] vdd gnd pinv_12
Xwl_driver_nand210 en_bar[210] in[210] net[210] vdd gnd pnand2_4
Xwl_driver_inv210 net[210] wl[210] vdd gnd pinv_11
Xwl_driver_inv_en211 en en_bar[211] vdd gnd pinv_12
Xwl_driver_nand211 en_bar[211] in[211] net[211] vdd gnd pnand2_4
Xwl_driver_inv211 net[211] wl[211] vdd gnd pinv_11
Xwl_driver_inv_en212 en en_bar[212] vdd gnd pinv_12
Xwl_driver_nand212 en_bar[212] in[212] net[212] vdd gnd pnand2_4
Xwl_driver_inv212 net[212] wl[212] vdd gnd pinv_11
Xwl_driver_inv_en213 en en_bar[213] vdd gnd pinv_12
Xwl_driver_nand213 en_bar[213] in[213] net[213] vdd gnd pnand2_4
Xwl_driver_inv213 net[213] wl[213] vdd gnd pinv_11
Xwl_driver_inv_en214 en en_bar[214] vdd gnd pinv_12
Xwl_driver_nand214 en_bar[214] in[214] net[214] vdd gnd pnand2_4
Xwl_driver_inv214 net[214] wl[214] vdd gnd pinv_11
Xwl_driver_inv_en215 en en_bar[215] vdd gnd pinv_12
Xwl_driver_nand215 en_bar[215] in[215] net[215] vdd gnd pnand2_4
Xwl_driver_inv215 net[215] wl[215] vdd gnd pinv_11
Xwl_driver_inv_en216 en en_bar[216] vdd gnd pinv_12
Xwl_driver_nand216 en_bar[216] in[216] net[216] vdd gnd pnand2_4
Xwl_driver_inv216 net[216] wl[216] vdd gnd pinv_11
Xwl_driver_inv_en217 en en_bar[217] vdd gnd pinv_12
Xwl_driver_nand217 en_bar[217] in[217] net[217] vdd gnd pnand2_4
Xwl_driver_inv217 net[217] wl[217] vdd gnd pinv_11
Xwl_driver_inv_en218 en en_bar[218] vdd gnd pinv_12
Xwl_driver_nand218 en_bar[218] in[218] net[218] vdd gnd pnand2_4
Xwl_driver_inv218 net[218] wl[218] vdd gnd pinv_11
Xwl_driver_inv_en219 en en_bar[219] vdd gnd pinv_12
Xwl_driver_nand219 en_bar[219] in[219] net[219] vdd gnd pnand2_4
Xwl_driver_inv219 net[219] wl[219] vdd gnd pinv_11
Xwl_driver_inv_en220 en en_bar[220] vdd gnd pinv_12
Xwl_driver_nand220 en_bar[220] in[220] net[220] vdd gnd pnand2_4
Xwl_driver_inv220 net[220] wl[220] vdd gnd pinv_11
Xwl_driver_inv_en221 en en_bar[221] vdd gnd pinv_12
Xwl_driver_nand221 en_bar[221] in[221] net[221] vdd gnd pnand2_4
Xwl_driver_inv221 net[221] wl[221] vdd gnd pinv_11
Xwl_driver_inv_en222 en en_bar[222] vdd gnd pinv_12
Xwl_driver_nand222 en_bar[222] in[222] net[222] vdd gnd pnand2_4
Xwl_driver_inv222 net[222] wl[222] vdd gnd pinv_11
Xwl_driver_inv_en223 en en_bar[223] vdd gnd pinv_12
Xwl_driver_nand223 en_bar[223] in[223] net[223] vdd gnd pnand2_4
Xwl_driver_inv223 net[223] wl[223] vdd gnd pinv_11
Xwl_driver_inv_en224 en en_bar[224] vdd gnd pinv_12
Xwl_driver_nand224 en_bar[224] in[224] net[224] vdd gnd pnand2_4
Xwl_driver_inv224 net[224] wl[224] vdd gnd pinv_11
Xwl_driver_inv_en225 en en_bar[225] vdd gnd pinv_12
Xwl_driver_nand225 en_bar[225] in[225] net[225] vdd gnd pnand2_4
Xwl_driver_inv225 net[225] wl[225] vdd gnd pinv_11
Xwl_driver_inv_en226 en en_bar[226] vdd gnd pinv_12
Xwl_driver_nand226 en_bar[226] in[226] net[226] vdd gnd pnand2_4
Xwl_driver_inv226 net[226] wl[226] vdd gnd pinv_11
Xwl_driver_inv_en227 en en_bar[227] vdd gnd pinv_12
Xwl_driver_nand227 en_bar[227] in[227] net[227] vdd gnd pnand2_4
Xwl_driver_inv227 net[227] wl[227] vdd gnd pinv_11
Xwl_driver_inv_en228 en en_bar[228] vdd gnd pinv_12
Xwl_driver_nand228 en_bar[228] in[228] net[228] vdd gnd pnand2_4
Xwl_driver_inv228 net[228] wl[228] vdd gnd pinv_11
Xwl_driver_inv_en229 en en_bar[229] vdd gnd pinv_12
Xwl_driver_nand229 en_bar[229] in[229] net[229] vdd gnd pnand2_4
Xwl_driver_inv229 net[229] wl[229] vdd gnd pinv_11
Xwl_driver_inv_en230 en en_bar[230] vdd gnd pinv_12
Xwl_driver_nand230 en_bar[230] in[230] net[230] vdd gnd pnand2_4
Xwl_driver_inv230 net[230] wl[230] vdd gnd pinv_11
Xwl_driver_inv_en231 en en_bar[231] vdd gnd pinv_12
Xwl_driver_nand231 en_bar[231] in[231] net[231] vdd gnd pnand2_4
Xwl_driver_inv231 net[231] wl[231] vdd gnd pinv_11
Xwl_driver_inv_en232 en en_bar[232] vdd gnd pinv_12
Xwl_driver_nand232 en_bar[232] in[232] net[232] vdd gnd pnand2_4
Xwl_driver_inv232 net[232] wl[232] vdd gnd pinv_11
Xwl_driver_inv_en233 en en_bar[233] vdd gnd pinv_12
Xwl_driver_nand233 en_bar[233] in[233] net[233] vdd gnd pnand2_4
Xwl_driver_inv233 net[233] wl[233] vdd gnd pinv_11
Xwl_driver_inv_en234 en en_bar[234] vdd gnd pinv_12
Xwl_driver_nand234 en_bar[234] in[234] net[234] vdd gnd pnand2_4
Xwl_driver_inv234 net[234] wl[234] vdd gnd pinv_11
Xwl_driver_inv_en235 en en_bar[235] vdd gnd pinv_12
Xwl_driver_nand235 en_bar[235] in[235] net[235] vdd gnd pnand2_4
Xwl_driver_inv235 net[235] wl[235] vdd gnd pinv_11
Xwl_driver_inv_en236 en en_bar[236] vdd gnd pinv_12
Xwl_driver_nand236 en_bar[236] in[236] net[236] vdd gnd pnand2_4
Xwl_driver_inv236 net[236] wl[236] vdd gnd pinv_11
Xwl_driver_inv_en237 en en_bar[237] vdd gnd pinv_12
Xwl_driver_nand237 en_bar[237] in[237] net[237] vdd gnd pnand2_4
Xwl_driver_inv237 net[237] wl[237] vdd gnd pinv_11
Xwl_driver_inv_en238 en en_bar[238] vdd gnd pinv_12
Xwl_driver_nand238 en_bar[238] in[238] net[238] vdd gnd pnand2_4
Xwl_driver_inv238 net[238] wl[238] vdd gnd pinv_11
Xwl_driver_inv_en239 en en_bar[239] vdd gnd pinv_12
Xwl_driver_nand239 en_bar[239] in[239] net[239] vdd gnd pnand2_4
Xwl_driver_inv239 net[239] wl[239] vdd gnd pinv_11
Xwl_driver_inv_en240 en en_bar[240] vdd gnd pinv_12
Xwl_driver_nand240 en_bar[240] in[240] net[240] vdd gnd pnand2_4
Xwl_driver_inv240 net[240] wl[240] vdd gnd pinv_11
Xwl_driver_inv_en241 en en_bar[241] vdd gnd pinv_12
Xwl_driver_nand241 en_bar[241] in[241] net[241] vdd gnd pnand2_4
Xwl_driver_inv241 net[241] wl[241] vdd gnd pinv_11
Xwl_driver_inv_en242 en en_bar[242] vdd gnd pinv_12
Xwl_driver_nand242 en_bar[242] in[242] net[242] vdd gnd pnand2_4
Xwl_driver_inv242 net[242] wl[242] vdd gnd pinv_11
Xwl_driver_inv_en243 en en_bar[243] vdd gnd pinv_12
Xwl_driver_nand243 en_bar[243] in[243] net[243] vdd gnd pnand2_4
Xwl_driver_inv243 net[243] wl[243] vdd gnd pinv_11
Xwl_driver_inv_en244 en en_bar[244] vdd gnd pinv_12
Xwl_driver_nand244 en_bar[244] in[244] net[244] vdd gnd pnand2_4
Xwl_driver_inv244 net[244] wl[244] vdd gnd pinv_11
Xwl_driver_inv_en245 en en_bar[245] vdd gnd pinv_12
Xwl_driver_nand245 en_bar[245] in[245] net[245] vdd gnd pnand2_4
Xwl_driver_inv245 net[245] wl[245] vdd gnd pinv_11
Xwl_driver_inv_en246 en en_bar[246] vdd gnd pinv_12
Xwl_driver_nand246 en_bar[246] in[246] net[246] vdd gnd pnand2_4
Xwl_driver_inv246 net[246] wl[246] vdd gnd pinv_11
Xwl_driver_inv_en247 en en_bar[247] vdd gnd pinv_12
Xwl_driver_nand247 en_bar[247] in[247] net[247] vdd gnd pnand2_4
Xwl_driver_inv247 net[247] wl[247] vdd gnd pinv_11
Xwl_driver_inv_en248 en en_bar[248] vdd gnd pinv_12
Xwl_driver_nand248 en_bar[248] in[248] net[248] vdd gnd pnand2_4
Xwl_driver_inv248 net[248] wl[248] vdd gnd pinv_11
Xwl_driver_inv_en249 en en_bar[249] vdd gnd pinv_12
Xwl_driver_nand249 en_bar[249] in[249] net[249] vdd gnd pnand2_4
Xwl_driver_inv249 net[249] wl[249] vdd gnd pinv_11
Xwl_driver_inv_en250 en en_bar[250] vdd gnd pinv_12
Xwl_driver_nand250 en_bar[250] in[250] net[250] vdd gnd pnand2_4
Xwl_driver_inv250 net[250] wl[250] vdd gnd pinv_11
Xwl_driver_inv_en251 en en_bar[251] vdd gnd pinv_12
Xwl_driver_nand251 en_bar[251] in[251] net[251] vdd gnd pnand2_4
Xwl_driver_inv251 net[251] wl[251] vdd gnd pinv_11
Xwl_driver_inv_en252 en en_bar[252] vdd gnd pinv_12
Xwl_driver_nand252 en_bar[252] in[252] net[252] vdd gnd pnand2_4
Xwl_driver_inv252 net[252] wl[252] vdd gnd pinv_11
Xwl_driver_inv_en253 en en_bar[253] vdd gnd pinv_12
Xwl_driver_nand253 en_bar[253] in[253] net[253] vdd gnd pnand2_4
Xwl_driver_inv253 net[253] wl[253] vdd gnd pinv_11
Xwl_driver_inv_en254 en en_bar[254] vdd gnd pinv_12
Xwl_driver_nand254 en_bar[254] in[254] net[254] vdd gnd pnand2_4
Xwl_driver_inv254 net[254] wl[254] vdd gnd pinv_11
Xwl_driver_inv_en255 en en_bar[255] vdd gnd pinv_12
Xwl_driver_nand255 en_bar[255] in[255] net[255] vdd gnd pnand2_4
Xwl_driver_inv255 net[255] wl[255] vdd gnd pinv_11
.ENDS wordline_driver

.SUBCKT pinv_13 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_13

.SUBCKT bank DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] ADDR[9] s_en w_en tri_en_bar tri_en clk_bar clk_buf vdd gnd
Xbitcell_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] vdd gnd bitcell_array
Xprecharge_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] clk_bar vdd precharge_array
Xcolumn_mux_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] sel[0] sel[1] sel[2] sel[3] bl_out[0] br_out[0] bl_out[1] br_out[1] bl_out[2] br_out[2] bl_out[3] br_out[3] bl_out[4] br_out[4] bl_out[5] br_out[5] bl_out[6] br_out[6] bl_out[7] br_out[7] bl_out[8] br_out[8] bl_out[9] br_out[9] bl_out[10] br_out[10] bl_out[11] br_out[11] bl_out[12] br_out[12] bl_out[13] br_out[13] bl_out[14] br_out[14] bl_out[15] br_out[15] bl_out[16] br_out[16] bl_out[17] br_out[17] bl_out[18] br_out[18] bl_out[19] br_out[19] bl_out[20] br_out[20] bl_out[21] br_out[21] bl_out[22] br_out[22] bl_out[23] br_out[23] bl_out[24] br_out[24] bl_out[25] br_out[25] bl_out[26] br_out[26] bl_out[27] br_out[27] bl_out[28] br_out[28] bl_out[29] br_out[29] bl_out[30] br_out[30] bl_out[31] br_out[31] gnd columnmux_array
Xcol_address_decoder A[8] A[9] sel[0] sel[1] sel[2] sel[3] vdd gnd pre2x4
Xsense_amp_array data_out[0] bl_out[0] br_out[0] data_out[1] bl_out[1] br_out[1] data_out[2] bl_out[2] br_out[2] data_out[3] bl_out[3] br_out[3] data_out[4] bl_out[4] br_out[4] data_out[5] bl_out[5] br_out[5] data_out[6] bl_out[6] br_out[6] data_out[7] bl_out[7] br_out[7] data_out[8] bl_out[8] br_out[8] data_out[9] bl_out[9] br_out[9] data_out[10] bl_out[10] br_out[10] data_out[11] bl_out[11] br_out[11] data_out[12] bl_out[12] br_out[12] data_out[13] bl_out[13] br_out[13] data_out[14] bl_out[14] br_out[14] data_out[15] bl_out[15] br_out[15] data_out[16] bl_out[16] br_out[16] data_out[17] bl_out[17] br_out[17] data_out[18] bl_out[18] br_out[18] data_out[19] bl_out[19] br_out[19] data_out[20] bl_out[20] br_out[20] data_out[21] bl_out[21] br_out[21] data_out[22] bl_out[22] br_out[22] data_out[23] bl_out[23] br_out[23] data_out[24] bl_out[24] br_out[24] data_out[25] bl_out[25] br_out[25] data_out[26] bl_out[26] br_out[26] data_out[27] bl_out[27] br_out[27] data_out[28] bl_out[28] br_out[28] data_out[29] bl_out[29] br_out[29] data_out[30] bl_out[30] br_out[30] data_out[31] bl_out[31] br_out[31] s_en vdd gnd sense_amp_array
Xwrite_driver_array data_in[0] data_in[1] data_in[2] data_in[3] data_in[4] data_in[5] data_in[6] data_in[7] data_in[8] data_in[9] data_in[10] data_in[11] data_in[12] data_in[13] data_in[14] data_in[15] data_in[16] data_in[17] data_in[18] data_in[19] data_in[20] data_in[21] data_in[22] data_in[23] data_in[24] data_in[25] data_in[26] data_in[27] data_in[28] data_in[29] data_in[30] data_in[31] bl_out[0] br_out[0] bl_out[1] br_out[1] bl_out[2] br_out[2] bl_out[3] br_out[3] bl_out[4] br_out[4] bl_out[5] br_out[5] bl_out[6] br_out[6] bl_out[7] br_out[7] bl_out[8] br_out[8] bl_out[9] br_out[9] bl_out[10] br_out[10] bl_out[11] br_out[11] bl_out[12] br_out[12] bl_out[13] br_out[13] bl_out[14] br_out[14] bl_out[15] br_out[15] bl_out[16] br_out[16] bl_out[17] br_out[17] bl_out[18] br_out[18] bl_out[19] br_out[19] bl_out[20] br_out[20] bl_out[21] br_out[21] bl_out[22] br_out[22] bl_out[23] br_out[23] bl_out[24] br_out[24] bl_out[25] br_out[25] bl_out[26] br_out[26] bl_out[27] br_out[27] bl_out[28] br_out[28] bl_out[29] br_out[29] bl_out[30] br_out[30] bl_out[31] br_out[31] w_en vdd gnd write_driver_array
Xdata_in_flop_array DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] data_in[0] data_in_bar[0] data_in[1] data_in_bar[1] data_in[2] data_in_bar[2] data_in[3] data_in_bar[3] data_in[4] data_in_bar[4] data_in[5] data_in_bar[5] data_in[6] data_in_bar[6] data_in[7] data_in_bar[7] data_in[8] data_in_bar[8] data_in[9] data_in_bar[9] data_in[10] data_in_bar[10] data_in[11] data_in_bar[11] data_in[12] data_in_bar[12] data_in[13] data_in_bar[13] data_in[14] data_in_bar[14] data_in[15] data_in_bar[15] data_in[16] data_in_bar[16] data_in[17] data_in_bar[17] data_in[18] data_in_bar[18] data_in[19] data_in_bar[19] data_in[20] data_in_bar[20] data_in[21] data_in_bar[21] data_in[22] data_in_bar[22] data_in[23] data_in_bar[23] data_in[24] data_in_bar[24] data_in[25] data_in_bar[25] data_in[26] data_in_bar[26] data_in[27] data_in_bar[27] data_in[28] data_in_bar[28] data_in[29] data_in_bar[29] data_in[30] data_in_bar[30] data_in[31] data_in_bar[31] clk_bar vdd gnd msf_data_in
Xtri_gate_array data_out[0] data_out[1] data_out[2] data_out[3] data_out[4] data_out[5] data_out[6] data_out[7] data_out[8] data_out[9] data_out[10] data_out[11] data_out[12] data_out[13] data_out[14] data_out[15] data_out[16] data_out[17] data_out[18] data_out[19] data_out[20] data_out[21] data_out[22] data_out[23] data_out[24] data_out[25] data_out[26] data_out[27] data_out[28] data_out[29] data_out[30] data_out[31] DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] tri_en tri_en_bar vdd gnd tri_gate_array
Xrow_decoder A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] dec_out[0] dec_out[1] dec_out[2] dec_out[3] dec_out[4] dec_out[5] dec_out[6] dec_out[7] dec_out[8] dec_out[9] dec_out[10] dec_out[11] dec_out[12] dec_out[13] dec_out[14] dec_out[15] dec_out[16] dec_out[17] dec_out[18] dec_out[19] dec_out[20] dec_out[21] dec_out[22] dec_out[23] dec_out[24] dec_out[25] dec_out[26] dec_out[27] dec_out[28] dec_out[29] dec_out[30] dec_out[31] dec_out[32] dec_out[33] dec_out[34] dec_out[35] dec_out[36] dec_out[37] dec_out[38] dec_out[39] dec_out[40] dec_out[41] dec_out[42] dec_out[43] dec_out[44] dec_out[45] dec_out[46] dec_out[47] dec_out[48] dec_out[49] dec_out[50] dec_out[51] dec_out[52] dec_out[53] dec_out[54] dec_out[55] dec_out[56] dec_out[57] dec_out[58] dec_out[59] dec_out[60] dec_out[61] dec_out[62] dec_out[63] dec_out[64] dec_out[65] dec_out[66] dec_out[67] dec_out[68] dec_out[69] dec_out[70] dec_out[71] dec_out[72] dec_out[73] dec_out[74] dec_out[75] dec_out[76] dec_out[77] dec_out[78] dec_out[79] dec_out[80] dec_out[81] dec_out[82] dec_out[83] dec_out[84] dec_out[85] dec_out[86] dec_out[87] dec_out[88] dec_out[89] dec_out[90] dec_out[91] dec_out[92] dec_out[93] dec_out[94] dec_out[95] dec_out[96] dec_out[97] dec_out[98] dec_out[99] dec_out[100] dec_out[101] dec_out[102] dec_out[103] dec_out[104] dec_out[105] dec_out[106] dec_out[107] dec_out[108] dec_out[109] dec_out[110] dec_out[111] dec_out[112] dec_out[113] dec_out[114] dec_out[115] dec_out[116] dec_out[117] dec_out[118] dec_out[119] dec_out[120] dec_out[121] dec_out[122] dec_out[123] dec_out[124] dec_out[125] dec_out[126] dec_out[127] dec_out[128] dec_out[129] dec_out[130] dec_out[131] dec_out[132] dec_out[133] dec_out[134] dec_out[135] dec_out[136] dec_out[137] dec_out[138] dec_out[139] dec_out[140] dec_out[141] dec_out[142] dec_out[143] dec_out[144] dec_out[145] dec_out[146] dec_out[147] dec_out[148] dec_out[149] dec_out[150] dec_out[151] dec_out[152] dec_out[153] dec_out[154] dec_out[155] dec_out[156] dec_out[157] dec_out[158] dec_out[159] dec_out[160] dec_out[161] dec_out[162] dec_out[163] dec_out[164] dec_out[165] dec_out[166] dec_out[167] dec_out[168] dec_out[169] dec_out[170] dec_out[171] dec_out[172] dec_out[173] dec_out[174] dec_out[175] dec_out[176] dec_out[177] dec_out[178] dec_out[179] dec_out[180] dec_out[181] dec_out[182] dec_out[183] dec_out[184] dec_out[185] dec_out[186] dec_out[187] dec_out[188] dec_out[189] dec_out[190] dec_out[191] dec_out[192] dec_out[193] dec_out[194] dec_out[195] dec_out[196] dec_out[197] dec_out[198] dec_out[199] dec_out[200] dec_out[201] dec_out[202] dec_out[203] dec_out[204] dec_out[205] dec_out[206] dec_out[207] dec_out[208] dec_out[209] dec_out[210] dec_out[211] dec_out[212] dec_out[213] dec_out[214] dec_out[215] dec_out[216] dec_out[217] dec_out[218] dec_out[219] dec_out[220] dec_out[221] dec_out[222] dec_out[223] dec_out[224] dec_out[225] dec_out[226] dec_out[227] dec_out[228] dec_out[229] dec_out[230] dec_out[231] dec_out[232] dec_out[233] dec_out[234] dec_out[235] dec_out[236] dec_out[237] dec_out[238] dec_out[239] dec_out[240] dec_out[241] dec_out[242] dec_out[243] dec_out[244] dec_out[245] dec_out[246] dec_out[247] dec_out[248] dec_out[249] dec_out[250] dec_out[251] dec_out[252] dec_out[253] dec_out[254] dec_out[255] vdd gnd hierarchical_decoder_256rows
Xwordline_driver dec_out[0] dec_out[1] dec_out[2] dec_out[3] dec_out[4] dec_out[5] dec_out[6] dec_out[7] dec_out[8] dec_out[9] dec_out[10] dec_out[11] dec_out[12] dec_out[13] dec_out[14] dec_out[15] dec_out[16] dec_out[17] dec_out[18] dec_out[19] dec_out[20] dec_out[21] dec_out[22] dec_out[23] dec_out[24] dec_out[25] dec_out[26] dec_out[27] dec_out[28] dec_out[29] dec_out[30] dec_out[31] dec_out[32] dec_out[33] dec_out[34] dec_out[35] dec_out[36] dec_out[37] dec_out[38] dec_out[39] dec_out[40] dec_out[41] dec_out[42] dec_out[43] dec_out[44] dec_out[45] dec_out[46] dec_out[47] dec_out[48] dec_out[49] dec_out[50] dec_out[51] dec_out[52] dec_out[53] dec_out[54] dec_out[55] dec_out[56] dec_out[57] dec_out[58] dec_out[59] dec_out[60] dec_out[61] dec_out[62] dec_out[63] dec_out[64] dec_out[65] dec_out[66] dec_out[67] dec_out[68] dec_out[69] dec_out[70] dec_out[71] dec_out[72] dec_out[73] dec_out[74] dec_out[75] dec_out[76] dec_out[77] dec_out[78] dec_out[79] dec_out[80] dec_out[81] dec_out[82] dec_out[83] dec_out[84] dec_out[85] dec_out[86] dec_out[87] dec_out[88] dec_out[89] dec_out[90] dec_out[91] dec_out[92] dec_out[93] dec_out[94] dec_out[95] dec_out[96] dec_out[97] dec_out[98] dec_out[99] dec_out[100] dec_out[101] dec_out[102] dec_out[103] dec_out[104] dec_out[105] dec_out[106] dec_out[107] dec_out[108] dec_out[109] dec_out[110] dec_out[111] dec_out[112] dec_out[113] dec_out[114] dec_out[115] dec_out[116] dec_out[117] dec_out[118] dec_out[119] dec_out[120] dec_out[121] dec_out[122] dec_out[123] dec_out[124] dec_out[125] dec_out[126] dec_out[127] dec_out[128] dec_out[129] dec_out[130] dec_out[131] dec_out[132] dec_out[133] dec_out[134] dec_out[135] dec_out[136] dec_out[137] dec_out[138] dec_out[139] dec_out[140] dec_out[141] dec_out[142] dec_out[143] dec_out[144] dec_out[145] dec_out[146] dec_out[147] dec_out[148] dec_out[149] dec_out[150] dec_out[151] dec_out[152] dec_out[153] dec_out[154] dec_out[155] dec_out[156] dec_out[157] dec_out[158] dec_out[159] dec_out[160] dec_out[161] dec_out[162] dec_out[163] dec_out[164] dec_out[165] dec_out[166] dec_out[167] dec_out[168] dec_out[169] dec_out[170] dec_out[171] dec_out[172] dec_out[173] dec_out[174] dec_out[175] dec_out[176] dec_out[177] dec_out[178] dec_out[179] dec_out[180] dec_out[181] dec_out[182] dec_out[183] dec_out[184] dec_out[185] dec_out[186] dec_out[187] dec_out[188] dec_out[189] dec_out[190] dec_out[191] dec_out[192] dec_out[193] dec_out[194] dec_out[195] dec_out[196] dec_out[197] dec_out[198] dec_out[199] dec_out[200] dec_out[201] dec_out[202] dec_out[203] dec_out[204] dec_out[205] dec_out[206] dec_out[207] dec_out[208] dec_out[209] dec_out[210] dec_out[211] dec_out[212] dec_out[213] dec_out[214] dec_out[215] dec_out[216] dec_out[217] dec_out[218] dec_out[219] dec_out[220] dec_out[221] dec_out[222] dec_out[223] dec_out[224] dec_out[225] dec_out[226] dec_out[227] dec_out[228] dec_out[229] dec_out[230] dec_out[231] dec_out[232] dec_out[233] dec_out[234] dec_out[235] dec_out[236] dec_out[237] dec_out[238] dec_out[239] dec_out[240] dec_out[241] dec_out[242] dec_out[243] dec_out[244] dec_out[245] dec_out[246] dec_out[247] dec_out[248] dec_out[249] dec_out[250] dec_out[251] dec_out[252] dec_out[253] dec_out[254] dec_out[255] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] clk_buf vdd gnd wordline_driver
Xaddress_flop_array ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] ADDR[9] A[0] A_bar[0] A[1] A_bar[1] A[2] A_bar[2] A[3] A_bar[3] A[4] A_bar[4] A[5] A_bar[5] A[6] A_bar[6] A[7] A_bar[7] A[8] A_bar[8] A[9] A_bar[9] clk_buf vdd gnd msf_address
.ENDS bank

.SUBCKT sram_1rw_32b_1024w_1bank_freepdk45 DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] ADDR[9] CSb WEb OEb clk vdd gnd
Xbank0 DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] ADDR[9] s_en w_en tri_en_bar tri_en clk_bar clk_buf vdd gnd bank
Xcontrol CSb WEb OEb clk s_en w_en tri_en tri_en_bar clk_bar clk_buf vdd gnd control_logic
.ENDS sram_1rw_32b_1024w_1bank_freepdk45
