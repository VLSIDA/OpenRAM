VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_2_16_scn4m_subm
   CLASS BLOCK ;
   SIZE 229.4 BY 372.8 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  193.4 56.6 194.2 57.4 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  215.2 56.6 216.0 57.4 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  72.4 301.4 73.2 302.2 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  72.4 323.4 73.2 324.2 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  72.4 341.4 73.2 342.2 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  72.4 363.4 73.2 364.2 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  10.4 10.8 11.2 11.6 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  10.4 32.8 11.2 33.6 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  51.5 2.2 52.1 12.0 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal2 ;
         RECT  200.0 119.8 200.8 122.8 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal2 ;
         RECT  206.8 119.8 207.6 122.8 ;
      END
   END dout0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  195.6 308.2 196.4 309.0 ;
         LAYER metal3 ;
         RECT  218.1 67.6 218.9 68.4 ;
         LAYER metal4 ;
         RECT  28.8 0.0 30.0 370.8 ;
         LAYER metal3 ;
         RECT  202.7 98.7 203.3 99.3 ;
         LAYER metal3 ;
         RECT  195.6 245.8 196.4 246.6 ;
         LAYER metal3 ;
         RECT  2.4 132.0 32.4 133.2 ;
         LAYER metal3 ;
         RECT  21.6 195.8 22.4 196.6 ;
         LAYER metal3 ;
         RECT  105.3 267.0 106.1 267.8 ;
         LAYER metal3 ;
         RECT  8.8 216.6 9.6 217.4 ;
         LAYER metal4 ;
         RECT  148.8 0.0 150.0 370.8 ;
         LAYER metal4 ;
         RECT  48.0 0.0 49.2 370.8 ;
         LAYER metal3 ;
         RECT  8.8 237.4 9.6 238.2 ;
         LAYER metal3 ;
         RECT  88.8 40.8 226.8 42.0 ;
         LAYER metal3 ;
         RECT  122.7 225.4 123.5 226.2 ;
         LAYER metal4 ;
         RECT  19.2 0.0 20.4 370.8 ;
         LAYER metal3 ;
         RECT  195.6 204.2 196.4 205.0 ;
         LAYER metal4 ;
         RECT  24.0 0.0 25.2 370.8 ;
         LAYER metal4 ;
         RECT  211.2 0.0 212.4 370.8 ;
         LAYER metal3 ;
         RECT  187.2 74.4 226.8 75.6 ;
         LAYER metal3 ;
         RECT  145.7 246.2 146.5 247.0 ;
         LAYER metal3 ;
         RECT  2.4 36.0 42.0 37.2 ;
         LAYER metal3 ;
         RECT  79.2 50.4 226.8 51.6 ;
         LAYER metal3 ;
         RECT  33.6 242.4 181.2 243.6 ;
         LAYER metal3 ;
         RECT  202.5 370.7 203.1 371.3 ;
         LAYER metal4 ;
         RECT  168.0 0.0 169.2 370.8 ;
         LAYER metal3 ;
         RECT  75.3 352.4 76.1 353.2 ;
         LAYER metal3 ;
         RECT  209.5 98.7 210.1 99.3 ;
         LAYER metal3 ;
         RECT  177.6 276.0 226.8 277.2 ;
         LAYER metal3 ;
         RECT  187.2 112.8 226.8 114.0 ;
         LAYER metal3 ;
         RECT  196.3 67.6 197.1 68.4 ;
         LAYER metal3 ;
         RECT  195.6 266.6 196.4 267.4 ;
         LAYER metal3 ;
         RECT  79.2 333.6 181.2 334.8 ;
         LAYER metal3 ;
         RECT  21.6 258.2 22.4 259.0 ;
         LAYER metal3 ;
         RECT  24.0 247.2 87.6 248.4 ;
         LAYER metal3 ;
         RECT  209.3 266.7 209.9 267.3 ;
         LAYER metal3 ;
         RECT  202.5 308.3 203.1 308.9 ;
         LAYER metal4 ;
         RECT  43.2 0.0 44.4 370.8 ;
         LAYER metal3 ;
         RECT  2.4 136.8 226.8 138.0 ;
         LAYER metal3 ;
         RECT  209.3 329.1 209.9 329.7 ;
         LAYER metal3 ;
         RECT  55.2 132.0 226.8 133.2 ;
         LAYER metal3 ;
         RECT  98.4 343.2 181.2 344.4 ;
         LAYER metal4 ;
         RECT  144.0 0.0 145.2 370.8 ;
         LAYER metal3 ;
         RECT  216.1 329.1 216.7 329.7 ;
         LAYER metal4 ;
         RECT  105.6 0.0 106.8 370.8 ;
         LAYER metal3 ;
         RECT  15.2 237.4 16.0 238.2 ;
         LAYER metal3 ;
         RECT  2.4 88.8 82.8 90.0 ;
         LAYER metal3 ;
         RECT  2.4 108.0 198.0 109.2 ;
         LAYER metal3 ;
         RECT  216.1 266.7 216.7 267.3 ;
         LAYER metal3 ;
         RECT  202.5 225.1 203.1 225.7 ;
         LAYER metal3 ;
         RECT  2.4 21.6 226.8 22.8 ;
         LAYER metal3 ;
         RECT  8.8 195.8 9.6 196.6 ;
         LAYER metal3 ;
         RECT  2.4 146.4 200.4 147.6 ;
         LAYER metal3 ;
         RECT  2.4 352.8 181.2 354.0 ;
         LAYER metal4 ;
         RECT  76.8 0.0 78.0 370.8 ;
         LAYER metal3 ;
         RECT  177.6 300.0 226.8 301.2 ;
         LAYER metal3 ;
         RECT  2.4 156.0 226.8 157.2 ;
         LAYER metal4 ;
         RECT  14.4 0.0 15.6 370.8 ;
         LAYER metal4 ;
         RECT  110.4 0.0 111.6 370.8 ;
         LAYER metal3 ;
         RECT  2.4 324.0 78.0 325.2 ;
         LAYER metal3 ;
         RECT  209.3 308.3 209.9 308.9 ;
         LAYER metal3 ;
         RECT  202.5 183.5 203.1 184.1 ;
         LAYER metal3 ;
         RECT  122.7 204.6 123.5 205.4 ;
         LAYER metal3 ;
         RECT  21.6 175.0 22.4 175.8 ;
         LAYER metal3 ;
         RECT  33.6 170.4 226.8 171.6 ;
         LAYER metal4 ;
         RECT  33.6 0.0 34.8 370.8 ;
         LAYER metal4 ;
         RECT  139.2 0.0 140.4 370.8 ;
         LAYER metal3 ;
         RECT  8.8 258.2 9.6 259.0 ;
         LAYER metal3 ;
         RECT  209.3 370.7 209.9 371.3 ;
         LAYER metal3 ;
         RECT  145.7 350.2 146.5 351.0 ;
         LAYER metal3 ;
         RECT  145.7 308.6 146.5 309.4 ;
         LAYER metal3 ;
         RECT  75.3 312.4 76.1 313.2 ;
         LAYER metal3 ;
         RECT  88.8 2.4 226.8 3.6 ;
         LAYER metal3 ;
         RECT  199.2 165.6 226.8 166.8 ;
         LAYER metal3 ;
         RECT  2.4 194.4 99.6 195.6 ;
         LAYER metal4 ;
         RECT  129.6 0.0 130.8 370.8 ;
         LAYER metal4 ;
         RECT  158.4 0.0 159.6 370.8 ;
         LAYER metal3 ;
         RECT  33.6 189.6 181.2 190.8 ;
         LAYER metal3 ;
         RECT  209.0 163.0 209.8 163.8 ;
         LAYER metal3 ;
         RECT  216.1 204.3 216.7 204.9 ;
         LAYER metal3 ;
         RECT  2.4 50.4 37.2 51.6 ;
         LAYER metal3 ;
         RECT  202.5 329.1 203.1 329.7 ;
         LAYER metal3 ;
         RECT  2.4 348.0 226.8 349.2 ;
         LAYER metal3 ;
         RECT  209.3 287.5 209.9 288.1 ;
         LAYER metal3 ;
         RECT  2.4 218.4 181.2 219.6 ;
         LAYER metal3 ;
         RECT  173.1 246.2 173.9 247.0 ;
         LAYER metal3 ;
         RECT  79.2 290.4 181.2 291.6 ;
         LAYER metal3 ;
         RECT  24.0 184.8 226.8 186.0 ;
         LAYER metal3 ;
         RECT  2.4 338.4 140.4 339.6 ;
         LAYER metal3 ;
         RECT  2.4 64.8 226.8 66.0 ;
         LAYER metal3 ;
         RECT  2.4 141.6 226.8 142.8 ;
         LAYER metal3 ;
         RECT  195.6 225.0 196.4 225.8 ;
         LAYER metal3 ;
         RECT  177.6 237.6 226.8 238.8 ;
         LAYER metal3 ;
         RECT  188.9 329.1 189.5 329.7 ;
         LAYER metal3 ;
         RECT  203.3 81.3 203.9 81.9 ;
         LAYER metal3 ;
         RECT  2.4 208.8 181.2 210.0 ;
         LAYER metal4 ;
         RECT  9.6 0.0 10.8 370.8 ;
         LAYER metal4 ;
         RECT  62.4 0.0 63.6 370.8 ;
         LAYER metal3 ;
         RECT  202.5 204.3 203.1 204.9 ;
         LAYER metal3 ;
         RECT  2.4 45.6 190.8 46.8 ;
         LAYER metal3 ;
         RECT  2.4 237.6 99.6 238.8 ;
         LAYER metal4 ;
         RECT  120.0 0.0 121.2 370.8 ;
         LAYER metal3 ;
         RECT  15.2 258.2 16.0 259.0 ;
         LAYER metal3 ;
         RECT  173.1 204.6 173.9 205.4 ;
         LAYER metal3 ;
         RECT  145.7 287.8 146.5 288.6 ;
         LAYER metal3 ;
         RECT  33.6 252.0 181.2 253.2 ;
         LAYER metal3 ;
         RECT  2.4 276.0 99.6 277.2 ;
         LAYER metal3 ;
         RECT  216.1 308.3 216.7 308.9 ;
         LAYER metal4 ;
         RECT  96.0 0.0 97.2 370.8 ;
         LAYER metal4 ;
         RECT  201.6 0.0 202.8 370.8 ;
         LAYER metal3 ;
         RECT  173.1 329.4 173.9 330.2 ;
         LAYER metal4 ;
         RECT  100.8 0.0 102.0 370.8 ;
         LAYER metal4 ;
         RECT  196.8 0.0 198.0 370.8 ;
         LAYER metal3 ;
         RECT  177.6 362.4 226.8 363.6 ;
         LAYER metal3 ;
         RECT  195.6 329.0 196.4 329.8 ;
         LAYER metal3 ;
         RECT  84.8 101.8 85.6 102.6 ;
         LAYER metal3 ;
         RECT  209.3 225.1 209.9 225.7 ;
         LAYER metal4 ;
         RECT  86.4 0.0 87.6 370.8 ;
         LAYER metal3 ;
         RECT  2.4 213.6 99.6 214.8 ;
         LAYER metal4 ;
         RECT  187.2 0.0 188.4 370.8 ;
         LAYER metal4 ;
         RECT  225.6 0.0 226.8 370.8 ;
         LAYER metal3 ;
         RECT  2.4 69.6 226.8 70.8 ;
         LAYER metal3 ;
         RECT  2.4 271.2 181.2 272.4 ;
         LAYER metal3 ;
         RECT  2.4 300.0 140.4 301.2 ;
         LAYER metal3 ;
         RECT  202.5 287.5 203.1 288.1 ;
         LAYER metal3 ;
         RECT  2.4 74.4 82.8 75.6 ;
         LAYER metal4 ;
         RECT  57.6 0.0 58.8 370.8 ;
         LAYER metal3 ;
         RECT  2.4 21.8 3.2 22.6 ;
         LAYER metal4 ;
         RECT  182.4 0.0 183.6 370.8 ;
         LAYER metal3 ;
         RECT  216.1 225.1 216.7 225.7 ;
         LAYER metal3 ;
         RECT  145.7 225.4 146.5 226.2 ;
         LAYER metal3 ;
         RECT  216.1 349.9 216.7 350.5 ;
         LAYER metal3 ;
         RECT  195.6 183.4 196.4 184.2 ;
         LAYER metal4 ;
         RECT  91.2 0.0 92.4 370.8 ;
         LAYER metal3 ;
         RECT  210.1 81.3 210.7 81.9 ;
         LAYER metal3 ;
         RECT  2.4 295.2 226.8 296.4 ;
         LAYER metal4 ;
         RECT  67.2 0.0 68.4 370.8 ;
         LAYER metal3 ;
         RECT  195.6 349.8 196.4 350.6 ;
         LAYER metal3 ;
         RECT  209.3 183.5 209.9 184.1 ;
         LAYER metal3 ;
         RECT  33.6 223.2 121.2 224.4 ;
         LAYER metal3 ;
         RECT  177.6 338.4 226.8 339.6 ;
         LAYER metal3 ;
         RECT  209.3 204.3 209.9 204.9 ;
         LAYER metal3 ;
         RECT  202.5 349.9 203.1 350.5 ;
         LAYER metal4 ;
         RECT  192.0 0.0 193.2 370.8 ;
         LAYER metal3 ;
         RECT  84.8 21.8 85.6 22.6 ;
         LAYER metal3 ;
         RECT  60.0 36.0 226.8 37.2 ;
         LAYER metal3 ;
         RECT  204.9 132.7 205.5 133.3 ;
         LAYER metal3 ;
         RECT  2.4 55.2 226.8 56.4 ;
         LAYER metal3 ;
         RECT  21.6 237.4 22.4 238.2 ;
         LAYER metal3 ;
         RECT  177.6 256.8 226.8 258.0 ;
         LAYER metal3 ;
         RECT  2.4 26.4 226.8 27.6 ;
         LAYER metal3 ;
         RECT  2.4 285.6 226.8 286.8 ;
         LAYER metal4 ;
         RECT  220.8 0.0 222.0 370.8 ;
         LAYER metal3 ;
         RECT  188.9 349.9 189.5 350.5 ;
         LAYER metal3 ;
         RECT  2.4 98.4 226.8 99.6 ;
         LAYER metal4 ;
         RECT  38.4 0.0 39.6 370.8 ;
         LAYER metal3 ;
         RECT  96.0 324.0 181.2 325.2 ;
         LAYER metal3 ;
         RECT  84.8 61.8 85.6 62.6 ;
         LAYER metal3 ;
         RECT  145.7 329.4 146.5 330.2 ;
         LAYER metal4 ;
         RECT  124.8 0.0 126.0 370.8 ;
         LAYER metal4 ;
         RECT  206.4 0.0 207.6 370.8 ;
         LAYER metal3 ;
         RECT  139.2 223.2 226.8 224.4 ;
         LAYER metal3 ;
         RECT  84.0 31.2 226.8 32.4 ;
         LAYER metal3 ;
         RECT  177.6 213.6 226.8 214.8 ;
         LAYER metal3 ;
         RECT  209.3 245.9 209.9 246.5 ;
         LAYER metal3 ;
         RECT  15.2 195.8 16.0 196.6 ;
         LAYER metal3 ;
         RECT  2.4 343.2 78.0 344.4 ;
         LAYER metal3 ;
         RECT  2.4 175.2 226.8 176.4 ;
         LAYER metal3 ;
         RECT  84.8 141.8 85.6 142.6 ;
         LAYER metal3 ;
         RECT  173.1 350.2 173.9 351.0 ;
         LAYER metal3 ;
         RECT  33.6 180.0 181.2 181.2 ;
         LAYER metal3 ;
         RECT  216.1 245.9 216.7 246.5 ;
         LAYER metal3 ;
         RECT  122.7 267.0 123.5 267.8 ;
         LAYER metal3 ;
         RECT  195.6 370.6 196.4 371.4 ;
         LAYER metal3 ;
         RECT  8.8 175.0 9.6 175.8 ;
         LAYER metal3 ;
         RECT  2.4 122.4 80.4 123.6 ;
         LAYER metal3 ;
         RECT  88.8 122.4 226.8 123.6 ;
         LAYER metal4 ;
         RECT  72.0 0.0 73.2 370.8 ;
         LAYER metal3 ;
         RECT  105.3 246.2 106.1 247.0 ;
         LAYER metal3 ;
         RECT  177.6 194.4 226.8 195.6 ;
         LAYER metal4 ;
         RECT  81.6 0.0 82.8 370.8 ;
         LAYER metal4 ;
         RECT  163.2 0.0 164.4 370.8 ;
         LAYER metal3 ;
         RECT  136.8 204.0 226.8 205.2 ;
         LAYER metal3 ;
         RECT  188.9 204.3 189.5 204.9 ;
         LAYER metal4 ;
         RECT  172.8 0.0 174.0 370.8 ;
         LAYER metal3 ;
         RECT  4.8 40.8 80.4 42.0 ;
         LAYER metal3 ;
         RECT  145.7 204.6 146.5 205.4 ;
         LAYER metal3 ;
         RECT  145.7 267.0 146.5 267.8 ;
         LAYER metal3 ;
         RECT  173.1 225.4 173.9 226.2 ;
         LAYER metal3 ;
         RECT  50.4 12.0 226.8 13.2 ;
         LAYER metal3 ;
         RECT  184.8 151.2 226.8 152.4 ;
         LAYER metal4 ;
         RECT  4.8 0.0 6.0 370.8 ;
         LAYER metal4 ;
         RECT  52.8 0.0 54.0 370.8 ;
         LAYER metal3 ;
         RECT  144.0 266.4 226.8 267.6 ;
         LAYER metal3 ;
         RECT  4.8 2.4 80.4 3.6 ;
         LAYER metal3 ;
         RECT  188.9 225.1 189.5 225.7 ;
         LAYER metal3 ;
         RECT  33.6 199.2 181.2 200.4 ;
         LAYER metal4 ;
         RECT  153.6 0.0 154.8 370.8 ;
         LAYER metal3 ;
         RECT  216.1 370.7 216.7 371.3 ;
         LAYER metal3 ;
         RECT  2.4 112.8 82.8 114.0 ;
         LAYER metal3 ;
         RECT  21.6 204.0 85.2 205.2 ;
         LAYER metal3 ;
         RECT  2.4 60.0 226.8 61.2 ;
         LAYER metal3 ;
         RECT  2.4 280.8 181.2 282.0 ;
         LAYER metal3 ;
         RECT  2.4 266.4 121.2 267.6 ;
         LAYER metal3 ;
         RECT  188.9 287.5 189.5 288.1 ;
         LAYER metal3 ;
         RECT  105.3 204.6 106.1 205.4 ;
         LAYER metal3 ;
         RECT  188.9 370.7 189.5 371.3 ;
         LAYER metal3 ;
         RECT  2.4 151.2 82.8 152.4 ;
         LAYER metal3 ;
         RECT  33.6 232.8 226.8 234.0 ;
         LAYER metal3 ;
         RECT  202.2 163.0 203.0 163.8 ;
         LAYER metal3 ;
         RECT  2.4 160.8 80.4 162.0 ;
         LAYER metal3 ;
         RECT  2.4 7.2 226.8 8.4 ;
         LAYER metal3 ;
         RECT  88.8 160.8 226.8 162.0 ;
         LAYER metal3 ;
         RECT  2.4 16.8 226.8 18.0 ;
         LAYER metal3 ;
         RECT  2.4 314.4 181.2 315.6 ;
         LAYER metal3 ;
         RECT  2.4 256.8 90.0 258.0 ;
         LAYER metal3 ;
         RECT  2.4 309.6 226.8 310.8 ;
         LAYER metal3 ;
         RECT  2.4 84.0 226.8 85.2 ;
         LAYER metal3 ;
         RECT  173.1 287.8 173.9 288.6 ;
         LAYER metal3 ;
         RECT  15.2 175.0 16.0 175.8 ;
         LAYER metal3 ;
         RECT  2.4 117.6 226.8 118.8 ;
         LAYER metal4 ;
         RECT  115.2 0.0 116.4 370.8 ;
         LAYER metal4 ;
         RECT  216.0 0.0 217.2 370.8 ;
         LAYER metal3 ;
         RECT  2.4 304.8 181.2 306.0 ;
         LAYER metal3 ;
         RECT  202.5 245.9 203.1 246.5 ;
         LAYER metal3 ;
         RECT  216.1 287.5 216.7 288.1 ;
         LAYER metal3 ;
         RECT  188.9 308.3 189.5 308.9 ;
         LAYER metal3 ;
         RECT  24.0 228.0 181.2 229.2 ;
         LAYER metal3 ;
         RECT  188.9 245.9 189.5 246.5 ;
         LAYER metal3 ;
         RECT  211.7 132.7 212.3 133.3 ;
         LAYER metal3 ;
         RECT  21.6 216.6 22.4 217.4 ;
         LAYER metal3 ;
         RECT  2.4 328.8 226.8 330.0 ;
         LAYER metal3 ;
         RECT  122.7 246.2 123.5 247.0 ;
         LAYER metal3 ;
         RECT  2.4 290.4 70.8 291.6 ;
         LAYER metal3 ;
         RECT  2.4 362.4 78.0 363.6 ;
         LAYER metal3 ;
         RECT  2.4 79.2 226.8 80.4 ;
         LAYER metal3 ;
         RECT  105.3 225.4 106.1 226.2 ;
         LAYER metal3 ;
         RECT  2.4 127.2 226.8 128.4 ;
         LAYER metal3 ;
         RECT  195.6 287.4 196.4 288.2 ;
         LAYER metal3 ;
         RECT  2.4 367.2 181.2 368.4 ;
         LAYER metal3 ;
         RECT  2.4 261.6 181.2 262.8 ;
         LAYER metal3 ;
         RECT  188.9 183.5 189.5 184.1 ;
         LAYER metal3 ;
         RECT  15.2 216.6 16.0 217.4 ;
         LAYER metal3 ;
         RECT  2.4 103.2 226.8 104.4 ;
         LAYER metal3 ;
         RECT  2.4 93.6 200.4 94.8 ;
         LAYER metal3 ;
         RECT  98.4 362.4 140.4 363.6 ;
         LAYER metal3 ;
         RECT  177.6 319.2 226.8 320.4 ;
         LAYER metal3 ;
         RECT  173.1 267.0 173.9 267.8 ;
         LAYER metal3 ;
         RECT  209.3 349.9 209.9 350.5 ;
         LAYER metal3 ;
         RECT  173.1 308.6 173.9 309.4 ;
         LAYER metal3 ;
         RECT  216.1 183.5 216.7 184.1 ;
         LAYER metal3 ;
         RECT  141.6 247.2 226.8 248.4 ;
         LAYER metal3 ;
         RECT  2.4 357.6 226.8 358.8 ;
         LAYER metal3 ;
         RECT  188.9 266.7 189.5 267.3 ;
         LAYER metal3 ;
         RECT  2.4 333.6 70.8 334.8 ;
         LAYER metal4 ;
         RECT  177.6 0.0 178.8 370.8 ;
         LAYER metal3 ;
         RECT  202.5 266.7 203.1 267.3 ;
         LAYER metal3 ;
         RECT  195.4 163.0 196.2 163.8 ;
         LAYER metal3 ;
         RECT  2.4 319.2 140.4 320.4 ;
         LAYER metal4 ;
         RECT  134.4 0.0 135.6 370.8 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  98.4 340.8 226.8 342.0 ;
         LAYER metal3 ;
         RECT  84.0 33.6 226.8 34.8 ;
         LAYER metal3 ;
         RECT  2.4 163.2 190.8 164.4 ;
         LAYER metal4 ;
         RECT  108.0 0.0 109.2 370.8 ;
         LAYER metal3 ;
         RECT  192.2 261.6 193.0 262.4 ;
         LAYER metal4 ;
         RECT  199.2 0.0 200.4 370.8 ;
         LAYER metal3 ;
         RECT  219.5 250.9 220.1 251.5 ;
         LAYER metal3 ;
         RECT  105.3 256.6 106.1 257.4 ;
         LAYER metal4 ;
         RECT  93.6 0.0 94.8 370.8 ;
         LAYER metal3 ;
         RECT  219.5 240.9 220.1 241.5 ;
         LAYER metal3 ;
         RECT  2.4 182.4 183.6 183.6 ;
         LAYER metal3 ;
         RECT  192.3 220.1 192.9 220.7 ;
         LAYER metal3 ;
         RECT  199.1 324.1 199.7 324.7 ;
         LAYER metal3 ;
         RECT  45.6 28.8 226.8 30.0 ;
         LAYER metal3 ;
         RECT  2.4 76.8 226.8 78.0 ;
         LAYER metal3 ;
         RECT  201.9 106.9 202.5 107.5 ;
         LAYER metal3 ;
         RECT  219.5 344.9 220.1 345.5 ;
         LAYER metal3 ;
         RECT  21.6 172.8 226.8 174.0 ;
         LAYER metal4 ;
         RECT  79.2 0.0 80.4 370.8 ;
         LAYER metal4 ;
         RECT  7.2 0.0 8.4 370.8 ;
         LAYER metal3 ;
         RECT  219.5 282.5 220.1 283.1 ;
         LAYER metal3 ;
         RECT  219.5 324.1 220.1 324.7 ;
         LAYER metal3 ;
         RECT  184.8 91.2 226.8 92.4 ;
         LAYER metal3 ;
         RECT  212.7 220.1 213.3 220.7 ;
         LAYER metal3 ;
         RECT  199.1 240.9 199.7 241.5 ;
         LAYER metal3 ;
         RECT  105.3 235.8 106.1 236.6 ;
         LAYER metal3 ;
         RECT  212.7 209.3 213.3 209.9 ;
         LAYER metal3 ;
         RECT  173.1 235.8 173.9 236.6 ;
         LAYER metal3 ;
         RECT  24.0 259.2 90.0 260.4 ;
         LAYER metal4 ;
         RECT  180.0 0.0 181.2 370.8 ;
         LAYER metal3 ;
         RECT  205.9 209.3 206.5 209.9 ;
         LAYER metal3 ;
         RECT  8.8 164.6 9.6 165.4 ;
         LAYER metal3 ;
         RECT  219.5 271.7 220.1 272.3 ;
         LAYER metal3 ;
         RECT  2.4 91.2 82.8 92.4 ;
         LAYER metal3 ;
         RECT  173.1 194.2 173.9 195.0 ;
         LAYER metal3 ;
         RECT  212.7 188.5 213.3 189.1 ;
         LAYER metal3 ;
         RECT  192.3 230.1 192.9 230.7 ;
         LAYER metal3 ;
         RECT  219.5 334.1 220.1 334.7 ;
         LAYER metal3 ;
         RECT  192.2 292.4 193.0 293.2 ;
         LAYER metal3 ;
         RECT  205.9 220.1 206.5 220.7 ;
         LAYER metal3 ;
         RECT  219.5 292.5 220.1 293.1 ;
         LAYER metal3 ;
         RECT  2.4 24.0 226.8 25.2 ;
         LAYER metal3 ;
         RECT  173.1 360.6 173.9 361.4 ;
         LAYER metal3 ;
         RECT  2.4 96.0 226.8 97.2 ;
         LAYER metal3 ;
         RECT  185.5 324.1 186.1 324.7 ;
         LAYER metal3 ;
         RECT  173.1 298.2 173.9 299.0 ;
         LAYER metal3 ;
         RECT  199.1 271.7 199.7 272.3 ;
         LAYER metal3 ;
         RECT  145.7 235.8 146.5 236.6 ;
         LAYER metal3 ;
         RECT  199.0 230.0 199.8 230.8 ;
         LAYER metal3 ;
         RECT  192.3 261.7 192.9 262.3 ;
         LAYER metal3 ;
         RECT  145.7 194.2 146.5 195.0 ;
         LAYER metal3 ;
         RECT  173.1 256.6 173.9 257.4 ;
         LAYER metal3 ;
         RECT  185.5 344.9 186.1 345.5 ;
         LAYER metal3 ;
         RECT  2.4 312.0 70.8 313.2 ;
         LAYER metal3 ;
         RECT  21.6 185.4 22.4 186.2 ;
         LAYER metal3 ;
         RECT  76.8 312.0 226.8 313.2 ;
         LAYER metal3 ;
         RECT  192.3 240.9 192.9 241.5 ;
         LAYER metal3 ;
         RECT  105.3 215.0 106.1 215.8 ;
         LAYER metal4 ;
         RECT  127.2 0.0 128.4 370.8 ;
         LAYER metal3 ;
         RECT  205.9 188.5 206.5 189.1 ;
         LAYER metal3 ;
         RECT  199.0 240.8 199.8 241.6 ;
         LAYER metal3 ;
         RECT  212.7 250.9 213.3 251.5 ;
         LAYER metal3 ;
         RECT  75.3 372.4 76.1 373.2 ;
         LAYER metal3 ;
         RECT  2.4 206.4 85.2 207.6 ;
         LAYER metal3 ;
         RECT  212.7 146.1 213.3 146.7 ;
         LAYER metal3 ;
         RECT  212.7 292.5 213.3 293.1 ;
         LAYER metal3 ;
         RECT  192.3 188.5 192.9 189.1 ;
         LAYER metal3 ;
         RECT  219.5 188.5 220.1 189.1 ;
         LAYER metal3 ;
         RECT  192.2 250.8 193.0 251.6 ;
         LAYER metal3 ;
         RECT  185.5 188.5 186.1 189.1 ;
         LAYER metal3 ;
         RECT  2.4 105.6 226.8 106.8 ;
         LAYER metal4 ;
         RECT  170.4 0.0 171.6 370.8 ;
         LAYER metal3 ;
         RECT  205.9 250.9 206.5 251.5 ;
         LAYER metal3 ;
         RECT  8.8 227.0 9.6 227.8 ;
         LAYER metal3 ;
         RECT  192.2 282.4 193.0 283.2 ;
         LAYER metal3 ;
         RECT  93.6 297.6 226.8 298.8 ;
         LAYER metal4 ;
         RECT  69.6 0.0 70.8 370.8 ;
         LAYER metal3 ;
         RECT  105.3 277.4 106.1 278.2 ;
         LAYER metal3 ;
         RECT  2.4 1.8 3.2 2.6 ;
         LAYER metal3 ;
         RECT  8.8 247.8 9.6 248.6 ;
         LAYER metal3 ;
         RECT  21.6 247.8 22.4 248.6 ;
         LAYER metal3 ;
         RECT  2.4 278.4 121.2 279.6 ;
         LAYER metal4 ;
         RECT  103.2 0.0 104.4 370.8 ;
         LAYER metal3 ;
         RECT  8.8 206.2 9.6 207.0 ;
         LAYER metal3 ;
         RECT  199.1 178.5 199.7 179.1 ;
         LAYER metal3 ;
         RECT  199.1 282.5 199.7 283.1 ;
         LAYER metal3 ;
         RECT  204.7 92.3 205.3 92.9 ;
         LAYER metal3 ;
         RECT  185.5 178.5 186.1 179.1 ;
         LAYER metal3 ;
         RECT  75.3 332.4 76.1 333.2 ;
         LAYER metal3 ;
         RECT  145.7 215.0 146.5 215.8 ;
         LAYER metal3 ;
         RECT  199.0 282.4 199.8 283.2 ;
         LAYER metal4 ;
         RECT  64.8 0.0 66.0 370.8 ;
         LAYER metal3 ;
         RECT  2.4 307.2 140.4 308.4 ;
         LAYER metal3 ;
         RECT  2.4 187.2 226.8 188.4 ;
         LAYER metal3 ;
         RECT  219.5 220.1 220.1 220.7 ;
         LAYER metal4 ;
         RECT  165.6 0.0 166.8 370.8 ;
         LAYER metal3 ;
         RECT  205.9 271.7 206.5 272.3 ;
         LAYER metal3 ;
         RECT  15.2 227.0 16.0 227.8 ;
         LAYER metal3 ;
         RECT  2.4 264.0 226.8 265.2 ;
         LAYER metal3 ;
         RECT  2.4 283.2 226.8 284.4 ;
         LAYER metal4 ;
         RECT  60.0 0.0 61.2 370.8 ;
         LAYER metal3 ;
         RECT  212.7 240.9 213.3 241.5 ;
         LAYER metal3 ;
         RECT  139.2 235.2 226.8 236.4 ;
         LAYER metal3 ;
         RECT  212.7 344.9 213.3 345.5 ;
         LAYER metal3 ;
         RECT  122.7 194.2 123.5 195.0 ;
         LAYER metal3 ;
         RECT  192.3 292.5 192.9 293.1 ;
         LAYER metal3 ;
         RECT  192.2 334.0 193.0 334.8 ;
         LAYER metal4 ;
         RECT  16.8 0.0 18.0 370.8 ;
         LAYER metal3 ;
         RECT  192.2 303.2 193.0 304.0 ;
         LAYER metal3 ;
         RECT  211.5 92.3 212.1 92.9 ;
         LAYER metal3 ;
         RECT  122.7 235.8 123.5 236.6 ;
         LAYER metal4 ;
         RECT  21.6 0.0 22.8 370.8 ;
         LAYER metal3 ;
         RECT  2.4 57.6 226.8 58.8 ;
         LAYER metal3 ;
         RECT  88.8 62.4 226.8 63.6 ;
         LAYER metal3 ;
         RECT  219.5 199.3 220.1 199.9 ;
         LAYER metal4 ;
         RECT  26.4 0.0 27.6 370.8 ;
         LAYER metal3 ;
         RECT  199.0 178.4 199.8 179.2 ;
         LAYER metal3 ;
         RECT  199.1 365.7 199.7 366.3 ;
         LAYER metal3 ;
         RECT  185.5 240.9 186.1 241.5 ;
         LAYER metal3 ;
         RECT  33.6 211.2 226.8 212.4 ;
         LAYER metal3 ;
         RECT  2.4 19.2 226.8 20.4 ;
         LAYER metal3 ;
         RECT  185.5 365.7 186.1 366.3 ;
         LAYER metal3 ;
         RECT  136.8 216.0 226.8 217.2 ;
         LAYER metal3 ;
         RECT  33.6 192.0 226.8 193.2 ;
         LAYER metal4 ;
         RECT  151.2 0.0 152.4 370.8 ;
         LAYER metal3 ;
         RECT  199.0 271.6 199.8 272.4 ;
         LAYER metal3 ;
         RECT  2.4 72.0 82.8 73.2 ;
         LAYER metal3 ;
         RECT  2.4 316.8 226.8 318.0 ;
         LAYER metal3 ;
         RECT  185.5 220.1 186.1 220.7 ;
         LAYER metal3 ;
         RECT  205.9 365.7 206.5 366.3 ;
         LAYER metal3 ;
         RECT  50.4 14.4 226.8 15.6 ;
         LAYER metal3 ;
         RECT  192.3 365.7 192.9 366.3 ;
         LAYER metal3 ;
         RECT  88.8 100.8 226.8 102.0 ;
         LAYER metal4 ;
         RECT  136.8 0.0 138.0 370.8 ;
         LAYER metal3 ;
         RECT  21.6 164.6 22.4 165.4 ;
         LAYER metal3 ;
         RECT  199.0 199.2 199.8 200.0 ;
         LAYER metal3 ;
         RECT  199.0 324.0 199.8 324.8 ;
         LAYER metal3 ;
         RECT  199.0 292.4 199.8 293.2 ;
         LAYER metal4 ;
         RECT  2.4 0.0 3.6 370.8 ;
         LAYER metal3 ;
         RECT  55.2 129.6 226.8 130.8 ;
         LAYER metal3 ;
         RECT  177.6 331.2 226.8 332.4 ;
         LAYER metal3 ;
         RECT  2.4 340.8 78.0 342.0 ;
         LAYER metal3 ;
         RECT  2.4 43.2 226.8 44.4 ;
         LAYER metal4 ;
         RECT  146.4 0.0 147.6 370.8 ;
         LAYER metal3 ;
         RECT  2.4 158.4 226.8 159.6 ;
         LAYER metal3 ;
         RECT  205.9 240.9 206.5 241.5 ;
         LAYER metal3 ;
         RECT  192.2 354.8 193.0 355.6 ;
         LAYER metal4 ;
         RECT  31.2 0.0 32.4 370.8 ;
         LAYER metal3 ;
         RECT  212.7 334.1 213.3 334.7 ;
         LAYER metal3 ;
         RECT  2.4 177.6 226.8 178.8 ;
         LAYER metal3 ;
         RECT  2.4 369.6 183.6 370.8 ;
         LAYER metal3 ;
         RECT  2.4 134.4 200.4 135.6 ;
         LAYER metal3 ;
         RECT  192.2 324.0 193.0 324.8 ;
         LAYER metal4 ;
         RECT  112.8 0.0 114.0 370.8 ;
         LAYER metal4 ;
         RECT  194.4 0.0 195.6 370.8 ;
         LAYER metal4 ;
         RECT  208.8 0.0 210.0 370.8 ;
         LAYER metal3 ;
         RECT  145.7 277.4 146.5 278.2 ;
         LAYER metal3 ;
         RECT  187.2 72.0 226.8 73.2 ;
         LAYER metal3 ;
         RECT  218.1 47.6 218.9 48.4 ;
         LAYER metal3 ;
         RECT  28.8 9.6 226.8 10.8 ;
         LAYER metal3 ;
         RECT  192.2 230.0 193.0 230.8 ;
         LAYER metal3 ;
         RECT  192.3 303.3 192.9 303.9 ;
         LAYER metal3 ;
         RECT  199.0 365.6 199.8 366.4 ;
         LAYER metal3 ;
         RECT  192.2 188.4 193.0 189.2 ;
         LAYER metal4 ;
         RECT  141.6 0.0 142.8 370.8 ;
         LAYER metal3 ;
         RECT  199.0 220.0 199.8 220.8 ;
         LAYER metal3 ;
         RECT  84.8 81.8 85.6 82.6 ;
         LAYER metal3 ;
         RECT  185.5 334.1 186.1 334.7 ;
         LAYER metal3 ;
         RECT  199.0 313.2 199.8 314.0 ;
         LAYER metal3 ;
         RECT  199.1 209.3 199.7 209.9 ;
         LAYER metal3 ;
         RECT  21.6 227.0 22.4 227.8 ;
         LAYER metal3 ;
         RECT  2.4 100.8 80.4 102.0 ;
         LAYER metal3 ;
         RECT  212.7 261.7 213.3 262.3 ;
         LAYER metal3 ;
         RECT  15.2 206.2 16.0 207.0 ;
         LAYER metal3 ;
         RECT  2.4 288.0 140.4 289.2 ;
         LAYER metal3 ;
         RECT  2.4 129.6 32.4 130.8 ;
         LAYER metal3 ;
         RECT  205.9 199.3 206.5 199.9 ;
         LAYER metal3 ;
         RECT  192.3 178.5 192.9 179.1 ;
         LAYER metal3 ;
         RECT  212.7 354.9 213.3 355.5 ;
         LAYER metal3 ;
         RECT  33.6 254.4 226.8 255.6 ;
         LAYER metal3 ;
         RECT  192.3 344.9 192.9 345.5 ;
         LAYER metal3 ;
         RECT  105.3 194.2 106.1 195.0 ;
         LAYER metal3 ;
         RECT  219.5 365.7 220.1 366.3 ;
         LAYER metal3 ;
         RECT  2.4 302.4 78.0 303.6 ;
         LAYER metal3 ;
         RECT  185.5 313.3 186.1 313.9 ;
         LAYER metal3 ;
         RECT  2.4 38.4 42.0 39.6 ;
         LAYER metal3 ;
         RECT  2.4 345.6 226.8 346.8 ;
         LAYER metal3 ;
         RECT  15.2 247.8 16.0 248.6 ;
         LAYER metal3 ;
         RECT  2.4 336.0 226.8 337.2 ;
         LAYER metal3 ;
         RECT  205.9 303.3 206.5 303.9 ;
         LAYER metal3 ;
         RECT  205.9 354.9 206.5 355.5 ;
         LAYER metal3 ;
         RECT  212.7 324.1 213.3 324.7 ;
         LAYER metal3 ;
         RECT  205.9 344.9 206.5 345.5 ;
         LAYER metal3 ;
         RECT  185.5 271.7 186.1 272.3 ;
         LAYER metal4 ;
         RECT  156.0 0.0 157.2 370.8 ;
         LAYER metal3 ;
         RECT  199.1 292.5 199.7 293.1 ;
         LAYER metal3 ;
         RECT  2.4 48.0 226.8 49.2 ;
         LAYER metal3 ;
         RECT  192.2 209.2 193.0 210.0 ;
         LAYER metal3 ;
         RECT  24.0 216.0 85.2 217.2 ;
         LAYER metal3 ;
         RECT  75.3 292.4 76.1 293.2 ;
         LAYER metal4 ;
         RECT  223.2 0.0 224.4 370.8 ;
         LAYER metal3 ;
         RECT  79.2 350.4 140.4 351.6 ;
         LAYER metal3 ;
         RECT  187.2 110.4 226.8 111.6 ;
         LAYER metal3 ;
         RECT  219.5 178.5 220.1 179.1 ;
         LAYER metal3 ;
         RECT  192.2 199.2 193.0 200.0 ;
         LAYER metal3 ;
         RECT  185.5 261.7 186.1 262.3 ;
         LAYER metal3 ;
         RECT  177.6 268.8 226.8 270.0 ;
         LAYER metal3 ;
         RECT  2.4 62.4 80.4 63.6 ;
         LAYER metal3 ;
         RECT  192.2 344.8 193.0 345.6 ;
         LAYER metal3 ;
         RECT  196.3 47.6 197.1 48.4 ;
         LAYER metal3 ;
         RECT  2.4 148.8 226.8 150.0 ;
         LAYER metal4 ;
         RECT  84.0 0.0 85.2 370.8 ;
         LAYER metal4 ;
         RECT  74.4 0.0 75.6 370.8 ;
         LAYER metal3 ;
         RECT  122.7 256.6 123.5 257.4 ;
         LAYER metal3 ;
         RECT  2.4 292.8 226.8 294.0 ;
         LAYER metal3 ;
         RECT  2.4 249.6 226.8 250.8 ;
         LAYER metal3 ;
         RECT  185.5 250.9 186.1 251.5 ;
         LAYER metal4 ;
         RECT  160.8 0.0 162.0 370.8 ;
         LAYER metal3 ;
         RECT  212.7 271.7 213.3 272.3 ;
         LAYER metal3 ;
         RECT  219.5 313.3 220.1 313.9 ;
         LAYER metal3 ;
         RECT  205.9 313.3 206.5 313.9 ;
         LAYER metal3 ;
         RECT  2.4 41.8 3.2 42.6 ;
         LAYER metal3 ;
         RECT  212.7 230.1 213.3 230.7 ;
         LAYER metal3 ;
         RECT  8.8 185.4 9.6 186.2 ;
         LAYER metal3 ;
         RECT  199.0 250.8 199.8 251.6 ;
         LAYER metal3 ;
         RECT  93.6 302.4 226.8 303.6 ;
         LAYER metal3 ;
         RECT  219.5 354.9 220.1 355.5 ;
         LAYER metal4 ;
         RECT  204.0 0.0 205.2 370.8 ;
         LAYER metal3 ;
         RECT  208.7 106.9 209.3 107.5 ;
         LAYER metal3 ;
         RECT  173.1 277.4 173.9 278.2 ;
         LAYER metal3 ;
         RECT  96.0 321.6 226.8 322.8 ;
         LAYER metal3 ;
         RECT  192.3 199.3 192.9 199.9 ;
         LAYER metal3 ;
         RECT  192.3 271.7 192.9 272.3 ;
         LAYER metal3 ;
         RECT  33.6 230.4 226.8 231.6 ;
         LAYER metal3 ;
         RECT  219.5 209.3 220.1 209.9 ;
         LAYER metal3 ;
         RECT  2.4 144.0 226.8 145.2 ;
         LAYER metal3 ;
         RECT  192.2 271.6 193.0 272.4 ;
         LAYER metal3 ;
         RECT  212.7 365.7 213.3 366.3 ;
         LAYER metal3 ;
         RECT  173.1 319.0 173.9 319.8 ;
         LAYER metal3 ;
         RECT  2.4 273.6 226.8 274.8 ;
         LAYER metal3 ;
         RECT  2.4 240.0 226.8 241.2 ;
         LAYER metal3 ;
         RECT  146.4 278.4 226.8 279.6 ;
         LAYER metal4 ;
         RECT  122.4 0.0 123.6 370.8 ;
         LAYER metal3 ;
         RECT  145.7 319.0 146.5 319.8 ;
         LAYER metal3 ;
         RECT  219.5 303.3 220.1 303.9 ;
         LAYER metal3 ;
         RECT  2.4 331.2 140.4 332.4 ;
         LAYER metal3 ;
         RECT  205.9 178.5 206.5 179.1 ;
         LAYER metal3 ;
         RECT  122.7 215.0 123.5 215.8 ;
         LAYER metal3 ;
         RECT  2.4 364.8 226.8 366.0 ;
         LAYER metal3 ;
         RECT  122.7 277.4 123.5 278.2 ;
         LAYER metal4 ;
         RECT  40.8 0.0 42.0 370.8 ;
         LAYER metal3 ;
         RECT  219.5 230.1 220.1 230.7 ;
         LAYER metal3 ;
         RECT  199.0 354.8 199.8 355.6 ;
         LAYER metal3 ;
         RECT  192.3 250.9 192.9 251.5 ;
         LAYER metal3 ;
         RECT  205.9 261.7 206.5 262.3 ;
         LAYER metal4 ;
         RECT  184.8 0.0 186.0 370.8 ;
         LAYER metal3 ;
         RECT  199.1 220.1 199.7 220.7 ;
         LAYER metal3 ;
         RECT  199.1 250.9 199.7 251.5 ;
         LAYER metal4 ;
         RECT  55.2 0.0 56.4 370.8 ;
         LAYER metal3 ;
         RECT  145.7 360.6 146.5 361.4 ;
         LAYER metal3 ;
         RECT  192.3 334.1 192.9 334.7 ;
         LAYER metal4 ;
         RECT  98.4 0.0 99.6 370.8 ;
         LAYER metal4 ;
         RECT  88.8 0.0 90.0 370.8 ;
         LAYER metal3 ;
         RECT  76.8 4.8 226.8 6.0 ;
         LAYER metal3 ;
         RECT  185.5 303.3 186.1 303.9 ;
         LAYER metal3 ;
         RECT  173.1 215.0 173.9 215.8 ;
         LAYER metal4 ;
         RECT  45.6 0.0 46.8 370.8 ;
         LAYER metal3 ;
         RECT  205.9 282.5 206.5 283.1 ;
         LAYER metal4 ;
         RECT  12.0 0.0 13.2 370.8 ;
         LAYER metal3 ;
         RECT  199.1 313.3 199.7 313.9 ;
         LAYER metal3 ;
         RECT  84.8 121.8 85.6 122.6 ;
         LAYER metal4 ;
         RECT  50.4 0.0 51.6 370.8 ;
         LAYER metal3 ;
         RECT  205.9 334.1 206.5 334.7 ;
         LAYER metal3 ;
         RECT  192.2 240.8 193.0 241.6 ;
         LAYER metal3 ;
         RECT  205.9 146.1 206.5 146.7 ;
         LAYER metal3 ;
         RECT  212.7 178.5 213.3 179.1 ;
         LAYER metal4 ;
         RECT  213.6 0.0 214.8 370.8 ;
         LAYER metal3 ;
         RECT  2.4 355.2 226.8 356.4 ;
         LAYER metal3 ;
         RECT  212.7 303.3 213.3 303.9 ;
         LAYER metal3 ;
         RECT  145.7 256.6 146.5 257.4 ;
         LAYER metal3 ;
         RECT  212.7 282.5 213.3 283.1 ;
         LAYER metal3 ;
         RECT  145.7 298.2 146.5 299.0 ;
         LAYER metal3 ;
         RECT  199.1 230.1 199.7 230.7 ;
         LAYER metal3 ;
         RECT  199.1 261.7 199.7 262.3 ;
         LAYER metal3 ;
         RECT  185.5 209.3 186.1 209.9 ;
         LAYER metal3 ;
         RECT  2.4 153.6 82.8 154.8 ;
         LAYER metal3 ;
         RECT  21.6 206.2 22.4 207.0 ;
         LAYER metal3 ;
         RECT  2.4 67.2 193.2 68.4 ;
         LAYER metal3 ;
         RECT  192.3 324.1 192.9 324.7 ;
         LAYER metal3 ;
         RECT  2.4 124.8 226.8 126.0 ;
         LAYER metal3 ;
         RECT  192.3 209.3 192.9 209.9 ;
         LAYER metal3 ;
         RECT  205.9 292.5 206.5 293.1 ;
         LAYER metal3 ;
         RECT  33.6 220.8 226.8 222.0 ;
         LAYER metal3 ;
         RECT  84.8 1.8 85.6 2.6 ;
         LAYER metal3 ;
         RECT  15.2 164.6 16.0 165.4 ;
         LAYER metal3 ;
         RECT  203.3 87.9 203.9 88.5 ;
         LAYER metal3 ;
         RECT  84.8 161.8 85.6 162.6 ;
         LAYER metal3 ;
         RECT  33.6 201.6 226.8 202.8 ;
         LAYER metal3 ;
         RECT  199.1 188.5 199.7 189.1 ;
         LAYER metal3 ;
         RECT  2.4 297.6 61.2 298.8 ;
         LAYER metal3 ;
         RECT  199.0 261.6 199.8 262.4 ;
         LAYER metal3 ;
         RECT  199.1 199.3 199.7 199.9 ;
         LAYER metal3 ;
         RECT  192.3 354.9 192.9 355.5 ;
         LAYER metal3 ;
         RECT  2.4 268.8 99.6 270.0 ;
         LAYER metal3 ;
         RECT  2.4 81.6 198.0 82.8 ;
         LAYER metal3 ;
         RECT  2.4 86.4 226.8 87.6 ;
         LAYER metal3 ;
         RECT  210.1 87.9 210.7 88.5 ;
         LAYER metal4 ;
         RECT  132.0 0.0 133.2 370.8 ;
         LAYER metal3 ;
         RECT  2.4 326.4 226.8 327.6 ;
         LAYER metal3 ;
         RECT  177.6 206.4 226.8 207.6 ;
         LAYER metal3 ;
         RECT  145.7 339.8 146.5 340.6 ;
         LAYER metal3 ;
         RECT  84.8 41.8 85.6 42.6 ;
         LAYER metal3 ;
         RECT  199.0 188.4 199.8 189.2 ;
         LAYER metal3 ;
         RECT  2.4 4.8 39.6 6.0 ;
         LAYER metal3 ;
         RECT  2.4 115.2 226.8 116.4 ;
         LAYER metal4 ;
         RECT  189.6 0.0 190.8 370.8 ;
         LAYER metal3 ;
         RECT  185.5 292.5 186.1 293.1 ;
         LAYER metal3 ;
         RECT  219.5 261.7 220.1 262.3 ;
         LAYER metal3 ;
         RECT  199.2 168.0 226.8 169.2 ;
         LAYER metal3 ;
         RECT  185.5 230.1 186.1 230.7 ;
         LAYER metal3 ;
         RECT  185.5 354.9 186.1 355.5 ;
         LAYER metal3 ;
         RECT  2.4 52.8 82.8 54.0 ;
         LAYER metal3 ;
         RECT  60.0 38.4 226.8 39.6 ;
         LAYER metal3 ;
         RECT  212.7 313.3 213.3 313.9 ;
         LAYER metal3 ;
         RECT  192.2 365.6 193.0 366.4 ;
         LAYER metal3 ;
         RECT  185.5 282.5 186.1 283.1 ;
         LAYER metal3 ;
         RECT  199.1 354.9 199.7 355.5 ;
         LAYER metal3 ;
         RECT  2.4 350.4 70.8 351.6 ;
         LAYER metal3 ;
         RECT  192.2 178.4 193.0 179.2 ;
         LAYER metal3 ;
         RECT  199.1 303.3 199.7 303.9 ;
         LAYER metal3 ;
         RECT  2.4 120.0 226.8 121.2 ;
         LAYER metal3 ;
         RECT  2.4 225.6 99.6 226.8 ;
         LAYER metal4 ;
         RECT  175.2 0.0 176.4 370.8 ;
         LAYER metal3 ;
         RECT  2.4 0.0 226.8 1.2 ;
         LAYER metal3 ;
         RECT  173.1 339.8 173.9 340.6 ;
         LAYER metal3 ;
         RECT  2.4 110.4 82.8 111.6 ;
         LAYER metal3 ;
         RECT  199.0 344.8 199.8 345.6 ;
         LAYER metal3 ;
         RECT  199.0 303.2 199.8 304.0 ;
         LAYER metal3 ;
         RECT  192.3 313.3 192.9 313.9 ;
         LAYER metal3 ;
         RECT  199.0 209.2 199.8 210.0 ;
         LAYER metal3 ;
         RECT  199.1 334.1 199.7 334.7 ;
         LAYER metal3 ;
         RECT  192.2 313.2 193.0 314.0 ;
         LAYER metal4 ;
         RECT  117.6 0.0 118.8 370.8 ;
         LAYER metal3 ;
         RECT  199.1 344.9 199.7 345.5 ;
         LAYER metal3 ;
         RECT  103.2 259.2 226.8 260.4 ;
         LAYER metal3 ;
         RECT  192.3 282.5 192.9 283.1 ;
         LAYER metal3 ;
         RECT  199.0 334.0 199.8 334.8 ;
         LAYER metal3 ;
         RECT  2.4 360.0 226.8 361.2 ;
         LAYER metal4 ;
         RECT  36.0 0.0 37.2 370.8 ;
         LAYER metal3 ;
         RECT  2.4 244.8 99.6 246.0 ;
         LAYER metal3 ;
         RECT  2.4 139.2 226.8 140.4 ;
         LAYER metal3 ;
         RECT  212.7 199.3 213.3 199.9 ;
         LAYER metal3 ;
         RECT  15.2 185.4 16.0 186.2 ;
         LAYER metal3 ;
         RECT  205.9 324.1 206.5 324.7 ;
         LAYER metal3 ;
         RECT  24.0 196.8 226.8 198.0 ;
         LAYER metal3 ;
         RECT  184.8 153.6 226.8 154.8 ;
         LAYER metal3 ;
         RECT  21.6 235.2 121.2 236.4 ;
         LAYER metal3 ;
         RECT  205.9 230.1 206.5 230.7 ;
         LAYER metal4 ;
         RECT  218.4 0.0 219.6 370.8 ;
         LAYER metal3 ;
         RECT  2.4 321.6 78.0 322.8 ;
         LAYER metal3 ;
         RECT  185.5 199.3 186.1 199.9 ;
         LAYER metal3 ;
         RECT  192.2 220.0 193.0 220.8 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  86.6 10.9 88.0 11.5 ;
      RECT  202.8 70.5 205.0 71.1 ;
      RECT  209.6 71.9 226.8 72.5 ;
      RECT  183.4 199.3 184.0 199.9 ;
      RECT  183.4 196.5 184.0 197.1 ;
      RECT  177.3 199.3 183.7 199.9 ;
      RECT  183.4 196.8 184.0 199.6 ;
      RECT  183.7 196.5 185.8 197.1 ;
      RECT  183.4 210.1 184.0 210.7 ;
      RECT  183.4 212.1 184.0 212.7 ;
      RECT  177.3 210.1 183.7 210.7 ;
      RECT  183.4 210.4 184.0 212.4 ;
      RECT  183.7 212.1 185.8 212.7 ;
      RECT  183.4 220.1 184.0 220.7 ;
      RECT  183.4 217.3 184.0 217.9 ;
      RECT  177.3 220.1 183.7 220.7 ;
      RECT  183.4 217.6 184.0 220.4 ;
      RECT  183.7 217.3 185.8 217.9 ;
      RECT  183.4 230.9 184.0 231.5 ;
      RECT  183.4 232.9 184.0 233.5 ;
      RECT  177.3 230.9 183.7 231.5 ;
      RECT  183.4 231.2 184.0 233.2 ;
      RECT  183.7 232.9 185.8 233.5 ;
      RECT  183.4 240.9 184.0 241.5 ;
      RECT  183.4 238.1 184.0 238.7 ;
      RECT  177.3 240.9 183.7 241.5 ;
      RECT  183.4 238.4 184.0 241.2 ;
      RECT  183.7 238.1 185.8 238.7 ;
      RECT  183.4 251.7 184.0 252.3 ;
      RECT  183.4 253.7 184.0 254.3 ;
      RECT  177.3 251.7 183.7 252.3 ;
      RECT  183.4 252.0 184.0 254.0 ;
      RECT  183.7 253.7 185.8 254.3 ;
      RECT  183.4 261.7 184.0 262.3 ;
      RECT  183.4 258.9 184.0 259.5 ;
      RECT  177.3 261.7 183.7 262.3 ;
      RECT  183.4 259.2 184.0 262.0 ;
      RECT  183.7 258.9 185.8 259.5 ;
      RECT  183.4 272.5 184.0 273.1 ;
      RECT  183.4 274.5 184.0 275.1 ;
      RECT  177.3 272.5 183.7 273.1 ;
      RECT  183.4 272.8 184.0 274.8 ;
      RECT  183.7 274.5 185.8 275.1 ;
      RECT  183.4 282.5 184.0 283.1 ;
      RECT  183.4 279.7 184.0 280.3 ;
      RECT  177.3 282.5 183.7 283.1 ;
      RECT  183.4 280.0 184.0 282.8 ;
      RECT  183.7 279.7 185.8 280.3 ;
      RECT  183.4 293.3 184.0 293.9 ;
      RECT  183.4 295.3 184.0 295.9 ;
      RECT  177.3 293.3 183.7 293.9 ;
      RECT  183.4 293.6 184.0 295.6 ;
      RECT  183.7 295.3 185.8 295.9 ;
      RECT  183.4 303.3 184.0 303.9 ;
      RECT  183.4 300.5 184.0 301.1 ;
      RECT  177.3 303.3 183.7 303.9 ;
      RECT  183.4 300.8 184.0 303.6 ;
      RECT  183.7 300.5 185.8 301.1 ;
      RECT  183.4 314.1 184.0 314.7 ;
      RECT  183.4 316.1 184.0 316.7 ;
      RECT  177.3 314.1 183.7 314.7 ;
      RECT  183.4 314.4 184.0 316.4 ;
      RECT  183.7 316.1 185.8 316.7 ;
      RECT  183.4 324.1 184.0 324.7 ;
      RECT  183.4 321.3 184.0 321.9 ;
      RECT  177.3 324.1 183.7 324.7 ;
      RECT  183.4 321.6 184.0 324.4 ;
      RECT  183.7 321.3 185.8 321.9 ;
      RECT  183.4 334.9 184.0 335.5 ;
      RECT  183.4 336.9 184.0 337.5 ;
      RECT  177.3 334.9 183.7 335.5 ;
      RECT  183.4 335.2 184.0 337.2 ;
      RECT  183.7 336.9 185.8 337.5 ;
      RECT  183.4 344.9 184.0 345.5 ;
      RECT  183.4 342.1 184.0 342.7 ;
      RECT  177.3 344.9 183.7 345.5 ;
      RECT  183.4 342.4 184.0 345.2 ;
      RECT  183.7 342.1 185.8 342.7 ;
      RECT  183.4 355.7 184.0 356.3 ;
      RECT  183.4 357.7 184.0 358.3 ;
      RECT  177.3 355.7 183.7 356.3 ;
      RECT  183.4 356.0 184.0 358.0 ;
      RECT  183.7 357.7 185.8 358.3 ;
      RECT  181.9 159.8 192.6 160.4 ;
      RECT  183.3 191.3 185.8 191.9 ;
      RECT  179.1 79.8 199.4 80.4 ;
      RECT  180.5 149.6 199.4 150.2 ;
      RECT  161.8 185.9 183.3 186.5 ;
      RECT  201.4 198.2 202.4 199.0 ;
      RECT  203.8 202.6 204.8 203.4 ;
      RECT  204.0 199.0 204.8 199.4 ;
      RECT  202.8 197.2 203.6 197.4 ;
      RECT  205.8 197.8 206.6 202.0 ;
      RECT  201.6 201.2 203.2 202.0 ;
      RECT  204.0 198.2 205.0 199.0 ;
      RECT  199.0 204.2 206.6 205.0 ;
      RECT  199.0 202.6 199.8 204.2 ;
      RECT  201.6 202.6 202.6 203.4 ;
      RECT  201.6 202.0 202.4 202.6 ;
      RECT  204.0 200.2 204.8 202.6 ;
      RECT  203.6 199.4 204.8 200.2 ;
      RECT  199.0 196.4 206.6 197.2 ;
      RECT  199.0 197.8 199.8 202.0 ;
      RECT  201.6 199.0 202.4 201.2 ;
      RECT  203.4 195.0 205.0 195.8 ;
      RECT  205.8 202.6 206.6 204.2 ;
      RECT  200.6 195.0 202.2 195.8 ;
      RECT  201.4 211.0 202.4 210.2 ;
      RECT  203.8 206.6 204.8 205.8 ;
      RECT  204.0 210.2 204.8 209.8 ;
      RECT  202.8 212.0 203.6 211.8 ;
      RECT  205.8 211.4 206.6 207.2 ;
      RECT  201.6 208.0 203.2 207.2 ;
      RECT  204.0 211.0 205.0 210.2 ;
      RECT  199.0 205.0 206.6 204.2 ;
      RECT  199.0 206.6 199.8 205.0 ;
      RECT  201.6 206.6 202.6 205.8 ;
      RECT  201.6 207.2 202.4 206.6 ;
      RECT  204.0 209.0 204.8 206.6 ;
      RECT  203.6 209.8 204.8 209.0 ;
      RECT  199.0 212.8 206.6 212.0 ;
      RECT  199.0 211.4 199.8 207.2 ;
      RECT  201.6 210.2 202.4 208.0 ;
      RECT  203.4 214.2 205.0 213.4 ;
      RECT  205.8 206.6 206.6 205.0 ;
      RECT  200.6 214.2 202.2 213.4 ;
      RECT  201.4 219.0 202.4 219.8 ;
      RECT  203.8 223.4 204.8 224.2 ;
      RECT  204.0 219.8 204.8 220.2 ;
      RECT  202.8 218.0 203.6 218.2 ;
      RECT  205.8 218.6 206.6 222.8 ;
      RECT  201.6 222.0 203.2 222.8 ;
      RECT  204.0 219.0 205.0 219.8 ;
      RECT  199.0 225.0 206.6 225.8 ;
      RECT  199.0 223.4 199.8 225.0 ;
      RECT  201.6 223.4 202.6 224.2 ;
      RECT  201.6 222.8 202.4 223.4 ;
      RECT  204.0 221.0 204.8 223.4 ;
      RECT  203.6 220.2 204.8 221.0 ;
      RECT  199.0 217.2 206.6 218.0 ;
      RECT  199.0 218.6 199.8 222.8 ;
      RECT  201.6 219.8 202.4 222.0 ;
      RECT  203.4 215.8 205.0 216.6 ;
      RECT  205.8 223.4 206.6 225.0 ;
      RECT  200.6 215.8 202.2 216.6 ;
      RECT  201.4 231.8 202.4 231.0 ;
      RECT  203.8 227.4 204.8 226.6 ;
      RECT  204.0 231.0 204.8 230.6 ;
      RECT  202.8 232.8 203.6 232.6 ;
      RECT  205.8 232.2 206.6 228.0 ;
      RECT  201.6 228.8 203.2 228.0 ;
      RECT  204.0 231.8 205.0 231.0 ;
      RECT  199.0 225.8 206.6 225.0 ;
      RECT  199.0 227.4 199.8 225.8 ;
      RECT  201.6 227.4 202.6 226.6 ;
      RECT  201.6 228.0 202.4 227.4 ;
      RECT  204.0 229.8 204.8 227.4 ;
      RECT  203.6 230.6 204.8 229.8 ;
      RECT  199.0 233.6 206.6 232.8 ;
      RECT  199.0 232.2 199.8 228.0 ;
      RECT  201.6 231.0 202.4 228.8 ;
      RECT  203.4 235.0 205.0 234.2 ;
      RECT  205.8 227.4 206.6 225.8 ;
      RECT  200.6 235.0 202.2 234.2 ;
      RECT  201.4 239.8 202.4 240.6 ;
      RECT  203.8 244.2 204.8 245.0 ;
      RECT  204.0 240.6 204.8 241.0 ;
      RECT  202.8 238.8 203.6 239.0 ;
      RECT  205.8 239.4 206.6 243.6 ;
      RECT  201.6 242.8 203.2 243.6 ;
      RECT  204.0 239.8 205.0 240.6 ;
      RECT  199.0 245.8 206.6 246.6 ;
      RECT  199.0 244.2 199.8 245.8 ;
      RECT  201.6 244.2 202.6 245.0 ;
      RECT  201.6 243.6 202.4 244.2 ;
      RECT  204.0 241.8 204.8 244.2 ;
      RECT  203.6 241.0 204.8 241.8 ;
      RECT  199.0 238.0 206.6 238.8 ;
      RECT  199.0 239.4 199.8 243.6 ;
      RECT  201.6 240.6 202.4 242.8 ;
      RECT  203.4 236.6 205.0 237.4 ;
      RECT  205.8 244.2 206.6 245.8 ;
      RECT  200.6 236.6 202.2 237.4 ;
      RECT  201.4 252.6 202.4 251.8 ;
      RECT  203.8 248.2 204.8 247.4 ;
      RECT  204.0 251.8 204.8 251.4 ;
      RECT  202.8 253.6 203.6 253.4 ;
      RECT  205.8 253.0 206.6 248.8 ;
      RECT  201.6 249.6 203.2 248.8 ;
      RECT  204.0 252.6 205.0 251.8 ;
      RECT  199.0 246.6 206.6 245.8 ;
      RECT  199.0 248.2 199.8 246.6 ;
      RECT  201.6 248.2 202.6 247.4 ;
      RECT  201.6 248.8 202.4 248.2 ;
      RECT  204.0 250.6 204.8 248.2 ;
      RECT  203.6 251.4 204.8 250.6 ;
      RECT  199.0 254.4 206.6 253.6 ;
      RECT  199.0 253.0 199.8 248.8 ;
      RECT  201.6 251.8 202.4 249.6 ;
      RECT  203.4 255.8 205.0 255.0 ;
      RECT  205.8 248.2 206.6 246.6 ;
      RECT  200.6 255.8 202.2 255.0 ;
      RECT  201.4 260.6 202.4 261.4 ;
      RECT  203.8 265.0 204.8 265.8 ;
      RECT  204.0 261.4 204.8 261.8 ;
      RECT  202.8 259.6 203.6 259.8 ;
      RECT  205.8 260.2 206.6 264.4 ;
      RECT  201.6 263.6 203.2 264.4 ;
      RECT  204.0 260.6 205.0 261.4 ;
      RECT  199.0 266.6 206.6 267.4 ;
      RECT  199.0 265.0 199.8 266.6 ;
      RECT  201.6 265.0 202.6 265.8 ;
      RECT  201.6 264.4 202.4 265.0 ;
      RECT  204.0 262.6 204.8 265.0 ;
      RECT  203.6 261.8 204.8 262.6 ;
      RECT  199.0 258.8 206.6 259.6 ;
      RECT  199.0 260.2 199.8 264.4 ;
      RECT  201.6 261.4 202.4 263.6 ;
      RECT  203.4 257.4 205.0 258.2 ;
      RECT  205.8 265.0 206.6 266.6 ;
      RECT  200.6 257.4 202.2 258.2 ;
      RECT  201.4 273.4 202.4 272.6 ;
      RECT  203.8 269.0 204.8 268.2 ;
      RECT  204.0 272.6 204.8 272.2 ;
      RECT  202.8 274.4 203.6 274.2 ;
      RECT  205.8 273.8 206.6 269.6 ;
      RECT  201.6 270.4 203.2 269.6 ;
      RECT  204.0 273.4 205.0 272.6 ;
      RECT  199.0 267.4 206.6 266.6 ;
      RECT  199.0 269.0 199.8 267.4 ;
      RECT  201.6 269.0 202.6 268.2 ;
      RECT  201.6 269.6 202.4 269.0 ;
      RECT  204.0 271.4 204.8 269.0 ;
      RECT  203.6 272.2 204.8 271.4 ;
      RECT  199.0 275.2 206.6 274.4 ;
      RECT  199.0 273.8 199.8 269.6 ;
      RECT  201.6 272.6 202.4 270.4 ;
      RECT  203.4 276.6 205.0 275.8 ;
      RECT  205.8 269.0 206.6 267.4 ;
      RECT  200.6 276.6 202.2 275.8 ;
      RECT  201.4 281.4 202.4 282.2 ;
      RECT  203.8 285.8 204.8 286.6 ;
      RECT  204.0 282.2 204.8 282.6 ;
      RECT  202.8 280.4 203.6 280.6 ;
      RECT  205.8 281.0 206.6 285.2 ;
      RECT  201.6 284.4 203.2 285.2 ;
      RECT  204.0 281.4 205.0 282.2 ;
      RECT  199.0 287.4 206.6 288.2 ;
      RECT  199.0 285.8 199.8 287.4 ;
      RECT  201.6 285.8 202.6 286.6 ;
      RECT  201.6 285.2 202.4 285.8 ;
      RECT  204.0 283.4 204.8 285.8 ;
      RECT  203.6 282.6 204.8 283.4 ;
      RECT  199.0 279.6 206.6 280.4 ;
      RECT  199.0 281.0 199.8 285.2 ;
      RECT  201.6 282.2 202.4 284.4 ;
      RECT  203.4 278.2 205.0 279.0 ;
      RECT  205.8 285.8 206.6 287.4 ;
      RECT  200.6 278.2 202.2 279.0 ;
      RECT  201.4 294.2 202.4 293.4 ;
      RECT  203.8 289.8 204.8 289.0 ;
      RECT  204.0 293.4 204.8 293.0 ;
      RECT  202.8 295.2 203.6 295.0 ;
      RECT  205.8 294.6 206.6 290.4 ;
      RECT  201.6 291.2 203.2 290.4 ;
      RECT  204.0 294.2 205.0 293.4 ;
      RECT  199.0 288.2 206.6 287.4 ;
      RECT  199.0 289.8 199.8 288.2 ;
      RECT  201.6 289.8 202.6 289.0 ;
      RECT  201.6 290.4 202.4 289.8 ;
      RECT  204.0 292.2 204.8 289.8 ;
      RECT  203.6 293.0 204.8 292.2 ;
      RECT  199.0 296.0 206.6 295.2 ;
      RECT  199.0 294.6 199.8 290.4 ;
      RECT  201.6 293.4 202.4 291.2 ;
      RECT  203.4 297.4 205.0 296.6 ;
      RECT  205.8 289.8 206.6 288.2 ;
      RECT  200.6 297.4 202.2 296.6 ;
      RECT  201.4 302.2 202.4 303.0 ;
      RECT  203.8 306.6 204.8 307.4 ;
      RECT  204.0 303.0 204.8 303.4 ;
      RECT  202.8 301.2 203.6 301.4 ;
      RECT  205.8 301.8 206.6 306.0 ;
      RECT  201.6 305.2 203.2 306.0 ;
      RECT  204.0 302.2 205.0 303.0 ;
      RECT  199.0 308.2 206.6 309.0 ;
      RECT  199.0 306.6 199.8 308.2 ;
      RECT  201.6 306.6 202.6 307.4 ;
      RECT  201.6 306.0 202.4 306.6 ;
      RECT  204.0 304.2 204.8 306.6 ;
      RECT  203.6 303.4 204.8 304.2 ;
      RECT  199.0 300.4 206.6 301.2 ;
      RECT  199.0 301.8 199.8 306.0 ;
      RECT  201.6 303.0 202.4 305.2 ;
      RECT  203.4 299.0 205.0 299.8 ;
      RECT  205.8 306.6 206.6 308.2 ;
      RECT  200.6 299.0 202.2 299.8 ;
      RECT  201.4 315.0 202.4 314.2 ;
      RECT  203.8 310.6 204.8 309.8 ;
      RECT  204.0 314.2 204.8 313.8 ;
      RECT  202.8 316.0 203.6 315.8 ;
      RECT  205.8 315.4 206.6 311.2 ;
      RECT  201.6 312.0 203.2 311.2 ;
      RECT  204.0 315.0 205.0 314.2 ;
      RECT  199.0 309.0 206.6 308.2 ;
      RECT  199.0 310.6 199.8 309.0 ;
      RECT  201.6 310.6 202.6 309.8 ;
      RECT  201.6 311.2 202.4 310.6 ;
      RECT  204.0 313.0 204.8 310.6 ;
      RECT  203.6 313.8 204.8 313.0 ;
      RECT  199.0 316.8 206.6 316.0 ;
      RECT  199.0 315.4 199.8 311.2 ;
      RECT  201.6 314.2 202.4 312.0 ;
      RECT  203.4 318.2 205.0 317.4 ;
      RECT  205.8 310.6 206.6 309.0 ;
      RECT  200.6 318.2 202.2 317.4 ;
      RECT  201.4 323.0 202.4 323.8 ;
      RECT  203.8 327.4 204.8 328.2 ;
      RECT  204.0 323.8 204.8 324.2 ;
      RECT  202.8 322.0 203.6 322.2 ;
      RECT  205.8 322.6 206.6 326.8 ;
      RECT  201.6 326.0 203.2 326.8 ;
      RECT  204.0 323.0 205.0 323.8 ;
      RECT  199.0 329.0 206.6 329.8 ;
      RECT  199.0 327.4 199.8 329.0 ;
      RECT  201.6 327.4 202.6 328.2 ;
      RECT  201.6 326.8 202.4 327.4 ;
      RECT  204.0 325.0 204.8 327.4 ;
      RECT  203.6 324.2 204.8 325.0 ;
      RECT  199.0 321.2 206.6 322.0 ;
      RECT  199.0 322.6 199.8 326.8 ;
      RECT  201.6 323.8 202.4 326.0 ;
      RECT  203.4 319.8 205.0 320.6 ;
      RECT  205.8 327.4 206.6 329.0 ;
      RECT  200.6 319.8 202.2 320.6 ;
      RECT  201.4 335.8 202.4 335.0 ;
      RECT  203.8 331.4 204.8 330.6 ;
      RECT  204.0 335.0 204.8 334.6 ;
      RECT  202.8 336.8 203.6 336.6 ;
      RECT  205.8 336.2 206.6 332.0 ;
      RECT  201.6 332.8 203.2 332.0 ;
      RECT  204.0 335.8 205.0 335.0 ;
      RECT  199.0 329.8 206.6 329.0 ;
      RECT  199.0 331.4 199.8 329.8 ;
      RECT  201.6 331.4 202.6 330.6 ;
      RECT  201.6 332.0 202.4 331.4 ;
      RECT  204.0 333.8 204.8 331.4 ;
      RECT  203.6 334.6 204.8 333.8 ;
      RECT  199.0 337.6 206.6 336.8 ;
      RECT  199.0 336.2 199.8 332.0 ;
      RECT  201.6 335.0 202.4 332.8 ;
      RECT  203.4 339.0 205.0 338.2 ;
      RECT  205.8 331.4 206.6 329.8 ;
      RECT  200.6 339.0 202.2 338.2 ;
      RECT  201.4 343.8 202.4 344.6 ;
      RECT  203.8 348.2 204.8 349.0 ;
      RECT  204.0 344.6 204.8 345.0 ;
      RECT  202.8 342.8 203.6 343.0 ;
      RECT  205.8 343.4 206.6 347.6 ;
      RECT  201.6 346.8 203.2 347.6 ;
      RECT  204.0 343.8 205.0 344.6 ;
      RECT  199.0 349.8 206.6 350.6 ;
      RECT  199.0 348.2 199.8 349.8 ;
      RECT  201.6 348.2 202.6 349.0 ;
      RECT  201.6 347.6 202.4 348.2 ;
      RECT  204.0 345.8 204.8 348.2 ;
      RECT  203.6 345.0 204.8 345.8 ;
      RECT  199.0 342.0 206.6 342.8 ;
      RECT  199.0 343.4 199.8 347.6 ;
      RECT  201.6 344.6 202.4 346.8 ;
      RECT  203.4 340.6 205.0 341.4 ;
      RECT  205.8 348.2 206.6 349.8 ;
      RECT  200.6 340.6 202.2 341.4 ;
      RECT  201.4 356.6 202.4 355.8 ;
      RECT  203.8 352.2 204.8 351.4 ;
      RECT  204.0 355.8 204.8 355.4 ;
      RECT  202.8 357.6 203.6 357.4 ;
      RECT  205.8 357.0 206.6 352.8 ;
      RECT  201.6 353.6 203.2 352.8 ;
      RECT  204.0 356.6 205.0 355.8 ;
      RECT  199.0 350.6 206.6 349.8 ;
      RECT  199.0 352.2 199.8 350.6 ;
      RECT  201.6 352.2 202.6 351.4 ;
      RECT  201.6 352.8 202.4 352.2 ;
      RECT  204.0 354.6 204.8 352.2 ;
      RECT  203.6 355.4 204.8 354.6 ;
      RECT  199.0 358.4 206.6 357.6 ;
      RECT  199.0 357.0 199.8 352.8 ;
      RECT  201.6 355.8 202.4 353.6 ;
      RECT  203.4 359.8 205.0 359.0 ;
      RECT  205.8 352.2 206.6 350.6 ;
      RECT  200.6 359.8 202.2 359.0 ;
      RECT  208.2 198.2 209.2 199.0 ;
      RECT  210.6 202.6 211.6 203.4 ;
      RECT  210.8 199.0 211.6 199.4 ;
      RECT  209.6 197.2 210.4 197.4 ;
      RECT  212.6 197.8 213.4 202.0 ;
      RECT  208.4 201.2 210.0 202.0 ;
      RECT  210.8 198.2 211.8 199.0 ;
      RECT  205.8 204.2 213.4 205.0 ;
      RECT  205.8 202.6 206.6 204.2 ;
      RECT  208.4 202.6 209.4 203.4 ;
      RECT  208.4 202.0 209.2 202.6 ;
      RECT  210.8 200.2 211.6 202.6 ;
      RECT  210.4 199.4 211.6 200.2 ;
      RECT  205.8 196.4 213.4 197.2 ;
      RECT  205.8 197.8 206.6 202.0 ;
      RECT  208.4 199.0 209.2 201.2 ;
      RECT  210.2 195.0 211.8 195.8 ;
      RECT  212.6 202.6 213.4 204.2 ;
      RECT  207.4 195.0 209.0 195.8 ;
      RECT  208.2 211.0 209.2 210.2 ;
      RECT  210.6 206.6 211.6 205.8 ;
      RECT  210.8 210.2 211.6 209.8 ;
      RECT  209.6 212.0 210.4 211.8 ;
      RECT  212.6 211.4 213.4 207.2 ;
      RECT  208.4 208.0 210.0 207.2 ;
      RECT  210.8 211.0 211.8 210.2 ;
      RECT  205.8 205.0 213.4 204.2 ;
      RECT  205.8 206.6 206.6 205.0 ;
      RECT  208.4 206.6 209.4 205.8 ;
      RECT  208.4 207.2 209.2 206.6 ;
      RECT  210.8 209.0 211.6 206.6 ;
      RECT  210.4 209.8 211.6 209.0 ;
      RECT  205.8 212.8 213.4 212.0 ;
      RECT  205.8 211.4 206.6 207.2 ;
      RECT  208.4 210.2 209.2 208.0 ;
      RECT  210.2 214.2 211.8 213.4 ;
      RECT  212.6 206.6 213.4 205.0 ;
      RECT  207.4 214.2 209.0 213.4 ;
      RECT  208.2 219.0 209.2 219.8 ;
      RECT  210.6 223.4 211.6 224.2 ;
      RECT  210.8 219.8 211.6 220.2 ;
      RECT  209.6 218.0 210.4 218.2 ;
      RECT  212.6 218.6 213.4 222.8 ;
      RECT  208.4 222.0 210.0 222.8 ;
      RECT  210.8 219.0 211.8 219.8 ;
      RECT  205.8 225.0 213.4 225.8 ;
      RECT  205.8 223.4 206.6 225.0 ;
      RECT  208.4 223.4 209.4 224.2 ;
      RECT  208.4 222.8 209.2 223.4 ;
      RECT  210.8 221.0 211.6 223.4 ;
      RECT  210.4 220.2 211.6 221.0 ;
      RECT  205.8 217.2 213.4 218.0 ;
      RECT  205.8 218.6 206.6 222.8 ;
      RECT  208.4 219.8 209.2 222.0 ;
      RECT  210.2 215.8 211.8 216.6 ;
      RECT  212.6 223.4 213.4 225.0 ;
      RECT  207.4 215.8 209.0 216.6 ;
      RECT  208.2 231.8 209.2 231.0 ;
      RECT  210.6 227.4 211.6 226.6 ;
      RECT  210.8 231.0 211.6 230.6 ;
      RECT  209.6 232.8 210.4 232.6 ;
      RECT  212.6 232.2 213.4 228.0 ;
      RECT  208.4 228.8 210.0 228.0 ;
      RECT  210.8 231.8 211.8 231.0 ;
      RECT  205.8 225.8 213.4 225.0 ;
      RECT  205.8 227.4 206.6 225.8 ;
      RECT  208.4 227.4 209.4 226.6 ;
      RECT  208.4 228.0 209.2 227.4 ;
      RECT  210.8 229.8 211.6 227.4 ;
      RECT  210.4 230.6 211.6 229.8 ;
      RECT  205.8 233.6 213.4 232.8 ;
      RECT  205.8 232.2 206.6 228.0 ;
      RECT  208.4 231.0 209.2 228.8 ;
      RECT  210.2 235.0 211.8 234.2 ;
      RECT  212.6 227.4 213.4 225.8 ;
      RECT  207.4 235.0 209.0 234.2 ;
      RECT  208.2 239.8 209.2 240.6 ;
      RECT  210.6 244.2 211.6 245.0 ;
      RECT  210.8 240.6 211.6 241.0 ;
      RECT  209.6 238.8 210.4 239.0 ;
      RECT  212.6 239.4 213.4 243.6 ;
      RECT  208.4 242.8 210.0 243.6 ;
      RECT  210.8 239.8 211.8 240.6 ;
      RECT  205.8 245.8 213.4 246.6 ;
      RECT  205.8 244.2 206.6 245.8 ;
      RECT  208.4 244.2 209.4 245.0 ;
      RECT  208.4 243.6 209.2 244.2 ;
      RECT  210.8 241.8 211.6 244.2 ;
      RECT  210.4 241.0 211.6 241.8 ;
      RECT  205.8 238.0 213.4 238.8 ;
      RECT  205.8 239.4 206.6 243.6 ;
      RECT  208.4 240.6 209.2 242.8 ;
      RECT  210.2 236.6 211.8 237.4 ;
      RECT  212.6 244.2 213.4 245.8 ;
      RECT  207.4 236.6 209.0 237.4 ;
      RECT  208.2 252.6 209.2 251.8 ;
      RECT  210.6 248.2 211.6 247.4 ;
      RECT  210.8 251.8 211.6 251.4 ;
      RECT  209.6 253.6 210.4 253.4 ;
      RECT  212.6 253.0 213.4 248.8 ;
      RECT  208.4 249.6 210.0 248.8 ;
      RECT  210.8 252.6 211.8 251.8 ;
      RECT  205.8 246.6 213.4 245.8 ;
      RECT  205.8 248.2 206.6 246.6 ;
      RECT  208.4 248.2 209.4 247.4 ;
      RECT  208.4 248.8 209.2 248.2 ;
      RECT  210.8 250.6 211.6 248.2 ;
      RECT  210.4 251.4 211.6 250.6 ;
      RECT  205.8 254.4 213.4 253.6 ;
      RECT  205.8 253.0 206.6 248.8 ;
      RECT  208.4 251.8 209.2 249.6 ;
      RECT  210.2 255.8 211.8 255.0 ;
      RECT  212.6 248.2 213.4 246.6 ;
      RECT  207.4 255.8 209.0 255.0 ;
      RECT  208.2 260.6 209.2 261.4 ;
      RECT  210.6 265.0 211.6 265.8 ;
      RECT  210.8 261.4 211.6 261.8 ;
      RECT  209.6 259.6 210.4 259.8 ;
      RECT  212.6 260.2 213.4 264.4 ;
      RECT  208.4 263.6 210.0 264.4 ;
      RECT  210.8 260.6 211.8 261.4 ;
      RECT  205.8 266.6 213.4 267.4 ;
      RECT  205.8 265.0 206.6 266.6 ;
      RECT  208.4 265.0 209.4 265.8 ;
      RECT  208.4 264.4 209.2 265.0 ;
      RECT  210.8 262.6 211.6 265.0 ;
      RECT  210.4 261.8 211.6 262.6 ;
      RECT  205.8 258.8 213.4 259.6 ;
      RECT  205.8 260.2 206.6 264.4 ;
      RECT  208.4 261.4 209.2 263.6 ;
      RECT  210.2 257.4 211.8 258.2 ;
      RECT  212.6 265.0 213.4 266.6 ;
      RECT  207.4 257.4 209.0 258.2 ;
      RECT  208.2 273.4 209.2 272.6 ;
      RECT  210.6 269.0 211.6 268.2 ;
      RECT  210.8 272.6 211.6 272.2 ;
      RECT  209.6 274.4 210.4 274.2 ;
      RECT  212.6 273.8 213.4 269.6 ;
      RECT  208.4 270.4 210.0 269.6 ;
      RECT  210.8 273.4 211.8 272.6 ;
      RECT  205.8 267.4 213.4 266.6 ;
      RECT  205.8 269.0 206.6 267.4 ;
      RECT  208.4 269.0 209.4 268.2 ;
      RECT  208.4 269.6 209.2 269.0 ;
      RECT  210.8 271.4 211.6 269.0 ;
      RECT  210.4 272.2 211.6 271.4 ;
      RECT  205.8 275.2 213.4 274.4 ;
      RECT  205.8 273.8 206.6 269.6 ;
      RECT  208.4 272.6 209.2 270.4 ;
      RECT  210.2 276.6 211.8 275.8 ;
      RECT  212.6 269.0 213.4 267.4 ;
      RECT  207.4 276.6 209.0 275.8 ;
      RECT  208.2 281.4 209.2 282.2 ;
      RECT  210.6 285.8 211.6 286.6 ;
      RECT  210.8 282.2 211.6 282.6 ;
      RECT  209.6 280.4 210.4 280.6 ;
      RECT  212.6 281.0 213.4 285.2 ;
      RECT  208.4 284.4 210.0 285.2 ;
      RECT  210.8 281.4 211.8 282.2 ;
      RECT  205.8 287.4 213.4 288.2 ;
      RECT  205.8 285.8 206.6 287.4 ;
      RECT  208.4 285.8 209.4 286.6 ;
      RECT  208.4 285.2 209.2 285.8 ;
      RECT  210.8 283.4 211.6 285.8 ;
      RECT  210.4 282.6 211.6 283.4 ;
      RECT  205.8 279.6 213.4 280.4 ;
      RECT  205.8 281.0 206.6 285.2 ;
      RECT  208.4 282.2 209.2 284.4 ;
      RECT  210.2 278.2 211.8 279.0 ;
      RECT  212.6 285.8 213.4 287.4 ;
      RECT  207.4 278.2 209.0 279.0 ;
      RECT  208.2 294.2 209.2 293.4 ;
      RECT  210.6 289.8 211.6 289.0 ;
      RECT  210.8 293.4 211.6 293.0 ;
      RECT  209.6 295.2 210.4 295.0 ;
      RECT  212.6 294.6 213.4 290.4 ;
      RECT  208.4 291.2 210.0 290.4 ;
      RECT  210.8 294.2 211.8 293.4 ;
      RECT  205.8 288.2 213.4 287.4 ;
      RECT  205.8 289.8 206.6 288.2 ;
      RECT  208.4 289.8 209.4 289.0 ;
      RECT  208.4 290.4 209.2 289.8 ;
      RECT  210.8 292.2 211.6 289.8 ;
      RECT  210.4 293.0 211.6 292.2 ;
      RECT  205.8 296.0 213.4 295.2 ;
      RECT  205.8 294.6 206.6 290.4 ;
      RECT  208.4 293.4 209.2 291.2 ;
      RECT  210.2 297.4 211.8 296.6 ;
      RECT  212.6 289.8 213.4 288.2 ;
      RECT  207.4 297.4 209.0 296.6 ;
      RECT  208.2 302.2 209.2 303.0 ;
      RECT  210.6 306.6 211.6 307.4 ;
      RECT  210.8 303.0 211.6 303.4 ;
      RECT  209.6 301.2 210.4 301.4 ;
      RECT  212.6 301.8 213.4 306.0 ;
      RECT  208.4 305.2 210.0 306.0 ;
      RECT  210.8 302.2 211.8 303.0 ;
      RECT  205.8 308.2 213.4 309.0 ;
      RECT  205.8 306.6 206.6 308.2 ;
      RECT  208.4 306.6 209.4 307.4 ;
      RECT  208.4 306.0 209.2 306.6 ;
      RECT  210.8 304.2 211.6 306.6 ;
      RECT  210.4 303.4 211.6 304.2 ;
      RECT  205.8 300.4 213.4 301.2 ;
      RECT  205.8 301.8 206.6 306.0 ;
      RECT  208.4 303.0 209.2 305.2 ;
      RECT  210.2 299.0 211.8 299.8 ;
      RECT  212.6 306.6 213.4 308.2 ;
      RECT  207.4 299.0 209.0 299.8 ;
      RECT  208.2 315.0 209.2 314.2 ;
      RECT  210.6 310.6 211.6 309.8 ;
      RECT  210.8 314.2 211.6 313.8 ;
      RECT  209.6 316.0 210.4 315.8 ;
      RECT  212.6 315.4 213.4 311.2 ;
      RECT  208.4 312.0 210.0 311.2 ;
      RECT  210.8 315.0 211.8 314.2 ;
      RECT  205.8 309.0 213.4 308.2 ;
      RECT  205.8 310.6 206.6 309.0 ;
      RECT  208.4 310.6 209.4 309.8 ;
      RECT  208.4 311.2 209.2 310.6 ;
      RECT  210.8 313.0 211.6 310.6 ;
      RECT  210.4 313.8 211.6 313.0 ;
      RECT  205.8 316.8 213.4 316.0 ;
      RECT  205.8 315.4 206.6 311.2 ;
      RECT  208.4 314.2 209.2 312.0 ;
      RECT  210.2 318.2 211.8 317.4 ;
      RECT  212.6 310.6 213.4 309.0 ;
      RECT  207.4 318.2 209.0 317.4 ;
      RECT  208.2 323.0 209.2 323.8 ;
      RECT  210.6 327.4 211.6 328.2 ;
      RECT  210.8 323.8 211.6 324.2 ;
      RECT  209.6 322.0 210.4 322.2 ;
      RECT  212.6 322.6 213.4 326.8 ;
      RECT  208.4 326.0 210.0 326.8 ;
      RECT  210.8 323.0 211.8 323.8 ;
      RECT  205.8 329.0 213.4 329.8 ;
      RECT  205.8 327.4 206.6 329.0 ;
      RECT  208.4 327.4 209.4 328.2 ;
      RECT  208.4 326.8 209.2 327.4 ;
      RECT  210.8 325.0 211.6 327.4 ;
      RECT  210.4 324.2 211.6 325.0 ;
      RECT  205.8 321.2 213.4 322.0 ;
      RECT  205.8 322.6 206.6 326.8 ;
      RECT  208.4 323.8 209.2 326.0 ;
      RECT  210.2 319.8 211.8 320.6 ;
      RECT  212.6 327.4 213.4 329.0 ;
      RECT  207.4 319.8 209.0 320.6 ;
      RECT  208.2 335.8 209.2 335.0 ;
      RECT  210.6 331.4 211.6 330.6 ;
      RECT  210.8 335.0 211.6 334.6 ;
      RECT  209.6 336.8 210.4 336.6 ;
      RECT  212.6 336.2 213.4 332.0 ;
      RECT  208.4 332.8 210.0 332.0 ;
      RECT  210.8 335.8 211.8 335.0 ;
      RECT  205.8 329.8 213.4 329.0 ;
      RECT  205.8 331.4 206.6 329.8 ;
      RECT  208.4 331.4 209.4 330.6 ;
      RECT  208.4 332.0 209.2 331.4 ;
      RECT  210.8 333.8 211.6 331.4 ;
      RECT  210.4 334.6 211.6 333.8 ;
      RECT  205.8 337.6 213.4 336.8 ;
      RECT  205.8 336.2 206.6 332.0 ;
      RECT  208.4 335.0 209.2 332.8 ;
      RECT  210.2 339.0 211.8 338.2 ;
      RECT  212.6 331.4 213.4 329.8 ;
      RECT  207.4 339.0 209.0 338.2 ;
      RECT  208.2 343.8 209.2 344.6 ;
      RECT  210.6 348.2 211.6 349.0 ;
      RECT  210.8 344.6 211.6 345.0 ;
      RECT  209.6 342.8 210.4 343.0 ;
      RECT  212.6 343.4 213.4 347.6 ;
      RECT  208.4 346.8 210.0 347.6 ;
      RECT  210.8 343.8 211.8 344.6 ;
      RECT  205.8 349.8 213.4 350.6 ;
      RECT  205.8 348.2 206.6 349.8 ;
      RECT  208.4 348.2 209.4 349.0 ;
      RECT  208.4 347.6 209.2 348.2 ;
      RECT  210.8 345.8 211.6 348.2 ;
      RECT  210.4 345.0 211.6 345.8 ;
      RECT  205.8 342.0 213.4 342.8 ;
      RECT  205.8 343.4 206.6 347.6 ;
      RECT  208.4 344.6 209.2 346.8 ;
      RECT  210.2 340.6 211.8 341.4 ;
      RECT  212.6 348.2 213.4 349.8 ;
      RECT  207.4 340.6 209.0 341.4 ;
      RECT  208.2 356.6 209.2 355.8 ;
      RECT  210.6 352.2 211.6 351.4 ;
      RECT  210.8 355.8 211.6 355.4 ;
      RECT  209.6 357.6 210.4 357.4 ;
      RECT  212.6 357.0 213.4 352.8 ;
      RECT  208.4 353.6 210.0 352.8 ;
      RECT  210.8 356.6 211.8 355.8 ;
      RECT  205.8 350.6 213.4 349.8 ;
      RECT  205.8 352.2 206.6 350.6 ;
      RECT  208.4 352.2 209.4 351.4 ;
      RECT  208.4 352.8 209.2 352.2 ;
      RECT  210.8 354.6 211.6 352.2 ;
      RECT  210.4 355.4 211.6 354.6 ;
      RECT  205.8 358.4 213.4 357.6 ;
      RECT  205.8 357.0 206.6 352.8 ;
      RECT  208.4 355.8 209.2 353.6 ;
      RECT  210.2 359.8 211.8 359.0 ;
      RECT  212.6 352.2 213.4 350.6 ;
      RECT  207.4 359.8 209.0 359.0 ;
      RECT  199.4 196.4 213.0 197.2 ;
      RECT  199.4 212.0 213.0 212.8 ;
      RECT  199.4 217.2 213.0 218.0 ;
      RECT  199.4 232.8 213.0 233.6 ;
      RECT  199.4 238.0 213.0 238.8 ;
      RECT  199.4 253.6 213.0 254.4 ;
      RECT  199.4 258.8 213.0 259.6 ;
      RECT  199.4 274.4 213.0 275.2 ;
      RECT  199.4 279.6 213.0 280.4 ;
      RECT  199.4 295.2 213.0 296.0 ;
      RECT  199.4 300.4 213.0 301.2 ;
      RECT  199.4 316.0 213.0 316.8 ;
      RECT  199.4 321.2 213.0 322.0 ;
      RECT  199.4 336.8 213.0 337.6 ;
      RECT  199.4 342.0 213.0 342.8 ;
      RECT  199.4 357.6 213.0 358.4 ;
      RECT  194.6 177.4 195.6 178.2 ;
      RECT  197.0 181.8 198.0 182.6 ;
      RECT  197.2 178.2 198.0 178.6 ;
      RECT  196.0 176.4 196.8 176.6 ;
      RECT  199.0 177.0 199.8 181.2 ;
      RECT  194.8 180.4 196.4 181.2 ;
      RECT  197.2 177.4 198.2 178.2 ;
      RECT  194.6 174.2 195.4 175.0 ;
      RECT  192.2 183.4 199.8 184.2 ;
      RECT  192.2 181.8 193.0 183.4 ;
      RECT  194.8 181.8 195.8 182.6 ;
      RECT  194.8 181.2 195.6 181.8 ;
      RECT  197.2 179.4 198.0 181.8 ;
      RECT  196.8 178.6 198.0 179.4 ;
      RECT  192.2 175.6 199.8 176.4 ;
      RECT  197.4 174.2 198.2 175.0 ;
      RECT  192.2 177.0 193.0 181.2 ;
      RECT  194.8 178.2 195.6 180.4 ;
      RECT  199.0 181.8 199.8 183.4 ;
      RECT  194.6 190.2 195.6 189.4 ;
      RECT  197.0 185.8 198.0 185.0 ;
      RECT  197.2 189.4 198.0 189.0 ;
      RECT  196.0 191.2 196.8 191.0 ;
      RECT  199.0 190.6 199.8 186.4 ;
      RECT  194.8 187.2 196.4 186.4 ;
      RECT  197.0 185.0 197.8 184.2 ;
      RECT  197.2 190.2 198.2 189.4 ;
      RECT  192.2 184.2 199.8 183.4 ;
      RECT  192.2 185.8 193.0 184.2 ;
      RECT  194.8 185.8 195.8 185.0 ;
      RECT  194.8 186.4 195.6 185.8 ;
      RECT  197.2 188.2 198.0 185.8 ;
      RECT  196.8 189.0 198.0 188.2 ;
      RECT  192.2 192.0 199.8 191.2 ;
      RECT  192.2 190.6 193.0 186.4 ;
      RECT  194.8 189.4 195.6 187.2 ;
      RECT  196.6 193.4 198.2 192.6 ;
      RECT  199.0 185.8 199.8 184.2 ;
      RECT  193.8 193.4 195.4 192.6 ;
      RECT  194.6 198.2 195.6 199.0 ;
      RECT  197.0 202.6 198.0 203.4 ;
      RECT  197.2 199.0 198.0 199.4 ;
      RECT  196.0 197.2 196.8 197.4 ;
      RECT  199.0 197.8 199.8 202.0 ;
      RECT  194.8 201.2 196.4 202.0 ;
      RECT  197.0 203.4 197.8 204.2 ;
      RECT  197.2 198.2 198.2 199.0 ;
      RECT  192.2 204.2 199.8 205.0 ;
      RECT  192.2 202.6 193.0 204.2 ;
      RECT  194.8 202.6 195.8 203.4 ;
      RECT  194.8 202.0 195.6 202.6 ;
      RECT  197.2 200.2 198.0 202.6 ;
      RECT  196.8 199.4 198.0 200.2 ;
      RECT  192.2 196.4 199.8 197.2 ;
      RECT  192.2 197.8 193.0 202.0 ;
      RECT  194.8 199.0 195.6 201.2 ;
      RECT  196.6 195.0 198.2 195.8 ;
      RECT  199.0 202.6 199.8 204.2 ;
      RECT  193.8 195.0 195.4 195.8 ;
      RECT  194.6 211.0 195.6 210.2 ;
      RECT  197.0 206.6 198.0 205.8 ;
      RECT  197.2 210.2 198.0 209.8 ;
      RECT  196.0 212.0 196.8 211.8 ;
      RECT  199.0 211.4 199.8 207.2 ;
      RECT  194.8 208.0 196.4 207.2 ;
      RECT  197.0 205.8 197.8 205.0 ;
      RECT  197.2 211.0 198.2 210.2 ;
      RECT  192.2 205.0 199.8 204.2 ;
      RECT  192.2 206.6 193.0 205.0 ;
      RECT  194.8 206.6 195.8 205.8 ;
      RECT  194.8 207.2 195.6 206.6 ;
      RECT  197.2 209.0 198.0 206.6 ;
      RECT  196.8 209.8 198.0 209.0 ;
      RECT  192.2 212.8 199.8 212.0 ;
      RECT  192.2 211.4 193.0 207.2 ;
      RECT  194.8 210.2 195.6 208.0 ;
      RECT  196.6 214.2 198.2 213.4 ;
      RECT  199.0 206.6 199.8 205.0 ;
      RECT  193.8 214.2 195.4 213.4 ;
      RECT  194.6 219.0 195.6 219.8 ;
      RECT  197.0 223.4 198.0 224.2 ;
      RECT  197.2 219.8 198.0 220.2 ;
      RECT  196.0 218.0 196.8 218.2 ;
      RECT  199.0 218.6 199.8 222.8 ;
      RECT  194.8 222.0 196.4 222.8 ;
      RECT  197.0 224.2 197.8 225.0 ;
      RECT  197.2 219.0 198.2 219.8 ;
      RECT  192.2 225.0 199.8 225.8 ;
      RECT  192.2 223.4 193.0 225.0 ;
      RECT  194.8 223.4 195.8 224.2 ;
      RECT  194.8 222.8 195.6 223.4 ;
      RECT  197.2 221.0 198.0 223.4 ;
      RECT  196.8 220.2 198.0 221.0 ;
      RECT  192.2 217.2 199.8 218.0 ;
      RECT  192.2 218.6 193.0 222.8 ;
      RECT  194.8 219.8 195.6 222.0 ;
      RECT  196.6 215.8 198.2 216.6 ;
      RECT  199.0 223.4 199.8 225.0 ;
      RECT  193.8 215.8 195.4 216.6 ;
      RECT  194.6 231.8 195.6 231.0 ;
      RECT  197.0 227.4 198.0 226.6 ;
      RECT  197.2 231.0 198.0 230.6 ;
      RECT  196.0 232.8 196.8 232.6 ;
      RECT  199.0 232.2 199.8 228.0 ;
      RECT  194.8 228.8 196.4 228.0 ;
      RECT  197.0 226.6 197.8 225.8 ;
      RECT  197.2 231.8 198.2 231.0 ;
      RECT  192.2 225.8 199.8 225.0 ;
      RECT  192.2 227.4 193.0 225.8 ;
      RECT  194.8 227.4 195.8 226.6 ;
      RECT  194.8 228.0 195.6 227.4 ;
      RECT  197.2 229.8 198.0 227.4 ;
      RECT  196.8 230.6 198.0 229.8 ;
      RECT  192.2 233.6 199.8 232.8 ;
      RECT  192.2 232.2 193.0 228.0 ;
      RECT  194.8 231.0 195.6 228.8 ;
      RECT  196.6 235.0 198.2 234.2 ;
      RECT  199.0 227.4 199.8 225.8 ;
      RECT  193.8 235.0 195.4 234.2 ;
      RECT  194.6 239.8 195.6 240.6 ;
      RECT  197.0 244.2 198.0 245.0 ;
      RECT  197.2 240.6 198.0 241.0 ;
      RECT  196.0 238.8 196.8 239.0 ;
      RECT  199.0 239.4 199.8 243.6 ;
      RECT  194.8 242.8 196.4 243.6 ;
      RECT  197.0 245.0 197.8 245.8 ;
      RECT  197.2 239.8 198.2 240.6 ;
      RECT  192.2 245.8 199.8 246.6 ;
      RECT  192.2 244.2 193.0 245.8 ;
      RECT  194.8 244.2 195.8 245.0 ;
      RECT  194.8 243.6 195.6 244.2 ;
      RECT  197.2 241.8 198.0 244.2 ;
      RECT  196.8 241.0 198.0 241.8 ;
      RECT  192.2 238.0 199.8 238.8 ;
      RECT  192.2 239.4 193.0 243.6 ;
      RECT  194.8 240.6 195.6 242.8 ;
      RECT  196.6 236.6 198.2 237.4 ;
      RECT  199.0 244.2 199.8 245.8 ;
      RECT  193.8 236.6 195.4 237.4 ;
      RECT  194.6 252.6 195.6 251.8 ;
      RECT  197.0 248.2 198.0 247.4 ;
      RECT  197.2 251.8 198.0 251.4 ;
      RECT  196.0 253.6 196.8 253.4 ;
      RECT  199.0 253.0 199.8 248.8 ;
      RECT  194.8 249.6 196.4 248.8 ;
      RECT  197.0 247.4 197.8 246.6 ;
      RECT  197.2 252.6 198.2 251.8 ;
      RECT  192.2 246.6 199.8 245.8 ;
      RECT  192.2 248.2 193.0 246.6 ;
      RECT  194.8 248.2 195.8 247.4 ;
      RECT  194.8 248.8 195.6 248.2 ;
      RECT  197.2 250.6 198.0 248.2 ;
      RECT  196.8 251.4 198.0 250.6 ;
      RECT  192.2 254.4 199.8 253.6 ;
      RECT  192.2 253.0 193.0 248.8 ;
      RECT  194.8 251.8 195.6 249.6 ;
      RECT  196.6 255.8 198.2 255.0 ;
      RECT  199.0 248.2 199.8 246.6 ;
      RECT  193.8 255.8 195.4 255.0 ;
      RECT  194.6 260.6 195.6 261.4 ;
      RECT  197.0 265.0 198.0 265.8 ;
      RECT  197.2 261.4 198.0 261.8 ;
      RECT  196.0 259.6 196.8 259.8 ;
      RECT  199.0 260.2 199.8 264.4 ;
      RECT  194.8 263.6 196.4 264.4 ;
      RECT  197.0 265.8 197.8 266.6 ;
      RECT  197.2 260.6 198.2 261.4 ;
      RECT  192.2 266.6 199.8 267.4 ;
      RECT  192.2 265.0 193.0 266.6 ;
      RECT  194.8 265.0 195.8 265.8 ;
      RECT  194.8 264.4 195.6 265.0 ;
      RECT  197.2 262.6 198.0 265.0 ;
      RECT  196.8 261.8 198.0 262.6 ;
      RECT  192.2 258.8 199.8 259.6 ;
      RECT  192.2 260.2 193.0 264.4 ;
      RECT  194.8 261.4 195.6 263.6 ;
      RECT  196.6 257.4 198.2 258.2 ;
      RECT  199.0 265.0 199.8 266.6 ;
      RECT  193.8 257.4 195.4 258.2 ;
      RECT  194.6 273.4 195.6 272.6 ;
      RECT  197.0 269.0 198.0 268.2 ;
      RECT  197.2 272.6 198.0 272.2 ;
      RECT  196.0 274.4 196.8 274.2 ;
      RECT  199.0 273.8 199.8 269.6 ;
      RECT  194.8 270.4 196.4 269.6 ;
      RECT  197.0 268.2 197.8 267.4 ;
      RECT  197.2 273.4 198.2 272.6 ;
      RECT  192.2 267.4 199.8 266.6 ;
      RECT  192.2 269.0 193.0 267.4 ;
      RECT  194.8 269.0 195.8 268.2 ;
      RECT  194.8 269.6 195.6 269.0 ;
      RECT  197.2 271.4 198.0 269.0 ;
      RECT  196.8 272.2 198.0 271.4 ;
      RECT  192.2 275.2 199.8 274.4 ;
      RECT  192.2 273.8 193.0 269.6 ;
      RECT  194.8 272.6 195.6 270.4 ;
      RECT  196.6 276.6 198.2 275.8 ;
      RECT  199.0 269.0 199.8 267.4 ;
      RECT  193.8 276.6 195.4 275.8 ;
      RECT  194.6 281.4 195.6 282.2 ;
      RECT  197.0 285.8 198.0 286.6 ;
      RECT  197.2 282.2 198.0 282.6 ;
      RECT  196.0 280.4 196.8 280.6 ;
      RECT  199.0 281.0 199.8 285.2 ;
      RECT  194.8 284.4 196.4 285.2 ;
      RECT  197.0 286.6 197.8 287.4 ;
      RECT  197.2 281.4 198.2 282.2 ;
      RECT  192.2 287.4 199.8 288.2 ;
      RECT  192.2 285.8 193.0 287.4 ;
      RECT  194.8 285.8 195.8 286.6 ;
      RECT  194.8 285.2 195.6 285.8 ;
      RECT  197.2 283.4 198.0 285.8 ;
      RECT  196.8 282.6 198.0 283.4 ;
      RECT  192.2 279.6 199.8 280.4 ;
      RECT  192.2 281.0 193.0 285.2 ;
      RECT  194.8 282.2 195.6 284.4 ;
      RECT  196.6 278.2 198.2 279.0 ;
      RECT  199.0 285.8 199.8 287.4 ;
      RECT  193.8 278.2 195.4 279.0 ;
      RECT  194.6 294.2 195.6 293.4 ;
      RECT  197.0 289.8 198.0 289.0 ;
      RECT  197.2 293.4 198.0 293.0 ;
      RECT  196.0 295.2 196.8 295.0 ;
      RECT  199.0 294.6 199.8 290.4 ;
      RECT  194.8 291.2 196.4 290.4 ;
      RECT  197.0 289.0 197.8 288.2 ;
      RECT  197.2 294.2 198.2 293.4 ;
      RECT  192.2 288.2 199.8 287.4 ;
      RECT  192.2 289.8 193.0 288.2 ;
      RECT  194.8 289.8 195.8 289.0 ;
      RECT  194.8 290.4 195.6 289.8 ;
      RECT  197.2 292.2 198.0 289.8 ;
      RECT  196.8 293.0 198.0 292.2 ;
      RECT  192.2 296.0 199.8 295.2 ;
      RECT  192.2 294.6 193.0 290.4 ;
      RECT  194.8 293.4 195.6 291.2 ;
      RECT  196.6 297.4 198.2 296.6 ;
      RECT  199.0 289.8 199.8 288.2 ;
      RECT  193.8 297.4 195.4 296.6 ;
      RECT  194.6 302.2 195.6 303.0 ;
      RECT  197.0 306.6 198.0 307.4 ;
      RECT  197.2 303.0 198.0 303.4 ;
      RECT  196.0 301.2 196.8 301.4 ;
      RECT  199.0 301.8 199.8 306.0 ;
      RECT  194.8 305.2 196.4 306.0 ;
      RECT  197.0 307.4 197.8 308.2 ;
      RECT  197.2 302.2 198.2 303.0 ;
      RECT  192.2 308.2 199.8 309.0 ;
      RECT  192.2 306.6 193.0 308.2 ;
      RECT  194.8 306.6 195.8 307.4 ;
      RECT  194.8 306.0 195.6 306.6 ;
      RECT  197.2 304.2 198.0 306.6 ;
      RECT  196.8 303.4 198.0 304.2 ;
      RECT  192.2 300.4 199.8 301.2 ;
      RECT  192.2 301.8 193.0 306.0 ;
      RECT  194.8 303.0 195.6 305.2 ;
      RECT  196.6 299.0 198.2 299.8 ;
      RECT  199.0 306.6 199.8 308.2 ;
      RECT  193.8 299.0 195.4 299.8 ;
      RECT  194.6 315.0 195.6 314.2 ;
      RECT  197.0 310.6 198.0 309.8 ;
      RECT  197.2 314.2 198.0 313.8 ;
      RECT  196.0 316.0 196.8 315.8 ;
      RECT  199.0 315.4 199.8 311.2 ;
      RECT  194.8 312.0 196.4 311.2 ;
      RECT  197.0 309.8 197.8 309.0 ;
      RECT  197.2 315.0 198.2 314.2 ;
      RECT  192.2 309.0 199.8 308.2 ;
      RECT  192.2 310.6 193.0 309.0 ;
      RECT  194.8 310.6 195.8 309.8 ;
      RECT  194.8 311.2 195.6 310.6 ;
      RECT  197.2 313.0 198.0 310.6 ;
      RECT  196.8 313.8 198.0 313.0 ;
      RECT  192.2 316.8 199.8 316.0 ;
      RECT  192.2 315.4 193.0 311.2 ;
      RECT  194.8 314.2 195.6 312.0 ;
      RECT  196.6 318.2 198.2 317.4 ;
      RECT  199.0 310.6 199.8 309.0 ;
      RECT  193.8 318.2 195.4 317.4 ;
      RECT  194.6 323.0 195.6 323.8 ;
      RECT  197.0 327.4 198.0 328.2 ;
      RECT  197.2 323.8 198.0 324.2 ;
      RECT  196.0 322.0 196.8 322.2 ;
      RECT  199.0 322.6 199.8 326.8 ;
      RECT  194.8 326.0 196.4 326.8 ;
      RECT  197.0 328.2 197.8 329.0 ;
      RECT  197.2 323.0 198.2 323.8 ;
      RECT  192.2 329.0 199.8 329.8 ;
      RECT  192.2 327.4 193.0 329.0 ;
      RECT  194.8 327.4 195.8 328.2 ;
      RECT  194.8 326.8 195.6 327.4 ;
      RECT  197.2 325.0 198.0 327.4 ;
      RECT  196.8 324.2 198.0 325.0 ;
      RECT  192.2 321.2 199.8 322.0 ;
      RECT  192.2 322.6 193.0 326.8 ;
      RECT  194.8 323.8 195.6 326.0 ;
      RECT  196.6 319.8 198.2 320.6 ;
      RECT  199.0 327.4 199.8 329.0 ;
      RECT  193.8 319.8 195.4 320.6 ;
      RECT  194.6 335.8 195.6 335.0 ;
      RECT  197.0 331.4 198.0 330.6 ;
      RECT  197.2 335.0 198.0 334.6 ;
      RECT  196.0 336.8 196.8 336.6 ;
      RECT  199.0 336.2 199.8 332.0 ;
      RECT  194.8 332.8 196.4 332.0 ;
      RECT  197.0 330.6 197.8 329.8 ;
      RECT  197.2 335.8 198.2 335.0 ;
      RECT  192.2 329.8 199.8 329.0 ;
      RECT  192.2 331.4 193.0 329.8 ;
      RECT  194.8 331.4 195.8 330.6 ;
      RECT  194.8 332.0 195.6 331.4 ;
      RECT  197.2 333.8 198.0 331.4 ;
      RECT  196.8 334.6 198.0 333.8 ;
      RECT  192.2 337.6 199.8 336.8 ;
      RECT  192.2 336.2 193.0 332.0 ;
      RECT  194.8 335.0 195.6 332.8 ;
      RECT  196.6 339.0 198.2 338.2 ;
      RECT  199.0 331.4 199.8 329.8 ;
      RECT  193.8 339.0 195.4 338.2 ;
      RECT  194.6 343.8 195.6 344.6 ;
      RECT  197.0 348.2 198.0 349.0 ;
      RECT  197.2 344.6 198.0 345.0 ;
      RECT  196.0 342.8 196.8 343.0 ;
      RECT  199.0 343.4 199.8 347.6 ;
      RECT  194.8 346.8 196.4 347.6 ;
      RECT  197.0 349.0 197.8 349.8 ;
      RECT  197.2 343.8 198.2 344.6 ;
      RECT  192.2 349.8 199.8 350.6 ;
      RECT  192.2 348.2 193.0 349.8 ;
      RECT  194.8 348.2 195.8 349.0 ;
      RECT  194.8 347.6 195.6 348.2 ;
      RECT  197.2 345.8 198.0 348.2 ;
      RECT  196.8 345.0 198.0 345.8 ;
      RECT  192.2 342.0 199.8 342.8 ;
      RECT  192.2 343.4 193.0 347.6 ;
      RECT  194.8 344.6 195.6 346.8 ;
      RECT  196.6 340.6 198.2 341.4 ;
      RECT  199.0 348.2 199.8 349.8 ;
      RECT  193.8 340.6 195.4 341.4 ;
      RECT  194.6 356.6 195.6 355.8 ;
      RECT  197.0 352.2 198.0 351.4 ;
      RECT  197.2 355.8 198.0 355.4 ;
      RECT  196.0 357.6 196.8 357.4 ;
      RECT  199.0 357.0 199.8 352.8 ;
      RECT  194.8 353.6 196.4 352.8 ;
      RECT  197.0 351.4 197.8 350.6 ;
      RECT  197.2 356.6 198.2 355.8 ;
      RECT  192.2 350.6 199.8 349.8 ;
      RECT  192.2 352.2 193.0 350.6 ;
      RECT  194.8 352.2 195.8 351.4 ;
      RECT  194.8 352.8 195.6 352.2 ;
      RECT  197.2 354.6 198.0 352.2 ;
      RECT  196.8 355.4 198.0 354.6 ;
      RECT  192.2 358.4 199.8 357.6 ;
      RECT  192.2 357.0 193.0 352.8 ;
      RECT  194.8 355.8 195.6 353.6 ;
      RECT  196.6 359.8 198.2 359.0 ;
      RECT  199.0 352.2 199.8 350.6 ;
      RECT  193.8 359.8 195.4 359.0 ;
      RECT  194.6 364.6 195.6 365.4 ;
      RECT  197.0 369.0 198.0 369.8 ;
      RECT  197.2 365.4 198.0 365.8 ;
      RECT  196.0 363.6 196.8 363.8 ;
      RECT  199.0 364.2 199.8 368.4 ;
      RECT  194.8 367.6 196.4 368.4 ;
      RECT  197.2 364.6 198.2 365.4 ;
      RECT  194.6 361.4 195.4 362.2 ;
      RECT  192.2 370.6 199.8 371.4 ;
      RECT  192.2 369.0 193.0 370.6 ;
      RECT  194.8 369.0 195.8 369.8 ;
      RECT  194.8 368.4 195.6 369.0 ;
      RECT  197.2 366.6 198.0 369.0 ;
      RECT  196.8 365.8 198.0 366.6 ;
      RECT  192.2 362.8 199.8 363.6 ;
      RECT  197.4 361.4 198.2 362.2 ;
      RECT  192.2 364.2 193.0 368.4 ;
      RECT  194.8 365.4 195.6 367.6 ;
      RECT  199.0 369.0 199.8 370.6 ;
      RECT  192.6 175.6 199.4 176.4 ;
      RECT  192.6 191.2 199.4 192.0 ;
      RECT  192.6 196.4 199.4 197.2 ;
      RECT  192.6 212.0 199.4 212.8 ;
      RECT  192.6 217.2 199.4 218.0 ;
      RECT  192.6 232.8 199.4 233.6 ;
      RECT  192.6 238.0 199.4 238.8 ;
      RECT  192.6 253.6 199.4 254.4 ;
      RECT  192.6 258.8 199.4 259.6 ;
      RECT  192.6 274.4 199.4 275.2 ;
      RECT  192.6 279.6 199.4 280.4 ;
      RECT  192.6 295.2 199.4 296.0 ;
      RECT  192.6 300.4 199.4 301.2 ;
      RECT  192.6 316.0 199.4 316.8 ;
      RECT  192.6 321.2 199.4 322.0 ;
      RECT  192.6 336.8 199.4 337.6 ;
      RECT  192.6 342.0 199.4 342.8 ;
      RECT  192.6 357.6 199.4 358.4 ;
      RECT  192.6 362.8 199.4 363.6 ;
      RECT  201.4 190.2 202.4 189.4 ;
      RECT  203.8 185.8 204.8 185.0 ;
      RECT  204.0 189.4 204.8 189.0 ;
      RECT  202.8 191.2 203.6 191.0 ;
      RECT  205.8 190.6 206.6 186.4 ;
      RECT  201.6 187.2 203.2 186.4 ;
      RECT  204.0 190.2 205.0 189.4 ;
      RECT  201.4 193.4 202.2 192.6 ;
      RECT  199.0 184.2 206.6 183.4 ;
      RECT  199.0 185.8 199.8 184.2 ;
      RECT  201.6 185.8 202.6 185.0 ;
      RECT  201.6 186.4 202.4 185.8 ;
      RECT  204.0 188.2 204.8 185.8 ;
      RECT  203.6 189.0 204.8 188.2 ;
      RECT  199.0 192.0 206.6 191.2 ;
      RECT  204.2 193.4 205.0 192.6 ;
      RECT  199.0 190.6 199.8 186.4 ;
      RECT  201.6 189.4 202.4 187.2 ;
      RECT  205.8 185.8 206.6 184.2 ;
      RECT  208.2 190.2 209.2 189.4 ;
      RECT  210.6 185.8 211.6 185.0 ;
      RECT  210.8 189.4 211.6 189.0 ;
      RECT  209.6 191.2 210.4 191.0 ;
      RECT  212.6 190.6 213.4 186.4 ;
      RECT  208.4 187.2 210.0 186.4 ;
      RECT  210.8 190.2 211.8 189.4 ;
      RECT  208.2 193.4 209.0 192.6 ;
      RECT  205.8 184.2 213.4 183.4 ;
      RECT  205.8 185.8 206.6 184.2 ;
      RECT  208.4 185.8 209.4 185.0 ;
      RECT  208.4 186.4 209.2 185.8 ;
      RECT  210.8 188.2 211.6 185.8 ;
      RECT  210.4 189.0 211.6 188.2 ;
      RECT  205.8 192.0 213.4 191.2 ;
      RECT  211.0 193.4 211.8 192.6 ;
      RECT  205.8 190.6 206.6 186.4 ;
      RECT  208.4 189.4 209.2 187.2 ;
      RECT  212.6 185.8 213.4 184.2 ;
      RECT  199.0 192.0 212.6 191.2 ;
      RECT  201.4 177.4 202.4 178.2 ;
      RECT  203.8 181.8 204.8 182.6 ;
      RECT  204.0 178.2 204.8 178.6 ;
      RECT  202.8 176.4 203.6 176.6 ;
      RECT  205.8 177.0 206.6 181.2 ;
      RECT  201.6 180.4 203.2 181.2 ;
      RECT  204.0 177.4 205.0 178.2 ;
      RECT  201.4 174.2 202.2 175.0 ;
      RECT  199.0 183.4 206.6 184.2 ;
      RECT  199.0 181.8 199.8 183.4 ;
      RECT  201.6 181.8 202.6 182.6 ;
      RECT  201.6 181.2 202.4 181.8 ;
      RECT  204.0 179.4 204.8 181.8 ;
      RECT  203.6 178.6 204.8 179.4 ;
      RECT  199.0 175.6 206.6 176.4 ;
      RECT  204.2 174.2 205.0 175.0 ;
      RECT  199.0 177.0 199.8 181.2 ;
      RECT  201.6 178.2 202.4 180.4 ;
      RECT  205.8 181.8 206.6 183.4 ;
      RECT  208.2 177.4 209.2 178.2 ;
      RECT  210.6 181.8 211.6 182.6 ;
      RECT  210.8 178.2 211.6 178.6 ;
      RECT  209.6 176.4 210.4 176.6 ;
      RECT  212.6 177.0 213.4 181.2 ;
      RECT  208.4 180.4 210.0 181.2 ;
      RECT  210.8 177.4 211.8 178.2 ;
      RECT  208.2 174.2 209.0 175.0 ;
      RECT  205.8 183.4 213.4 184.2 ;
      RECT  205.8 181.8 206.6 183.4 ;
      RECT  208.4 181.8 209.4 182.6 ;
      RECT  208.4 181.2 209.2 181.8 ;
      RECT  210.8 179.4 211.6 181.8 ;
      RECT  210.4 178.6 211.6 179.4 ;
      RECT  205.8 175.6 213.4 176.4 ;
      RECT  211.0 174.2 211.8 175.0 ;
      RECT  205.8 177.0 206.6 181.2 ;
      RECT  208.4 178.2 209.2 180.4 ;
      RECT  212.6 181.8 213.4 183.4 ;
      RECT  199.0 175.6 212.6 176.4 ;
      RECT  201.4 364.6 202.4 365.4 ;
      RECT  203.8 369.0 204.8 369.8 ;
      RECT  204.0 365.4 204.8 365.8 ;
      RECT  202.8 363.6 203.6 363.8 ;
      RECT  205.8 364.2 206.6 368.4 ;
      RECT  201.6 367.6 203.2 368.4 ;
      RECT  204.0 364.6 205.0 365.4 ;
      RECT  201.4 361.4 202.2 362.2 ;
      RECT  199.0 370.6 206.6 371.4 ;
      RECT  199.0 369.0 199.8 370.6 ;
      RECT  201.6 369.0 202.6 369.8 ;
      RECT  201.6 368.4 202.4 369.0 ;
      RECT  204.0 366.6 204.8 369.0 ;
      RECT  203.6 365.8 204.8 366.6 ;
      RECT  199.0 362.8 206.6 363.6 ;
      RECT  204.2 361.4 205.0 362.2 ;
      RECT  199.0 364.2 199.8 368.4 ;
      RECT  201.6 365.4 202.4 367.6 ;
      RECT  205.8 369.0 206.6 370.6 ;
      RECT  208.2 364.6 209.2 365.4 ;
      RECT  210.6 369.0 211.6 369.8 ;
      RECT  210.8 365.4 211.6 365.8 ;
      RECT  209.6 363.6 210.4 363.8 ;
      RECT  212.6 364.2 213.4 368.4 ;
      RECT  208.4 367.6 210.0 368.4 ;
      RECT  210.8 364.6 211.8 365.4 ;
      RECT  208.2 361.4 209.0 362.2 ;
      RECT  205.8 370.6 213.4 371.4 ;
      RECT  205.8 369.0 206.6 370.6 ;
      RECT  208.4 369.0 209.4 369.8 ;
      RECT  208.4 368.4 209.2 369.0 ;
      RECT  210.8 366.6 211.6 369.0 ;
      RECT  210.4 365.8 211.6 366.6 ;
      RECT  205.8 362.8 213.4 363.6 ;
      RECT  211.0 361.4 211.8 362.2 ;
      RECT  205.8 364.2 206.6 368.4 ;
      RECT  208.4 365.4 209.2 367.6 ;
      RECT  212.6 369.0 213.4 370.6 ;
      RECT  199.0 362.8 212.6 363.6 ;
      RECT  187.8 177.4 188.8 178.2 ;
      RECT  190.2 181.8 191.2 182.6 ;
      RECT  190.4 178.2 191.2 178.6 ;
      RECT  189.2 176.4 190.0 176.6 ;
      RECT  192.2 177.0 193.0 181.2 ;
      RECT  188.0 180.4 189.6 181.2 ;
      RECT  190.4 177.4 191.4 178.2 ;
      RECT  187.8 174.2 188.6 175.0 ;
      RECT  185.4 183.4 193.0 184.2 ;
      RECT  185.4 181.8 186.2 183.4 ;
      RECT  188.0 181.8 189.0 182.6 ;
      RECT  188.0 181.2 188.8 181.8 ;
      RECT  190.4 179.4 191.2 181.8 ;
      RECT  190.0 178.6 191.2 179.4 ;
      RECT  185.4 175.6 193.0 176.4 ;
      RECT  190.6 174.2 191.4 175.0 ;
      RECT  185.4 177.0 186.2 181.2 ;
      RECT  188.0 178.2 188.8 180.4 ;
      RECT  192.2 181.8 193.0 183.4 ;
      RECT  187.8 190.2 188.8 189.4 ;
      RECT  190.2 185.8 191.2 185.0 ;
      RECT  190.4 189.4 191.2 189.0 ;
      RECT  189.2 191.2 190.0 191.0 ;
      RECT  192.2 190.6 193.0 186.4 ;
      RECT  188.0 187.2 189.6 186.4 ;
      RECT  190.4 190.2 191.4 189.4 ;
      RECT  187.8 193.4 188.6 192.6 ;
      RECT  185.4 184.2 193.0 183.4 ;
      RECT  185.4 185.8 186.2 184.2 ;
      RECT  188.0 185.8 189.0 185.0 ;
      RECT  188.0 186.4 188.8 185.8 ;
      RECT  190.4 188.2 191.2 185.8 ;
      RECT  190.0 189.0 191.2 188.2 ;
      RECT  185.4 192.0 193.0 191.2 ;
      RECT  190.6 193.4 191.4 192.6 ;
      RECT  185.4 190.6 186.2 186.4 ;
      RECT  188.0 189.4 188.8 187.2 ;
      RECT  192.2 185.8 193.0 184.2 ;
      RECT  187.8 198.2 188.8 199.0 ;
      RECT  190.2 202.6 191.2 203.4 ;
      RECT  190.4 199.0 191.2 199.4 ;
      RECT  189.2 197.2 190.0 197.4 ;
      RECT  192.2 197.8 193.0 202.0 ;
      RECT  188.0 201.2 189.6 202.0 ;
      RECT  190.4 198.2 191.4 199.0 ;
      RECT  187.8 195.0 188.6 195.8 ;
      RECT  185.4 204.2 193.0 205.0 ;
      RECT  185.4 202.6 186.2 204.2 ;
      RECT  188.0 202.6 189.0 203.4 ;
      RECT  188.0 202.0 188.8 202.6 ;
      RECT  190.4 200.2 191.2 202.6 ;
      RECT  190.0 199.4 191.2 200.2 ;
      RECT  185.4 196.4 193.0 197.2 ;
      RECT  190.6 195.0 191.4 195.8 ;
      RECT  185.4 197.8 186.2 202.0 ;
      RECT  188.0 199.0 188.8 201.2 ;
      RECT  192.2 202.6 193.0 204.2 ;
      RECT  187.8 211.0 188.8 210.2 ;
      RECT  190.2 206.6 191.2 205.8 ;
      RECT  190.4 210.2 191.2 209.8 ;
      RECT  189.2 212.0 190.0 211.8 ;
      RECT  192.2 211.4 193.0 207.2 ;
      RECT  188.0 208.0 189.6 207.2 ;
      RECT  190.4 211.0 191.4 210.2 ;
      RECT  187.8 214.2 188.6 213.4 ;
      RECT  185.4 205.0 193.0 204.2 ;
      RECT  185.4 206.6 186.2 205.0 ;
      RECT  188.0 206.6 189.0 205.8 ;
      RECT  188.0 207.2 188.8 206.6 ;
      RECT  190.4 209.0 191.2 206.6 ;
      RECT  190.0 209.8 191.2 209.0 ;
      RECT  185.4 212.8 193.0 212.0 ;
      RECT  190.6 214.2 191.4 213.4 ;
      RECT  185.4 211.4 186.2 207.2 ;
      RECT  188.0 210.2 188.8 208.0 ;
      RECT  192.2 206.6 193.0 205.0 ;
      RECT  187.8 219.0 188.8 219.8 ;
      RECT  190.2 223.4 191.2 224.2 ;
      RECT  190.4 219.8 191.2 220.2 ;
      RECT  189.2 218.0 190.0 218.2 ;
      RECT  192.2 218.6 193.0 222.8 ;
      RECT  188.0 222.0 189.6 222.8 ;
      RECT  190.4 219.0 191.4 219.8 ;
      RECT  187.8 215.8 188.6 216.6 ;
      RECT  185.4 225.0 193.0 225.8 ;
      RECT  185.4 223.4 186.2 225.0 ;
      RECT  188.0 223.4 189.0 224.2 ;
      RECT  188.0 222.8 188.8 223.4 ;
      RECT  190.4 221.0 191.2 223.4 ;
      RECT  190.0 220.2 191.2 221.0 ;
      RECT  185.4 217.2 193.0 218.0 ;
      RECT  190.6 215.8 191.4 216.6 ;
      RECT  185.4 218.6 186.2 222.8 ;
      RECT  188.0 219.8 188.8 222.0 ;
      RECT  192.2 223.4 193.0 225.0 ;
      RECT  187.8 231.8 188.8 231.0 ;
      RECT  190.2 227.4 191.2 226.6 ;
      RECT  190.4 231.0 191.2 230.6 ;
      RECT  189.2 232.8 190.0 232.6 ;
      RECT  192.2 232.2 193.0 228.0 ;
      RECT  188.0 228.8 189.6 228.0 ;
      RECT  190.4 231.8 191.4 231.0 ;
      RECT  187.8 235.0 188.6 234.2 ;
      RECT  185.4 225.8 193.0 225.0 ;
      RECT  185.4 227.4 186.2 225.8 ;
      RECT  188.0 227.4 189.0 226.6 ;
      RECT  188.0 228.0 188.8 227.4 ;
      RECT  190.4 229.8 191.2 227.4 ;
      RECT  190.0 230.6 191.2 229.8 ;
      RECT  185.4 233.6 193.0 232.8 ;
      RECT  190.6 235.0 191.4 234.2 ;
      RECT  185.4 232.2 186.2 228.0 ;
      RECT  188.0 231.0 188.8 228.8 ;
      RECT  192.2 227.4 193.0 225.8 ;
      RECT  187.8 239.8 188.8 240.6 ;
      RECT  190.2 244.2 191.2 245.0 ;
      RECT  190.4 240.6 191.2 241.0 ;
      RECT  189.2 238.8 190.0 239.0 ;
      RECT  192.2 239.4 193.0 243.6 ;
      RECT  188.0 242.8 189.6 243.6 ;
      RECT  190.4 239.8 191.4 240.6 ;
      RECT  187.8 236.6 188.6 237.4 ;
      RECT  185.4 245.8 193.0 246.6 ;
      RECT  185.4 244.2 186.2 245.8 ;
      RECT  188.0 244.2 189.0 245.0 ;
      RECT  188.0 243.6 188.8 244.2 ;
      RECT  190.4 241.8 191.2 244.2 ;
      RECT  190.0 241.0 191.2 241.8 ;
      RECT  185.4 238.0 193.0 238.8 ;
      RECT  190.6 236.6 191.4 237.4 ;
      RECT  185.4 239.4 186.2 243.6 ;
      RECT  188.0 240.6 188.8 242.8 ;
      RECT  192.2 244.2 193.0 245.8 ;
      RECT  187.8 252.6 188.8 251.8 ;
      RECT  190.2 248.2 191.2 247.4 ;
      RECT  190.4 251.8 191.2 251.4 ;
      RECT  189.2 253.6 190.0 253.4 ;
      RECT  192.2 253.0 193.0 248.8 ;
      RECT  188.0 249.6 189.6 248.8 ;
      RECT  190.4 252.6 191.4 251.8 ;
      RECT  187.8 255.8 188.6 255.0 ;
      RECT  185.4 246.6 193.0 245.8 ;
      RECT  185.4 248.2 186.2 246.6 ;
      RECT  188.0 248.2 189.0 247.4 ;
      RECT  188.0 248.8 188.8 248.2 ;
      RECT  190.4 250.6 191.2 248.2 ;
      RECT  190.0 251.4 191.2 250.6 ;
      RECT  185.4 254.4 193.0 253.6 ;
      RECT  190.6 255.8 191.4 255.0 ;
      RECT  185.4 253.0 186.2 248.8 ;
      RECT  188.0 251.8 188.8 249.6 ;
      RECT  192.2 248.2 193.0 246.6 ;
      RECT  187.8 260.6 188.8 261.4 ;
      RECT  190.2 265.0 191.2 265.8 ;
      RECT  190.4 261.4 191.2 261.8 ;
      RECT  189.2 259.6 190.0 259.8 ;
      RECT  192.2 260.2 193.0 264.4 ;
      RECT  188.0 263.6 189.6 264.4 ;
      RECT  190.4 260.6 191.4 261.4 ;
      RECT  187.8 257.4 188.6 258.2 ;
      RECT  185.4 266.6 193.0 267.4 ;
      RECT  185.4 265.0 186.2 266.6 ;
      RECT  188.0 265.0 189.0 265.8 ;
      RECT  188.0 264.4 188.8 265.0 ;
      RECT  190.4 262.6 191.2 265.0 ;
      RECT  190.0 261.8 191.2 262.6 ;
      RECT  185.4 258.8 193.0 259.6 ;
      RECT  190.6 257.4 191.4 258.2 ;
      RECT  185.4 260.2 186.2 264.4 ;
      RECT  188.0 261.4 188.8 263.6 ;
      RECT  192.2 265.0 193.0 266.6 ;
      RECT  187.8 273.4 188.8 272.6 ;
      RECT  190.2 269.0 191.2 268.2 ;
      RECT  190.4 272.6 191.2 272.2 ;
      RECT  189.2 274.4 190.0 274.2 ;
      RECT  192.2 273.8 193.0 269.6 ;
      RECT  188.0 270.4 189.6 269.6 ;
      RECT  190.4 273.4 191.4 272.6 ;
      RECT  187.8 276.6 188.6 275.8 ;
      RECT  185.4 267.4 193.0 266.6 ;
      RECT  185.4 269.0 186.2 267.4 ;
      RECT  188.0 269.0 189.0 268.2 ;
      RECT  188.0 269.6 188.8 269.0 ;
      RECT  190.4 271.4 191.2 269.0 ;
      RECT  190.0 272.2 191.2 271.4 ;
      RECT  185.4 275.2 193.0 274.4 ;
      RECT  190.6 276.6 191.4 275.8 ;
      RECT  185.4 273.8 186.2 269.6 ;
      RECT  188.0 272.6 188.8 270.4 ;
      RECT  192.2 269.0 193.0 267.4 ;
      RECT  187.8 281.4 188.8 282.2 ;
      RECT  190.2 285.8 191.2 286.6 ;
      RECT  190.4 282.2 191.2 282.6 ;
      RECT  189.2 280.4 190.0 280.6 ;
      RECT  192.2 281.0 193.0 285.2 ;
      RECT  188.0 284.4 189.6 285.2 ;
      RECT  190.4 281.4 191.4 282.2 ;
      RECT  187.8 278.2 188.6 279.0 ;
      RECT  185.4 287.4 193.0 288.2 ;
      RECT  185.4 285.8 186.2 287.4 ;
      RECT  188.0 285.8 189.0 286.6 ;
      RECT  188.0 285.2 188.8 285.8 ;
      RECT  190.4 283.4 191.2 285.8 ;
      RECT  190.0 282.6 191.2 283.4 ;
      RECT  185.4 279.6 193.0 280.4 ;
      RECT  190.6 278.2 191.4 279.0 ;
      RECT  185.4 281.0 186.2 285.2 ;
      RECT  188.0 282.2 188.8 284.4 ;
      RECT  192.2 285.8 193.0 287.4 ;
      RECT  187.8 294.2 188.8 293.4 ;
      RECT  190.2 289.8 191.2 289.0 ;
      RECT  190.4 293.4 191.2 293.0 ;
      RECT  189.2 295.2 190.0 295.0 ;
      RECT  192.2 294.6 193.0 290.4 ;
      RECT  188.0 291.2 189.6 290.4 ;
      RECT  190.4 294.2 191.4 293.4 ;
      RECT  187.8 297.4 188.6 296.6 ;
      RECT  185.4 288.2 193.0 287.4 ;
      RECT  185.4 289.8 186.2 288.2 ;
      RECT  188.0 289.8 189.0 289.0 ;
      RECT  188.0 290.4 188.8 289.8 ;
      RECT  190.4 292.2 191.2 289.8 ;
      RECT  190.0 293.0 191.2 292.2 ;
      RECT  185.4 296.0 193.0 295.2 ;
      RECT  190.6 297.4 191.4 296.6 ;
      RECT  185.4 294.6 186.2 290.4 ;
      RECT  188.0 293.4 188.8 291.2 ;
      RECT  192.2 289.8 193.0 288.2 ;
      RECT  187.8 302.2 188.8 303.0 ;
      RECT  190.2 306.6 191.2 307.4 ;
      RECT  190.4 303.0 191.2 303.4 ;
      RECT  189.2 301.2 190.0 301.4 ;
      RECT  192.2 301.8 193.0 306.0 ;
      RECT  188.0 305.2 189.6 306.0 ;
      RECT  190.4 302.2 191.4 303.0 ;
      RECT  187.8 299.0 188.6 299.8 ;
      RECT  185.4 308.2 193.0 309.0 ;
      RECT  185.4 306.6 186.2 308.2 ;
      RECT  188.0 306.6 189.0 307.4 ;
      RECT  188.0 306.0 188.8 306.6 ;
      RECT  190.4 304.2 191.2 306.6 ;
      RECT  190.0 303.4 191.2 304.2 ;
      RECT  185.4 300.4 193.0 301.2 ;
      RECT  190.6 299.0 191.4 299.8 ;
      RECT  185.4 301.8 186.2 306.0 ;
      RECT  188.0 303.0 188.8 305.2 ;
      RECT  192.2 306.6 193.0 308.2 ;
      RECT  187.8 315.0 188.8 314.2 ;
      RECT  190.2 310.6 191.2 309.8 ;
      RECT  190.4 314.2 191.2 313.8 ;
      RECT  189.2 316.0 190.0 315.8 ;
      RECT  192.2 315.4 193.0 311.2 ;
      RECT  188.0 312.0 189.6 311.2 ;
      RECT  190.4 315.0 191.4 314.2 ;
      RECT  187.8 318.2 188.6 317.4 ;
      RECT  185.4 309.0 193.0 308.2 ;
      RECT  185.4 310.6 186.2 309.0 ;
      RECT  188.0 310.6 189.0 309.8 ;
      RECT  188.0 311.2 188.8 310.6 ;
      RECT  190.4 313.0 191.2 310.6 ;
      RECT  190.0 313.8 191.2 313.0 ;
      RECT  185.4 316.8 193.0 316.0 ;
      RECT  190.6 318.2 191.4 317.4 ;
      RECT  185.4 315.4 186.2 311.2 ;
      RECT  188.0 314.2 188.8 312.0 ;
      RECT  192.2 310.6 193.0 309.0 ;
      RECT  187.8 323.0 188.8 323.8 ;
      RECT  190.2 327.4 191.2 328.2 ;
      RECT  190.4 323.8 191.2 324.2 ;
      RECT  189.2 322.0 190.0 322.2 ;
      RECT  192.2 322.6 193.0 326.8 ;
      RECT  188.0 326.0 189.6 326.8 ;
      RECT  190.4 323.0 191.4 323.8 ;
      RECT  187.8 319.8 188.6 320.6 ;
      RECT  185.4 329.0 193.0 329.8 ;
      RECT  185.4 327.4 186.2 329.0 ;
      RECT  188.0 327.4 189.0 328.2 ;
      RECT  188.0 326.8 188.8 327.4 ;
      RECT  190.4 325.0 191.2 327.4 ;
      RECT  190.0 324.2 191.2 325.0 ;
      RECT  185.4 321.2 193.0 322.0 ;
      RECT  190.6 319.8 191.4 320.6 ;
      RECT  185.4 322.6 186.2 326.8 ;
      RECT  188.0 323.8 188.8 326.0 ;
      RECT  192.2 327.4 193.0 329.0 ;
      RECT  187.8 335.8 188.8 335.0 ;
      RECT  190.2 331.4 191.2 330.6 ;
      RECT  190.4 335.0 191.2 334.6 ;
      RECT  189.2 336.8 190.0 336.6 ;
      RECT  192.2 336.2 193.0 332.0 ;
      RECT  188.0 332.8 189.6 332.0 ;
      RECT  190.4 335.8 191.4 335.0 ;
      RECT  187.8 339.0 188.6 338.2 ;
      RECT  185.4 329.8 193.0 329.0 ;
      RECT  185.4 331.4 186.2 329.8 ;
      RECT  188.0 331.4 189.0 330.6 ;
      RECT  188.0 332.0 188.8 331.4 ;
      RECT  190.4 333.8 191.2 331.4 ;
      RECT  190.0 334.6 191.2 333.8 ;
      RECT  185.4 337.6 193.0 336.8 ;
      RECT  190.6 339.0 191.4 338.2 ;
      RECT  185.4 336.2 186.2 332.0 ;
      RECT  188.0 335.0 188.8 332.8 ;
      RECT  192.2 331.4 193.0 329.8 ;
      RECT  187.8 343.8 188.8 344.6 ;
      RECT  190.2 348.2 191.2 349.0 ;
      RECT  190.4 344.6 191.2 345.0 ;
      RECT  189.2 342.8 190.0 343.0 ;
      RECT  192.2 343.4 193.0 347.6 ;
      RECT  188.0 346.8 189.6 347.6 ;
      RECT  190.4 343.8 191.4 344.6 ;
      RECT  187.8 340.6 188.6 341.4 ;
      RECT  185.4 349.8 193.0 350.6 ;
      RECT  185.4 348.2 186.2 349.8 ;
      RECT  188.0 348.2 189.0 349.0 ;
      RECT  188.0 347.6 188.8 348.2 ;
      RECT  190.4 345.8 191.2 348.2 ;
      RECT  190.0 345.0 191.2 345.8 ;
      RECT  185.4 342.0 193.0 342.8 ;
      RECT  190.6 340.6 191.4 341.4 ;
      RECT  185.4 343.4 186.2 347.6 ;
      RECT  188.0 344.6 188.8 346.8 ;
      RECT  192.2 348.2 193.0 349.8 ;
      RECT  187.8 356.6 188.8 355.8 ;
      RECT  190.2 352.2 191.2 351.4 ;
      RECT  190.4 355.8 191.2 355.4 ;
      RECT  189.2 357.6 190.0 357.4 ;
      RECT  192.2 357.0 193.0 352.8 ;
      RECT  188.0 353.6 189.6 352.8 ;
      RECT  190.4 356.6 191.4 355.8 ;
      RECT  187.8 359.8 188.6 359.0 ;
      RECT  185.4 350.6 193.0 349.8 ;
      RECT  185.4 352.2 186.2 350.6 ;
      RECT  188.0 352.2 189.0 351.4 ;
      RECT  188.0 352.8 188.8 352.2 ;
      RECT  190.4 354.6 191.2 352.2 ;
      RECT  190.0 355.4 191.2 354.6 ;
      RECT  185.4 358.4 193.0 357.6 ;
      RECT  190.6 359.8 191.4 359.0 ;
      RECT  185.4 357.0 186.2 352.8 ;
      RECT  188.0 355.8 188.8 353.6 ;
      RECT  192.2 352.2 193.0 350.6 ;
      RECT  187.8 364.6 188.8 365.4 ;
      RECT  190.2 369.0 191.2 369.8 ;
      RECT  190.4 365.4 191.2 365.8 ;
      RECT  189.2 363.6 190.0 363.8 ;
      RECT  192.2 364.2 193.0 368.4 ;
      RECT  188.0 367.6 189.6 368.4 ;
      RECT  190.4 364.6 191.4 365.4 ;
      RECT  187.8 361.4 188.6 362.2 ;
      RECT  185.4 370.6 193.0 371.4 ;
      RECT  185.4 369.0 186.2 370.6 ;
      RECT  188.0 369.0 189.0 369.8 ;
      RECT  188.0 368.4 188.8 369.0 ;
      RECT  190.4 366.6 191.2 369.0 ;
      RECT  190.0 365.8 191.2 366.6 ;
      RECT  185.4 362.8 193.0 363.6 ;
      RECT  190.6 361.4 191.4 362.2 ;
      RECT  185.4 364.2 186.2 368.4 ;
      RECT  188.0 365.4 188.8 367.6 ;
      RECT  192.2 369.0 193.0 370.6 ;
      RECT  185.4 175.6 192.2 176.4 ;
      RECT  185.4 191.2 192.2 192.0 ;
      RECT  185.4 196.4 192.2 197.2 ;
      RECT  185.4 212.0 192.2 212.8 ;
      RECT  185.4 217.2 192.2 218.0 ;
      RECT  185.4 232.8 192.2 233.6 ;
      RECT  185.4 238.0 192.2 238.8 ;
      RECT  185.4 253.6 192.2 254.4 ;
      RECT  185.4 258.8 192.2 259.6 ;
      RECT  185.4 274.4 192.2 275.2 ;
      RECT  185.4 279.6 192.2 280.4 ;
      RECT  185.4 295.2 192.2 296.0 ;
      RECT  185.4 300.4 192.2 301.2 ;
      RECT  185.4 316.0 192.2 316.8 ;
      RECT  185.4 321.2 192.2 322.0 ;
      RECT  185.4 336.8 192.2 337.6 ;
      RECT  185.4 342.0 192.2 342.8 ;
      RECT  185.4 357.6 192.2 358.4 ;
      RECT  185.4 362.8 192.2 363.6 ;
      RECT  215.0 177.4 216.0 178.2 ;
      RECT  217.4 181.8 218.4 182.6 ;
      RECT  217.6 178.2 218.4 178.6 ;
      RECT  216.4 176.4 217.2 176.6 ;
      RECT  219.4 177.0 220.2 181.2 ;
      RECT  215.2 180.4 216.8 181.2 ;
      RECT  217.6 177.4 218.6 178.2 ;
      RECT  215.0 174.2 215.8 175.0 ;
      RECT  212.6 183.4 220.2 184.2 ;
      RECT  212.6 181.8 213.4 183.4 ;
      RECT  215.2 181.8 216.2 182.6 ;
      RECT  215.2 181.2 216.0 181.8 ;
      RECT  217.6 179.4 218.4 181.8 ;
      RECT  217.2 178.6 218.4 179.4 ;
      RECT  212.6 175.6 220.2 176.4 ;
      RECT  217.8 174.2 218.6 175.0 ;
      RECT  212.6 177.0 213.4 181.2 ;
      RECT  215.2 178.2 216.0 180.4 ;
      RECT  219.4 181.8 220.2 183.4 ;
      RECT  215.0 190.2 216.0 189.4 ;
      RECT  217.4 185.8 218.4 185.0 ;
      RECT  217.6 189.4 218.4 189.0 ;
      RECT  216.4 191.2 217.2 191.0 ;
      RECT  219.4 190.6 220.2 186.4 ;
      RECT  215.2 187.2 216.8 186.4 ;
      RECT  217.6 190.2 218.6 189.4 ;
      RECT  215.0 193.4 215.8 192.6 ;
      RECT  212.6 184.2 220.2 183.4 ;
      RECT  212.6 185.8 213.4 184.2 ;
      RECT  215.2 185.8 216.2 185.0 ;
      RECT  215.2 186.4 216.0 185.8 ;
      RECT  217.6 188.2 218.4 185.8 ;
      RECT  217.2 189.0 218.4 188.2 ;
      RECT  212.6 192.0 220.2 191.2 ;
      RECT  217.8 193.4 218.6 192.6 ;
      RECT  212.6 190.6 213.4 186.4 ;
      RECT  215.2 189.4 216.0 187.2 ;
      RECT  219.4 185.8 220.2 184.2 ;
      RECT  215.0 198.2 216.0 199.0 ;
      RECT  217.4 202.6 218.4 203.4 ;
      RECT  217.6 199.0 218.4 199.4 ;
      RECT  216.4 197.2 217.2 197.4 ;
      RECT  219.4 197.8 220.2 202.0 ;
      RECT  215.2 201.2 216.8 202.0 ;
      RECT  217.6 198.2 218.6 199.0 ;
      RECT  215.0 195.0 215.8 195.8 ;
      RECT  212.6 204.2 220.2 205.0 ;
      RECT  212.6 202.6 213.4 204.2 ;
      RECT  215.2 202.6 216.2 203.4 ;
      RECT  215.2 202.0 216.0 202.6 ;
      RECT  217.6 200.2 218.4 202.6 ;
      RECT  217.2 199.4 218.4 200.2 ;
      RECT  212.6 196.4 220.2 197.2 ;
      RECT  217.8 195.0 218.6 195.8 ;
      RECT  212.6 197.8 213.4 202.0 ;
      RECT  215.2 199.0 216.0 201.2 ;
      RECT  219.4 202.6 220.2 204.2 ;
      RECT  215.0 211.0 216.0 210.2 ;
      RECT  217.4 206.6 218.4 205.8 ;
      RECT  217.6 210.2 218.4 209.8 ;
      RECT  216.4 212.0 217.2 211.8 ;
      RECT  219.4 211.4 220.2 207.2 ;
      RECT  215.2 208.0 216.8 207.2 ;
      RECT  217.6 211.0 218.6 210.2 ;
      RECT  215.0 214.2 215.8 213.4 ;
      RECT  212.6 205.0 220.2 204.2 ;
      RECT  212.6 206.6 213.4 205.0 ;
      RECT  215.2 206.6 216.2 205.8 ;
      RECT  215.2 207.2 216.0 206.6 ;
      RECT  217.6 209.0 218.4 206.6 ;
      RECT  217.2 209.8 218.4 209.0 ;
      RECT  212.6 212.8 220.2 212.0 ;
      RECT  217.8 214.2 218.6 213.4 ;
      RECT  212.6 211.4 213.4 207.2 ;
      RECT  215.2 210.2 216.0 208.0 ;
      RECT  219.4 206.6 220.2 205.0 ;
      RECT  215.0 219.0 216.0 219.8 ;
      RECT  217.4 223.4 218.4 224.2 ;
      RECT  217.6 219.8 218.4 220.2 ;
      RECT  216.4 218.0 217.2 218.2 ;
      RECT  219.4 218.6 220.2 222.8 ;
      RECT  215.2 222.0 216.8 222.8 ;
      RECT  217.6 219.0 218.6 219.8 ;
      RECT  215.0 215.8 215.8 216.6 ;
      RECT  212.6 225.0 220.2 225.8 ;
      RECT  212.6 223.4 213.4 225.0 ;
      RECT  215.2 223.4 216.2 224.2 ;
      RECT  215.2 222.8 216.0 223.4 ;
      RECT  217.6 221.0 218.4 223.4 ;
      RECT  217.2 220.2 218.4 221.0 ;
      RECT  212.6 217.2 220.2 218.0 ;
      RECT  217.8 215.8 218.6 216.6 ;
      RECT  212.6 218.6 213.4 222.8 ;
      RECT  215.2 219.8 216.0 222.0 ;
      RECT  219.4 223.4 220.2 225.0 ;
      RECT  215.0 231.8 216.0 231.0 ;
      RECT  217.4 227.4 218.4 226.6 ;
      RECT  217.6 231.0 218.4 230.6 ;
      RECT  216.4 232.8 217.2 232.6 ;
      RECT  219.4 232.2 220.2 228.0 ;
      RECT  215.2 228.8 216.8 228.0 ;
      RECT  217.6 231.8 218.6 231.0 ;
      RECT  215.0 235.0 215.8 234.2 ;
      RECT  212.6 225.8 220.2 225.0 ;
      RECT  212.6 227.4 213.4 225.8 ;
      RECT  215.2 227.4 216.2 226.6 ;
      RECT  215.2 228.0 216.0 227.4 ;
      RECT  217.6 229.8 218.4 227.4 ;
      RECT  217.2 230.6 218.4 229.8 ;
      RECT  212.6 233.6 220.2 232.8 ;
      RECT  217.8 235.0 218.6 234.2 ;
      RECT  212.6 232.2 213.4 228.0 ;
      RECT  215.2 231.0 216.0 228.8 ;
      RECT  219.4 227.4 220.2 225.8 ;
      RECT  215.0 239.8 216.0 240.6 ;
      RECT  217.4 244.2 218.4 245.0 ;
      RECT  217.6 240.6 218.4 241.0 ;
      RECT  216.4 238.8 217.2 239.0 ;
      RECT  219.4 239.4 220.2 243.6 ;
      RECT  215.2 242.8 216.8 243.6 ;
      RECT  217.6 239.8 218.6 240.6 ;
      RECT  215.0 236.6 215.8 237.4 ;
      RECT  212.6 245.8 220.2 246.6 ;
      RECT  212.6 244.2 213.4 245.8 ;
      RECT  215.2 244.2 216.2 245.0 ;
      RECT  215.2 243.6 216.0 244.2 ;
      RECT  217.6 241.8 218.4 244.2 ;
      RECT  217.2 241.0 218.4 241.8 ;
      RECT  212.6 238.0 220.2 238.8 ;
      RECT  217.8 236.6 218.6 237.4 ;
      RECT  212.6 239.4 213.4 243.6 ;
      RECT  215.2 240.6 216.0 242.8 ;
      RECT  219.4 244.2 220.2 245.8 ;
      RECT  215.0 252.6 216.0 251.8 ;
      RECT  217.4 248.2 218.4 247.4 ;
      RECT  217.6 251.8 218.4 251.4 ;
      RECT  216.4 253.6 217.2 253.4 ;
      RECT  219.4 253.0 220.2 248.8 ;
      RECT  215.2 249.6 216.8 248.8 ;
      RECT  217.6 252.6 218.6 251.8 ;
      RECT  215.0 255.8 215.8 255.0 ;
      RECT  212.6 246.6 220.2 245.8 ;
      RECT  212.6 248.2 213.4 246.6 ;
      RECT  215.2 248.2 216.2 247.4 ;
      RECT  215.2 248.8 216.0 248.2 ;
      RECT  217.6 250.6 218.4 248.2 ;
      RECT  217.2 251.4 218.4 250.6 ;
      RECT  212.6 254.4 220.2 253.6 ;
      RECT  217.8 255.8 218.6 255.0 ;
      RECT  212.6 253.0 213.4 248.8 ;
      RECT  215.2 251.8 216.0 249.6 ;
      RECT  219.4 248.2 220.2 246.6 ;
      RECT  215.0 260.6 216.0 261.4 ;
      RECT  217.4 265.0 218.4 265.8 ;
      RECT  217.6 261.4 218.4 261.8 ;
      RECT  216.4 259.6 217.2 259.8 ;
      RECT  219.4 260.2 220.2 264.4 ;
      RECT  215.2 263.6 216.8 264.4 ;
      RECT  217.6 260.6 218.6 261.4 ;
      RECT  215.0 257.4 215.8 258.2 ;
      RECT  212.6 266.6 220.2 267.4 ;
      RECT  212.6 265.0 213.4 266.6 ;
      RECT  215.2 265.0 216.2 265.8 ;
      RECT  215.2 264.4 216.0 265.0 ;
      RECT  217.6 262.6 218.4 265.0 ;
      RECT  217.2 261.8 218.4 262.6 ;
      RECT  212.6 258.8 220.2 259.6 ;
      RECT  217.8 257.4 218.6 258.2 ;
      RECT  212.6 260.2 213.4 264.4 ;
      RECT  215.2 261.4 216.0 263.6 ;
      RECT  219.4 265.0 220.2 266.6 ;
      RECT  215.0 273.4 216.0 272.6 ;
      RECT  217.4 269.0 218.4 268.2 ;
      RECT  217.6 272.6 218.4 272.2 ;
      RECT  216.4 274.4 217.2 274.2 ;
      RECT  219.4 273.8 220.2 269.6 ;
      RECT  215.2 270.4 216.8 269.6 ;
      RECT  217.6 273.4 218.6 272.6 ;
      RECT  215.0 276.6 215.8 275.8 ;
      RECT  212.6 267.4 220.2 266.6 ;
      RECT  212.6 269.0 213.4 267.4 ;
      RECT  215.2 269.0 216.2 268.2 ;
      RECT  215.2 269.6 216.0 269.0 ;
      RECT  217.6 271.4 218.4 269.0 ;
      RECT  217.2 272.2 218.4 271.4 ;
      RECT  212.6 275.2 220.2 274.4 ;
      RECT  217.8 276.6 218.6 275.8 ;
      RECT  212.6 273.8 213.4 269.6 ;
      RECT  215.2 272.6 216.0 270.4 ;
      RECT  219.4 269.0 220.2 267.4 ;
      RECT  215.0 281.4 216.0 282.2 ;
      RECT  217.4 285.8 218.4 286.6 ;
      RECT  217.6 282.2 218.4 282.6 ;
      RECT  216.4 280.4 217.2 280.6 ;
      RECT  219.4 281.0 220.2 285.2 ;
      RECT  215.2 284.4 216.8 285.2 ;
      RECT  217.6 281.4 218.6 282.2 ;
      RECT  215.0 278.2 215.8 279.0 ;
      RECT  212.6 287.4 220.2 288.2 ;
      RECT  212.6 285.8 213.4 287.4 ;
      RECT  215.2 285.8 216.2 286.6 ;
      RECT  215.2 285.2 216.0 285.8 ;
      RECT  217.6 283.4 218.4 285.8 ;
      RECT  217.2 282.6 218.4 283.4 ;
      RECT  212.6 279.6 220.2 280.4 ;
      RECT  217.8 278.2 218.6 279.0 ;
      RECT  212.6 281.0 213.4 285.2 ;
      RECT  215.2 282.2 216.0 284.4 ;
      RECT  219.4 285.8 220.2 287.4 ;
      RECT  215.0 294.2 216.0 293.4 ;
      RECT  217.4 289.8 218.4 289.0 ;
      RECT  217.6 293.4 218.4 293.0 ;
      RECT  216.4 295.2 217.2 295.0 ;
      RECT  219.4 294.6 220.2 290.4 ;
      RECT  215.2 291.2 216.8 290.4 ;
      RECT  217.6 294.2 218.6 293.4 ;
      RECT  215.0 297.4 215.8 296.6 ;
      RECT  212.6 288.2 220.2 287.4 ;
      RECT  212.6 289.8 213.4 288.2 ;
      RECT  215.2 289.8 216.2 289.0 ;
      RECT  215.2 290.4 216.0 289.8 ;
      RECT  217.6 292.2 218.4 289.8 ;
      RECT  217.2 293.0 218.4 292.2 ;
      RECT  212.6 296.0 220.2 295.2 ;
      RECT  217.8 297.4 218.6 296.6 ;
      RECT  212.6 294.6 213.4 290.4 ;
      RECT  215.2 293.4 216.0 291.2 ;
      RECT  219.4 289.8 220.2 288.2 ;
      RECT  215.0 302.2 216.0 303.0 ;
      RECT  217.4 306.6 218.4 307.4 ;
      RECT  217.6 303.0 218.4 303.4 ;
      RECT  216.4 301.2 217.2 301.4 ;
      RECT  219.4 301.8 220.2 306.0 ;
      RECT  215.2 305.2 216.8 306.0 ;
      RECT  217.6 302.2 218.6 303.0 ;
      RECT  215.0 299.0 215.8 299.8 ;
      RECT  212.6 308.2 220.2 309.0 ;
      RECT  212.6 306.6 213.4 308.2 ;
      RECT  215.2 306.6 216.2 307.4 ;
      RECT  215.2 306.0 216.0 306.6 ;
      RECT  217.6 304.2 218.4 306.6 ;
      RECT  217.2 303.4 218.4 304.2 ;
      RECT  212.6 300.4 220.2 301.2 ;
      RECT  217.8 299.0 218.6 299.8 ;
      RECT  212.6 301.8 213.4 306.0 ;
      RECT  215.2 303.0 216.0 305.2 ;
      RECT  219.4 306.6 220.2 308.2 ;
      RECT  215.0 315.0 216.0 314.2 ;
      RECT  217.4 310.6 218.4 309.8 ;
      RECT  217.6 314.2 218.4 313.8 ;
      RECT  216.4 316.0 217.2 315.8 ;
      RECT  219.4 315.4 220.2 311.2 ;
      RECT  215.2 312.0 216.8 311.2 ;
      RECT  217.6 315.0 218.6 314.2 ;
      RECT  215.0 318.2 215.8 317.4 ;
      RECT  212.6 309.0 220.2 308.2 ;
      RECT  212.6 310.6 213.4 309.0 ;
      RECT  215.2 310.6 216.2 309.8 ;
      RECT  215.2 311.2 216.0 310.6 ;
      RECT  217.6 313.0 218.4 310.6 ;
      RECT  217.2 313.8 218.4 313.0 ;
      RECT  212.6 316.8 220.2 316.0 ;
      RECT  217.8 318.2 218.6 317.4 ;
      RECT  212.6 315.4 213.4 311.2 ;
      RECT  215.2 314.2 216.0 312.0 ;
      RECT  219.4 310.6 220.2 309.0 ;
      RECT  215.0 323.0 216.0 323.8 ;
      RECT  217.4 327.4 218.4 328.2 ;
      RECT  217.6 323.8 218.4 324.2 ;
      RECT  216.4 322.0 217.2 322.2 ;
      RECT  219.4 322.6 220.2 326.8 ;
      RECT  215.2 326.0 216.8 326.8 ;
      RECT  217.6 323.0 218.6 323.8 ;
      RECT  215.0 319.8 215.8 320.6 ;
      RECT  212.6 329.0 220.2 329.8 ;
      RECT  212.6 327.4 213.4 329.0 ;
      RECT  215.2 327.4 216.2 328.2 ;
      RECT  215.2 326.8 216.0 327.4 ;
      RECT  217.6 325.0 218.4 327.4 ;
      RECT  217.2 324.2 218.4 325.0 ;
      RECT  212.6 321.2 220.2 322.0 ;
      RECT  217.8 319.8 218.6 320.6 ;
      RECT  212.6 322.6 213.4 326.8 ;
      RECT  215.2 323.8 216.0 326.0 ;
      RECT  219.4 327.4 220.2 329.0 ;
      RECT  215.0 335.8 216.0 335.0 ;
      RECT  217.4 331.4 218.4 330.6 ;
      RECT  217.6 335.0 218.4 334.6 ;
      RECT  216.4 336.8 217.2 336.6 ;
      RECT  219.4 336.2 220.2 332.0 ;
      RECT  215.2 332.8 216.8 332.0 ;
      RECT  217.6 335.8 218.6 335.0 ;
      RECT  215.0 339.0 215.8 338.2 ;
      RECT  212.6 329.8 220.2 329.0 ;
      RECT  212.6 331.4 213.4 329.8 ;
      RECT  215.2 331.4 216.2 330.6 ;
      RECT  215.2 332.0 216.0 331.4 ;
      RECT  217.6 333.8 218.4 331.4 ;
      RECT  217.2 334.6 218.4 333.8 ;
      RECT  212.6 337.6 220.2 336.8 ;
      RECT  217.8 339.0 218.6 338.2 ;
      RECT  212.6 336.2 213.4 332.0 ;
      RECT  215.2 335.0 216.0 332.8 ;
      RECT  219.4 331.4 220.2 329.8 ;
      RECT  215.0 343.8 216.0 344.6 ;
      RECT  217.4 348.2 218.4 349.0 ;
      RECT  217.6 344.6 218.4 345.0 ;
      RECT  216.4 342.8 217.2 343.0 ;
      RECT  219.4 343.4 220.2 347.6 ;
      RECT  215.2 346.8 216.8 347.6 ;
      RECT  217.6 343.8 218.6 344.6 ;
      RECT  215.0 340.6 215.8 341.4 ;
      RECT  212.6 349.8 220.2 350.6 ;
      RECT  212.6 348.2 213.4 349.8 ;
      RECT  215.2 348.2 216.2 349.0 ;
      RECT  215.2 347.6 216.0 348.2 ;
      RECT  217.6 345.8 218.4 348.2 ;
      RECT  217.2 345.0 218.4 345.8 ;
      RECT  212.6 342.0 220.2 342.8 ;
      RECT  217.8 340.6 218.6 341.4 ;
      RECT  212.6 343.4 213.4 347.6 ;
      RECT  215.2 344.6 216.0 346.8 ;
      RECT  219.4 348.2 220.2 349.8 ;
      RECT  215.0 356.6 216.0 355.8 ;
      RECT  217.4 352.2 218.4 351.4 ;
      RECT  217.6 355.8 218.4 355.4 ;
      RECT  216.4 357.6 217.2 357.4 ;
      RECT  219.4 357.0 220.2 352.8 ;
      RECT  215.2 353.6 216.8 352.8 ;
      RECT  217.6 356.6 218.6 355.8 ;
      RECT  215.0 359.8 215.8 359.0 ;
      RECT  212.6 350.6 220.2 349.8 ;
      RECT  212.6 352.2 213.4 350.6 ;
      RECT  215.2 352.2 216.2 351.4 ;
      RECT  215.2 352.8 216.0 352.2 ;
      RECT  217.6 354.6 218.4 352.2 ;
      RECT  217.2 355.4 218.4 354.6 ;
      RECT  212.6 358.4 220.2 357.6 ;
      RECT  217.8 359.8 218.6 359.0 ;
      RECT  212.6 357.0 213.4 352.8 ;
      RECT  215.2 355.8 216.0 353.6 ;
      RECT  219.4 352.2 220.2 350.6 ;
      RECT  215.0 364.6 216.0 365.4 ;
      RECT  217.4 369.0 218.4 369.8 ;
      RECT  217.6 365.4 218.4 365.8 ;
      RECT  216.4 363.6 217.2 363.8 ;
      RECT  219.4 364.2 220.2 368.4 ;
      RECT  215.2 367.6 216.8 368.4 ;
      RECT  217.6 364.6 218.6 365.4 ;
      RECT  215.0 361.4 215.8 362.2 ;
      RECT  212.6 370.6 220.2 371.4 ;
      RECT  212.6 369.0 213.4 370.6 ;
      RECT  215.2 369.0 216.2 369.8 ;
      RECT  215.2 368.4 216.0 369.0 ;
      RECT  217.6 366.6 218.4 369.0 ;
      RECT  217.2 365.8 218.4 366.6 ;
      RECT  212.6 362.8 220.2 363.6 ;
      RECT  217.8 361.4 218.6 362.2 ;
      RECT  212.6 364.2 213.4 368.4 ;
      RECT  215.2 365.4 216.0 367.6 ;
      RECT  219.4 369.0 220.2 370.6 ;
      RECT  212.6 175.6 219.4 176.4 ;
      RECT  212.6 191.2 219.4 192.0 ;
      RECT  212.6 196.4 219.4 197.2 ;
      RECT  212.6 212.0 219.4 212.8 ;
      RECT  212.6 217.2 219.4 218.0 ;
      RECT  212.6 232.8 219.4 233.6 ;
      RECT  212.6 238.0 219.4 238.8 ;
      RECT  212.6 253.6 219.4 254.4 ;
      RECT  212.6 258.8 219.4 259.6 ;
      RECT  212.6 274.4 219.4 275.2 ;
      RECT  212.6 279.6 219.4 280.4 ;
      RECT  212.6 295.2 219.4 296.0 ;
      RECT  212.6 300.4 219.4 301.2 ;
      RECT  212.6 316.0 219.4 316.8 ;
      RECT  212.6 321.2 219.4 322.0 ;
      RECT  212.6 336.8 219.4 337.6 ;
      RECT  212.6 342.0 219.4 342.8 ;
      RECT  212.6 357.6 219.4 358.4 ;
      RECT  212.6 362.8 219.4 363.6 ;
      RECT  185.8 196.4 219.8 197.2 ;
      RECT  185.8 212.0 219.8 212.8 ;
      RECT  185.8 217.2 219.8 218.0 ;
      RECT  185.8 232.8 219.8 233.6 ;
      RECT  185.8 238.0 219.8 238.8 ;
      RECT  185.8 253.6 219.8 254.4 ;
      RECT  185.8 258.8 219.8 259.6 ;
      RECT  185.8 274.4 219.8 275.2 ;
      RECT  185.8 279.6 219.8 280.4 ;
      RECT  185.8 295.2 219.8 296.0 ;
      RECT  185.8 300.4 219.8 301.2 ;
      RECT  185.8 316.0 219.8 316.8 ;
      RECT  185.8 321.2 219.8 322.0 ;
      RECT  185.8 336.8 219.8 337.6 ;
      RECT  185.8 342.0 219.8 342.8 ;
      RECT  185.8 357.6 219.8 358.4 ;
      RECT  185.8 191.2 219.8 192.0 ;
      RECT  192.6 168.9 199.4 169.5 ;
      RECT  195.5 163.8 196.1 169.2 ;
      RECT  195.8 158.3 197.8 158.9 ;
      RECT  197.4 163.1 197.8 163.7 ;
      RECT  193.8 158.2 194.6 159.0 ;
      RECT  195.4 158.2 196.2 159.0 ;
      RECT  195.4 158.2 196.2 159.0 ;
      RECT  193.8 158.2 194.6 159.0 ;
      RECT  193.8 163.0 194.6 163.8 ;
      RECT  195.4 163.0 196.2 163.8 ;
      RECT  195.4 163.0 196.2 163.8 ;
      RECT  193.8 163.0 194.6 163.8 ;
      RECT  195.4 163.0 196.2 163.8 ;
      RECT  197.0 163.0 197.8 163.8 ;
      RECT  197.0 163.0 197.8 163.8 ;
      RECT  195.4 163.0 196.2 163.8 ;
      RECT  194.4 159.7 195.2 160.5 ;
      RECT  195.4 166.6 196.2 167.4 ;
      RECT  195.4 163.0 196.2 163.8 ;
      RECT  193.8 163.0 194.6 163.8 ;
      RECT  193.8 158.2 194.6 159.0 ;
      RECT  197.4 163.0 198.2 163.8 ;
      RECT  197.4 158.2 198.2 159.0 ;
      RECT  192.6 159.8 199.4 160.4 ;
      RECT  199.4 168.9 206.2 169.5 ;
      RECT  202.3 163.8 202.9 169.2 ;
      RECT  202.6 158.3 204.6 158.9 ;
      RECT  204.2 163.1 204.6 163.7 ;
      RECT  200.6 158.2 201.4 159.0 ;
      RECT  202.2 158.2 203.0 159.0 ;
      RECT  202.2 158.2 203.0 159.0 ;
      RECT  200.6 158.2 201.4 159.0 ;
      RECT  200.6 163.0 201.4 163.8 ;
      RECT  202.2 163.0 203.0 163.8 ;
      RECT  202.2 163.0 203.0 163.8 ;
      RECT  200.6 163.0 201.4 163.8 ;
      RECT  202.2 163.0 203.0 163.8 ;
      RECT  203.8 163.0 204.6 163.8 ;
      RECT  203.8 163.0 204.6 163.8 ;
      RECT  202.2 163.0 203.0 163.8 ;
      RECT  201.2 159.7 202.0 160.5 ;
      RECT  202.2 166.6 203.0 167.4 ;
      RECT  202.2 163.0 203.0 163.8 ;
      RECT  200.6 163.0 201.4 163.8 ;
      RECT  200.6 158.2 201.4 159.0 ;
      RECT  204.2 163.0 205.0 163.8 ;
      RECT  204.2 158.2 205.0 159.0 ;
      RECT  199.4 159.8 206.2 160.4 ;
      RECT  206.2 168.9 213.0 169.5 ;
      RECT  209.1 163.8 209.7 169.2 ;
      RECT  209.4 158.3 211.4 158.9 ;
      RECT  211.0 163.1 211.4 163.7 ;
      RECT  207.4 158.2 208.2 159.0 ;
      RECT  209.0 158.2 209.8 159.0 ;
      RECT  209.0 158.2 209.8 159.0 ;
      RECT  207.4 158.2 208.2 159.0 ;
      RECT  207.4 163.0 208.2 163.8 ;
      RECT  209.0 163.0 209.8 163.8 ;
      RECT  209.0 163.0 209.8 163.8 ;
      RECT  207.4 163.0 208.2 163.8 ;
      RECT  209.0 163.0 209.8 163.8 ;
      RECT  210.6 163.0 211.4 163.8 ;
      RECT  210.6 163.0 211.4 163.8 ;
      RECT  209.0 163.0 209.8 163.8 ;
      RECT  208.0 159.7 208.8 160.5 ;
      RECT  209.0 166.6 209.8 167.4 ;
      RECT  209.0 163.0 209.8 163.8 ;
      RECT  207.4 163.0 208.2 163.8 ;
      RECT  207.4 158.2 208.2 159.0 ;
      RECT  211.0 163.0 211.8 163.8 ;
      RECT  211.0 158.2 211.8 159.0 ;
      RECT  206.2 159.8 213.0 160.4 ;
      RECT  192.6 159.8 213.0 160.4 ;
      RECT  202.2 123.8 203.0 128.6 ;
      RECT  204.8 133.0 205.6 134.2 ;
      RECT  204.0 140.8 204.8 143.2 ;
      RECT  202.4 141.4 203.2 143.2 ;
      RECT  205.8 147.2 206.6 148.0 ;
      RECT  200.6 124.4 201.4 128.6 ;
      RECT  202.4 134.2 205.6 134.8 ;
      RECT  200.8 133.6 201.6 143.2 ;
      RECT  205.6 128.6 206.2 130.0 ;
      RECT  199.0 149.6 206.6 150.4 ;
      RECT  200.8 132.8 202.0 133.6 ;
      RECT  200.6 130.0 202.0 130.6 ;
      RECT  201.2 130.6 202.0 130.8 ;
      RECT  204.2 147.2 205.0 147.6 ;
      RECT  203.8 123.8 204.6 129.4 ;
      RECT  202.0 128.6 202.8 129.4 ;
      RECT  200.6 128.6 201.2 130.0 ;
      RECT  202.6 143.2 203.2 145.8 ;
      RECT  205.4 123.8 206.2 128.6 ;
      RECT  202.6 145.8 203.4 147.6 ;
      RECT  200.0 122.0 200.8 123.8 ;
      RECT  204.0 135.4 204.8 140.0 ;
      RECT  200.0 123.8 201.4 124.4 ;
      RECT  205.2 130.0 206.2 130.8 ;
      RECT  202.4 135.4 203.2 139.0 ;
      RECT  204.2 146.4 206.6 147.2 ;
      RECT  202.4 134.8 203.0 135.4 ;
      RECT  204.0 140.0 205.4 140.8 ;
      RECT  204.2 145.8 205.0 146.4 ;
      RECT  209.0 123.8 209.8 128.6 ;
      RECT  211.6 133.0 212.4 134.2 ;
      RECT  210.8 140.8 211.6 143.2 ;
      RECT  209.2 141.4 210.0 143.2 ;
      RECT  212.6 147.2 213.4 148.0 ;
      RECT  207.4 124.4 208.2 128.6 ;
      RECT  209.2 134.2 212.4 134.8 ;
      RECT  207.6 133.6 208.4 143.2 ;
      RECT  212.4 128.6 213.0 130.0 ;
      RECT  205.8 149.6 213.4 150.4 ;
      RECT  207.6 132.8 208.8 133.6 ;
      RECT  207.4 130.0 208.8 130.6 ;
      RECT  208.0 130.6 208.8 130.8 ;
      RECT  211.0 147.2 211.8 147.6 ;
      RECT  210.6 123.8 211.4 129.4 ;
      RECT  208.8 128.6 209.6 129.4 ;
      RECT  207.4 128.6 208.0 130.0 ;
      RECT  209.4 143.2 210.0 145.8 ;
      RECT  212.2 123.8 213.0 128.6 ;
      RECT  209.4 145.8 210.2 147.6 ;
      RECT  206.8 122.0 207.6 123.8 ;
      RECT  210.8 135.4 211.6 140.0 ;
      RECT  206.8 123.8 208.2 124.4 ;
      RECT  212.0 130.0 213.0 130.8 ;
      RECT  209.2 135.4 210.0 139.0 ;
      RECT  211.0 146.4 213.4 147.2 ;
      RECT  209.2 134.8 209.8 135.4 ;
      RECT  210.8 140.0 212.2 140.8 ;
      RECT  211.0 145.8 211.8 146.4 ;
      RECT  199.4 149.6 213.0 150.2 ;
      RECT  200.4 91.4 201.2 95.2 ;
      RECT  203.6 94.2 204.8 95.0 ;
      RECT  200.0 79.8 205.6 80.6 ;
      RECT  200.4 113.6 202.2 114.4 ;
      RECT  200.0 82.0 200.8 84.0 ;
      RECT  203.4 100.0 204.2 102.6 ;
      RECT  202.0 96.4 202.8 98.6 ;
      RECT  200.0 81.2 204.0 82.0 ;
      RECT  202.0 91.4 202.8 92.8 ;
      RECT  200.4 95.8 201.2 97.8 ;
      RECT  201.6 82.6 202.4 84.6 ;
      RECT  200.0 85.2 200.8 87.8 ;
      RECT  203.4 103.4 204.2 104.6 ;
      RECT  200.2 100.0 201.0 108.6 ;
      RECT  200.4 95.2 204.4 95.8 ;
      RECT  201.8 98.6 203.4 99.4 ;
      RECT  203.2 82.0 204.0 84.0 ;
      RECT  203.6 95.8 204.4 97.8 ;
      RECT  201.6 86.4 202.4 87.8 ;
      RECT  203.6 95.0 204.4 95.2 ;
      RECT  203.4 110.6 204.2 113.8 ;
      RECT  201.8 99.4 202.6 101.4 ;
      RECT  203.4 102.6 206.0 103.4 ;
      RECT  200.0 89.2 200.8 90.0 ;
      RECT  204.4 92.8 205.4 93.0 ;
      RECT  200.4 113.0 201.0 113.6 ;
      RECT  201.8 103.8 202.6 113.0 ;
      RECT  200.2 110.6 201.0 113.0 ;
      RECT  200.0 84.6 202.4 85.2 ;
      RECT  205.0 111.4 206.0 112.2 ;
      RECT  200.2 87.8 200.8 89.2 ;
      RECT  202.4 76.2 203.2 77.8 ;
      RECT  203.2 86.4 204.0 88.6 ;
      RECT  205.4 103.4 206.0 111.4 ;
      RECT  204.0 90.0 205.6 90.8 ;
      RECT  203.6 91.4 205.4 92.8 ;
      RECT  204.8 82.6 205.6 90.0 ;
      RECT  207.2 91.4 208.0 95.2 ;
      RECT  210.4 94.2 211.6 95.0 ;
      RECT  206.8 79.8 212.4 80.6 ;
      RECT  207.2 113.6 209.0 114.4 ;
      RECT  206.8 82.0 207.6 84.0 ;
      RECT  210.2 100.0 211.0 102.6 ;
      RECT  208.8 96.4 209.6 98.6 ;
      RECT  206.8 81.2 210.8 82.0 ;
      RECT  208.8 91.4 209.6 92.8 ;
      RECT  207.2 95.8 208.0 97.8 ;
      RECT  208.4 82.6 209.2 84.6 ;
      RECT  206.8 85.2 207.6 87.8 ;
      RECT  210.2 103.4 211.0 104.6 ;
      RECT  207.0 100.0 207.8 108.6 ;
      RECT  207.2 95.2 211.2 95.8 ;
      RECT  208.6 98.6 210.2 99.4 ;
      RECT  210.0 82.0 210.8 84.0 ;
      RECT  210.4 95.8 211.2 97.8 ;
      RECT  208.4 86.4 209.2 87.8 ;
      RECT  210.4 95.0 211.2 95.2 ;
      RECT  210.2 110.6 211.0 113.8 ;
      RECT  208.6 99.4 209.4 101.4 ;
      RECT  210.2 102.6 212.8 103.4 ;
      RECT  206.8 89.2 207.6 90.0 ;
      RECT  211.2 92.8 212.2 93.0 ;
      RECT  207.2 113.0 207.8 113.6 ;
      RECT  208.6 103.8 209.4 113.0 ;
      RECT  207.0 110.6 207.8 113.0 ;
      RECT  206.8 84.6 209.2 85.2 ;
      RECT  211.8 111.4 212.8 112.2 ;
      RECT  207.0 87.8 207.6 89.2 ;
      RECT  209.2 76.2 210.0 77.8 ;
      RECT  210.0 86.4 210.8 88.6 ;
      RECT  212.2 103.4 212.8 111.4 ;
      RECT  210.8 90.0 212.4 90.8 ;
      RECT  210.4 91.4 212.2 92.8 ;
      RECT  211.6 82.6 212.4 90.0 ;
      RECT  199.4 79.8 213.0 80.4 ;
      RECT  199.4 150.2 213.0 149.6 ;
      RECT  192.6 160.4 213.0 159.8 ;
      RECT  199.4 80.4 213.0 79.8 ;
      RECT  156.9 199.3 157.5 199.9 ;
      RECT  156.9 197.1 157.5 197.7 ;
      RECT  154.7 199.3 157.2 199.9 ;
      RECT  156.9 197.4 157.5 199.6 ;
      RECT  157.2 197.1 159.7 197.7 ;
      RECT  156.9 210.1 157.5 210.7 ;
      RECT  156.9 212.3 157.5 212.9 ;
      RECT  154.7 210.1 157.2 210.7 ;
      RECT  156.9 210.4 157.5 212.6 ;
      RECT  157.2 212.3 159.7 212.9 ;
      RECT  156.9 220.1 157.5 220.7 ;
      RECT  156.9 217.9 157.5 218.5 ;
      RECT  154.7 220.1 157.2 220.7 ;
      RECT  156.9 218.2 157.5 220.4 ;
      RECT  157.2 217.9 159.7 218.5 ;
      RECT  156.9 230.9 157.5 231.5 ;
      RECT  156.9 233.1 157.5 233.7 ;
      RECT  154.7 230.9 157.2 231.5 ;
      RECT  156.9 231.2 157.5 233.4 ;
      RECT  157.2 233.1 159.7 233.7 ;
      RECT  156.9 240.9 157.5 241.5 ;
      RECT  156.9 238.7 157.5 239.3 ;
      RECT  154.7 240.9 157.2 241.5 ;
      RECT  156.9 239.0 157.5 241.2 ;
      RECT  157.2 238.7 159.7 239.3 ;
      RECT  156.9 251.7 157.5 252.3 ;
      RECT  156.9 253.9 157.5 254.5 ;
      RECT  154.7 251.7 157.2 252.3 ;
      RECT  156.9 252.0 157.5 254.2 ;
      RECT  157.2 253.9 159.7 254.5 ;
      RECT  156.9 261.7 157.5 262.3 ;
      RECT  156.9 259.5 157.5 260.1 ;
      RECT  154.7 261.7 157.2 262.3 ;
      RECT  156.9 259.8 157.5 262.0 ;
      RECT  157.2 259.5 159.7 260.1 ;
      RECT  156.9 272.5 157.5 273.1 ;
      RECT  156.9 274.7 157.5 275.3 ;
      RECT  154.7 272.5 157.2 273.1 ;
      RECT  156.9 272.8 157.5 275.0 ;
      RECT  157.2 274.7 159.7 275.3 ;
      RECT  156.9 282.5 157.5 283.1 ;
      RECT  156.9 280.3 157.5 280.9 ;
      RECT  154.7 282.5 157.2 283.1 ;
      RECT  156.9 280.6 157.5 282.8 ;
      RECT  157.2 280.3 159.7 280.9 ;
      RECT  156.9 293.3 157.5 293.9 ;
      RECT  156.9 295.5 157.5 296.1 ;
      RECT  154.7 293.3 157.2 293.9 ;
      RECT  156.9 293.6 157.5 295.8 ;
      RECT  157.2 295.5 159.7 296.1 ;
      RECT  156.9 303.3 157.5 303.9 ;
      RECT  156.9 301.1 157.5 301.7 ;
      RECT  154.7 303.3 157.2 303.9 ;
      RECT  156.9 301.4 157.5 303.6 ;
      RECT  157.2 301.1 159.7 301.7 ;
      RECT  156.9 314.1 157.5 314.7 ;
      RECT  156.9 316.3 157.5 316.9 ;
      RECT  154.7 314.1 157.2 314.7 ;
      RECT  156.9 314.4 157.5 316.6 ;
      RECT  157.2 316.3 159.7 316.9 ;
      RECT  156.9 324.1 157.5 324.7 ;
      RECT  156.9 321.9 157.5 322.5 ;
      RECT  154.7 324.1 157.2 324.7 ;
      RECT  156.9 322.2 157.5 324.4 ;
      RECT  157.2 321.9 159.7 322.5 ;
      RECT  156.9 334.9 157.5 335.5 ;
      RECT  156.9 337.1 157.5 337.7 ;
      RECT  154.7 334.9 157.2 335.5 ;
      RECT  156.9 335.2 157.5 337.4 ;
      RECT  157.2 337.1 159.7 337.7 ;
      RECT  156.9 344.9 157.5 345.5 ;
      RECT  156.9 342.7 157.5 343.3 ;
      RECT  154.7 344.9 157.2 345.5 ;
      RECT  156.9 343.0 157.5 345.2 ;
      RECT  157.2 342.7 159.7 343.3 ;
      RECT  156.9 355.7 157.5 356.3 ;
      RECT  156.9 357.9 157.5 358.5 ;
      RECT  154.7 355.7 157.2 356.3 ;
      RECT  156.9 356.0 157.5 358.2 ;
      RECT  157.2 357.9 159.7 358.5 ;
      RECT  149.8 199.1 150.4 199.7 ;
      RECT  149.8 199.3 150.4 199.9 ;
      RECT  147.9 199.1 150.1 199.7 ;
      RECT  149.8 199.4 150.4 199.6 ;
      RECT  150.1 199.3 152.3 199.9 ;
      RECT  149.8 210.3 150.4 210.9 ;
      RECT  149.8 210.1 150.4 210.7 ;
      RECT  147.9 210.3 150.1 210.9 ;
      RECT  149.8 210.4 150.4 210.6 ;
      RECT  150.1 210.1 152.3 210.7 ;
      RECT  149.8 219.9 150.4 220.5 ;
      RECT  149.8 220.1 150.4 220.7 ;
      RECT  147.9 219.9 150.1 220.5 ;
      RECT  149.8 220.2 150.4 220.4 ;
      RECT  150.1 220.1 152.3 220.7 ;
      RECT  149.8 231.1 150.4 231.7 ;
      RECT  149.8 230.9 150.4 231.5 ;
      RECT  147.9 231.1 150.1 231.7 ;
      RECT  149.8 231.2 150.4 231.4 ;
      RECT  150.1 230.9 152.3 231.5 ;
      RECT  149.8 240.7 150.4 241.3 ;
      RECT  149.8 240.9 150.4 241.5 ;
      RECT  147.9 240.7 150.1 241.3 ;
      RECT  149.8 241.0 150.4 241.2 ;
      RECT  150.1 240.9 152.3 241.5 ;
      RECT  149.8 251.9 150.4 252.5 ;
      RECT  149.8 251.7 150.4 252.3 ;
      RECT  147.9 251.9 150.1 252.5 ;
      RECT  149.8 252.0 150.4 252.2 ;
      RECT  150.1 251.7 152.3 252.3 ;
      RECT  149.8 261.5 150.4 262.1 ;
      RECT  149.8 261.7 150.4 262.3 ;
      RECT  147.9 261.5 150.1 262.1 ;
      RECT  149.8 261.8 150.4 262.0 ;
      RECT  150.1 261.7 152.3 262.3 ;
      RECT  149.8 272.7 150.4 273.3 ;
      RECT  149.8 272.5 150.4 273.1 ;
      RECT  147.9 272.7 150.1 273.3 ;
      RECT  149.8 272.8 150.4 273.0 ;
      RECT  150.1 272.5 152.3 273.1 ;
      RECT  149.8 282.3 150.4 282.9 ;
      RECT  149.8 282.5 150.4 283.1 ;
      RECT  147.9 282.3 150.1 282.9 ;
      RECT  149.8 282.6 150.4 282.8 ;
      RECT  150.1 282.5 152.3 283.1 ;
      RECT  149.8 293.5 150.4 294.1 ;
      RECT  149.8 293.3 150.4 293.9 ;
      RECT  147.9 293.5 150.1 294.1 ;
      RECT  149.8 293.6 150.4 293.8 ;
      RECT  150.1 293.3 152.3 293.9 ;
      RECT  149.8 303.1 150.4 303.7 ;
      RECT  149.8 303.3 150.4 303.9 ;
      RECT  147.9 303.1 150.1 303.7 ;
      RECT  149.8 303.4 150.4 303.6 ;
      RECT  150.1 303.3 152.3 303.9 ;
      RECT  149.8 314.3 150.4 314.9 ;
      RECT  149.8 314.1 150.4 314.7 ;
      RECT  147.9 314.3 150.1 314.9 ;
      RECT  149.8 314.4 150.4 314.6 ;
      RECT  150.1 314.1 152.3 314.7 ;
      RECT  149.8 323.9 150.4 324.5 ;
      RECT  149.8 324.1 150.4 324.7 ;
      RECT  147.9 323.9 150.1 324.5 ;
      RECT  149.8 324.2 150.4 324.4 ;
      RECT  150.1 324.1 152.3 324.7 ;
      RECT  149.8 335.1 150.4 335.7 ;
      RECT  149.8 334.9 150.4 335.5 ;
      RECT  147.9 335.1 150.1 335.7 ;
      RECT  149.8 335.2 150.4 335.4 ;
      RECT  150.1 334.9 152.3 335.5 ;
      RECT  149.8 344.7 150.4 345.3 ;
      RECT  149.8 344.9 150.4 345.5 ;
      RECT  147.9 344.7 150.1 345.3 ;
      RECT  149.8 345.0 150.4 345.2 ;
      RECT  150.1 344.9 152.3 345.5 ;
      RECT  149.8 355.9 150.4 356.5 ;
      RECT  149.8 355.7 150.4 356.3 ;
      RECT  147.9 355.9 150.1 356.5 ;
      RECT  149.8 356.0 150.4 356.2 ;
      RECT  150.1 355.7 152.3 356.3 ;
      RECT  130.7 199.1 142.9 199.7 ;
      RECT  136.3 197.7 144.9 198.3 ;
      RECT  132.1 210.3 142.9 210.9 ;
      RECT  136.3 211.7 144.9 212.3 ;
      RECT  133.5 219.9 142.9 220.5 ;
      RECT  136.3 218.5 144.9 219.1 ;
      RECT  134.9 231.1 142.9 231.7 ;
      RECT  136.3 232.5 144.9 233.1 ;
      RECT  130.7 240.7 142.9 241.3 ;
      RECT  137.7 239.3 144.9 239.9 ;
      RECT  132.1 251.9 142.9 252.5 ;
      RECT  137.7 253.3 144.9 253.9 ;
      RECT  133.5 261.5 142.9 262.1 ;
      RECT  137.7 260.1 144.9 260.7 ;
      RECT  134.9 272.7 142.9 273.3 ;
      RECT  137.7 274.1 144.9 274.7 ;
      RECT  130.7 282.3 142.9 282.9 ;
      RECT  139.1 280.9 144.9 281.5 ;
      RECT  132.1 293.5 142.9 294.1 ;
      RECT  139.1 294.9 144.9 295.5 ;
      RECT  133.5 303.1 142.9 303.7 ;
      RECT  139.1 301.7 144.9 302.3 ;
      RECT  134.9 314.3 142.9 314.9 ;
      RECT  139.1 315.7 144.9 316.3 ;
      RECT  130.7 323.9 142.9 324.5 ;
      RECT  140.5 322.5 144.9 323.1 ;
      RECT  132.1 335.1 142.9 335.7 ;
      RECT  140.5 336.5 144.9 337.1 ;
      RECT  133.5 344.7 142.9 345.3 ;
      RECT  140.5 343.3 144.9 343.9 ;
      RECT  134.9 355.9 142.9 356.5 ;
      RECT  140.5 357.3 144.9 357.9 ;
      RECT  141.3 204.7 157.3 205.3 ;
      RECT  141.3 194.3 157.3 194.9 ;
      RECT  141.3 225.5 157.3 226.1 ;
      RECT  141.3 215.1 157.3 215.7 ;
      RECT  141.3 246.3 157.3 246.9 ;
      RECT  141.3 235.9 157.3 236.5 ;
      RECT  141.3 267.1 157.3 267.7 ;
      RECT  141.3 256.7 157.3 257.3 ;
      RECT  141.3 287.9 157.3 288.5 ;
      RECT  141.3 277.5 157.3 278.1 ;
      RECT  141.3 308.7 157.3 309.3 ;
      RECT  141.3 298.3 157.3 298.9 ;
      RECT  141.3 329.5 157.3 330.1 ;
      RECT  141.3 319.1 157.3 319.7 ;
      RECT  141.3 350.3 157.3 350.9 ;
      RECT  141.3 339.9 157.3 340.5 ;
      RECT  106.0 199.3 106.6 199.9 ;
      RECT  106.0 202.9 106.6 203.5 ;
      RECT  103.1 199.3 106.3 199.9 ;
      RECT  106.0 199.6 106.6 203.2 ;
      RECT  106.3 202.9 108.8 203.5 ;
      RECT  97.1 199.3 100.7 199.9 ;
      RECT  106.0 210.1 106.6 210.7 ;
      RECT  106.0 213.3 106.6 213.9 ;
      RECT  103.1 210.1 106.3 210.7 ;
      RECT  106.0 210.4 106.6 213.6 ;
      RECT  106.3 213.3 110.2 213.9 ;
      RECT  98.5 210.1 100.7 210.7 ;
      RECT  97.1 216.5 111.6 217.1 ;
      RECT  98.5 226.9 113.0 227.5 ;
      RECT  108.8 199.1 115.7 199.7 ;
      RECT  110.2 197.7 117.7 198.3 ;
      RECT  111.6 210.3 115.7 210.9 ;
      RECT  110.2 211.7 117.7 212.3 ;
      RECT  108.8 219.9 115.7 220.5 ;
      RECT  113.0 218.5 117.7 219.1 ;
      RECT  111.6 231.1 115.7 231.7 ;
      RECT  113.0 232.5 117.7 233.1 ;
      RECT  122.6 199.1 123.2 199.7 ;
      RECT  122.6 199.3 123.2 199.9 ;
      RECT  120.7 199.1 122.9 199.7 ;
      RECT  122.6 199.4 123.2 199.6 ;
      RECT  122.9 199.3 125.1 199.9 ;
      RECT  122.6 210.3 123.2 210.9 ;
      RECT  122.6 210.1 123.2 210.7 ;
      RECT  120.7 210.3 122.9 210.9 ;
      RECT  122.6 210.4 123.2 210.6 ;
      RECT  122.9 210.1 125.1 210.7 ;
      RECT  122.6 219.9 123.2 220.5 ;
      RECT  122.6 220.1 123.2 220.7 ;
      RECT  120.7 219.9 122.9 220.5 ;
      RECT  122.6 220.2 123.2 220.4 ;
      RECT  122.9 220.1 125.1 220.7 ;
      RECT  122.6 231.1 123.2 231.7 ;
      RECT  122.6 230.9 123.2 231.5 ;
      RECT  120.7 231.1 122.9 231.7 ;
      RECT  122.6 231.2 123.2 231.4 ;
      RECT  122.9 230.9 125.1 231.5 ;
      RECT  96.5 204.7 130.1 205.3 ;
      RECT  96.5 194.3 130.1 194.9 ;
      RECT  96.5 204.7 130.1 205.3 ;
      RECT  96.5 215.1 130.1 215.7 ;
      RECT  96.5 225.5 130.1 226.1 ;
      RECT  96.5 215.1 130.1 215.7 ;
      RECT  96.5 225.5 130.1 226.1 ;
      RECT  96.5 235.9 130.1 236.5 ;
      RECT  103.7 203.7 104.5 205.0 ;
      RECT  103.7 194.6 104.5 195.9 ;
      RECT  100.5 195.5 101.3 194.3 ;
      RECT  100.5 202.9 101.3 205.3 ;
      RECT  102.2 195.5 102.8 203.7 ;
      RECT  100.5 202.9 101.3 203.7 ;
      RECT  102.1 202.9 102.9 203.7 ;
      RECT  102.1 202.9 102.9 203.7 ;
      RECT  100.5 202.9 101.3 203.7 ;
      RECT  100.5 195.5 101.3 196.3 ;
      RECT  102.1 195.5 102.9 196.3 ;
      RECT  102.1 195.5 102.9 196.3 ;
      RECT  100.5 195.5 101.3 196.3 ;
      RECT  103.7 203.3 104.5 204.1 ;
      RECT  103.7 195.5 104.5 196.3 ;
      RECT  100.7 199.2 101.5 200.0 ;
      RECT  100.7 199.2 101.5 200.0 ;
      RECT  102.5 199.3 103.1 199.9 ;
      RECT  99.3 204.7 105.7 205.3 ;
      RECT  99.3 194.3 105.7 194.9 ;
      RECT  103.7 206.3 104.5 205.0 ;
      RECT  103.7 215.4 104.5 214.1 ;
      RECT  100.5 214.5 101.3 215.7 ;
      RECT  100.5 207.1 101.3 204.7 ;
      RECT  102.2 214.5 102.8 206.3 ;
      RECT  100.5 207.1 101.3 206.3 ;
      RECT  102.1 207.1 102.9 206.3 ;
      RECT  102.1 207.1 102.9 206.3 ;
      RECT  100.5 207.1 101.3 206.3 ;
      RECT  100.5 214.5 101.3 213.7 ;
      RECT  102.1 214.5 102.9 213.7 ;
      RECT  102.1 214.5 102.9 213.7 ;
      RECT  100.5 214.5 101.3 213.7 ;
      RECT  103.7 206.7 104.5 205.9 ;
      RECT  103.7 214.5 104.5 213.7 ;
      RECT  100.7 210.8 101.5 210.0 ;
      RECT  100.7 210.8 101.5 210.0 ;
      RECT  102.5 210.7 103.1 210.1 ;
      RECT  99.3 205.3 105.7 204.7 ;
      RECT  99.3 215.7 105.7 215.1 ;
      RECT  128.1 203.7 128.9 205.0 ;
      RECT  128.1 194.6 128.9 195.9 ;
      RECT  124.9 195.5 125.7 194.3 ;
      RECT  124.9 202.9 125.7 205.3 ;
      RECT  126.6 195.5 127.2 203.7 ;
      RECT  124.9 202.9 125.7 203.7 ;
      RECT  126.5 202.9 127.3 203.7 ;
      RECT  126.5 202.9 127.3 203.7 ;
      RECT  124.9 202.9 125.7 203.7 ;
      RECT  124.9 195.5 125.7 196.3 ;
      RECT  126.5 195.5 127.3 196.3 ;
      RECT  126.5 195.5 127.3 196.3 ;
      RECT  124.9 195.5 125.7 196.3 ;
      RECT  128.1 203.3 128.9 204.1 ;
      RECT  128.1 195.5 128.9 196.3 ;
      RECT  125.1 199.2 125.9 200.0 ;
      RECT  125.1 199.2 125.9 200.0 ;
      RECT  126.9 199.3 127.5 199.9 ;
      RECT  123.7 204.7 130.1 205.3 ;
      RECT  123.7 194.3 130.1 194.9 ;
      RECT  128.1 206.3 128.9 205.0 ;
      RECT  128.1 215.4 128.9 214.1 ;
      RECT  124.9 214.5 125.7 215.7 ;
      RECT  124.9 207.1 125.7 204.7 ;
      RECT  126.6 214.5 127.2 206.3 ;
      RECT  124.9 207.1 125.7 206.3 ;
      RECT  126.5 207.1 127.3 206.3 ;
      RECT  126.5 207.1 127.3 206.3 ;
      RECT  124.9 207.1 125.7 206.3 ;
      RECT  124.9 214.5 125.7 213.7 ;
      RECT  126.5 214.5 127.3 213.7 ;
      RECT  126.5 214.5 127.3 213.7 ;
      RECT  124.9 214.5 125.7 213.7 ;
      RECT  128.1 206.7 128.9 205.9 ;
      RECT  128.1 214.5 128.9 213.7 ;
      RECT  125.1 210.8 125.9 210.0 ;
      RECT  125.1 210.8 125.9 210.0 ;
      RECT  126.9 210.7 127.5 210.1 ;
      RECT  123.7 205.3 130.1 204.7 ;
      RECT  123.7 215.7 130.1 215.1 ;
      RECT  128.1 224.5 128.9 225.8 ;
      RECT  128.1 215.4 128.9 216.7 ;
      RECT  124.9 216.3 125.7 215.1 ;
      RECT  124.9 223.7 125.7 226.1 ;
      RECT  126.6 216.3 127.2 224.5 ;
      RECT  124.9 223.7 125.7 224.5 ;
      RECT  126.5 223.7 127.3 224.5 ;
      RECT  126.5 223.7 127.3 224.5 ;
      RECT  124.9 223.7 125.7 224.5 ;
      RECT  124.9 216.3 125.7 217.1 ;
      RECT  126.5 216.3 127.3 217.1 ;
      RECT  126.5 216.3 127.3 217.1 ;
      RECT  124.9 216.3 125.7 217.1 ;
      RECT  128.1 224.1 128.9 224.9 ;
      RECT  128.1 216.3 128.9 217.1 ;
      RECT  125.1 220.0 125.9 220.8 ;
      RECT  125.1 220.0 125.9 220.8 ;
      RECT  126.9 220.1 127.5 220.7 ;
      RECT  123.7 225.5 130.1 226.1 ;
      RECT  123.7 215.1 130.1 215.7 ;
      RECT  128.1 227.1 128.9 225.8 ;
      RECT  128.1 236.2 128.9 234.9 ;
      RECT  124.9 235.3 125.7 236.5 ;
      RECT  124.9 227.9 125.7 225.5 ;
      RECT  126.6 235.3 127.2 227.1 ;
      RECT  124.9 227.9 125.7 227.1 ;
      RECT  126.5 227.9 127.3 227.1 ;
      RECT  126.5 227.9 127.3 227.1 ;
      RECT  124.9 227.9 125.7 227.1 ;
      RECT  124.9 235.3 125.7 234.5 ;
      RECT  126.5 235.3 127.3 234.5 ;
      RECT  126.5 235.3 127.3 234.5 ;
      RECT  124.9 235.3 125.7 234.5 ;
      RECT  128.1 227.5 128.9 226.7 ;
      RECT  128.1 235.3 128.9 234.5 ;
      RECT  125.1 231.6 125.9 230.8 ;
      RECT  125.1 231.6 125.9 230.8 ;
      RECT  126.9 231.5 127.5 230.9 ;
      RECT  123.7 226.1 130.1 225.5 ;
      RECT  123.7 236.5 130.1 235.9 ;
      RECT  115.3 195.9 116.1 194.3 ;
      RECT  115.3 202.9 116.1 205.3 ;
      RECT  118.5 202.9 119.3 205.3 ;
      RECT  120.1 203.7 120.9 205.0 ;
      RECT  120.1 194.6 120.9 195.9 ;
      RECT  115.3 202.9 116.1 203.7 ;
      RECT  116.9 202.9 117.7 203.7 ;
      RECT  116.9 202.9 117.7 203.7 ;
      RECT  115.3 202.9 116.1 203.7 ;
      RECT  116.9 202.9 117.7 203.7 ;
      RECT  118.5 202.9 119.3 203.7 ;
      RECT  118.5 202.9 119.3 203.7 ;
      RECT  116.9 202.9 117.7 203.7 ;
      RECT  115.3 195.9 116.1 196.7 ;
      RECT  116.9 195.9 117.7 196.7 ;
      RECT  116.9 195.9 117.7 196.7 ;
      RECT  115.3 195.9 116.1 196.7 ;
      RECT  116.9 195.9 117.7 196.7 ;
      RECT  118.5 195.9 119.3 196.7 ;
      RECT  118.5 195.9 119.3 196.7 ;
      RECT  116.9 195.9 117.7 196.7 ;
      RECT  120.1 203.3 120.9 204.1 ;
      RECT  120.1 195.5 120.9 196.3 ;
      RECT  117.7 197.6 118.5 198.4 ;
      RECT  115.7 199.0 116.5 199.8 ;
      RECT  116.9 202.9 117.7 203.7 ;
      RECT  118.5 195.9 119.3 196.7 ;
      RECT  119.9 199.0 120.7 199.8 ;
      RECT  115.7 199.0 116.5 199.8 ;
      RECT  117.7 197.6 118.5 198.4 ;
      RECT  119.9 199.0 120.7 199.8 ;
      RECT  114.1 204.7 123.7 205.3 ;
      RECT  114.1 194.3 123.7 194.9 ;
      RECT  115.3 214.1 116.1 215.7 ;
      RECT  115.3 207.1 116.1 204.7 ;
      RECT  118.5 207.1 119.3 204.7 ;
      RECT  120.1 206.3 120.9 205.0 ;
      RECT  120.1 215.4 120.9 214.1 ;
      RECT  115.3 207.1 116.1 206.3 ;
      RECT  116.9 207.1 117.7 206.3 ;
      RECT  116.9 207.1 117.7 206.3 ;
      RECT  115.3 207.1 116.1 206.3 ;
      RECT  116.9 207.1 117.7 206.3 ;
      RECT  118.5 207.1 119.3 206.3 ;
      RECT  118.5 207.1 119.3 206.3 ;
      RECT  116.9 207.1 117.7 206.3 ;
      RECT  115.3 214.1 116.1 213.3 ;
      RECT  116.9 214.1 117.7 213.3 ;
      RECT  116.9 214.1 117.7 213.3 ;
      RECT  115.3 214.1 116.1 213.3 ;
      RECT  116.9 214.1 117.7 213.3 ;
      RECT  118.5 214.1 119.3 213.3 ;
      RECT  118.5 214.1 119.3 213.3 ;
      RECT  116.9 214.1 117.7 213.3 ;
      RECT  120.1 206.7 120.9 205.9 ;
      RECT  120.1 214.5 120.9 213.7 ;
      RECT  117.7 212.4 118.5 211.6 ;
      RECT  115.7 211.0 116.5 210.2 ;
      RECT  116.9 207.1 117.7 206.3 ;
      RECT  118.5 214.1 119.3 213.3 ;
      RECT  119.9 211.0 120.7 210.2 ;
      RECT  115.7 211.0 116.5 210.2 ;
      RECT  117.7 212.4 118.5 211.6 ;
      RECT  119.9 211.0 120.7 210.2 ;
      RECT  114.1 205.3 123.7 204.7 ;
      RECT  114.1 215.7 123.7 215.1 ;
      RECT  115.3 216.7 116.1 215.1 ;
      RECT  115.3 223.7 116.1 226.1 ;
      RECT  118.5 223.7 119.3 226.1 ;
      RECT  120.1 224.5 120.9 225.8 ;
      RECT  120.1 215.4 120.9 216.7 ;
      RECT  115.3 223.7 116.1 224.5 ;
      RECT  116.9 223.7 117.7 224.5 ;
      RECT  116.9 223.7 117.7 224.5 ;
      RECT  115.3 223.7 116.1 224.5 ;
      RECT  116.9 223.7 117.7 224.5 ;
      RECT  118.5 223.7 119.3 224.5 ;
      RECT  118.5 223.7 119.3 224.5 ;
      RECT  116.9 223.7 117.7 224.5 ;
      RECT  115.3 216.7 116.1 217.5 ;
      RECT  116.9 216.7 117.7 217.5 ;
      RECT  116.9 216.7 117.7 217.5 ;
      RECT  115.3 216.7 116.1 217.5 ;
      RECT  116.9 216.7 117.7 217.5 ;
      RECT  118.5 216.7 119.3 217.5 ;
      RECT  118.5 216.7 119.3 217.5 ;
      RECT  116.9 216.7 117.7 217.5 ;
      RECT  120.1 224.1 120.9 224.9 ;
      RECT  120.1 216.3 120.9 217.1 ;
      RECT  117.7 218.4 118.5 219.2 ;
      RECT  115.7 219.8 116.5 220.6 ;
      RECT  116.9 223.7 117.7 224.5 ;
      RECT  118.5 216.7 119.3 217.5 ;
      RECT  119.9 219.8 120.7 220.6 ;
      RECT  115.7 219.8 116.5 220.6 ;
      RECT  117.7 218.4 118.5 219.2 ;
      RECT  119.9 219.8 120.7 220.6 ;
      RECT  114.1 225.5 123.7 226.1 ;
      RECT  114.1 215.1 123.7 215.7 ;
      RECT  115.3 234.9 116.1 236.5 ;
      RECT  115.3 227.9 116.1 225.5 ;
      RECT  118.5 227.9 119.3 225.5 ;
      RECT  120.1 227.1 120.9 225.8 ;
      RECT  120.1 236.2 120.9 234.9 ;
      RECT  115.3 227.9 116.1 227.1 ;
      RECT  116.9 227.9 117.7 227.1 ;
      RECT  116.9 227.9 117.7 227.1 ;
      RECT  115.3 227.9 116.1 227.1 ;
      RECT  116.9 227.9 117.7 227.1 ;
      RECT  118.5 227.9 119.3 227.1 ;
      RECT  118.5 227.9 119.3 227.1 ;
      RECT  116.9 227.9 117.7 227.1 ;
      RECT  115.3 234.9 116.1 234.1 ;
      RECT  116.9 234.9 117.7 234.1 ;
      RECT  116.9 234.9 117.7 234.1 ;
      RECT  115.3 234.9 116.1 234.1 ;
      RECT  116.9 234.9 117.7 234.1 ;
      RECT  118.5 234.9 119.3 234.1 ;
      RECT  118.5 234.9 119.3 234.1 ;
      RECT  116.9 234.9 117.7 234.1 ;
      RECT  120.1 227.5 120.9 226.7 ;
      RECT  120.1 235.3 120.9 234.5 ;
      RECT  117.7 233.2 118.5 232.4 ;
      RECT  115.7 231.8 116.5 231.0 ;
      RECT  116.9 227.9 117.7 227.1 ;
      RECT  118.5 234.9 119.3 234.1 ;
      RECT  119.9 231.8 120.7 231.0 ;
      RECT  115.7 231.8 116.5 231.0 ;
      RECT  117.7 233.2 118.5 232.4 ;
      RECT  119.9 231.8 120.7 231.0 ;
      RECT  114.1 226.1 123.7 225.5 ;
      RECT  114.1 236.5 123.7 235.9 ;
      RECT  108.4 202.8 109.2 203.6 ;
      RECT  96.7 199.2 97.5 200.0 ;
      RECT  109.8 213.2 110.6 214.0 ;
      RECT  98.1 210.0 98.9 210.8 ;
      RECT  96.7 216.4 97.5 217.2 ;
      RECT  111.2 216.4 112.0 217.2 ;
      RECT  98.1 226.8 98.9 227.6 ;
      RECT  112.6 226.8 113.4 227.6 ;
      RECT  108.4 199.0 109.2 199.8 ;
      RECT  109.8 197.6 110.6 198.4 ;
      RECT  111.2 210.2 112.0 211.0 ;
      RECT  109.8 211.6 110.6 212.4 ;
      RECT  108.4 219.8 109.2 220.6 ;
      RECT  112.6 218.4 113.4 219.2 ;
      RECT  111.2 231.0 112.0 231.8 ;
      RECT  112.6 232.4 113.4 233.2 ;
      RECT  105.3 204.6 106.1 205.4 ;
      RECT  122.7 204.6 123.5 205.4 ;
      RECT  105.3 194.2 106.1 195.0 ;
      RECT  122.7 194.2 123.5 195.0 ;
      RECT  105.3 204.6 106.1 205.4 ;
      RECT  122.7 204.6 123.5 205.4 ;
      RECT  105.3 215.0 106.1 215.8 ;
      RECT  122.7 215.0 123.5 215.8 ;
      RECT  105.3 225.4 106.1 226.2 ;
      RECT  122.7 225.4 123.5 226.2 ;
      RECT  105.3 215.0 106.1 215.8 ;
      RECT  122.7 215.0 123.5 215.8 ;
      RECT  105.3 225.4 106.1 226.2 ;
      RECT  122.7 225.4 123.5 226.2 ;
      RECT  105.3 235.8 106.1 236.6 ;
      RECT  122.7 235.8 123.5 236.6 ;
      RECT  126.9 199.3 127.5 199.9 ;
      RECT  126.9 210.1 127.5 210.7 ;
      RECT  126.9 220.1 127.5 220.7 ;
      RECT  126.9 230.9 127.5 231.5 ;
      RECT  106.0 240.9 106.6 241.5 ;
      RECT  106.0 244.5 106.6 245.1 ;
      RECT  103.1 240.9 106.3 241.5 ;
      RECT  106.0 241.2 106.6 244.8 ;
      RECT  106.3 244.5 108.8 245.1 ;
      RECT  97.1 240.9 100.7 241.5 ;
      RECT  106.0 251.7 106.6 252.3 ;
      RECT  106.0 254.9 106.6 255.5 ;
      RECT  103.1 251.7 106.3 252.3 ;
      RECT  106.0 252.0 106.6 255.2 ;
      RECT  106.3 254.9 110.2 255.5 ;
      RECT  98.5 251.7 100.7 252.3 ;
      RECT  97.1 258.1 111.6 258.7 ;
      RECT  98.5 268.5 113.0 269.1 ;
      RECT  108.8 240.7 115.7 241.3 ;
      RECT  110.2 239.3 117.7 239.9 ;
      RECT  111.6 251.9 115.7 252.5 ;
      RECT  110.2 253.3 117.7 253.9 ;
      RECT  108.8 261.5 115.7 262.1 ;
      RECT  113.0 260.1 117.7 260.7 ;
      RECT  111.6 272.7 115.7 273.3 ;
      RECT  113.0 274.1 117.7 274.7 ;
      RECT  122.6 240.7 123.2 241.3 ;
      RECT  122.6 240.9 123.2 241.5 ;
      RECT  120.7 240.7 122.9 241.3 ;
      RECT  122.6 241.0 123.2 241.2 ;
      RECT  122.9 240.9 125.1 241.5 ;
      RECT  122.6 251.9 123.2 252.5 ;
      RECT  122.6 251.7 123.2 252.3 ;
      RECT  120.7 251.9 122.9 252.5 ;
      RECT  122.6 252.0 123.2 252.2 ;
      RECT  122.9 251.7 125.1 252.3 ;
      RECT  122.6 261.5 123.2 262.1 ;
      RECT  122.6 261.7 123.2 262.3 ;
      RECT  120.7 261.5 122.9 262.1 ;
      RECT  122.6 261.8 123.2 262.0 ;
      RECT  122.9 261.7 125.1 262.3 ;
      RECT  122.6 272.7 123.2 273.3 ;
      RECT  122.6 272.5 123.2 273.1 ;
      RECT  120.7 272.7 122.9 273.3 ;
      RECT  122.6 272.8 123.2 273.0 ;
      RECT  122.9 272.5 125.1 273.1 ;
      RECT  96.5 246.3 130.1 246.9 ;
      RECT  96.5 235.9 130.1 236.5 ;
      RECT  96.5 246.3 130.1 246.9 ;
      RECT  96.5 256.7 130.1 257.3 ;
      RECT  96.5 267.1 130.1 267.7 ;
      RECT  96.5 256.7 130.1 257.3 ;
      RECT  96.5 267.1 130.1 267.7 ;
      RECT  96.5 277.5 130.1 278.1 ;
      RECT  103.7 245.3 104.5 246.6 ;
      RECT  103.7 236.2 104.5 237.5 ;
      RECT  100.5 237.1 101.3 235.9 ;
      RECT  100.5 244.5 101.3 246.9 ;
      RECT  102.2 237.1 102.8 245.3 ;
      RECT  100.5 244.5 101.3 245.3 ;
      RECT  102.1 244.5 102.9 245.3 ;
      RECT  102.1 244.5 102.9 245.3 ;
      RECT  100.5 244.5 101.3 245.3 ;
      RECT  100.5 237.1 101.3 237.9 ;
      RECT  102.1 237.1 102.9 237.9 ;
      RECT  102.1 237.1 102.9 237.9 ;
      RECT  100.5 237.1 101.3 237.9 ;
      RECT  103.7 244.9 104.5 245.7 ;
      RECT  103.7 237.1 104.5 237.9 ;
      RECT  100.7 240.8 101.5 241.6 ;
      RECT  100.7 240.8 101.5 241.6 ;
      RECT  102.5 240.9 103.1 241.5 ;
      RECT  99.3 246.3 105.7 246.9 ;
      RECT  99.3 235.9 105.7 236.5 ;
      RECT  103.7 247.9 104.5 246.6 ;
      RECT  103.7 257.0 104.5 255.7 ;
      RECT  100.5 256.1 101.3 257.3 ;
      RECT  100.5 248.7 101.3 246.3 ;
      RECT  102.2 256.1 102.8 247.9 ;
      RECT  100.5 248.7 101.3 247.9 ;
      RECT  102.1 248.7 102.9 247.9 ;
      RECT  102.1 248.7 102.9 247.9 ;
      RECT  100.5 248.7 101.3 247.9 ;
      RECT  100.5 256.1 101.3 255.3 ;
      RECT  102.1 256.1 102.9 255.3 ;
      RECT  102.1 256.1 102.9 255.3 ;
      RECT  100.5 256.1 101.3 255.3 ;
      RECT  103.7 248.3 104.5 247.5 ;
      RECT  103.7 256.1 104.5 255.3 ;
      RECT  100.7 252.4 101.5 251.6 ;
      RECT  100.7 252.4 101.5 251.6 ;
      RECT  102.5 252.3 103.1 251.7 ;
      RECT  99.3 246.9 105.7 246.3 ;
      RECT  99.3 257.3 105.7 256.7 ;
      RECT  128.1 245.3 128.9 246.6 ;
      RECT  128.1 236.2 128.9 237.5 ;
      RECT  124.9 237.1 125.7 235.9 ;
      RECT  124.9 244.5 125.7 246.9 ;
      RECT  126.6 237.1 127.2 245.3 ;
      RECT  124.9 244.5 125.7 245.3 ;
      RECT  126.5 244.5 127.3 245.3 ;
      RECT  126.5 244.5 127.3 245.3 ;
      RECT  124.9 244.5 125.7 245.3 ;
      RECT  124.9 237.1 125.7 237.9 ;
      RECT  126.5 237.1 127.3 237.9 ;
      RECT  126.5 237.1 127.3 237.9 ;
      RECT  124.9 237.1 125.7 237.9 ;
      RECT  128.1 244.9 128.9 245.7 ;
      RECT  128.1 237.1 128.9 237.9 ;
      RECT  125.1 240.8 125.9 241.6 ;
      RECT  125.1 240.8 125.9 241.6 ;
      RECT  126.9 240.9 127.5 241.5 ;
      RECT  123.7 246.3 130.1 246.9 ;
      RECT  123.7 235.9 130.1 236.5 ;
      RECT  128.1 247.9 128.9 246.6 ;
      RECT  128.1 257.0 128.9 255.7 ;
      RECT  124.9 256.1 125.7 257.3 ;
      RECT  124.9 248.7 125.7 246.3 ;
      RECT  126.6 256.1 127.2 247.9 ;
      RECT  124.9 248.7 125.7 247.9 ;
      RECT  126.5 248.7 127.3 247.9 ;
      RECT  126.5 248.7 127.3 247.9 ;
      RECT  124.9 248.7 125.7 247.9 ;
      RECT  124.9 256.1 125.7 255.3 ;
      RECT  126.5 256.1 127.3 255.3 ;
      RECT  126.5 256.1 127.3 255.3 ;
      RECT  124.9 256.1 125.7 255.3 ;
      RECT  128.1 248.3 128.9 247.5 ;
      RECT  128.1 256.1 128.9 255.3 ;
      RECT  125.1 252.4 125.9 251.6 ;
      RECT  125.1 252.4 125.9 251.6 ;
      RECT  126.9 252.3 127.5 251.7 ;
      RECT  123.7 246.9 130.1 246.3 ;
      RECT  123.7 257.3 130.1 256.7 ;
      RECT  128.1 266.1 128.9 267.4 ;
      RECT  128.1 257.0 128.9 258.3 ;
      RECT  124.9 257.9 125.7 256.7 ;
      RECT  124.9 265.3 125.7 267.7 ;
      RECT  126.6 257.9 127.2 266.1 ;
      RECT  124.9 265.3 125.7 266.1 ;
      RECT  126.5 265.3 127.3 266.1 ;
      RECT  126.5 265.3 127.3 266.1 ;
      RECT  124.9 265.3 125.7 266.1 ;
      RECT  124.9 257.9 125.7 258.7 ;
      RECT  126.5 257.9 127.3 258.7 ;
      RECT  126.5 257.9 127.3 258.7 ;
      RECT  124.9 257.9 125.7 258.7 ;
      RECT  128.1 265.7 128.9 266.5 ;
      RECT  128.1 257.9 128.9 258.7 ;
      RECT  125.1 261.6 125.9 262.4 ;
      RECT  125.1 261.6 125.9 262.4 ;
      RECT  126.9 261.7 127.5 262.3 ;
      RECT  123.7 267.1 130.1 267.7 ;
      RECT  123.7 256.7 130.1 257.3 ;
      RECT  128.1 268.7 128.9 267.4 ;
      RECT  128.1 277.8 128.9 276.5 ;
      RECT  124.9 276.9 125.7 278.1 ;
      RECT  124.9 269.5 125.7 267.1 ;
      RECT  126.6 276.9 127.2 268.7 ;
      RECT  124.9 269.5 125.7 268.7 ;
      RECT  126.5 269.5 127.3 268.7 ;
      RECT  126.5 269.5 127.3 268.7 ;
      RECT  124.9 269.5 125.7 268.7 ;
      RECT  124.9 276.9 125.7 276.1 ;
      RECT  126.5 276.9 127.3 276.1 ;
      RECT  126.5 276.9 127.3 276.1 ;
      RECT  124.9 276.9 125.7 276.1 ;
      RECT  128.1 269.1 128.9 268.3 ;
      RECT  128.1 276.9 128.9 276.1 ;
      RECT  125.1 273.2 125.9 272.4 ;
      RECT  125.1 273.2 125.9 272.4 ;
      RECT  126.9 273.1 127.5 272.5 ;
      RECT  123.7 267.7 130.1 267.1 ;
      RECT  123.7 278.1 130.1 277.5 ;
      RECT  115.3 237.5 116.1 235.9 ;
      RECT  115.3 244.5 116.1 246.9 ;
      RECT  118.5 244.5 119.3 246.9 ;
      RECT  120.1 245.3 120.9 246.6 ;
      RECT  120.1 236.2 120.9 237.5 ;
      RECT  115.3 244.5 116.1 245.3 ;
      RECT  116.9 244.5 117.7 245.3 ;
      RECT  116.9 244.5 117.7 245.3 ;
      RECT  115.3 244.5 116.1 245.3 ;
      RECT  116.9 244.5 117.7 245.3 ;
      RECT  118.5 244.5 119.3 245.3 ;
      RECT  118.5 244.5 119.3 245.3 ;
      RECT  116.9 244.5 117.7 245.3 ;
      RECT  115.3 237.5 116.1 238.3 ;
      RECT  116.9 237.5 117.7 238.3 ;
      RECT  116.9 237.5 117.7 238.3 ;
      RECT  115.3 237.5 116.1 238.3 ;
      RECT  116.9 237.5 117.7 238.3 ;
      RECT  118.5 237.5 119.3 238.3 ;
      RECT  118.5 237.5 119.3 238.3 ;
      RECT  116.9 237.5 117.7 238.3 ;
      RECT  120.1 244.9 120.9 245.7 ;
      RECT  120.1 237.1 120.9 237.9 ;
      RECT  117.7 239.2 118.5 240.0 ;
      RECT  115.7 240.6 116.5 241.4 ;
      RECT  116.9 244.5 117.7 245.3 ;
      RECT  118.5 237.5 119.3 238.3 ;
      RECT  119.9 240.6 120.7 241.4 ;
      RECT  115.7 240.6 116.5 241.4 ;
      RECT  117.7 239.2 118.5 240.0 ;
      RECT  119.9 240.6 120.7 241.4 ;
      RECT  114.1 246.3 123.7 246.9 ;
      RECT  114.1 235.9 123.7 236.5 ;
      RECT  115.3 255.7 116.1 257.3 ;
      RECT  115.3 248.7 116.1 246.3 ;
      RECT  118.5 248.7 119.3 246.3 ;
      RECT  120.1 247.9 120.9 246.6 ;
      RECT  120.1 257.0 120.9 255.7 ;
      RECT  115.3 248.7 116.1 247.9 ;
      RECT  116.9 248.7 117.7 247.9 ;
      RECT  116.9 248.7 117.7 247.9 ;
      RECT  115.3 248.7 116.1 247.9 ;
      RECT  116.9 248.7 117.7 247.9 ;
      RECT  118.5 248.7 119.3 247.9 ;
      RECT  118.5 248.7 119.3 247.9 ;
      RECT  116.9 248.7 117.7 247.9 ;
      RECT  115.3 255.7 116.1 254.9 ;
      RECT  116.9 255.7 117.7 254.9 ;
      RECT  116.9 255.7 117.7 254.9 ;
      RECT  115.3 255.7 116.1 254.9 ;
      RECT  116.9 255.7 117.7 254.9 ;
      RECT  118.5 255.7 119.3 254.9 ;
      RECT  118.5 255.7 119.3 254.9 ;
      RECT  116.9 255.7 117.7 254.9 ;
      RECT  120.1 248.3 120.9 247.5 ;
      RECT  120.1 256.1 120.9 255.3 ;
      RECT  117.7 254.0 118.5 253.2 ;
      RECT  115.7 252.6 116.5 251.8 ;
      RECT  116.9 248.7 117.7 247.9 ;
      RECT  118.5 255.7 119.3 254.9 ;
      RECT  119.9 252.6 120.7 251.8 ;
      RECT  115.7 252.6 116.5 251.8 ;
      RECT  117.7 254.0 118.5 253.2 ;
      RECT  119.9 252.6 120.7 251.8 ;
      RECT  114.1 246.9 123.7 246.3 ;
      RECT  114.1 257.3 123.7 256.7 ;
      RECT  115.3 258.3 116.1 256.7 ;
      RECT  115.3 265.3 116.1 267.7 ;
      RECT  118.5 265.3 119.3 267.7 ;
      RECT  120.1 266.1 120.9 267.4 ;
      RECT  120.1 257.0 120.9 258.3 ;
      RECT  115.3 265.3 116.1 266.1 ;
      RECT  116.9 265.3 117.7 266.1 ;
      RECT  116.9 265.3 117.7 266.1 ;
      RECT  115.3 265.3 116.1 266.1 ;
      RECT  116.9 265.3 117.7 266.1 ;
      RECT  118.5 265.3 119.3 266.1 ;
      RECT  118.5 265.3 119.3 266.1 ;
      RECT  116.9 265.3 117.7 266.1 ;
      RECT  115.3 258.3 116.1 259.1 ;
      RECT  116.9 258.3 117.7 259.1 ;
      RECT  116.9 258.3 117.7 259.1 ;
      RECT  115.3 258.3 116.1 259.1 ;
      RECT  116.9 258.3 117.7 259.1 ;
      RECT  118.5 258.3 119.3 259.1 ;
      RECT  118.5 258.3 119.3 259.1 ;
      RECT  116.9 258.3 117.7 259.1 ;
      RECT  120.1 265.7 120.9 266.5 ;
      RECT  120.1 257.9 120.9 258.7 ;
      RECT  117.7 260.0 118.5 260.8 ;
      RECT  115.7 261.4 116.5 262.2 ;
      RECT  116.9 265.3 117.7 266.1 ;
      RECT  118.5 258.3 119.3 259.1 ;
      RECT  119.9 261.4 120.7 262.2 ;
      RECT  115.7 261.4 116.5 262.2 ;
      RECT  117.7 260.0 118.5 260.8 ;
      RECT  119.9 261.4 120.7 262.2 ;
      RECT  114.1 267.1 123.7 267.7 ;
      RECT  114.1 256.7 123.7 257.3 ;
      RECT  115.3 276.5 116.1 278.1 ;
      RECT  115.3 269.5 116.1 267.1 ;
      RECT  118.5 269.5 119.3 267.1 ;
      RECT  120.1 268.7 120.9 267.4 ;
      RECT  120.1 277.8 120.9 276.5 ;
      RECT  115.3 269.5 116.1 268.7 ;
      RECT  116.9 269.5 117.7 268.7 ;
      RECT  116.9 269.5 117.7 268.7 ;
      RECT  115.3 269.5 116.1 268.7 ;
      RECT  116.9 269.5 117.7 268.7 ;
      RECT  118.5 269.5 119.3 268.7 ;
      RECT  118.5 269.5 119.3 268.7 ;
      RECT  116.9 269.5 117.7 268.7 ;
      RECT  115.3 276.5 116.1 275.7 ;
      RECT  116.9 276.5 117.7 275.7 ;
      RECT  116.9 276.5 117.7 275.7 ;
      RECT  115.3 276.5 116.1 275.7 ;
      RECT  116.9 276.5 117.7 275.7 ;
      RECT  118.5 276.5 119.3 275.7 ;
      RECT  118.5 276.5 119.3 275.7 ;
      RECT  116.9 276.5 117.7 275.7 ;
      RECT  120.1 269.1 120.9 268.3 ;
      RECT  120.1 276.9 120.9 276.1 ;
      RECT  117.7 274.8 118.5 274.0 ;
      RECT  115.7 273.4 116.5 272.6 ;
      RECT  116.9 269.5 117.7 268.7 ;
      RECT  118.5 276.5 119.3 275.7 ;
      RECT  119.9 273.4 120.7 272.6 ;
      RECT  115.7 273.4 116.5 272.6 ;
      RECT  117.7 274.8 118.5 274.0 ;
      RECT  119.9 273.4 120.7 272.6 ;
      RECT  114.1 267.7 123.7 267.1 ;
      RECT  114.1 278.1 123.7 277.5 ;
      RECT  108.4 244.4 109.2 245.2 ;
      RECT  96.7 240.8 97.5 241.6 ;
      RECT  109.8 254.8 110.6 255.6 ;
      RECT  98.1 251.6 98.9 252.4 ;
      RECT  96.7 258.0 97.5 258.8 ;
      RECT  111.2 258.0 112.0 258.8 ;
      RECT  98.1 268.4 98.9 269.2 ;
      RECT  112.6 268.4 113.4 269.2 ;
      RECT  108.4 240.6 109.2 241.4 ;
      RECT  109.8 239.2 110.6 240.0 ;
      RECT  111.2 251.8 112.0 252.6 ;
      RECT  109.8 253.2 110.6 254.0 ;
      RECT  108.4 261.4 109.2 262.2 ;
      RECT  112.6 260.0 113.4 260.8 ;
      RECT  111.2 272.6 112.0 273.4 ;
      RECT  112.6 274.0 113.4 274.8 ;
      RECT  105.3 246.2 106.1 247.0 ;
      RECT  122.7 246.2 123.5 247.0 ;
      RECT  105.3 235.8 106.1 236.6 ;
      RECT  122.7 235.8 123.5 236.6 ;
      RECT  105.3 246.2 106.1 247.0 ;
      RECT  122.7 246.2 123.5 247.0 ;
      RECT  105.3 256.6 106.1 257.4 ;
      RECT  122.7 256.6 123.5 257.4 ;
      RECT  105.3 267.0 106.1 267.8 ;
      RECT  122.7 267.0 123.5 267.8 ;
      RECT  105.3 256.6 106.1 257.4 ;
      RECT  122.7 256.6 123.5 257.4 ;
      RECT  105.3 267.0 106.1 267.8 ;
      RECT  122.7 267.0 123.5 267.8 ;
      RECT  105.3 277.4 106.1 278.2 ;
      RECT  122.7 277.4 123.5 278.2 ;
      RECT  126.9 240.9 127.5 241.5 ;
      RECT  126.9 251.7 127.5 252.3 ;
      RECT  126.9 261.7 127.5 262.3 ;
      RECT  126.9 272.5 127.5 273.1 ;
      RECT  142.5 195.9 143.3 194.3 ;
      RECT  142.5 202.9 143.3 205.3 ;
      RECT  145.7 202.9 146.5 205.3 ;
      RECT  147.3 203.7 148.1 205.0 ;
      RECT  147.3 194.6 148.1 195.9 ;
      RECT  142.5 202.9 143.3 203.7 ;
      RECT  144.1 202.9 144.9 203.7 ;
      RECT  144.1 202.9 144.9 203.7 ;
      RECT  142.5 202.9 143.3 203.7 ;
      RECT  144.1 202.9 144.9 203.7 ;
      RECT  145.7 202.9 146.5 203.7 ;
      RECT  145.7 202.9 146.5 203.7 ;
      RECT  144.1 202.9 144.9 203.7 ;
      RECT  142.5 195.9 143.3 196.7 ;
      RECT  144.1 195.9 144.9 196.7 ;
      RECT  144.1 195.9 144.9 196.7 ;
      RECT  142.5 195.9 143.3 196.7 ;
      RECT  144.1 195.9 144.9 196.7 ;
      RECT  145.7 195.9 146.5 196.7 ;
      RECT  145.7 195.9 146.5 196.7 ;
      RECT  144.1 195.9 144.9 196.7 ;
      RECT  147.3 203.3 148.1 204.1 ;
      RECT  147.3 195.5 148.1 196.3 ;
      RECT  144.9 197.6 145.7 198.4 ;
      RECT  142.9 199.0 143.7 199.8 ;
      RECT  144.1 202.9 144.9 203.7 ;
      RECT  145.7 195.9 146.5 196.7 ;
      RECT  147.1 199.0 147.9 199.8 ;
      RECT  142.9 199.0 143.7 199.8 ;
      RECT  144.9 197.6 145.7 198.4 ;
      RECT  147.1 199.0 147.9 199.8 ;
      RECT  141.3 204.7 150.9 205.3 ;
      RECT  141.3 194.3 150.9 194.9 ;
      RECT  142.5 214.1 143.3 215.7 ;
      RECT  142.5 207.1 143.3 204.7 ;
      RECT  145.7 207.1 146.5 204.7 ;
      RECT  147.3 206.3 148.1 205.0 ;
      RECT  147.3 215.4 148.1 214.1 ;
      RECT  142.5 207.1 143.3 206.3 ;
      RECT  144.1 207.1 144.9 206.3 ;
      RECT  144.1 207.1 144.9 206.3 ;
      RECT  142.5 207.1 143.3 206.3 ;
      RECT  144.1 207.1 144.9 206.3 ;
      RECT  145.7 207.1 146.5 206.3 ;
      RECT  145.7 207.1 146.5 206.3 ;
      RECT  144.1 207.1 144.9 206.3 ;
      RECT  142.5 214.1 143.3 213.3 ;
      RECT  144.1 214.1 144.9 213.3 ;
      RECT  144.1 214.1 144.9 213.3 ;
      RECT  142.5 214.1 143.3 213.3 ;
      RECT  144.1 214.1 144.9 213.3 ;
      RECT  145.7 214.1 146.5 213.3 ;
      RECT  145.7 214.1 146.5 213.3 ;
      RECT  144.1 214.1 144.9 213.3 ;
      RECT  147.3 206.7 148.1 205.9 ;
      RECT  147.3 214.5 148.1 213.7 ;
      RECT  144.9 212.4 145.7 211.6 ;
      RECT  142.9 211.0 143.7 210.2 ;
      RECT  144.1 207.1 144.9 206.3 ;
      RECT  145.7 214.1 146.5 213.3 ;
      RECT  147.1 211.0 147.9 210.2 ;
      RECT  142.9 211.0 143.7 210.2 ;
      RECT  144.9 212.4 145.7 211.6 ;
      RECT  147.1 211.0 147.9 210.2 ;
      RECT  141.3 205.3 150.9 204.7 ;
      RECT  141.3 215.7 150.9 215.1 ;
      RECT  142.5 216.7 143.3 215.1 ;
      RECT  142.5 223.7 143.3 226.1 ;
      RECT  145.7 223.7 146.5 226.1 ;
      RECT  147.3 224.5 148.1 225.8 ;
      RECT  147.3 215.4 148.1 216.7 ;
      RECT  142.5 223.7 143.3 224.5 ;
      RECT  144.1 223.7 144.9 224.5 ;
      RECT  144.1 223.7 144.9 224.5 ;
      RECT  142.5 223.7 143.3 224.5 ;
      RECT  144.1 223.7 144.9 224.5 ;
      RECT  145.7 223.7 146.5 224.5 ;
      RECT  145.7 223.7 146.5 224.5 ;
      RECT  144.1 223.7 144.9 224.5 ;
      RECT  142.5 216.7 143.3 217.5 ;
      RECT  144.1 216.7 144.9 217.5 ;
      RECT  144.1 216.7 144.9 217.5 ;
      RECT  142.5 216.7 143.3 217.5 ;
      RECT  144.1 216.7 144.9 217.5 ;
      RECT  145.7 216.7 146.5 217.5 ;
      RECT  145.7 216.7 146.5 217.5 ;
      RECT  144.1 216.7 144.9 217.5 ;
      RECT  147.3 224.1 148.1 224.9 ;
      RECT  147.3 216.3 148.1 217.1 ;
      RECT  144.9 218.4 145.7 219.2 ;
      RECT  142.9 219.8 143.7 220.6 ;
      RECT  144.1 223.7 144.9 224.5 ;
      RECT  145.7 216.7 146.5 217.5 ;
      RECT  147.1 219.8 147.9 220.6 ;
      RECT  142.9 219.8 143.7 220.6 ;
      RECT  144.9 218.4 145.7 219.2 ;
      RECT  147.1 219.8 147.9 220.6 ;
      RECT  141.3 225.5 150.9 226.1 ;
      RECT  141.3 215.1 150.9 215.7 ;
      RECT  142.5 234.9 143.3 236.5 ;
      RECT  142.5 227.9 143.3 225.5 ;
      RECT  145.7 227.9 146.5 225.5 ;
      RECT  147.3 227.1 148.1 225.8 ;
      RECT  147.3 236.2 148.1 234.9 ;
      RECT  142.5 227.9 143.3 227.1 ;
      RECT  144.1 227.9 144.9 227.1 ;
      RECT  144.1 227.9 144.9 227.1 ;
      RECT  142.5 227.9 143.3 227.1 ;
      RECT  144.1 227.9 144.9 227.1 ;
      RECT  145.7 227.9 146.5 227.1 ;
      RECT  145.7 227.9 146.5 227.1 ;
      RECT  144.1 227.9 144.9 227.1 ;
      RECT  142.5 234.9 143.3 234.1 ;
      RECT  144.1 234.9 144.9 234.1 ;
      RECT  144.1 234.9 144.9 234.1 ;
      RECT  142.5 234.9 143.3 234.1 ;
      RECT  144.1 234.9 144.9 234.1 ;
      RECT  145.7 234.9 146.5 234.1 ;
      RECT  145.7 234.9 146.5 234.1 ;
      RECT  144.1 234.9 144.9 234.1 ;
      RECT  147.3 227.5 148.1 226.7 ;
      RECT  147.3 235.3 148.1 234.5 ;
      RECT  144.9 233.2 145.7 232.4 ;
      RECT  142.9 231.8 143.7 231.0 ;
      RECT  144.1 227.9 144.9 227.1 ;
      RECT  145.7 234.9 146.5 234.1 ;
      RECT  147.1 231.8 147.9 231.0 ;
      RECT  142.9 231.8 143.7 231.0 ;
      RECT  144.9 233.2 145.7 232.4 ;
      RECT  147.1 231.8 147.9 231.0 ;
      RECT  141.3 226.1 150.9 225.5 ;
      RECT  141.3 236.5 150.9 235.9 ;
      RECT  142.5 237.5 143.3 235.9 ;
      RECT  142.5 244.5 143.3 246.9 ;
      RECT  145.7 244.5 146.5 246.9 ;
      RECT  147.3 245.3 148.1 246.6 ;
      RECT  147.3 236.2 148.1 237.5 ;
      RECT  142.5 244.5 143.3 245.3 ;
      RECT  144.1 244.5 144.9 245.3 ;
      RECT  144.1 244.5 144.9 245.3 ;
      RECT  142.5 244.5 143.3 245.3 ;
      RECT  144.1 244.5 144.9 245.3 ;
      RECT  145.7 244.5 146.5 245.3 ;
      RECT  145.7 244.5 146.5 245.3 ;
      RECT  144.1 244.5 144.9 245.3 ;
      RECT  142.5 237.5 143.3 238.3 ;
      RECT  144.1 237.5 144.9 238.3 ;
      RECT  144.1 237.5 144.9 238.3 ;
      RECT  142.5 237.5 143.3 238.3 ;
      RECT  144.1 237.5 144.9 238.3 ;
      RECT  145.7 237.5 146.5 238.3 ;
      RECT  145.7 237.5 146.5 238.3 ;
      RECT  144.1 237.5 144.9 238.3 ;
      RECT  147.3 244.9 148.1 245.7 ;
      RECT  147.3 237.1 148.1 237.9 ;
      RECT  144.9 239.2 145.7 240.0 ;
      RECT  142.9 240.6 143.7 241.4 ;
      RECT  144.1 244.5 144.9 245.3 ;
      RECT  145.7 237.5 146.5 238.3 ;
      RECT  147.1 240.6 147.9 241.4 ;
      RECT  142.9 240.6 143.7 241.4 ;
      RECT  144.9 239.2 145.7 240.0 ;
      RECT  147.1 240.6 147.9 241.4 ;
      RECT  141.3 246.3 150.9 246.9 ;
      RECT  141.3 235.9 150.9 236.5 ;
      RECT  142.5 255.7 143.3 257.3 ;
      RECT  142.5 248.7 143.3 246.3 ;
      RECT  145.7 248.7 146.5 246.3 ;
      RECT  147.3 247.9 148.1 246.6 ;
      RECT  147.3 257.0 148.1 255.7 ;
      RECT  142.5 248.7 143.3 247.9 ;
      RECT  144.1 248.7 144.9 247.9 ;
      RECT  144.1 248.7 144.9 247.9 ;
      RECT  142.5 248.7 143.3 247.9 ;
      RECT  144.1 248.7 144.9 247.9 ;
      RECT  145.7 248.7 146.5 247.9 ;
      RECT  145.7 248.7 146.5 247.9 ;
      RECT  144.1 248.7 144.9 247.9 ;
      RECT  142.5 255.7 143.3 254.9 ;
      RECT  144.1 255.7 144.9 254.9 ;
      RECT  144.1 255.7 144.9 254.9 ;
      RECT  142.5 255.7 143.3 254.9 ;
      RECT  144.1 255.7 144.9 254.9 ;
      RECT  145.7 255.7 146.5 254.9 ;
      RECT  145.7 255.7 146.5 254.9 ;
      RECT  144.1 255.7 144.9 254.9 ;
      RECT  147.3 248.3 148.1 247.5 ;
      RECT  147.3 256.1 148.1 255.3 ;
      RECT  144.9 254.0 145.7 253.2 ;
      RECT  142.9 252.6 143.7 251.8 ;
      RECT  144.1 248.7 144.9 247.9 ;
      RECT  145.7 255.7 146.5 254.9 ;
      RECT  147.1 252.6 147.9 251.8 ;
      RECT  142.9 252.6 143.7 251.8 ;
      RECT  144.9 254.0 145.7 253.2 ;
      RECT  147.1 252.6 147.9 251.8 ;
      RECT  141.3 246.9 150.9 246.3 ;
      RECT  141.3 257.3 150.9 256.7 ;
      RECT  142.5 258.3 143.3 256.7 ;
      RECT  142.5 265.3 143.3 267.7 ;
      RECT  145.7 265.3 146.5 267.7 ;
      RECT  147.3 266.1 148.1 267.4 ;
      RECT  147.3 257.0 148.1 258.3 ;
      RECT  142.5 265.3 143.3 266.1 ;
      RECT  144.1 265.3 144.9 266.1 ;
      RECT  144.1 265.3 144.9 266.1 ;
      RECT  142.5 265.3 143.3 266.1 ;
      RECT  144.1 265.3 144.9 266.1 ;
      RECT  145.7 265.3 146.5 266.1 ;
      RECT  145.7 265.3 146.5 266.1 ;
      RECT  144.1 265.3 144.9 266.1 ;
      RECT  142.5 258.3 143.3 259.1 ;
      RECT  144.1 258.3 144.9 259.1 ;
      RECT  144.1 258.3 144.9 259.1 ;
      RECT  142.5 258.3 143.3 259.1 ;
      RECT  144.1 258.3 144.9 259.1 ;
      RECT  145.7 258.3 146.5 259.1 ;
      RECT  145.7 258.3 146.5 259.1 ;
      RECT  144.1 258.3 144.9 259.1 ;
      RECT  147.3 265.7 148.1 266.5 ;
      RECT  147.3 257.9 148.1 258.7 ;
      RECT  144.9 260.0 145.7 260.8 ;
      RECT  142.9 261.4 143.7 262.2 ;
      RECT  144.1 265.3 144.9 266.1 ;
      RECT  145.7 258.3 146.5 259.1 ;
      RECT  147.1 261.4 147.9 262.2 ;
      RECT  142.9 261.4 143.7 262.2 ;
      RECT  144.9 260.0 145.7 260.8 ;
      RECT  147.1 261.4 147.9 262.2 ;
      RECT  141.3 267.1 150.9 267.7 ;
      RECT  141.3 256.7 150.9 257.3 ;
      RECT  142.5 276.5 143.3 278.1 ;
      RECT  142.5 269.5 143.3 267.1 ;
      RECT  145.7 269.5 146.5 267.1 ;
      RECT  147.3 268.7 148.1 267.4 ;
      RECT  147.3 277.8 148.1 276.5 ;
      RECT  142.5 269.5 143.3 268.7 ;
      RECT  144.1 269.5 144.9 268.7 ;
      RECT  144.1 269.5 144.9 268.7 ;
      RECT  142.5 269.5 143.3 268.7 ;
      RECT  144.1 269.5 144.9 268.7 ;
      RECT  145.7 269.5 146.5 268.7 ;
      RECT  145.7 269.5 146.5 268.7 ;
      RECT  144.1 269.5 144.9 268.7 ;
      RECT  142.5 276.5 143.3 275.7 ;
      RECT  144.1 276.5 144.9 275.7 ;
      RECT  144.1 276.5 144.9 275.7 ;
      RECT  142.5 276.5 143.3 275.7 ;
      RECT  144.1 276.5 144.9 275.7 ;
      RECT  145.7 276.5 146.5 275.7 ;
      RECT  145.7 276.5 146.5 275.7 ;
      RECT  144.1 276.5 144.9 275.7 ;
      RECT  147.3 269.1 148.1 268.3 ;
      RECT  147.3 276.9 148.1 276.1 ;
      RECT  144.9 274.8 145.7 274.0 ;
      RECT  142.9 273.4 143.7 272.6 ;
      RECT  144.1 269.5 144.9 268.7 ;
      RECT  145.7 276.5 146.5 275.7 ;
      RECT  147.1 273.4 147.9 272.6 ;
      RECT  142.9 273.4 143.7 272.6 ;
      RECT  144.9 274.8 145.7 274.0 ;
      RECT  147.1 273.4 147.9 272.6 ;
      RECT  141.3 267.7 150.9 267.1 ;
      RECT  141.3 278.1 150.9 277.5 ;
      RECT  142.5 279.1 143.3 277.5 ;
      RECT  142.5 286.1 143.3 288.5 ;
      RECT  145.7 286.1 146.5 288.5 ;
      RECT  147.3 286.9 148.1 288.2 ;
      RECT  147.3 277.8 148.1 279.1 ;
      RECT  142.5 286.1 143.3 286.9 ;
      RECT  144.1 286.1 144.9 286.9 ;
      RECT  144.1 286.1 144.9 286.9 ;
      RECT  142.5 286.1 143.3 286.9 ;
      RECT  144.1 286.1 144.9 286.9 ;
      RECT  145.7 286.1 146.5 286.9 ;
      RECT  145.7 286.1 146.5 286.9 ;
      RECT  144.1 286.1 144.9 286.9 ;
      RECT  142.5 279.1 143.3 279.9 ;
      RECT  144.1 279.1 144.9 279.9 ;
      RECT  144.1 279.1 144.9 279.9 ;
      RECT  142.5 279.1 143.3 279.9 ;
      RECT  144.1 279.1 144.9 279.9 ;
      RECT  145.7 279.1 146.5 279.9 ;
      RECT  145.7 279.1 146.5 279.9 ;
      RECT  144.1 279.1 144.9 279.9 ;
      RECT  147.3 286.5 148.1 287.3 ;
      RECT  147.3 278.7 148.1 279.5 ;
      RECT  144.9 280.8 145.7 281.6 ;
      RECT  142.9 282.2 143.7 283.0 ;
      RECT  144.1 286.1 144.9 286.9 ;
      RECT  145.7 279.1 146.5 279.9 ;
      RECT  147.1 282.2 147.9 283.0 ;
      RECT  142.9 282.2 143.7 283.0 ;
      RECT  144.9 280.8 145.7 281.6 ;
      RECT  147.1 282.2 147.9 283.0 ;
      RECT  141.3 287.9 150.9 288.5 ;
      RECT  141.3 277.5 150.9 278.1 ;
      RECT  142.5 297.3 143.3 298.9 ;
      RECT  142.5 290.3 143.3 287.9 ;
      RECT  145.7 290.3 146.5 287.9 ;
      RECT  147.3 289.5 148.1 288.2 ;
      RECT  147.3 298.6 148.1 297.3 ;
      RECT  142.5 290.3 143.3 289.5 ;
      RECT  144.1 290.3 144.9 289.5 ;
      RECT  144.1 290.3 144.9 289.5 ;
      RECT  142.5 290.3 143.3 289.5 ;
      RECT  144.1 290.3 144.9 289.5 ;
      RECT  145.7 290.3 146.5 289.5 ;
      RECT  145.7 290.3 146.5 289.5 ;
      RECT  144.1 290.3 144.9 289.5 ;
      RECT  142.5 297.3 143.3 296.5 ;
      RECT  144.1 297.3 144.9 296.5 ;
      RECT  144.1 297.3 144.9 296.5 ;
      RECT  142.5 297.3 143.3 296.5 ;
      RECT  144.1 297.3 144.9 296.5 ;
      RECT  145.7 297.3 146.5 296.5 ;
      RECT  145.7 297.3 146.5 296.5 ;
      RECT  144.1 297.3 144.9 296.5 ;
      RECT  147.3 289.9 148.1 289.1 ;
      RECT  147.3 297.7 148.1 296.9 ;
      RECT  144.9 295.6 145.7 294.8 ;
      RECT  142.9 294.2 143.7 293.4 ;
      RECT  144.1 290.3 144.9 289.5 ;
      RECT  145.7 297.3 146.5 296.5 ;
      RECT  147.1 294.2 147.9 293.4 ;
      RECT  142.9 294.2 143.7 293.4 ;
      RECT  144.9 295.6 145.7 294.8 ;
      RECT  147.1 294.2 147.9 293.4 ;
      RECT  141.3 288.5 150.9 287.9 ;
      RECT  141.3 298.9 150.9 298.3 ;
      RECT  142.5 299.9 143.3 298.3 ;
      RECT  142.5 306.9 143.3 309.3 ;
      RECT  145.7 306.9 146.5 309.3 ;
      RECT  147.3 307.7 148.1 309.0 ;
      RECT  147.3 298.6 148.1 299.9 ;
      RECT  142.5 306.9 143.3 307.7 ;
      RECT  144.1 306.9 144.9 307.7 ;
      RECT  144.1 306.9 144.9 307.7 ;
      RECT  142.5 306.9 143.3 307.7 ;
      RECT  144.1 306.9 144.9 307.7 ;
      RECT  145.7 306.9 146.5 307.7 ;
      RECT  145.7 306.9 146.5 307.7 ;
      RECT  144.1 306.9 144.9 307.7 ;
      RECT  142.5 299.9 143.3 300.7 ;
      RECT  144.1 299.9 144.9 300.7 ;
      RECT  144.1 299.9 144.9 300.7 ;
      RECT  142.5 299.9 143.3 300.7 ;
      RECT  144.1 299.9 144.9 300.7 ;
      RECT  145.7 299.9 146.5 300.7 ;
      RECT  145.7 299.9 146.5 300.7 ;
      RECT  144.1 299.9 144.9 300.7 ;
      RECT  147.3 307.3 148.1 308.1 ;
      RECT  147.3 299.5 148.1 300.3 ;
      RECT  144.9 301.6 145.7 302.4 ;
      RECT  142.9 303.0 143.7 303.8 ;
      RECT  144.1 306.9 144.9 307.7 ;
      RECT  145.7 299.9 146.5 300.7 ;
      RECT  147.1 303.0 147.9 303.8 ;
      RECT  142.9 303.0 143.7 303.8 ;
      RECT  144.9 301.6 145.7 302.4 ;
      RECT  147.1 303.0 147.9 303.8 ;
      RECT  141.3 308.7 150.9 309.3 ;
      RECT  141.3 298.3 150.9 298.9 ;
      RECT  142.5 318.1 143.3 319.7 ;
      RECT  142.5 311.1 143.3 308.7 ;
      RECT  145.7 311.1 146.5 308.7 ;
      RECT  147.3 310.3 148.1 309.0 ;
      RECT  147.3 319.4 148.1 318.1 ;
      RECT  142.5 311.1 143.3 310.3 ;
      RECT  144.1 311.1 144.9 310.3 ;
      RECT  144.1 311.1 144.9 310.3 ;
      RECT  142.5 311.1 143.3 310.3 ;
      RECT  144.1 311.1 144.9 310.3 ;
      RECT  145.7 311.1 146.5 310.3 ;
      RECT  145.7 311.1 146.5 310.3 ;
      RECT  144.1 311.1 144.9 310.3 ;
      RECT  142.5 318.1 143.3 317.3 ;
      RECT  144.1 318.1 144.9 317.3 ;
      RECT  144.1 318.1 144.9 317.3 ;
      RECT  142.5 318.1 143.3 317.3 ;
      RECT  144.1 318.1 144.9 317.3 ;
      RECT  145.7 318.1 146.5 317.3 ;
      RECT  145.7 318.1 146.5 317.3 ;
      RECT  144.1 318.1 144.9 317.3 ;
      RECT  147.3 310.7 148.1 309.9 ;
      RECT  147.3 318.5 148.1 317.7 ;
      RECT  144.9 316.4 145.7 315.6 ;
      RECT  142.9 315.0 143.7 314.2 ;
      RECT  144.1 311.1 144.9 310.3 ;
      RECT  145.7 318.1 146.5 317.3 ;
      RECT  147.1 315.0 147.9 314.2 ;
      RECT  142.9 315.0 143.7 314.2 ;
      RECT  144.9 316.4 145.7 315.6 ;
      RECT  147.1 315.0 147.9 314.2 ;
      RECT  141.3 309.3 150.9 308.7 ;
      RECT  141.3 319.7 150.9 319.1 ;
      RECT  142.5 320.7 143.3 319.1 ;
      RECT  142.5 327.7 143.3 330.1 ;
      RECT  145.7 327.7 146.5 330.1 ;
      RECT  147.3 328.5 148.1 329.8 ;
      RECT  147.3 319.4 148.1 320.7 ;
      RECT  142.5 327.7 143.3 328.5 ;
      RECT  144.1 327.7 144.9 328.5 ;
      RECT  144.1 327.7 144.9 328.5 ;
      RECT  142.5 327.7 143.3 328.5 ;
      RECT  144.1 327.7 144.9 328.5 ;
      RECT  145.7 327.7 146.5 328.5 ;
      RECT  145.7 327.7 146.5 328.5 ;
      RECT  144.1 327.7 144.9 328.5 ;
      RECT  142.5 320.7 143.3 321.5 ;
      RECT  144.1 320.7 144.9 321.5 ;
      RECT  144.1 320.7 144.9 321.5 ;
      RECT  142.5 320.7 143.3 321.5 ;
      RECT  144.1 320.7 144.9 321.5 ;
      RECT  145.7 320.7 146.5 321.5 ;
      RECT  145.7 320.7 146.5 321.5 ;
      RECT  144.1 320.7 144.9 321.5 ;
      RECT  147.3 328.1 148.1 328.9 ;
      RECT  147.3 320.3 148.1 321.1 ;
      RECT  144.9 322.4 145.7 323.2 ;
      RECT  142.9 323.8 143.7 324.6 ;
      RECT  144.1 327.7 144.9 328.5 ;
      RECT  145.7 320.7 146.5 321.5 ;
      RECT  147.1 323.8 147.9 324.6 ;
      RECT  142.9 323.8 143.7 324.6 ;
      RECT  144.9 322.4 145.7 323.2 ;
      RECT  147.1 323.8 147.9 324.6 ;
      RECT  141.3 329.5 150.9 330.1 ;
      RECT  141.3 319.1 150.9 319.7 ;
      RECT  142.5 338.9 143.3 340.5 ;
      RECT  142.5 331.9 143.3 329.5 ;
      RECT  145.7 331.9 146.5 329.5 ;
      RECT  147.3 331.1 148.1 329.8 ;
      RECT  147.3 340.2 148.1 338.9 ;
      RECT  142.5 331.9 143.3 331.1 ;
      RECT  144.1 331.9 144.9 331.1 ;
      RECT  144.1 331.9 144.9 331.1 ;
      RECT  142.5 331.9 143.3 331.1 ;
      RECT  144.1 331.9 144.9 331.1 ;
      RECT  145.7 331.9 146.5 331.1 ;
      RECT  145.7 331.9 146.5 331.1 ;
      RECT  144.1 331.9 144.9 331.1 ;
      RECT  142.5 338.9 143.3 338.1 ;
      RECT  144.1 338.9 144.9 338.1 ;
      RECT  144.1 338.9 144.9 338.1 ;
      RECT  142.5 338.9 143.3 338.1 ;
      RECT  144.1 338.9 144.9 338.1 ;
      RECT  145.7 338.9 146.5 338.1 ;
      RECT  145.7 338.9 146.5 338.1 ;
      RECT  144.1 338.9 144.9 338.1 ;
      RECT  147.3 331.5 148.1 330.7 ;
      RECT  147.3 339.3 148.1 338.5 ;
      RECT  144.9 337.2 145.7 336.4 ;
      RECT  142.9 335.8 143.7 335.0 ;
      RECT  144.1 331.9 144.9 331.1 ;
      RECT  145.7 338.9 146.5 338.1 ;
      RECT  147.1 335.8 147.9 335.0 ;
      RECT  142.9 335.8 143.7 335.0 ;
      RECT  144.9 337.2 145.7 336.4 ;
      RECT  147.1 335.8 147.9 335.0 ;
      RECT  141.3 330.1 150.9 329.5 ;
      RECT  141.3 340.5 150.9 339.9 ;
      RECT  142.5 341.5 143.3 339.9 ;
      RECT  142.5 348.5 143.3 350.9 ;
      RECT  145.7 348.5 146.5 350.9 ;
      RECT  147.3 349.3 148.1 350.6 ;
      RECT  147.3 340.2 148.1 341.5 ;
      RECT  142.5 348.5 143.3 349.3 ;
      RECT  144.1 348.5 144.9 349.3 ;
      RECT  144.1 348.5 144.9 349.3 ;
      RECT  142.5 348.5 143.3 349.3 ;
      RECT  144.1 348.5 144.9 349.3 ;
      RECT  145.7 348.5 146.5 349.3 ;
      RECT  145.7 348.5 146.5 349.3 ;
      RECT  144.1 348.5 144.9 349.3 ;
      RECT  142.5 341.5 143.3 342.3 ;
      RECT  144.1 341.5 144.9 342.3 ;
      RECT  144.1 341.5 144.9 342.3 ;
      RECT  142.5 341.5 143.3 342.3 ;
      RECT  144.1 341.5 144.9 342.3 ;
      RECT  145.7 341.5 146.5 342.3 ;
      RECT  145.7 341.5 146.5 342.3 ;
      RECT  144.1 341.5 144.9 342.3 ;
      RECT  147.3 348.9 148.1 349.7 ;
      RECT  147.3 341.1 148.1 341.9 ;
      RECT  144.9 343.2 145.7 344.0 ;
      RECT  142.9 344.6 143.7 345.4 ;
      RECT  144.1 348.5 144.9 349.3 ;
      RECT  145.7 341.5 146.5 342.3 ;
      RECT  147.1 344.6 147.9 345.4 ;
      RECT  142.9 344.6 143.7 345.4 ;
      RECT  144.9 343.2 145.7 344.0 ;
      RECT  147.1 344.6 147.9 345.4 ;
      RECT  141.3 350.3 150.9 350.9 ;
      RECT  141.3 339.9 150.9 340.5 ;
      RECT  142.5 359.7 143.3 361.3 ;
      RECT  142.5 352.7 143.3 350.3 ;
      RECT  145.7 352.7 146.5 350.3 ;
      RECT  147.3 351.9 148.1 350.6 ;
      RECT  147.3 361.0 148.1 359.7 ;
      RECT  142.5 352.7 143.3 351.9 ;
      RECT  144.1 352.7 144.9 351.9 ;
      RECT  144.1 352.7 144.9 351.9 ;
      RECT  142.5 352.7 143.3 351.9 ;
      RECT  144.1 352.7 144.9 351.9 ;
      RECT  145.7 352.7 146.5 351.9 ;
      RECT  145.7 352.7 146.5 351.9 ;
      RECT  144.1 352.7 144.9 351.9 ;
      RECT  142.5 359.7 143.3 358.9 ;
      RECT  144.1 359.7 144.9 358.9 ;
      RECT  144.1 359.7 144.9 358.9 ;
      RECT  142.5 359.7 143.3 358.9 ;
      RECT  144.1 359.7 144.9 358.9 ;
      RECT  145.7 359.7 146.5 358.9 ;
      RECT  145.7 359.7 146.5 358.9 ;
      RECT  144.1 359.7 144.9 358.9 ;
      RECT  147.3 352.3 148.1 351.5 ;
      RECT  147.3 360.1 148.1 359.3 ;
      RECT  144.9 358.0 145.7 357.2 ;
      RECT  142.9 356.6 143.7 355.8 ;
      RECT  144.1 352.7 144.9 351.9 ;
      RECT  145.7 359.7 146.5 358.9 ;
      RECT  147.1 356.6 147.9 355.8 ;
      RECT  142.9 356.6 143.7 355.8 ;
      RECT  144.9 358.0 145.7 357.2 ;
      RECT  147.1 356.6 147.9 355.8 ;
      RECT  141.3 350.9 150.9 350.3 ;
      RECT  141.3 361.3 150.9 360.7 ;
      RECT  155.3 203.7 156.1 205.0 ;
      RECT  155.3 194.6 156.1 195.9 ;
      RECT  152.1 195.5 152.9 194.3 ;
      RECT  152.1 202.9 152.9 205.3 ;
      RECT  153.8 195.5 154.4 203.7 ;
      RECT  152.1 202.9 152.9 203.7 ;
      RECT  153.7 202.9 154.5 203.7 ;
      RECT  153.7 202.9 154.5 203.7 ;
      RECT  152.1 202.9 152.9 203.7 ;
      RECT  152.1 195.5 152.9 196.3 ;
      RECT  153.7 195.5 154.5 196.3 ;
      RECT  153.7 195.5 154.5 196.3 ;
      RECT  152.1 195.5 152.9 196.3 ;
      RECT  155.3 203.3 156.1 204.1 ;
      RECT  155.3 195.5 156.1 196.3 ;
      RECT  152.3 199.2 153.1 200.0 ;
      RECT  152.3 199.2 153.1 200.0 ;
      RECT  154.1 199.3 154.7 199.9 ;
      RECT  150.9 204.7 157.3 205.3 ;
      RECT  150.9 194.3 157.3 194.9 ;
      RECT  155.3 206.3 156.1 205.0 ;
      RECT  155.3 215.4 156.1 214.1 ;
      RECT  152.1 214.5 152.9 215.7 ;
      RECT  152.1 207.1 152.9 204.7 ;
      RECT  153.8 214.5 154.4 206.3 ;
      RECT  152.1 207.1 152.9 206.3 ;
      RECT  153.7 207.1 154.5 206.3 ;
      RECT  153.7 207.1 154.5 206.3 ;
      RECT  152.1 207.1 152.9 206.3 ;
      RECT  152.1 214.5 152.9 213.7 ;
      RECT  153.7 214.5 154.5 213.7 ;
      RECT  153.7 214.5 154.5 213.7 ;
      RECT  152.1 214.5 152.9 213.7 ;
      RECT  155.3 206.7 156.1 205.9 ;
      RECT  155.3 214.5 156.1 213.7 ;
      RECT  152.3 210.8 153.1 210.0 ;
      RECT  152.3 210.8 153.1 210.0 ;
      RECT  154.1 210.7 154.7 210.1 ;
      RECT  150.9 205.3 157.3 204.7 ;
      RECT  150.9 215.7 157.3 215.1 ;
      RECT  155.3 224.5 156.1 225.8 ;
      RECT  155.3 215.4 156.1 216.7 ;
      RECT  152.1 216.3 152.9 215.1 ;
      RECT  152.1 223.7 152.9 226.1 ;
      RECT  153.8 216.3 154.4 224.5 ;
      RECT  152.1 223.7 152.9 224.5 ;
      RECT  153.7 223.7 154.5 224.5 ;
      RECT  153.7 223.7 154.5 224.5 ;
      RECT  152.1 223.7 152.9 224.5 ;
      RECT  152.1 216.3 152.9 217.1 ;
      RECT  153.7 216.3 154.5 217.1 ;
      RECT  153.7 216.3 154.5 217.1 ;
      RECT  152.1 216.3 152.9 217.1 ;
      RECT  155.3 224.1 156.1 224.9 ;
      RECT  155.3 216.3 156.1 217.1 ;
      RECT  152.3 220.0 153.1 220.8 ;
      RECT  152.3 220.0 153.1 220.8 ;
      RECT  154.1 220.1 154.7 220.7 ;
      RECT  150.9 225.5 157.3 226.1 ;
      RECT  150.9 215.1 157.3 215.7 ;
      RECT  155.3 227.1 156.1 225.8 ;
      RECT  155.3 236.2 156.1 234.9 ;
      RECT  152.1 235.3 152.9 236.5 ;
      RECT  152.1 227.9 152.9 225.5 ;
      RECT  153.8 235.3 154.4 227.1 ;
      RECT  152.1 227.9 152.9 227.1 ;
      RECT  153.7 227.9 154.5 227.1 ;
      RECT  153.7 227.9 154.5 227.1 ;
      RECT  152.1 227.9 152.9 227.1 ;
      RECT  152.1 235.3 152.9 234.5 ;
      RECT  153.7 235.3 154.5 234.5 ;
      RECT  153.7 235.3 154.5 234.5 ;
      RECT  152.1 235.3 152.9 234.5 ;
      RECT  155.3 227.5 156.1 226.7 ;
      RECT  155.3 235.3 156.1 234.5 ;
      RECT  152.3 231.6 153.1 230.8 ;
      RECT  152.3 231.6 153.1 230.8 ;
      RECT  154.1 231.5 154.7 230.9 ;
      RECT  150.9 226.1 157.3 225.5 ;
      RECT  150.9 236.5 157.3 235.9 ;
      RECT  155.3 245.3 156.1 246.6 ;
      RECT  155.3 236.2 156.1 237.5 ;
      RECT  152.1 237.1 152.9 235.9 ;
      RECT  152.1 244.5 152.9 246.9 ;
      RECT  153.8 237.1 154.4 245.3 ;
      RECT  152.1 244.5 152.9 245.3 ;
      RECT  153.7 244.5 154.5 245.3 ;
      RECT  153.7 244.5 154.5 245.3 ;
      RECT  152.1 244.5 152.9 245.3 ;
      RECT  152.1 237.1 152.9 237.9 ;
      RECT  153.7 237.1 154.5 237.9 ;
      RECT  153.7 237.1 154.5 237.9 ;
      RECT  152.1 237.1 152.9 237.9 ;
      RECT  155.3 244.9 156.1 245.7 ;
      RECT  155.3 237.1 156.1 237.9 ;
      RECT  152.3 240.8 153.1 241.6 ;
      RECT  152.3 240.8 153.1 241.6 ;
      RECT  154.1 240.9 154.7 241.5 ;
      RECT  150.9 246.3 157.3 246.9 ;
      RECT  150.9 235.9 157.3 236.5 ;
      RECT  155.3 247.9 156.1 246.6 ;
      RECT  155.3 257.0 156.1 255.7 ;
      RECT  152.1 256.1 152.9 257.3 ;
      RECT  152.1 248.7 152.9 246.3 ;
      RECT  153.8 256.1 154.4 247.9 ;
      RECT  152.1 248.7 152.9 247.9 ;
      RECT  153.7 248.7 154.5 247.9 ;
      RECT  153.7 248.7 154.5 247.9 ;
      RECT  152.1 248.7 152.9 247.9 ;
      RECT  152.1 256.1 152.9 255.3 ;
      RECT  153.7 256.1 154.5 255.3 ;
      RECT  153.7 256.1 154.5 255.3 ;
      RECT  152.1 256.1 152.9 255.3 ;
      RECT  155.3 248.3 156.1 247.5 ;
      RECT  155.3 256.1 156.1 255.3 ;
      RECT  152.3 252.4 153.1 251.6 ;
      RECT  152.3 252.4 153.1 251.6 ;
      RECT  154.1 252.3 154.7 251.7 ;
      RECT  150.9 246.9 157.3 246.3 ;
      RECT  150.9 257.3 157.3 256.7 ;
      RECT  155.3 266.1 156.1 267.4 ;
      RECT  155.3 257.0 156.1 258.3 ;
      RECT  152.1 257.9 152.9 256.7 ;
      RECT  152.1 265.3 152.9 267.7 ;
      RECT  153.8 257.9 154.4 266.1 ;
      RECT  152.1 265.3 152.9 266.1 ;
      RECT  153.7 265.3 154.5 266.1 ;
      RECT  153.7 265.3 154.5 266.1 ;
      RECT  152.1 265.3 152.9 266.1 ;
      RECT  152.1 257.9 152.9 258.7 ;
      RECT  153.7 257.9 154.5 258.7 ;
      RECT  153.7 257.9 154.5 258.7 ;
      RECT  152.1 257.9 152.9 258.7 ;
      RECT  155.3 265.7 156.1 266.5 ;
      RECT  155.3 257.9 156.1 258.7 ;
      RECT  152.3 261.6 153.1 262.4 ;
      RECT  152.3 261.6 153.1 262.4 ;
      RECT  154.1 261.7 154.7 262.3 ;
      RECT  150.9 267.1 157.3 267.7 ;
      RECT  150.9 256.7 157.3 257.3 ;
      RECT  155.3 268.7 156.1 267.4 ;
      RECT  155.3 277.8 156.1 276.5 ;
      RECT  152.1 276.9 152.9 278.1 ;
      RECT  152.1 269.5 152.9 267.1 ;
      RECT  153.8 276.9 154.4 268.7 ;
      RECT  152.1 269.5 152.9 268.7 ;
      RECT  153.7 269.5 154.5 268.7 ;
      RECT  153.7 269.5 154.5 268.7 ;
      RECT  152.1 269.5 152.9 268.7 ;
      RECT  152.1 276.9 152.9 276.1 ;
      RECT  153.7 276.9 154.5 276.1 ;
      RECT  153.7 276.9 154.5 276.1 ;
      RECT  152.1 276.9 152.9 276.1 ;
      RECT  155.3 269.1 156.1 268.3 ;
      RECT  155.3 276.9 156.1 276.1 ;
      RECT  152.3 273.2 153.1 272.4 ;
      RECT  152.3 273.2 153.1 272.4 ;
      RECT  154.1 273.1 154.7 272.5 ;
      RECT  150.9 267.7 157.3 267.1 ;
      RECT  150.9 278.1 157.3 277.5 ;
      RECT  155.3 286.9 156.1 288.2 ;
      RECT  155.3 277.8 156.1 279.1 ;
      RECT  152.1 278.7 152.9 277.5 ;
      RECT  152.1 286.1 152.9 288.5 ;
      RECT  153.8 278.7 154.4 286.9 ;
      RECT  152.1 286.1 152.9 286.9 ;
      RECT  153.7 286.1 154.5 286.9 ;
      RECT  153.7 286.1 154.5 286.9 ;
      RECT  152.1 286.1 152.9 286.9 ;
      RECT  152.1 278.7 152.9 279.5 ;
      RECT  153.7 278.7 154.5 279.5 ;
      RECT  153.7 278.7 154.5 279.5 ;
      RECT  152.1 278.7 152.9 279.5 ;
      RECT  155.3 286.5 156.1 287.3 ;
      RECT  155.3 278.7 156.1 279.5 ;
      RECT  152.3 282.4 153.1 283.2 ;
      RECT  152.3 282.4 153.1 283.2 ;
      RECT  154.1 282.5 154.7 283.1 ;
      RECT  150.9 287.9 157.3 288.5 ;
      RECT  150.9 277.5 157.3 278.1 ;
      RECT  155.3 289.5 156.1 288.2 ;
      RECT  155.3 298.6 156.1 297.3 ;
      RECT  152.1 297.7 152.9 298.9 ;
      RECT  152.1 290.3 152.9 287.9 ;
      RECT  153.8 297.7 154.4 289.5 ;
      RECT  152.1 290.3 152.9 289.5 ;
      RECT  153.7 290.3 154.5 289.5 ;
      RECT  153.7 290.3 154.5 289.5 ;
      RECT  152.1 290.3 152.9 289.5 ;
      RECT  152.1 297.7 152.9 296.9 ;
      RECT  153.7 297.7 154.5 296.9 ;
      RECT  153.7 297.7 154.5 296.9 ;
      RECT  152.1 297.7 152.9 296.9 ;
      RECT  155.3 289.9 156.1 289.1 ;
      RECT  155.3 297.7 156.1 296.9 ;
      RECT  152.3 294.0 153.1 293.2 ;
      RECT  152.3 294.0 153.1 293.2 ;
      RECT  154.1 293.9 154.7 293.3 ;
      RECT  150.9 288.5 157.3 287.9 ;
      RECT  150.9 298.9 157.3 298.3 ;
      RECT  155.3 307.7 156.1 309.0 ;
      RECT  155.3 298.6 156.1 299.9 ;
      RECT  152.1 299.5 152.9 298.3 ;
      RECT  152.1 306.9 152.9 309.3 ;
      RECT  153.8 299.5 154.4 307.7 ;
      RECT  152.1 306.9 152.9 307.7 ;
      RECT  153.7 306.9 154.5 307.7 ;
      RECT  153.7 306.9 154.5 307.7 ;
      RECT  152.1 306.9 152.9 307.7 ;
      RECT  152.1 299.5 152.9 300.3 ;
      RECT  153.7 299.5 154.5 300.3 ;
      RECT  153.7 299.5 154.5 300.3 ;
      RECT  152.1 299.5 152.9 300.3 ;
      RECT  155.3 307.3 156.1 308.1 ;
      RECT  155.3 299.5 156.1 300.3 ;
      RECT  152.3 303.2 153.1 304.0 ;
      RECT  152.3 303.2 153.1 304.0 ;
      RECT  154.1 303.3 154.7 303.9 ;
      RECT  150.9 308.7 157.3 309.3 ;
      RECT  150.9 298.3 157.3 298.9 ;
      RECT  155.3 310.3 156.1 309.0 ;
      RECT  155.3 319.4 156.1 318.1 ;
      RECT  152.1 318.5 152.9 319.7 ;
      RECT  152.1 311.1 152.9 308.7 ;
      RECT  153.8 318.5 154.4 310.3 ;
      RECT  152.1 311.1 152.9 310.3 ;
      RECT  153.7 311.1 154.5 310.3 ;
      RECT  153.7 311.1 154.5 310.3 ;
      RECT  152.1 311.1 152.9 310.3 ;
      RECT  152.1 318.5 152.9 317.7 ;
      RECT  153.7 318.5 154.5 317.7 ;
      RECT  153.7 318.5 154.5 317.7 ;
      RECT  152.1 318.5 152.9 317.7 ;
      RECT  155.3 310.7 156.1 309.9 ;
      RECT  155.3 318.5 156.1 317.7 ;
      RECT  152.3 314.8 153.1 314.0 ;
      RECT  152.3 314.8 153.1 314.0 ;
      RECT  154.1 314.7 154.7 314.1 ;
      RECT  150.9 309.3 157.3 308.7 ;
      RECT  150.9 319.7 157.3 319.1 ;
      RECT  155.3 328.5 156.1 329.8 ;
      RECT  155.3 319.4 156.1 320.7 ;
      RECT  152.1 320.3 152.9 319.1 ;
      RECT  152.1 327.7 152.9 330.1 ;
      RECT  153.8 320.3 154.4 328.5 ;
      RECT  152.1 327.7 152.9 328.5 ;
      RECT  153.7 327.7 154.5 328.5 ;
      RECT  153.7 327.7 154.5 328.5 ;
      RECT  152.1 327.7 152.9 328.5 ;
      RECT  152.1 320.3 152.9 321.1 ;
      RECT  153.7 320.3 154.5 321.1 ;
      RECT  153.7 320.3 154.5 321.1 ;
      RECT  152.1 320.3 152.9 321.1 ;
      RECT  155.3 328.1 156.1 328.9 ;
      RECT  155.3 320.3 156.1 321.1 ;
      RECT  152.3 324.0 153.1 324.8 ;
      RECT  152.3 324.0 153.1 324.8 ;
      RECT  154.1 324.1 154.7 324.7 ;
      RECT  150.9 329.5 157.3 330.1 ;
      RECT  150.9 319.1 157.3 319.7 ;
      RECT  155.3 331.1 156.1 329.8 ;
      RECT  155.3 340.2 156.1 338.9 ;
      RECT  152.1 339.3 152.9 340.5 ;
      RECT  152.1 331.9 152.9 329.5 ;
      RECT  153.8 339.3 154.4 331.1 ;
      RECT  152.1 331.9 152.9 331.1 ;
      RECT  153.7 331.9 154.5 331.1 ;
      RECT  153.7 331.9 154.5 331.1 ;
      RECT  152.1 331.9 152.9 331.1 ;
      RECT  152.1 339.3 152.9 338.5 ;
      RECT  153.7 339.3 154.5 338.5 ;
      RECT  153.7 339.3 154.5 338.5 ;
      RECT  152.1 339.3 152.9 338.5 ;
      RECT  155.3 331.5 156.1 330.7 ;
      RECT  155.3 339.3 156.1 338.5 ;
      RECT  152.3 335.6 153.1 334.8 ;
      RECT  152.3 335.6 153.1 334.8 ;
      RECT  154.1 335.5 154.7 334.9 ;
      RECT  150.9 330.1 157.3 329.5 ;
      RECT  150.9 340.5 157.3 339.9 ;
      RECT  155.3 349.3 156.1 350.6 ;
      RECT  155.3 340.2 156.1 341.5 ;
      RECT  152.1 341.1 152.9 339.9 ;
      RECT  152.1 348.5 152.9 350.9 ;
      RECT  153.8 341.1 154.4 349.3 ;
      RECT  152.1 348.5 152.9 349.3 ;
      RECT  153.7 348.5 154.5 349.3 ;
      RECT  153.7 348.5 154.5 349.3 ;
      RECT  152.1 348.5 152.9 349.3 ;
      RECT  152.1 341.1 152.9 341.9 ;
      RECT  153.7 341.1 154.5 341.9 ;
      RECT  153.7 341.1 154.5 341.9 ;
      RECT  152.1 341.1 152.9 341.9 ;
      RECT  155.3 348.9 156.1 349.7 ;
      RECT  155.3 341.1 156.1 341.9 ;
      RECT  152.3 344.8 153.1 345.6 ;
      RECT  152.3 344.8 153.1 345.6 ;
      RECT  154.1 344.9 154.7 345.5 ;
      RECT  150.9 350.3 157.3 350.9 ;
      RECT  150.9 339.9 157.3 340.5 ;
      RECT  155.3 351.9 156.1 350.6 ;
      RECT  155.3 361.0 156.1 359.7 ;
      RECT  152.1 360.1 152.9 361.3 ;
      RECT  152.1 352.7 152.9 350.3 ;
      RECT  153.8 360.1 154.4 351.9 ;
      RECT  152.1 352.7 152.9 351.9 ;
      RECT  153.7 352.7 154.5 351.9 ;
      RECT  153.7 352.7 154.5 351.9 ;
      RECT  152.1 352.7 152.9 351.9 ;
      RECT  152.1 360.1 152.9 359.3 ;
      RECT  153.7 360.1 154.5 359.3 ;
      RECT  153.7 360.1 154.5 359.3 ;
      RECT  152.1 360.1 152.9 359.3 ;
      RECT  155.3 352.3 156.1 351.5 ;
      RECT  155.3 360.1 156.1 359.3 ;
      RECT  152.3 356.4 153.1 355.6 ;
      RECT  152.3 356.4 153.1 355.6 ;
      RECT  154.1 356.3 154.7 355.7 ;
      RECT  150.9 350.9 157.3 350.3 ;
      RECT  150.9 361.3 157.3 360.7 ;
      RECT  126.8 199.2 127.6 200.0 ;
      RECT  126.8 210.0 127.6 210.8 ;
      RECT  126.8 220.0 127.6 220.8 ;
      RECT  126.8 230.8 127.6 231.6 ;
      RECT  126.8 240.8 127.6 241.6 ;
      RECT  126.8 251.6 127.6 252.4 ;
      RECT  126.8 261.6 127.6 262.4 ;
      RECT  126.8 272.4 127.6 273.2 ;
      RECT  130.3 199.0 131.1 199.8 ;
      RECT  135.9 197.6 136.7 198.4 ;
      RECT  131.7 210.2 132.5 211.0 ;
      RECT  135.9 211.6 136.7 212.4 ;
      RECT  133.1 219.8 133.9 220.6 ;
      RECT  135.9 218.4 136.7 219.2 ;
      RECT  134.5 231.0 135.3 231.8 ;
      RECT  135.9 232.4 136.7 233.2 ;
      RECT  130.3 240.6 131.1 241.4 ;
      RECT  137.3 239.2 138.1 240.0 ;
      RECT  131.7 251.8 132.5 252.6 ;
      RECT  137.3 253.2 138.1 254.0 ;
      RECT  133.1 261.4 133.9 262.2 ;
      RECT  137.3 260.0 138.1 260.8 ;
      RECT  134.5 272.6 135.3 273.4 ;
      RECT  137.3 274.0 138.1 274.8 ;
      RECT  130.3 282.2 131.1 283.0 ;
      RECT  138.7 280.8 139.5 281.6 ;
      RECT  131.7 293.4 132.5 294.2 ;
      RECT  138.7 294.8 139.5 295.6 ;
      RECT  133.1 303.0 133.9 303.8 ;
      RECT  138.7 301.6 139.5 302.4 ;
      RECT  134.5 314.2 135.3 315.0 ;
      RECT  138.7 315.6 139.5 316.4 ;
      RECT  130.3 323.8 131.1 324.6 ;
      RECT  140.1 322.4 140.9 323.2 ;
      RECT  131.7 335.0 132.5 335.8 ;
      RECT  140.1 336.4 140.9 337.2 ;
      RECT  133.1 344.6 133.9 345.4 ;
      RECT  140.1 343.2 140.9 344.0 ;
      RECT  134.5 355.8 135.3 356.6 ;
      RECT  140.1 357.2 140.9 358.0 ;
      RECT  145.7 204.6 146.5 205.4 ;
      RECT  145.7 194.2 146.5 195.0 ;
      RECT  145.7 204.6 146.5 205.4 ;
      RECT  145.7 215.0 146.5 215.8 ;
      RECT  145.7 225.4 146.5 226.2 ;
      RECT  145.7 215.0 146.5 215.8 ;
      RECT  145.7 225.4 146.5 226.2 ;
      RECT  145.7 235.8 146.5 236.6 ;
      RECT  145.7 246.2 146.5 247.0 ;
      RECT  145.7 235.8 146.5 236.6 ;
      RECT  145.7 246.2 146.5 247.0 ;
      RECT  145.7 256.6 146.5 257.4 ;
      RECT  145.7 267.0 146.5 267.8 ;
      RECT  145.7 256.6 146.5 257.4 ;
      RECT  145.7 267.0 146.5 267.8 ;
      RECT  145.7 277.4 146.5 278.2 ;
      RECT  145.7 287.8 146.5 288.6 ;
      RECT  145.7 277.4 146.5 278.2 ;
      RECT  145.7 287.8 146.5 288.6 ;
      RECT  145.7 298.2 146.5 299.0 ;
      RECT  145.7 308.6 146.5 309.4 ;
      RECT  145.7 298.2 146.5 299.0 ;
      RECT  145.7 308.6 146.5 309.4 ;
      RECT  145.7 319.0 146.5 319.8 ;
      RECT  145.7 329.4 146.5 330.2 ;
      RECT  145.7 319.0 146.5 319.8 ;
      RECT  145.7 329.4 146.5 330.2 ;
      RECT  145.7 339.8 146.5 340.6 ;
      RECT  145.7 350.2 146.5 351.0 ;
      RECT  145.7 339.8 146.5 340.6 ;
      RECT  145.7 350.2 146.5 351.0 ;
      RECT  145.7 360.6 146.5 361.4 ;
      RECT  154.1 199.3 154.7 199.9 ;
      RECT  154.1 210.1 154.7 210.7 ;
      RECT  154.1 220.1 154.7 220.7 ;
      RECT  154.1 230.9 154.7 231.5 ;
      RECT  154.1 240.9 154.7 241.5 ;
      RECT  154.1 251.7 154.7 252.3 ;
      RECT  154.1 261.7 154.7 262.3 ;
      RECT  154.1 272.5 154.7 273.1 ;
      RECT  154.1 282.5 154.7 283.1 ;
      RECT  154.1 293.3 154.7 293.9 ;
      RECT  154.1 303.3 154.7 303.9 ;
      RECT  154.1 314.1 154.7 314.7 ;
      RECT  154.1 324.1 154.7 324.7 ;
      RECT  154.1 334.9 154.7 335.5 ;
      RECT  154.1 344.9 154.7 345.5 ;
      RECT  154.1 355.7 154.7 356.3 ;
      RECT  161.8 199.1 165.5 199.7 ;
      RECT  172.4 199.1 173.0 199.7 ;
      RECT  172.4 199.3 173.0 199.9 ;
      RECT  170.5 199.1 172.7 199.7 ;
      RECT  172.4 199.4 173.0 199.6 ;
      RECT  172.7 199.3 174.9 199.9 ;
      RECT  161.8 210.3 165.5 210.9 ;
      RECT  172.4 210.3 173.0 210.9 ;
      RECT  172.4 210.1 173.0 210.7 ;
      RECT  170.5 210.3 172.7 210.9 ;
      RECT  172.4 210.4 173.0 210.6 ;
      RECT  172.7 210.1 174.9 210.7 ;
      RECT  161.8 219.9 165.5 220.5 ;
      RECT  172.4 219.9 173.0 220.5 ;
      RECT  172.4 220.1 173.0 220.7 ;
      RECT  170.5 219.9 172.7 220.5 ;
      RECT  172.4 220.2 173.0 220.4 ;
      RECT  172.7 220.1 174.9 220.7 ;
      RECT  161.8 231.1 165.5 231.7 ;
      RECT  172.4 231.1 173.0 231.7 ;
      RECT  172.4 230.9 173.0 231.5 ;
      RECT  170.5 231.1 172.7 231.7 ;
      RECT  172.4 231.2 173.0 231.4 ;
      RECT  172.7 230.9 174.9 231.5 ;
      RECT  161.8 240.7 165.5 241.3 ;
      RECT  172.4 240.7 173.0 241.3 ;
      RECT  172.4 240.9 173.0 241.5 ;
      RECT  170.5 240.7 172.7 241.3 ;
      RECT  172.4 241.0 173.0 241.2 ;
      RECT  172.7 240.9 174.9 241.5 ;
      RECT  161.8 251.9 165.5 252.5 ;
      RECT  172.4 251.9 173.0 252.5 ;
      RECT  172.4 251.7 173.0 252.3 ;
      RECT  170.5 251.9 172.7 252.5 ;
      RECT  172.4 252.0 173.0 252.2 ;
      RECT  172.7 251.7 174.9 252.3 ;
      RECT  161.8 261.5 165.5 262.1 ;
      RECT  172.4 261.5 173.0 262.1 ;
      RECT  172.4 261.7 173.0 262.3 ;
      RECT  170.5 261.5 172.7 262.1 ;
      RECT  172.4 261.8 173.0 262.0 ;
      RECT  172.7 261.7 174.9 262.3 ;
      RECT  161.8 272.7 165.5 273.3 ;
      RECT  172.4 272.7 173.0 273.3 ;
      RECT  172.4 272.5 173.0 273.1 ;
      RECT  170.5 272.7 172.7 273.3 ;
      RECT  172.4 272.8 173.0 273.0 ;
      RECT  172.7 272.5 174.9 273.1 ;
      RECT  161.8 282.3 165.5 282.9 ;
      RECT  172.4 282.3 173.0 282.9 ;
      RECT  172.4 282.5 173.0 283.1 ;
      RECT  170.5 282.3 172.7 282.9 ;
      RECT  172.4 282.6 173.0 282.8 ;
      RECT  172.7 282.5 174.9 283.1 ;
      RECT  161.8 293.5 165.5 294.1 ;
      RECT  172.4 293.5 173.0 294.1 ;
      RECT  172.4 293.3 173.0 293.9 ;
      RECT  170.5 293.5 172.7 294.1 ;
      RECT  172.4 293.6 173.0 293.8 ;
      RECT  172.7 293.3 174.9 293.9 ;
      RECT  161.8 303.1 165.5 303.7 ;
      RECT  172.4 303.1 173.0 303.7 ;
      RECT  172.4 303.3 173.0 303.9 ;
      RECT  170.5 303.1 172.7 303.7 ;
      RECT  172.4 303.4 173.0 303.6 ;
      RECT  172.7 303.3 174.9 303.9 ;
      RECT  161.8 314.3 165.5 314.9 ;
      RECT  172.4 314.3 173.0 314.9 ;
      RECT  172.4 314.1 173.0 314.7 ;
      RECT  170.5 314.3 172.7 314.9 ;
      RECT  172.4 314.4 173.0 314.6 ;
      RECT  172.7 314.1 174.9 314.7 ;
      RECT  161.8 323.9 165.5 324.5 ;
      RECT  172.4 323.9 173.0 324.5 ;
      RECT  172.4 324.1 173.0 324.7 ;
      RECT  170.5 323.9 172.7 324.5 ;
      RECT  172.4 324.2 173.0 324.4 ;
      RECT  172.7 324.1 174.9 324.7 ;
      RECT  161.8 335.1 165.5 335.7 ;
      RECT  172.4 335.1 173.0 335.7 ;
      RECT  172.4 334.9 173.0 335.5 ;
      RECT  170.5 335.1 172.7 335.7 ;
      RECT  172.4 335.2 173.0 335.4 ;
      RECT  172.7 334.9 174.9 335.5 ;
      RECT  161.8 344.7 165.5 345.3 ;
      RECT  172.4 344.7 173.0 345.3 ;
      RECT  172.4 344.9 173.0 345.5 ;
      RECT  170.5 344.7 172.7 345.3 ;
      RECT  172.4 345.0 173.0 345.2 ;
      RECT  172.7 344.9 174.9 345.5 ;
      RECT  161.8 355.9 165.5 356.5 ;
      RECT  172.4 355.9 173.0 356.5 ;
      RECT  172.4 355.7 173.0 356.3 ;
      RECT  170.5 355.9 172.7 356.5 ;
      RECT  172.4 356.0 173.0 356.2 ;
      RECT  172.7 355.7 174.9 356.3 ;
      RECT  165.1 195.9 165.9 194.3 ;
      RECT  165.1 202.9 165.9 205.3 ;
      RECT  168.3 202.9 169.1 205.3 ;
      RECT  169.9 203.7 170.7 205.0 ;
      RECT  169.9 194.6 170.7 195.9 ;
      RECT  165.1 202.9 165.9 203.7 ;
      RECT  166.7 202.9 167.5 203.7 ;
      RECT  166.7 202.9 167.5 203.7 ;
      RECT  165.1 202.9 165.9 203.7 ;
      RECT  166.7 202.9 167.5 203.7 ;
      RECT  168.3 202.9 169.1 203.7 ;
      RECT  168.3 202.9 169.1 203.7 ;
      RECT  166.7 202.9 167.5 203.7 ;
      RECT  165.1 195.9 165.9 196.7 ;
      RECT  166.7 195.9 167.5 196.7 ;
      RECT  166.7 195.9 167.5 196.7 ;
      RECT  165.1 195.9 165.9 196.7 ;
      RECT  166.7 195.9 167.5 196.7 ;
      RECT  168.3 195.9 169.1 196.7 ;
      RECT  168.3 195.9 169.1 196.7 ;
      RECT  166.7 195.9 167.5 196.7 ;
      RECT  169.9 203.3 170.7 204.1 ;
      RECT  169.9 195.5 170.7 196.3 ;
      RECT  167.5 197.6 168.3 198.4 ;
      RECT  165.5 199.0 166.3 199.8 ;
      RECT  166.7 202.9 167.5 203.7 ;
      RECT  168.3 195.9 169.1 196.7 ;
      RECT  169.7 199.0 170.5 199.8 ;
      RECT  165.5 199.0 166.3 199.8 ;
      RECT  167.5 197.6 168.3 198.4 ;
      RECT  169.7 199.0 170.5 199.8 ;
      RECT  163.9 204.7 173.5 205.3 ;
      RECT  163.9 194.3 173.5 194.9 ;
      RECT  177.9 203.7 178.7 205.0 ;
      RECT  177.9 194.6 178.7 195.9 ;
      RECT  174.7 195.5 175.5 194.3 ;
      RECT  174.7 202.9 175.5 205.3 ;
      RECT  176.4 195.5 177.0 203.7 ;
      RECT  174.7 202.9 175.5 203.7 ;
      RECT  176.3 202.9 177.1 203.7 ;
      RECT  176.3 202.9 177.1 203.7 ;
      RECT  174.7 202.9 175.5 203.7 ;
      RECT  174.7 195.5 175.5 196.3 ;
      RECT  176.3 195.5 177.1 196.3 ;
      RECT  176.3 195.5 177.1 196.3 ;
      RECT  174.7 195.5 175.5 196.3 ;
      RECT  177.9 203.3 178.7 204.1 ;
      RECT  177.9 195.5 178.7 196.3 ;
      RECT  174.9 199.2 175.7 200.0 ;
      RECT  174.9 199.2 175.7 200.0 ;
      RECT  176.7 199.3 177.3 199.9 ;
      RECT  173.5 204.7 179.9 205.3 ;
      RECT  173.5 194.3 179.9 194.9 ;
      RECT  174.9 199.2 175.7 200.0 ;
      RECT  176.7 199.3 177.3 199.9 ;
      RECT  173.5 204.7 174.1 205.3 ;
      RECT  173.5 194.3 174.1 194.9 ;
      RECT  165.1 214.1 165.9 215.7 ;
      RECT  165.1 207.1 165.9 204.7 ;
      RECT  168.3 207.1 169.1 204.7 ;
      RECT  169.9 206.3 170.7 205.0 ;
      RECT  169.9 215.4 170.7 214.1 ;
      RECT  165.1 207.1 165.9 206.3 ;
      RECT  166.7 207.1 167.5 206.3 ;
      RECT  166.7 207.1 167.5 206.3 ;
      RECT  165.1 207.1 165.9 206.3 ;
      RECT  166.7 207.1 167.5 206.3 ;
      RECT  168.3 207.1 169.1 206.3 ;
      RECT  168.3 207.1 169.1 206.3 ;
      RECT  166.7 207.1 167.5 206.3 ;
      RECT  165.1 214.1 165.9 213.3 ;
      RECT  166.7 214.1 167.5 213.3 ;
      RECT  166.7 214.1 167.5 213.3 ;
      RECT  165.1 214.1 165.9 213.3 ;
      RECT  166.7 214.1 167.5 213.3 ;
      RECT  168.3 214.1 169.1 213.3 ;
      RECT  168.3 214.1 169.1 213.3 ;
      RECT  166.7 214.1 167.5 213.3 ;
      RECT  169.9 206.7 170.7 205.9 ;
      RECT  169.9 214.5 170.7 213.7 ;
      RECT  167.5 212.4 168.3 211.6 ;
      RECT  165.5 211.0 166.3 210.2 ;
      RECT  166.7 207.1 167.5 206.3 ;
      RECT  168.3 214.1 169.1 213.3 ;
      RECT  169.7 211.0 170.5 210.2 ;
      RECT  165.5 211.0 166.3 210.2 ;
      RECT  167.5 212.4 168.3 211.6 ;
      RECT  169.7 211.0 170.5 210.2 ;
      RECT  163.9 205.3 173.5 204.7 ;
      RECT  163.9 215.7 173.5 215.1 ;
      RECT  177.9 206.3 178.7 205.0 ;
      RECT  177.9 215.4 178.7 214.1 ;
      RECT  174.7 214.5 175.5 215.7 ;
      RECT  174.7 207.1 175.5 204.7 ;
      RECT  176.4 214.5 177.0 206.3 ;
      RECT  174.7 207.1 175.5 206.3 ;
      RECT  176.3 207.1 177.1 206.3 ;
      RECT  176.3 207.1 177.1 206.3 ;
      RECT  174.7 207.1 175.5 206.3 ;
      RECT  174.7 214.5 175.5 213.7 ;
      RECT  176.3 214.5 177.1 213.7 ;
      RECT  176.3 214.5 177.1 213.7 ;
      RECT  174.7 214.5 175.5 213.7 ;
      RECT  177.9 206.7 178.7 205.9 ;
      RECT  177.9 214.5 178.7 213.7 ;
      RECT  174.9 210.8 175.7 210.0 ;
      RECT  174.9 210.8 175.7 210.0 ;
      RECT  176.7 210.7 177.3 210.1 ;
      RECT  173.5 205.3 179.9 204.7 ;
      RECT  173.5 215.7 179.9 215.1 ;
      RECT  174.9 210.8 175.7 210.0 ;
      RECT  176.7 210.7 177.3 210.1 ;
      RECT  173.5 205.3 174.1 204.7 ;
      RECT  173.5 215.7 174.1 215.1 ;
      RECT  165.1 216.7 165.9 215.1 ;
      RECT  165.1 223.7 165.9 226.1 ;
      RECT  168.3 223.7 169.1 226.1 ;
      RECT  169.9 224.5 170.7 225.8 ;
      RECT  169.9 215.4 170.7 216.7 ;
      RECT  165.1 223.7 165.9 224.5 ;
      RECT  166.7 223.7 167.5 224.5 ;
      RECT  166.7 223.7 167.5 224.5 ;
      RECT  165.1 223.7 165.9 224.5 ;
      RECT  166.7 223.7 167.5 224.5 ;
      RECT  168.3 223.7 169.1 224.5 ;
      RECT  168.3 223.7 169.1 224.5 ;
      RECT  166.7 223.7 167.5 224.5 ;
      RECT  165.1 216.7 165.9 217.5 ;
      RECT  166.7 216.7 167.5 217.5 ;
      RECT  166.7 216.7 167.5 217.5 ;
      RECT  165.1 216.7 165.9 217.5 ;
      RECT  166.7 216.7 167.5 217.5 ;
      RECT  168.3 216.7 169.1 217.5 ;
      RECT  168.3 216.7 169.1 217.5 ;
      RECT  166.7 216.7 167.5 217.5 ;
      RECT  169.9 224.1 170.7 224.9 ;
      RECT  169.9 216.3 170.7 217.1 ;
      RECT  167.5 218.4 168.3 219.2 ;
      RECT  165.5 219.8 166.3 220.6 ;
      RECT  166.7 223.7 167.5 224.5 ;
      RECT  168.3 216.7 169.1 217.5 ;
      RECT  169.7 219.8 170.5 220.6 ;
      RECT  165.5 219.8 166.3 220.6 ;
      RECT  167.5 218.4 168.3 219.2 ;
      RECT  169.7 219.8 170.5 220.6 ;
      RECT  163.9 225.5 173.5 226.1 ;
      RECT  163.9 215.1 173.5 215.7 ;
      RECT  177.9 224.5 178.7 225.8 ;
      RECT  177.9 215.4 178.7 216.7 ;
      RECT  174.7 216.3 175.5 215.1 ;
      RECT  174.7 223.7 175.5 226.1 ;
      RECT  176.4 216.3 177.0 224.5 ;
      RECT  174.7 223.7 175.5 224.5 ;
      RECT  176.3 223.7 177.1 224.5 ;
      RECT  176.3 223.7 177.1 224.5 ;
      RECT  174.7 223.7 175.5 224.5 ;
      RECT  174.7 216.3 175.5 217.1 ;
      RECT  176.3 216.3 177.1 217.1 ;
      RECT  176.3 216.3 177.1 217.1 ;
      RECT  174.7 216.3 175.5 217.1 ;
      RECT  177.9 224.1 178.7 224.9 ;
      RECT  177.9 216.3 178.7 217.1 ;
      RECT  174.9 220.0 175.7 220.8 ;
      RECT  174.9 220.0 175.7 220.8 ;
      RECT  176.7 220.1 177.3 220.7 ;
      RECT  173.5 225.5 179.9 226.1 ;
      RECT  173.5 215.1 179.9 215.7 ;
      RECT  174.9 220.0 175.7 220.8 ;
      RECT  176.7 220.1 177.3 220.7 ;
      RECT  173.5 225.5 174.1 226.1 ;
      RECT  173.5 215.1 174.1 215.7 ;
      RECT  165.1 234.9 165.9 236.5 ;
      RECT  165.1 227.9 165.9 225.5 ;
      RECT  168.3 227.9 169.1 225.5 ;
      RECT  169.9 227.1 170.7 225.8 ;
      RECT  169.9 236.2 170.7 234.9 ;
      RECT  165.1 227.9 165.9 227.1 ;
      RECT  166.7 227.9 167.5 227.1 ;
      RECT  166.7 227.9 167.5 227.1 ;
      RECT  165.1 227.9 165.9 227.1 ;
      RECT  166.7 227.9 167.5 227.1 ;
      RECT  168.3 227.9 169.1 227.1 ;
      RECT  168.3 227.9 169.1 227.1 ;
      RECT  166.7 227.9 167.5 227.1 ;
      RECT  165.1 234.9 165.9 234.1 ;
      RECT  166.7 234.9 167.5 234.1 ;
      RECT  166.7 234.9 167.5 234.1 ;
      RECT  165.1 234.9 165.9 234.1 ;
      RECT  166.7 234.9 167.5 234.1 ;
      RECT  168.3 234.9 169.1 234.1 ;
      RECT  168.3 234.9 169.1 234.1 ;
      RECT  166.7 234.9 167.5 234.1 ;
      RECT  169.9 227.5 170.7 226.7 ;
      RECT  169.9 235.3 170.7 234.5 ;
      RECT  167.5 233.2 168.3 232.4 ;
      RECT  165.5 231.8 166.3 231.0 ;
      RECT  166.7 227.9 167.5 227.1 ;
      RECT  168.3 234.9 169.1 234.1 ;
      RECT  169.7 231.8 170.5 231.0 ;
      RECT  165.5 231.8 166.3 231.0 ;
      RECT  167.5 233.2 168.3 232.4 ;
      RECT  169.7 231.8 170.5 231.0 ;
      RECT  163.9 226.1 173.5 225.5 ;
      RECT  163.9 236.5 173.5 235.9 ;
      RECT  177.9 227.1 178.7 225.8 ;
      RECT  177.9 236.2 178.7 234.9 ;
      RECT  174.7 235.3 175.5 236.5 ;
      RECT  174.7 227.9 175.5 225.5 ;
      RECT  176.4 235.3 177.0 227.1 ;
      RECT  174.7 227.9 175.5 227.1 ;
      RECT  176.3 227.9 177.1 227.1 ;
      RECT  176.3 227.9 177.1 227.1 ;
      RECT  174.7 227.9 175.5 227.1 ;
      RECT  174.7 235.3 175.5 234.5 ;
      RECT  176.3 235.3 177.1 234.5 ;
      RECT  176.3 235.3 177.1 234.5 ;
      RECT  174.7 235.3 175.5 234.5 ;
      RECT  177.9 227.5 178.7 226.7 ;
      RECT  177.9 235.3 178.7 234.5 ;
      RECT  174.9 231.6 175.7 230.8 ;
      RECT  174.9 231.6 175.7 230.8 ;
      RECT  176.7 231.5 177.3 230.9 ;
      RECT  173.5 226.1 179.9 225.5 ;
      RECT  173.5 236.5 179.9 235.9 ;
      RECT  174.9 231.6 175.7 230.8 ;
      RECT  176.7 231.5 177.3 230.9 ;
      RECT  173.5 226.1 174.1 225.5 ;
      RECT  173.5 236.5 174.1 235.9 ;
      RECT  165.1 237.5 165.9 235.9 ;
      RECT  165.1 244.5 165.9 246.9 ;
      RECT  168.3 244.5 169.1 246.9 ;
      RECT  169.9 245.3 170.7 246.6 ;
      RECT  169.9 236.2 170.7 237.5 ;
      RECT  165.1 244.5 165.9 245.3 ;
      RECT  166.7 244.5 167.5 245.3 ;
      RECT  166.7 244.5 167.5 245.3 ;
      RECT  165.1 244.5 165.9 245.3 ;
      RECT  166.7 244.5 167.5 245.3 ;
      RECT  168.3 244.5 169.1 245.3 ;
      RECT  168.3 244.5 169.1 245.3 ;
      RECT  166.7 244.5 167.5 245.3 ;
      RECT  165.1 237.5 165.9 238.3 ;
      RECT  166.7 237.5 167.5 238.3 ;
      RECT  166.7 237.5 167.5 238.3 ;
      RECT  165.1 237.5 165.9 238.3 ;
      RECT  166.7 237.5 167.5 238.3 ;
      RECT  168.3 237.5 169.1 238.3 ;
      RECT  168.3 237.5 169.1 238.3 ;
      RECT  166.7 237.5 167.5 238.3 ;
      RECT  169.9 244.9 170.7 245.7 ;
      RECT  169.9 237.1 170.7 237.9 ;
      RECT  167.5 239.2 168.3 240.0 ;
      RECT  165.5 240.6 166.3 241.4 ;
      RECT  166.7 244.5 167.5 245.3 ;
      RECT  168.3 237.5 169.1 238.3 ;
      RECT  169.7 240.6 170.5 241.4 ;
      RECT  165.5 240.6 166.3 241.4 ;
      RECT  167.5 239.2 168.3 240.0 ;
      RECT  169.7 240.6 170.5 241.4 ;
      RECT  163.9 246.3 173.5 246.9 ;
      RECT  163.9 235.9 173.5 236.5 ;
      RECT  177.9 245.3 178.7 246.6 ;
      RECT  177.9 236.2 178.7 237.5 ;
      RECT  174.7 237.1 175.5 235.9 ;
      RECT  174.7 244.5 175.5 246.9 ;
      RECT  176.4 237.1 177.0 245.3 ;
      RECT  174.7 244.5 175.5 245.3 ;
      RECT  176.3 244.5 177.1 245.3 ;
      RECT  176.3 244.5 177.1 245.3 ;
      RECT  174.7 244.5 175.5 245.3 ;
      RECT  174.7 237.1 175.5 237.9 ;
      RECT  176.3 237.1 177.1 237.9 ;
      RECT  176.3 237.1 177.1 237.9 ;
      RECT  174.7 237.1 175.5 237.9 ;
      RECT  177.9 244.9 178.7 245.7 ;
      RECT  177.9 237.1 178.7 237.9 ;
      RECT  174.9 240.8 175.7 241.6 ;
      RECT  174.9 240.8 175.7 241.6 ;
      RECT  176.7 240.9 177.3 241.5 ;
      RECT  173.5 246.3 179.9 246.9 ;
      RECT  173.5 235.9 179.9 236.5 ;
      RECT  174.9 240.8 175.7 241.6 ;
      RECT  176.7 240.9 177.3 241.5 ;
      RECT  173.5 246.3 174.1 246.9 ;
      RECT  173.5 235.9 174.1 236.5 ;
      RECT  165.1 255.7 165.9 257.3 ;
      RECT  165.1 248.7 165.9 246.3 ;
      RECT  168.3 248.7 169.1 246.3 ;
      RECT  169.9 247.9 170.7 246.6 ;
      RECT  169.9 257.0 170.7 255.7 ;
      RECT  165.1 248.7 165.9 247.9 ;
      RECT  166.7 248.7 167.5 247.9 ;
      RECT  166.7 248.7 167.5 247.9 ;
      RECT  165.1 248.7 165.9 247.9 ;
      RECT  166.7 248.7 167.5 247.9 ;
      RECT  168.3 248.7 169.1 247.9 ;
      RECT  168.3 248.7 169.1 247.9 ;
      RECT  166.7 248.7 167.5 247.9 ;
      RECT  165.1 255.7 165.9 254.9 ;
      RECT  166.7 255.7 167.5 254.9 ;
      RECT  166.7 255.7 167.5 254.9 ;
      RECT  165.1 255.7 165.9 254.9 ;
      RECT  166.7 255.7 167.5 254.9 ;
      RECT  168.3 255.7 169.1 254.9 ;
      RECT  168.3 255.7 169.1 254.9 ;
      RECT  166.7 255.7 167.5 254.9 ;
      RECT  169.9 248.3 170.7 247.5 ;
      RECT  169.9 256.1 170.7 255.3 ;
      RECT  167.5 254.0 168.3 253.2 ;
      RECT  165.5 252.6 166.3 251.8 ;
      RECT  166.7 248.7 167.5 247.9 ;
      RECT  168.3 255.7 169.1 254.9 ;
      RECT  169.7 252.6 170.5 251.8 ;
      RECT  165.5 252.6 166.3 251.8 ;
      RECT  167.5 254.0 168.3 253.2 ;
      RECT  169.7 252.6 170.5 251.8 ;
      RECT  163.9 246.9 173.5 246.3 ;
      RECT  163.9 257.3 173.5 256.7 ;
      RECT  177.9 247.9 178.7 246.6 ;
      RECT  177.9 257.0 178.7 255.7 ;
      RECT  174.7 256.1 175.5 257.3 ;
      RECT  174.7 248.7 175.5 246.3 ;
      RECT  176.4 256.1 177.0 247.9 ;
      RECT  174.7 248.7 175.5 247.9 ;
      RECT  176.3 248.7 177.1 247.9 ;
      RECT  176.3 248.7 177.1 247.9 ;
      RECT  174.7 248.7 175.5 247.9 ;
      RECT  174.7 256.1 175.5 255.3 ;
      RECT  176.3 256.1 177.1 255.3 ;
      RECT  176.3 256.1 177.1 255.3 ;
      RECT  174.7 256.1 175.5 255.3 ;
      RECT  177.9 248.3 178.7 247.5 ;
      RECT  177.9 256.1 178.7 255.3 ;
      RECT  174.9 252.4 175.7 251.6 ;
      RECT  174.9 252.4 175.7 251.6 ;
      RECT  176.7 252.3 177.3 251.7 ;
      RECT  173.5 246.9 179.9 246.3 ;
      RECT  173.5 257.3 179.9 256.7 ;
      RECT  174.9 252.4 175.7 251.6 ;
      RECT  176.7 252.3 177.3 251.7 ;
      RECT  173.5 246.9 174.1 246.3 ;
      RECT  173.5 257.3 174.1 256.7 ;
      RECT  165.1 258.3 165.9 256.7 ;
      RECT  165.1 265.3 165.9 267.7 ;
      RECT  168.3 265.3 169.1 267.7 ;
      RECT  169.9 266.1 170.7 267.4 ;
      RECT  169.9 257.0 170.7 258.3 ;
      RECT  165.1 265.3 165.9 266.1 ;
      RECT  166.7 265.3 167.5 266.1 ;
      RECT  166.7 265.3 167.5 266.1 ;
      RECT  165.1 265.3 165.9 266.1 ;
      RECT  166.7 265.3 167.5 266.1 ;
      RECT  168.3 265.3 169.1 266.1 ;
      RECT  168.3 265.3 169.1 266.1 ;
      RECT  166.7 265.3 167.5 266.1 ;
      RECT  165.1 258.3 165.9 259.1 ;
      RECT  166.7 258.3 167.5 259.1 ;
      RECT  166.7 258.3 167.5 259.1 ;
      RECT  165.1 258.3 165.9 259.1 ;
      RECT  166.7 258.3 167.5 259.1 ;
      RECT  168.3 258.3 169.1 259.1 ;
      RECT  168.3 258.3 169.1 259.1 ;
      RECT  166.7 258.3 167.5 259.1 ;
      RECT  169.9 265.7 170.7 266.5 ;
      RECT  169.9 257.9 170.7 258.7 ;
      RECT  167.5 260.0 168.3 260.8 ;
      RECT  165.5 261.4 166.3 262.2 ;
      RECT  166.7 265.3 167.5 266.1 ;
      RECT  168.3 258.3 169.1 259.1 ;
      RECT  169.7 261.4 170.5 262.2 ;
      RECT  165.5 261.4 166.3 262.2 ;
      RECT  167.5 260.0 168.3 260.8 ;
      RECT  169.7 261.4 170.5 262.2 ;
      RECT  163.9 267.1 173.5 267.7 ;
      RECT  163.9 256.7 173.5 257.3 ;
      RECT  177.9 266.1 178.7 267.4 ;
      RECT  177.9 257.0 178.7 258.3 ;
      RECT  174.7 257.9 175.5 256.7 ;
      RECT  174.7 265.3 175.5 267.7 ;
      RECT  176.4 257.9 177.0 266.1 ;
      RECT  174.7 265.3 175.5 266.1 ;
      RECT  176.3 265.3 177.1 266.1 ;
      RECT  176.3 265.3 177.1 266.1 ;
      RECT  174.7 265.3 175.5 266.1 ;
      RECT  174.7 257.9 175.5 258.7 ;
      RECT  176.3 257.9 177.1 258.7 ;
      RECT  176.3 257.9 177.1 258.7 ;
      RECT  174.7 257.9 175.5 258.7 ;
      RECT  177.9 265.7 178.7 266.5 ;
      RECT  177.9 257.9 178.7 258.7 ;
      RECT  174.9 261.6 175.7 262.4 ;
      RECT  174.9 261.6 175.7 262.4 ;
      RECT  176.7 261.7 177.3 262.3 ;
      RECT  173.5 267.1 179.9 267.7 ;
      RECT  173.5 256.7 179.9 257.3 ;
      RECT  174.9 261.6 175.7 262.4 ;
      RECT  176.7 261.7 177.3 262.3 ;
      RECT  173.5 267.1 174.1 267.7 ;
      RECT  173.5 256.7 174.1 257.3 ;
      RECT  165.1 276.5 165.9 278.1 ;
      RECT  165.1 269.5 165.9 267.1 ;
      RECT  168.3 269.5 169.1 267.1 ;
      RECT  169.9 268.7 170.7 267.4 ;
      RECT  169.9 277.8 170.7 276.5 ;
      RECT  165.1 269.5 165.9 268.7 ;
      RECT  166.7 269.5 167.5 268.7 ;
      RECT  166.7 269.5 167.5 268.7 ;
      RECT  165.1 269.5 165.9 268.7 ;
      RECT  166.7 269.5 167.5 268.7 ;
      RECT  168.3 269.5 169.1 268.7 ;
      RECT  168.3 269.5 169.1 268.7 ;
      RECT  166.7 269.5 167.5 268.7 ;
      RECT  165.1 276.5 165.9 275.7 ;
      RECT  166.7 276.5 167.5 275.7 ;
      RECT  166.7 276.5 167.5 275.7 ;
      RECT  165.1 276.5 165.9 275.7 ;
      RECT  166.7 276.5 167.5 275.7 ;
      RECT  168.3 276.5 169.1 275.7 ;
      RECT  168.3 276.5 169.1 275.7 ;
      RECT  166.7 276.5 167.5 275.7 ;
      RECT  169.9 269.1 170.7 268.3 ;
      RECT  169.9 276.9 170.7 276.1 ;
      RECT  167.5 274.8 168.3 274.0 ;
      RECT  165.5 273.4 166.3 272.6 ;
      RECT  166.7 269.5 167.5 268.7 ;
      RECT  168.3 276.5 169.1 275.7 ;
      RECT  169.7 273.4 170.5 272.6 ;
      RECT  165.5 273.4 166.3 272.6 ;
      RECT  167.5 274.8 168.3 274.0 ;
      RECT  169.7 273.4 170.5 272.6 ;
      RECT  163.9 267.7 173.5 267.1 ;
      RECT  163.9 278.1 173.5 277.5 ;
      RECT  177.9 268.7 178.7 267.4 ;
      RECT  177.9 277.8 178.7 276.5 ;
      RECT  174.7 276.9 175.5 278.1 ;
      RECT  174.7 269.5 175.5 267.1 ;
      RECT  176.4 276.9 177.0 268.7 ;
      RECT  174.7 269.5 175.5 268.7 ;
      RECT  176.3 269.5 177.1 268.7 ;
      RECT  176.3 269.5 177.1 268.7 ;
      RECT  174.7 269.5 175.5 268.7 ;
      RECT  174.7 276.9 175.5 276.1 ;
      RECT  176.3 276.9 177.1 276.1 ;
      RECT  176.3 276.9 177.1 276.1 ;
      RECT  174.7 276.9 175.5 276.1 ;
      RECT  177.9 269.1 178.7 268.3 ;
      RECT  177.9 276.9 178.7 276.1 ;
      RECT  174.9 273.2 175.7 272.4 ;
      RECT  174.9 273.2 175.7 272.4 ;
      RECT  176.7 273.1 177.3 272.5 ;
      RECT  173.5 267.7 179.9 267.1 ;
      RECT  173.5 278.1 179.9 277.5 ;
      RECT  174.9 273.2 175.7 272.4 ;
      RECT  176.7 273.1 177.3 272.5 ;
      RECT  173.5 267.7 174.1 267.1 ;
      RECT  173.5 278.1 174.1 277.5 ;
      RECT  165.1 279.1 165.9 277.5 ;
      RECT  165.1 286.1 165.9 288.5 ;
      RECT  168.3 286.1 169.1 288.5 ;
      RECT  169.9 286.9 170.7 288.2 ;
      RECT  169.9 277.8 170.7 279.1 ;
      RECT  165.1 286.1 165.9 286.9 ;
      RECT  166.7 286.1 167.5 286.9 ;
      RECT  166.7 286.1 167.5 286.9 ;
      RECT  165.1 286.1 165.9 286.9 ;
      RECT  166.7 286.1 167.5 286.9 ;
      RECT  168.3 286.1 169.1 286.9 ;
      RECT  168.3 286.1 169.1 286.9 ;
      RECT  166.7 286.1 167.5 286.9 ;
      RECT  165.1 279.1 165.9 279.9 ;
      RECT  166.7 279.1 167.5 279.9 ;
      RECT  166.7 279.1 167.5 279.9 ;
      RECT  165.1 279.1 165.9 279.9 ;
      RECT  166.7 279.1 167.5 279.9 ;
      RECT  168.3 279.1 169.1 279.9 ;
      RECT  168.3 279.1 169.1 279.9 ;
      RECT  166.7 279.1 167.5 279.9 ;
      RECT  169.9 286.5 170.7 287.3 ;
      RECT  169.9 278.7 170.7 279.5 ;
      RECT  167.5 280.8 168.3 281.6 ;
      RECT  165.5 282.2 166.3 283.0 ;
      RECT  166.7 286.1 167.5 286.9 ;
      RECT  168.3 279.1 169.1 279.9 ;
      RECT  169.7 282.2 170.5 283.0 ;
      RECT  165.5 282.2 166.3 283.0 ;
      RECT  167.5 280.8 168.3 281.6 ;
      RECT  169.7 282.2 170.5 283.0 ;
      RECT  163.9 287.9 173.5 288.5 ;
      RECT  163.9 277.5 173.5 278.1 ;
      RECT  177.9 286.9 178.7 288.2 ;
      RECT  177.9 277.8 178.7 279.1 ;
      RECT  174.7 278.7 175.5 277.5 ;
      RECT  174.7 286.1 175.5 288.5 ;
      RECT  176.4 278.7 177.0 286.9 ;
      RECT  174.7 286.1 175.5 286.9 ;
      RECT  176.3 286.1 177.1 286.9 ;
      RECT  176.3 286.1 177.1 286.9 ;
      RECT  174.7 286.1 175.5 286.9 ;
      RECT  174.7 278.7 175.5 279.5 ;
      RECT  176.3 278.7 177.1 279.5 ;
      RECT  176.3 278.7 177.1 279.5 ;
      RECT  174.7 278.7 175.5 279.5 ;
      RECT  177.9 286.5 178.7 287.3 ;
      RECT  177.9 278.7 178.7 279.5 ;
      RECT  174.9 282.4 175.7 283.2 ;
      RECT  174.9 282.4 175.7 283.2 ;
      RECT  176.7 282.5 177.3 283.1 ;
      RECT  173.5 287.9 179.9 288.5 ;
      RECT  173.5 277.5 179.9 278.1 ;
      RECT  174.9 282.4 175.7 283.2 ;
      RECT  176.7 282.5 177.3 283.1 ;
      RECT  173.5 287.9 174.1 288.5 ;
      RECT  173.5 277.5 174.1 278.1 ;
      RECT  165.1 297.3 165.9 298.9 ;
      RECT  165.1 290.3 165.9 287.9 ;
      RECT  168.3 290.3 169.1 287.9 ;
      RECT  169.9 289.5 170.7 288.2 ;
      RECT  169.9 298.6 170.7 297.3 ;
      RECT  165.1 290.3 165.9 289.5 ;
      RECT  166.7 290.3 167.5 289.5 ;
      RECT  166.7 290.3 167.5 289.5 ;
      RECT  165.1 290.3 165.9 289.5 ;
      RECT  166.7 290.3 167.5 289.5 ;
      RECT  168.3 290.3 169.1 289.5 ;
      RECT  168.3 290.3 169.1 289.5 ;
      RECT  166.7 290.3 167.5 289.5 ;
      RECT  165.1 297.3 165.9 296.5 ;
      RECT  166.7 297.3 167.5 296.5 ;
      RECT  166.7 297.3 167.5 296.5 ;
      RECT  165.1 297.3 165.9 296.5 ;
      RECT  166.7 297.3 167.5 296.5 ;
      RECT  168.3 297.3 169.1 296.5 ;
      RECT  168.3 297.3 169.1 296.5 ;
      RECT  166.7 297.3 167.5 296.5 ;
      RECT  169.9 289.9 170.7 289.1 ;
      RECT  169.9 297.7 170.7 296.9 ;
      RECT  167.5 295.6 168.3 294.8 ;
      RECT  165.5 294.2 166.3 293.4 ;
      RECT  166.7 290.3 167.5 289.5 ;
      RECT  168.3 297.3 169.1 296.5 ;
      RECT  169.7 294.2 170.5 293.4 ;
      RECT  165.5 294.2 166.3 293.4 ;
      RECT  167.5 295.6 168.3 294.8 ;
      RECT  169.7 294.2 170.5 293.4 ;
      RECT  163.9 288.5 173.5 287.9 ;
      RECT  163.9 298.9 173.5 298.3 ;
      RECT  177.9 289.5 178.7 288.2 ;
      RECT  177.9 298.6 178.7 297.3 ;
      RECT  174.7 297.7 175.5 298.9 ;
      RECT  174.7 290.3 175.5 287.9 ;
      RECT  176.4 297.7 177.0 289.5 ;
      RECT  174.7 290.3 175.5 289.5 ;
      RECT  176.3 290.3 177.1 289.5 ;
      RECT  176.3 290.3 177.1 289.5 ;
      RECT  174.7 290.3 175.5 289.5 ;
      RECT  174.7 297.7 175.5 296.9 ;
      RECT  176.3 297.7 177.1 296.9 ;
      RECT  176.3 297.7 177.1 296.9 ;
      RECT  174.7 297.7 175.5 296.9 ;
      RECT  177.9 289.9 178.7 289.1 ;
      RECT  177.9 297.7 178.7 296.9 ;
      RECT  174.9 294.0 175.7 293.2 ;
      RECT  174.9 294.0 175.7 293.2 ;
      RECT  176.7 293.9 177.3 293.3 ;
      RECT  173.5 288.5 179.9 287.9 ;
      RECT  173.5 298.9 179.9 298.3 ;
      RECT  174.9 294.0 175.7 293.2 ;
      RECT  176.7 293.9 177.3 293.3 ;
      RECT  173.5 288.5 174.1 287.9 ;
      RECT  173.5 298.9 174.1 298.3 ;
      RECT  165.1 299.9 165.9 298.3 ;
      RECT  165.1 306.9 165.9 309.3 ;
      RECT  168.3 306.9 169.1 309.3 ;
      RECT  169.9 307.7 170.7 309.0 ;
      RECT  169.9 298.6 170.7 299.9 ;
      RECT  165.1 306.9 165.9 307.7 ;
      RECT  166.7 306.9 167.5 307.7 ;
      RECT  166.7 306.9 167.5 307.7 ;
      RECT  165.1 306.9 165.9 307.7 ;
      RECT  166.7 306.9 167.5 307.7 ;
      RECT  168.3 306.9 169.1 307.7 ;
      RECT  168.3 306.9 169.1 307.7 ;
      RECT  166.7 306.9 167.5 307.7 ;
      RECT  165.1 299.9 165.9 300.7 ;
      RECT  166.7 299.9 167.5 300.7 ;
      RECT  166.7 299.9 167.5 300.7 ;
      RECT  165.1 299.9 165.9 300.7 ;
      RECT  166.7 299.9 167.5 300.7 ;
      RECT  168.3 299.9 169.1 300.7 ;
      RECT  168.3 299.9 169.1 300.7 ;
      RECT  166.7 299.9 167.5 300.7 ;
      RECT  169.9 307.3 170.7 308.1 ;
      RECT  169.9 299.5 170.7 300.3 ;
      RECT  167.5 301.6 168.3 302.4 ;
      RECT  165.5 303.0 166.3 303.8 ;
      RECT  166.7 306.9 167.5 307.7 ;
      RECT  168.3 299.9 169.1 300.7 ;
      RECT  169.7 303.0 170.5 303.8 ;
      RECT  165.5 303.0 166.3 303.8 ;
      RECT  167.5 301.6 168.3 302.4 ;
      RECT  169.7 303.0 170.5 303.8 ;
      RECT  163.9 308.7 173.5 309.3 ;
      RECT  163.9 298.3 173.5 298.9 ;
      RECT  177.9 307.7 178.7 309.0 ;
      RECT  177.9 298.6 178.7 299.9 ;
      RECT  174.7 299.5 175.5 298.3 ;
      RECT  174.7 306.9 175.5 309.3 ;
      RECT  176.4 299.5 177.0 307.7 ;
      RECT  174.7 306.9 175.5 307.7 ;
      RECT  176.3 306.9 177.1 307.7 ;
      RECT  176.3 306.9 177.1 307.7 ;
      RECT  174.7 306.9 175.5 307.7 ;
      RECT  174.7 299.5 175.5 300.3 ;
      RECT  176.3 299.5 177.1 300.3 ;
      RECT  176.3 299.5 177.1 300.3 ;
      RECT  174.7 299.5 175.5 300.3 ;
      RECT  177.9 307.3 178.7 308.1 ;
      RECT  177.9 299.5 178.7 300.3 ;
      RECT  174.9 303.2 175.7 304.0 ;
      RECT  174.9 303.2 175.7 304.0 ;
      RECT  176.7 303.3 177.3 303.9 ;
      RECT  173.5 308.7 179.9 309.3 ;
      RECT  173.5 298.3 179.9 298.9 ;
      RECT  174.9 303.2 175.7 304.0 ;
      RECT  176.7 303.3 177.3 303.9 ;
      RECT  173.5 308.7 174.1 309.3 ;
      RECT  173.5 298.3 174.1 298.9 ;
      RECT  165.1 318.1 165.9 319.7 ;
      RECT  165.1 311.1 165.9 308.7 ;
      RECT  168.3 311.1 169.1 308.7 ;
      RECT  169.9 310.3 170.7 309.0 ;
      RECT  169.9 319.4 170.7 318.1 ;
      RECT  165.1 311.1 165.9 310.3 ;
      RECT  166.7 311.1 167.5 310.3 ;
      RECT  166.7 311.1 167.5 310.3 ;
      RECT  165.1 311.1 165.9 310.3 ;
      RECT  166.7 311.1 167.5 310.3 ;
      RECT  168.3 311.1 169.1 310.3 ;
      RECT  168.3 311.1 169.1 310.3 ;
      RECT  166.7 311.1 167.5 310.3 ;
      RECT  165.1 318.1 165.9 317.3 ;
      RECT  166.7 318.1 167.5 317.3 ;
      RECT  166.7 318.1 167.5 317.3 ;
      RECT  165.1 318.1 165.9 317.3 ;
      RECT  166.7 318.1 167.5 317.3 ;
      RECT  168.3 318.1 169.1 317.3 ;
      RECT  168.3 318.1 169.1 317.3 ;
      RECT  166.7 318.1 167.5 317.3 ;
      RECT  169.9 310.7 170.7 309.9 ;
      RECT  169.9 318.5 170.7 317.7 ;
      RECT  167.5 316.4 168.3 315.6 ;
      RECT  165.5 315.0 166.3 314.2 ;
      RECT  166.7 311.1 167.5 310.3 ;
      RECT  168.3 318.1 169.1 317.3 ;
      RECT  169.7 315.0 170.5 314.2 ;
      RECT  165.5 315.0 166.3 314.2 ;
      RECT  167.5 316.4 168.3 315.6 ;
      RECT  169.7 315.0 170.5 314.2 ;
      RECT  163.9 309.3 173.5 308.7 ;
      RECT  163.9 319.7 173.5 319.1 ;
      RECT  177.9 310.3 178.7 309.0 ;
      RECT  177.9 319.4 178.7 318.1 ;
      RECT  174.7 318.5 175.5 319.7 ;
      RECT  174.7 311.1 175.5 308.7 ;
      RECT  176.4 318.5 177.0 310.3 ;
      RECT  174.7 311.1 175.5 310.3 ;
      RECT  176.3 311.1 177.1 310.3 ;
      RECT  176.3 311.1 177.1 310.3 ;
      RECT  174.7 311.1 175.5 310.3 ;
      RECT  174.7 318.5 175.5 317.7 ;
      RECT  176.3 318.5 177.1 317.7 ;
      RECT  176.3 318.5 177.1 317.7 ;
      RECT  174.7 318.5 175.5 317.7 ;
      RECT  177.9 310.7 178.7 309.9 ;
      RECT  177.9 318.5 178.7 317.7 ;
      RECT  174.9 314.8 175.7 314.0 ;
      RECT  174.9 314.8 175.7 314.0 ;
      RECT  176.7 314.7 177.3 314.1 ;
      RECT  173.5 309.3 179.9 308.7 ;
      RECT  173.5 319.7 179.9 319.1 ;
      RECT  174.9 314.8 175.7 314.0 ;
      RECT  176.7 314.7 177.3 314.1 ;
      RECT  173.5 309.3 174.1 308.7 ;
      RECT  173.5 319.7 174.1 319.1 ;
      RECT  165.1 320.7 165.9 319.1 ;
      RECT  165.1 327.7 165.9 330.1 ;
      RECT  168.3 327.7 169.1 330.1 ;
      RECT  169.9 328.5 170.7 329.8 ;
      RECT  169.9 319.4 170.7 320.7 ;
      RECT  165.1 327.7 165.9 328.5 ;
      RECT  166.7 327.7 167.5 328.5 ;
      RECT  166.7 327.7 167.5 328.5 ;
      RECT  165.1 327.7 165.9 328.5 ;
      RECT  166.7 327.7 167.5 328.5 ;
      RECT  168.3 327.7 169.1 328.5 ;
      RECT  168.3 327.7 169.1 328.5 ;
      RECT  166.7 327.7 167.5 328.5 ;
      RECT  165.1 320.7 165.9 321.5 ;
      RECT  166.7 320.7 167.5 321.5 ;
      RECT  166.7 320.7 167.5 321.5 ;
      RECT  165.1 320.7 165.9 321.5 ;
      RECT  166.7 320.7 167.5 321.5 ;
      RECT  168.3 320.7 169.1 321.5 ;
      RECT  168.3 320.7 169.1 321.5 ;
      RECT  166.7 320.7 167.5 321.5 ;
      RECT  169.9 328.1 170.7 328.9 ;
      RECT  169.9 320.3 170.7 321.1 ;
      RECT  167.5 322.4 168.3 323.2 ;
      RECT  165.5 323.8 166.3 324.6 ;
      RECT  166.7 327.7 167.5 328.5 ;
      RECT  168.3 320.7 169.1 321.5 ;
      RECT  169.7 323.8 170.5 324.6 ;
      RECT  165.5 323.8 166.3 324.6 ;
      RECT  167.5 322.4 168.3 323.2 ;
      RECT  169.7 323.8 170.5 324.6 ;
      RECT  163.9 329.5 173.5 330.1 ;
      RECT  163.9 319.1 173.5 319.7 ;
      RECT  177.9 328.5 178.7 329.8 ;
      RECT  177.9 319.4 178.7 320.7 ;
      RECT  174.7 320.3 175.5 319.1 ;
      RECT  174.7 327.7 175.5 330.1 ;
      RECT  176.4 320.3 177.0 328.5 ;
      RECT  174.7 327.7 175.5 328.5 ;
      RECT  176.3 327.7 177.1 328.5 ;
      RECT  176.3 327.7 177.1 328.5 ;
      RECT  174.7 327.7 175.5 328.5 ;
      RECT  174.7 320.3 175.5 321.1 ;
      RECT  176.3 320.3 177.1 321.1 ;
      RECT  176.3 320.3 177.1 321.1 ;
      RECT  174.7 320.3 175.5 321.1 ;
      RECT  177.9 328.1 178.7 328.9 ;
      RECT  177.9 320.3 178.7 321.1 ;
      RECT  174.9 324.0 175.7 324.8 ;
      RECT  174.9 324.0 175.7 324.8 ;
      RECT  176.7 324.1 177.3 324.7 ;
      RECT  173.5 329.5 179.9 330.1 ;
      RECT  173.5 319.1 179.9 319.7 ;
      RECT  174.9 324.0 175.7 324.8 ;
      RECT  176.7 324.1 177.3 324.7 ;
      RECT  173.5 329.5 174.1 330.1 ;
      RECT  173.5 319.1 174.1 319.7 ;
      RECT  165.1 338.9 165.9 340.5 ;
      RECT  165.1 331.9 165.9 329.5 ;
      RECT  168.3 331.9 169.1 329.5 ;
      RECT  169.9 331.1 170.7 329.8 ;
      RECT  169.9 340.2 170.7 338.9 ;
      RECT  165.1 331.9 165.9 331.1 ;
      RECT  166.7 331.9 167.5 331.1 ;
      RECT  166.7 331.9 167.5 331.1 ;
      RECT  165.1 331.9 165.9 331.1 ;
      RECT  166.7 331.9 167.5 331.1 ;
      RECT  168.3 331.9 169.1 331.1 ;
      RECT  168.3 331.9 169.1 331.1 ;
      RECT  166.7 331.9 167.5 331.1 ;
      RECT  165.1 338.9 165.9 338.1 ;
      RECT  166.7 338.9 167.5 338.1 ;
      RECT  166.7 338.9 167.5 338.1 ;
      RECT  165.1 338.9 165.9 338.1 ;
      RECT  166.7 338.9 167.5 338.1 ;
      RECT  168.3 338.9 169.1 338.1 ;
      RECT  168.3 338.9 169.1 338.1 ;
      RECT  166.7 338.9 167.5 338.1 ;
      RECT  169.9 331.5 170.7 330.7 ;
      RECT  169.9 339.3 170.7 338.5 ;
      RECT  167.5 337.2 168.3 336.4 ;
      RECT  165.5 335.8 166.3 335.0 ;
      RECT  166.7 331.9 167.5 331.1 ;
      RECT  168.3 338.9 169.1 338.1 ;
      RECT  169.7 335.8 170.5 335.0 ;
      RECT  165.5 335.8 166.3 335.0 ;
      RECT  167.5 337.2 168.3 336.4 ;
      RECT  169.7 335.8 170.5 335.0 ;
      RECT  163.9 330.1 173.5 329.5 ;
      RECT  163.9 340.5 173.5 339.9 ;
      RECT  177.9 331.1 178.7 329.8 ;
      RECT  177.9 340.2 178.7 338.9 ;
      RECT  174.7 339.3 175.5 340.5 ;
      RECT  174.7 331.9 175.5 329.5 ;
      RECT  176.4 339.3 177.0 331.1 ;
      RECT  174.7 331.9 175.5 331.1 ;
      RECT  176.3 331.9 177.1 331.1 ;
      RECT  176.3 331.9 177.1 331.1 ;
      RECT  174.7 331.9 175.5 331.1 ;
      RECT  174.7 339.3 175.5 338.5 ;
      RECT  176.3 339.3 177.1 338.5 ;
      RECT  176.3 339.3 177.1 338.5 ;
      RECT  174.7 339.3 175.5 338.5 ;
      RECT  177.9 331.5 178.7 330.7 ;
      RECT  177.9 339.3 178.7 338.5 ;
      RECT  174.9 335.6 175.7 334.8 ;
      RECT  174.9 335.6 175.7 334.8 ;
      RECT  176.7 335.5 177.3 334.9 ;
      RECT  173.5 330.1 179.9 329.5 ;
      RECT  173.5 340.5 179.9 339.9 ;
      RECT  174.9 335.6 175.7 334.8 ;
      RECT  176.7 335.5 177.3 334.9 ;
      RECT  173.5 330.1 174.1 329.5 ;
      RECT  173.5 340.5 174.1 339.9 ;
      RECT  165.1 341.5 165.9 339.9 ;
      RECT  165.1 348.5 165.9 350.9 ;
      RECT  168.3 348.5 169.1 350.9 ;
      RECT  169.9 349.3 170.7 350.6 ;
      RECT  169.9 340.2 170.7 341.5 ;
      RECT  165.1 348.5 165.9 349.3 ;
      RECT  166.7 348.5 167.5 349.3 ;
      RECT  166.7 348.5 167.5 349.3 ;
      RECT  165.1 348.5 165.9 349.3 ;
      RECT  166.7 348.5 167.5 349.3 ;
      RECT  168.3 348.5 169.1 349.3 ;
      RECT  168.3 348.5 169.1 349.3 ;
      RECT  166.7 348.5 167.5 349.3 ;
      RECT  165.1 341.5 165.9 342.3 ;
      RECT  166.7 341.5 167.5 342.3 ;
      RECT  166.7 341.5 167.5 342.3 ;
      RECT  165.1 341.5 165.9 342.3 ;
      RECT  166.7 341.5 167.5 342.3 ;
      RECT  168.3 341.5 169.1 342.3 ;
      RECT  168.3 341.5 169.1 342.3 ;
      RECT  166.7 341.5 167.5 342.3 ;
      RECT  169.9 348.9 170.7 349.7 ;
      RECT  169.9 341.1 170.7 341.9 ;
      RECT  167.5 343.2 168.3 344.0 ;
      RECT  165.5 344.6 166.3 345.4 ;
      RECT  166.7 348.5 167.5 349.3 ;
      RECT  168.3 341.5 169.1 342.3 ;
      RECT  169.7 344.6 170.5 345.4 ;
      RECT  165.5 344.6 166.3 345.4 ;
      RECT  167.5 343.2 168.3 344.0 ;
      RECT  169.7 344.6 170.5 345.4 ;
      RECT  163.9 350.3 173.5 350.9 ;
      RECT  163.9 339.9 173.5 340.5 ;
      RECT  177.9 349.3 178.7 350.6 ;
      RECT  177.9 340.2 178.7 341.5 ;
      RECT  174.7 341.1 175.5 339.9 ;
      RECT  174.7 348.5 175.5 350.9 ;
      RECT  176.4 341.1 177.0 349.3 ;
      RECT  174.7 348.5 175.5 349.3 ;
      RECT  176.3 348.5 177.1 349.3 ;
      RECT  176.3 348.5 177.1 349.3 ;
      RECT  174.7 348.5 175.5 349.3 ;
      RECT  174.7 341.1 175.5 341.9 ;
      RECT  176.3 341.1 177.1 341.9 ;
      RECT  176.3 341.1 177.1 341.9 ;
      RECT  174.7 341.1 175.5 341.9 ;
      RECT  177.9 348.9 178.7 349.7 ;
      RECT  177.9 341.1 178.7 341.9 ;
      RECT  174.9 344.8 175.7 345.6 ;
      RECT  174.9 344.8 175.7 345.6 ;
      RECT  176.7 344.9 177.3 345.5 ;
      RECT  173.5 350.3 179.9 350.9 ;
      RECT  173.5 339.9 179.9 340.5 ;
      RECT  174.9 344.8 175.7 345.6 ;
      RECT  176.7 344.9 177.3 345.5 ;
      RECT  173.5 350.3 174.1 350.9 ;
      RECT  173.5 339.9 174.1 340.5 ;
      RECT  165.1 359.7 165.9 361.3 ;
      RECT  165.1 352.7 165.9 350.3 ;
      RECT  168.3 352.7 169.1 350.3 ;
      RECT  169.9 351.9 170.7 350.6 ;
      RECT  169.9 361.0 170.7 359.7 ;
      RECT  165.1 352.7 165.9 351.9 ;
      RECT  166.7 352.7 167.5 351.9 ;
      RECT  166.7 352.7 167.5 351.9 ;
      RECT  165.1 352.7 165.9 351.9 ;
      RECT  166.7 352.7 167.5 351.9 ;
      RECT  168.3 352.7 169.1 351.9 ;
      RECT  168.3 352.7 169.1 351.9 ;
      RECT  166.7 352.7 167.5 351.9 ;
      RECT  165.1 359.7 165.9 358.9 ;
      RECT  166.7 359.7 167.5 358.9 ;
      RECT  166.7 359.7 167.5 358.9 ;
      RECT  165.1 359.7 165.9 358.9 ;
      RECT  166.7 359.7 167.5 358.9 ;
      RECT  168.3 359.7 169.1 358.9 ;
      RECT  168.3 359.7 169.1 358.9 ;
      RECT  166.7 359.7 167.5 358.9 ;
      RECT  169.9 352.3 170.7 351.5 ;
      RECT  169.9 360.1 170.7 359.3 ;
      RECT  167.5 358.0 168.3 357.2 ;
      RECT  165.5 356.6 166.3 355.8 ;
      RECT  166.7 352.7 167.5 351.9 ;
      RECT  168.3 359.7 169.1 358.9 ;
      RECT  169.7 356.6 170.5 355.8 ;
      RECT  165.5 356.6 166.3 355.8 ;
      RECT  167.5 358.0 168.3 357.2 ;
      RECT  169.7 356.6 170.5 355.8 ;
      RECT  163.9 350.9 173.5 350.3 ;
      RECT  163.9 361.3 173.5 360.7 ;
      RECT  177.9 351.9 178.7 350.6 ;
      RECT  177.9 361.0 178.7 359.7 ;
      RECT  174.7 360.1 175.5 361.3 ;
      RECT  174.7 352.7 175.5 350.3 ;
      RECT  176.4 360.1 177.0 351.9 ;
      RECT  174.7 352.7 175.5 351.9 ;
      RECT  176.3 352.7 177.1 351.9 ;
      RECT  176.3 352.7 177.1 351.9 ;
      RECT  174.7 352.7 175.5 351.9 ;
      RECT  174.7 360.1 175.5 359.3 ;
      RECT  176.3 360.1 177.1 359.3 ;
      RECT  176.3 360.1 177.1 359.3 ;
      RECT  174.7 360.1 175.5 359.3 ;
      RECT  177.9 352.3 178.7 351.5 ;
      RECT  177.9 360.1 178.7 359.3 ;
      RECT  174.9 356.4 175.7 355.6 ;
      RECT  174.9 356.4 175.7 355.6 ;
      RECT  176.7 356.3 177.3 355.7 ;
      RECT  173.5 350.9 179.9 350.3 ;
      RECT  173.5 361.3 179.9 360.7 ;
      RECT  174.9 356.4 175.7 355.6 ;
      RECT  176.7 356.3 177.3 355.7 ;
      RECT  173.5 350.9 174.1 350.3 ;
      RECT  173.5 361.3 174.1 360.7 ;
      RECT  161.4 199.0 162.2 199.8 ;
      RECT  162.7 197.0 163.5 197.8 ;
      RECT  166.7 197.6 167.5 198.4 ;
      RECT  161.4 210.2 162.2 211.0 ;
      RECT  162.7 212.2 163.5 213.0 ;
      RECT  166.7 211.6 167.5 212.4 ;
      RECT  161.4 219.8 162.2 220.6 ;
      RECT  162.7 217.8 163.5 218.6 ;
      RECT  166.7 218.4 167.5 219.2 ;
      RECT  161.4 231.0 162.2 231.8 ;
      RECT  162.7 233.0 163.5 233.8 ;
      RECT  166.7 232.4 167.5 233.2 ;
      RECT  161.4 240.6 162.2 241.4 ;
      RECT  162.7 238.6 163.5 239.4 ;
      RECT  166.7 239.2 167.5 240.0 ;
      RECT  161.4 251.8 162.2 252.6 ;
      RECT  162.7 253.8 163.5 254.6 ;
      RECT  166.7 253.2 167.5 254.0 ;
      RECT  161.4 261.4 162.2 262.2 ;
      RECT  162.7 259.4 163.5 260.2 ;
      RECT  166.7 260.0 167.5 260.8 ;
      RECT  161.4 272.6 162.2 273.4 ;
      RECT  162.7 274.6 163.5 275.4 ;
      RECT  166.7 274.0 167.5 274.8 ;
      RECT  161.4 282.2 162.2 283.0 ;
      RECT  162.7 280.2 163.5 281.0 ;
      RECT  166.7 280.8 167.5 281.6 ;
      RECT  161.4 293.4 162.2 294.2 ;
      RECT  162.7 295.4 163.5 296.2 ;
      RECT  166.7 294.8 167.5 295.6 ;
      RECT  161.4 303.0 162.2 303.8 ;
      RECT  162.7 301.0 163.5 301.8 ;
      RECT  166.7 301.6 167.5 302.4 ;
      RECT  161.4 314.2 162.2 315.0 ;
      RECT  162.7 316.2 163.5 317.0 ;
      RECT  166.7 315.6 167.5 316.4 ;
      RECT  161.4 323.8 162.2 324.6 ;
      RECT  162.7 321.8 163.5 322.6 ;
      RECT  166.7 322.4 167.5 323.2 ;
      RECT  161.4 335.0 162.2 335.8 ;
      RECT  162.7 337.0 163.5 337.8 ;
      RECT  166.7 336.4 167.5 337.2 ;
      RECT  161.4 344.6 162.2 345.4 ;
      RECT  162.7 342.6 163.5 343.4 ;
      RECT  166.7 343.2 167.5 344.0 ;
      RECT  161.4 355.8 162.2 356.6 ;
      RECT  162.7 357.8 163.5 358.6 ;
      RECT  166.7 357.2 167.5 358.0 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 194.2 173.9 195.0 ;
      RECT  173.1 194.2 173.9 195.0 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 360.6 173.9 361.4 ;
      RECT  173.1 360.6 173.9 361.4 ;
      RECT  159.7 197.1 163.1 197.7 ;
      RECT  159.7 212.3 163.1 212.9 ;
      RECT  159.7 217.9 163.1 218.5 ;
      RECT  159.7 233.1 163.1 233.7 ;
      RECT  159.7 238.7 163.1 239.3 ;
      RECT  159.7 253.9 163.1 254.5 ;
      RECT  159.7 259.5 163.1 260.1 ;
      RECT  159.7 274.7 163.1 275.3 ;
      RECT  159.7 280.3 163.1 280.9 ;
      RECT  159.7 295.5 163.1 296.1 ;
      RECT  159.7 301.1 163.1 301.7 ;
      RECT  159.7 316.3 163.1 316.9 ;
      RECT  159.7 321.9 163.1 322.5 ;
      RECT  159.7 337.1 163.1 337.7 ;
      RECT  159.7 342.7 163.1 343.3 ;
      RECT  159.7 357.9 163.1 358.5 ;
      RECT  176.7 199.3 177.3 199.9 ;
      RECT  176.7 210.1 177.3 210.7 ;
      RECT  176.7 220.1 177.3 220.7 ;
      RECT  176.7 230.9 177.3 231.5 ;
      RECT  176.7 240.9 177.3 241.5 ;
      RECT  176.7 251.7 177.3 252.3 ;
      RECT  176.7 261.7 177.3 262.3 ;
      RECT  176.7 272.5 177.3 273.1 ;
      RECT  176.7 282.5 177.3 283.1 ;
      RECT  176.7 293.3 177.3 293.9 ;
      RECT  176.7 303.3 177.3 303.9 ;
      RECT  176.7 314.1 177.3 314.7 ;
      RECT  176.7 324.1 177.3 324.7 ;
      RECT  176.7 334.9 177.3 335.5 ;
      RECT  176.7 344.9 177.3 345.5 ;
      RECT  176.7 355.7 177.3 356.3 ;
      RECT  176.7 199.3 177.3 199.9 ;
      RECT  176.7 210.1 177.3 210.7 ;
      RECT  176.7 220.1 177.3 220.7 ;
      RECT  176.7 230.9 177.3 231.5 ;
      RECT  176.7 240.9 177.3 241.5 ;
      RECT  176.7 251.7 177.3 252.3 ;
      RECT  176.7 261.7 177.3 262.3 ;
      RECT  176.7 272.5 177.3 273.1 ;
      RECT  176.7 282.5 177.3 283.1 ;
      RECT  176.7 293.3 177.3 293.9 ;
      RECT  176.7 303.3 177.3 303.9 ;
      RECT  176.7 314.1 177.3 314.7 ;
      RECT  176.7 324.1 177.3 324.7 ;
      RECT  176.7 334.9 177.3 335.5 ;
      RECT  176.7 344.9 177.3 345.5 ;
      RECT  176.7 355.7 177.3 356.3 ;
      RECT  181.5 159.7 182.3 160.5 ;
      RECT  181.5 159.7 182.3 160.5 ;
      RECT  182.9 191.2 183.7 192.0 ;
      RECT  182.9 191.2 183.7 192.0 ;
      RECT  178.7 79.7 179.5 80.5 ;
      RECT  178.7 79.7 179.5 80.5 ;
      RECT  180.1 149.5 180.9 150.3 ;
      RECT  180.1 149.5 180.9 150.3 ;
      RECT  161.4 185.8 162.2 186.6 ;
      RECT  182.9 185.8 183.7 186.6 ;
      RECT  5.9 44.7 44.7 45.3 ;
      RECT  40.5 72.1 51.8 72.7 ;
      RECT  39.1 131.7 51.8 132.3 ;
      RECT  43.3 87.6 52.4 88.2 ;
      RECT  37.7 86.3 54.0 86.9 ;
      RECT  40.5 85.0 55.6 85.6 ;
      RECT  39.1 156.2 52.4 156.8 ;
      RECT  40.5 157.5 54.0 158.1 ;
      RECT  46.1 158.8 55.6 159.4 ;
      RECT  5.6 101.6 39.1 102.2 ;
      RECT  41.9 117.1 52.0 117.7 ;
      RECT  39.1 118.5 54.0 119.1 ;
      RECT  56.6 112.1 61.0 112.7 ;
      RECT  44.7 32.1 51.8 32.7 ;
      RECT  60.1 32.1 60.7 32.7 ;
      RECT  53.5 32.1 60.4 32.7 ;
      RECT  60.1 32.4 60.7 38.8 ;
      RECT  44.7 46.7 52.0 47.3 ;
      RECT  47.5 45.3 54.0 45.9 ;
      RECT  50.6 21.9 85.2 22.5 ;
      RECT  50.6 1.9 85.2 2.5 ;
      RECT  78.8 61.9 85.2 62.5 ;
      RECT  78.8 41.9 85.2 42.5 ;
      RECT  50.6 61.9 85.2 62.5 ;
      RECT  50.6 81.9 85.2 82.5 ;
      RECT  68.4 101.9 85.2 102.5 ;
      RECT  68.4 81.9 85.2 82.5 ;
      RECT  60.2 101.9 85.2 102.5 ;
      RECT  60.2 121.9 85.2 122.5 ;
      RECT  56.4 141.9 85.2 142.5 ;
      RECT  56.4 121.9 85.2 122.5 ;
      RECT  66.8 141.9 85.2 142.5 ;
      RECT  66.8 161.9 85.2 162.5 ;
      RECT  30.1 11.5 30.7 12.1 ;
      RECT  30.1 11.1 30.7 11.7 ;
      RECT  28.1 11.5 30.4 12.1 ;
      RECT  30.1 11.4 30.7 11.8 ;
      RECT  30.4 11.1 32.8 11.7 ;
      RECT  35.6 11.1 36.2 11.7 ;
      RECT  34.5 11.1 35.9 11.7 ;
      RECT  35.6 10.0 36.2 11.4 ;
      RECT  30.1 11.8 30.7 13.2 ;
      RECT  16.8 10.2 17.6 10.4 ;
      RECT  4.0 3.4 4.8 8.2 ;
      RECT  12.8 16.4 13.4 17.0 ;
      RECT  10.6 15.8 14.2 16.4 ;
      RECT  4.0 12.0 9.6 12.2 ;
      RECT  4.8 9.0 15.8 9.6 ;
      RECT  21.6 12.4 22.4 21.0 ;
      RECT  12.8 5.4 13.4 6.0 ;
      RECT  8.4 3.4 9.2 4.8 ;
      RECT  10.6 15.6 11.4 15.8 ;
      RECT  16.8 16.2 17.6 17.0 ;
      RECT  13.2 13.0 13.8 14.2 ;
      RECT  7.2 17.0 9.2 17.6 ;
      RECT  14.4 2.8 15.2 5.4 ;
      RECT  10.6 6.0 13.4 6.6 ;
      RECT  7.2 4.8 9.2 5.4 ;
      RECT  21.6 8.4 22.4 11.8 ;
      RECT  17.0 17.0 18.2 21.0 ;
      RECT  5.6 13.2 6.4 21.6 ;
      RECT  7.2 13.6 12.6 14.2 ;
      RECT  15.2 9.6 15.8 12.8 ;
      RECT  2.8 21.6 24.6 22.8 ;
      RECT  18.2 11.8 22.4 12.4 ;
      RECT  20.0 13.0 20.8 21.6 ;
      RECT  23.2 2.8 24.0 4.2 ;
      RECT  17.0 13.4 17.6 14.4 ;
      RECT  15.2 12.8 17.6 13.4 ;
      RECT  4.0 12.6 4.8 21.0 ;
      RECT  16.8 4.8 18.2 5.4 ;
      RECT  13.2 14.2 15.4 14.8 ;
      RECT  8.4 17.6 9.2 21.0 ;
      RECT  6.2 10.8 11.2 11.4 ;
      RECT  23.2 20.0 24.0 21.6 ;
      RECT  16.8 10.4 20.6 11.0 ;
      RECT  16.8 5.4 17.6 6.2 ;
      RECT  2.8 1.6 24.6 2.8 ;
      RECT  10.4 11.4 11.2 11.6 ;
      RECT  7.8 9.6 8.6 9.8 ;
      RECT  13.4 15.6 14.2 15.8 ;
      RECT  21.6 3.4 22.4 7.8 ;
      RECT  4.8 8.8 6.4 9.0 ;
      RECT  7.2 16.2 8.0 17.0 ;
      RECT  12.8 3.4 13.6 5.4 ;
      RECT  6.2 10.6 7.0 10.8 ;
      RECT  7.2 14.2 8.0 14.4 ;
      RECT  18.6 7.6 19.4 7.8 ;
      RECT  8.8 6.0 9.6 6.8 ;
      RECT  20.0 2.8 20.8 7.2 ;
      RECT  14.6 14.0 15.4 14.2 ;
      RECT  11.0 2.8 12.0 5.4 ;
      RECT  9.0 6.8 9.6 9.0 ;
      RECT  14.4 17.0 15.2 21.6 ;
      RECT  11.2 17.0 12.0 21.6 ;
      RECT  14.6 8.8 15.4 9.0 ;
      RECT  9.0 12.6 13.8 13.0 ;
      RECT  4.0 12.2 9.8 12.4 ;
      RECT  12.8 17.0 13.6 21.0 ;
      RECT  19.8 11.0 20.6 11.2 ;
      RECT  4.0 12.4 13.8 12.6 ;
      RECT  11.8 14.2 12.6 14.4 ;
      RECT  17.0 3.4 18.2 4.8 ;
      RECT  10.6 6.6 11.4 6.8 ;
      RECT  17.0 14.4 18.4 15.2 ;
      RECT  18.2 11.6 19.0 11.8 ;
      RECT  7.2 5.4 8.0 6.2 ;
      RECT  5.6 2.8 6.4 7.4 ;
      RECT  18.6 7.8 22.4 8.4 ;
      RECT  29.0 20.9 29.8 22.2 ;
      RECT  29.0 2.2 29.8 3.5 ;
      RECT  25.8 3.5 26.6 1.9 ;
      RECT  25.8 19.3 26.6 22.5 ;
      RECT  27.5 3.5 28.1 20.1 ;
      RECT  25.8 19.3 26.6 20.1 ;
      RECT  27.4 19.3 28.2 20.1 ;
      RECT  27.4 19.3 28.2 20.1 ;
      RECT  25.8 19.3 26.6 20.1 ;
      RECT  25.8 3.5 26.6 4.3 ;
      RECT  27.4 3.5 28.2 4.3 ;
      RECT  27.4 3.5 28.2 4.3 ;
      RECT  25.8 3.5 26.6 4.3 ;
      RECT  29.0 20.5 29.8 21.3 ;
      RECT  29.0 3.1 29.8 3.9 ;
      RECT  26.0 11.4 26.8 12.2 ;
      RECT  26.0 11.4 26.8 12.2 ;
      RECT  27.8 11.5 28.4 12.1 ;
      RECT  24.6 21.9 31.0 22.5 ;
      RECT  24.6 1.9 31.0 2.5 ;
      RECT  35.4 20.9 36.2 22.2 ;
      RECT  35.4 2.2 36.2 3.5 ;
      RECT  32.2 4.3 33.0 1.9 ;
      RECT  32.2 17.7 33.0 22.5 ;
      RECT  33.9 4.3 34.5 18.5 ;
      RECT  32.2 17.7 33.0 18.5 ;
      RECT  33.8 17.7 34.6 18.5 ;
      RECT  33.8 17.7 34.6 18.5 ;
      RECT  32.2 17.7 33.0 18.5 ;
      RECT  32.2 4.3 33.0 5.1 ;
      RECT  33.8 4.3 34.6 5.1 ;
      RECT  33.8 4.3 34.6 5.1 ;
      RECT  32.2 4.3 33.0 5.1 ;
      RECT  35.4 20.5 36.2 21.3 ;
      RECT  35.4 3.1 36.2 3.9 ;
      RECT  32.4 11.0 33.2 11.8 ;
      RECT  32.4 11.0 33.2 11.8 ;
      RECT  34.2 11.1 34.8 11.7 ;
      RECT  31.0 21.9 37.4 22.5 ;
      RECT  31.0 1.9 37.4 2.5 ;
      RECT  26.0 11.4 26.8 12.2 ;
      RECT  35.5 9.6 36.3 10.4 ;
      RECT  30.0 12.8 30.8 13.6 ;
      RECT  2.8 21.6 37.4 22.8 ;
      RECT  2.8 1.6 37.4 2.8 ;
      RECT  30.1 32.9 30.7 32.3 ;
      RECT  30.1 33.3 30.7 32.7 ;
      RECT  28.1 32.9 30.4 32.3 ;
      RECT  30.1 33.0 30.7 32.6 ;
      RECT  30.4 33.3 32.8 32.7 ;
      RECT  35.6 33.3 36.2 32.7 ;
      RECT  34.5 33.3 35.9 32.7 ;
      RECT  35.6 34.4 36.2 33.0 ;
      RECT  30.1 32.6 30.7 31.2 ;
      RECT  16.8 34.2 17.6 34.0 ;
      RECT  4.0 41.0 4.8 36.2 ;
      RECT  12.8 28.0 13.4 27.4 ;
      RECT  10.6 28.6 14.2 28.0 ;
      RECT  4.0 32.4 9.6 32.2 ;
      RECT  4.8 35.4 15.8 34.8 ;
      RECT  21.6 32.0 22.4 23.4 ;
      RECT  12.8 39.0 13.4 38.4 ;
      RECT  8.4 41.0 9.2 39.6 ;
      RECT  10.6 28.8 11.4 28.6 ;
      RECT  16.8 28.2 17.6 27.4 ;
      RECT  13.2 31.4 13.8 30.2 ;
      RECT  7.2 27.4 9.2 26.8 ;
      RECT  14.4 41.6 15.2 39.0 ;
      RECT  10.6 38.4 13.4 37.8 ;
      RECT  7.2 39.6 9.2 39.0 ;
      RECT  21.6 36.0 22.4 32.6 ;
      RECT  17.0 27.4 18.2 23.4 ;
      RECT  5.6 31.2 6.4 22.8 ;
      RECT  7.2 30.8 12.6 30.2 ;
      RECT  15.2 34.8 15.8 31.6 ;
      RECT  2.8 22.8 24.6 21.6 ;
      RECT  18.2 32.6 22.4 32.0 ;
      RECT  20.0 31.4 20.8 22.8 ;
      RECT  23.2 41.6 24.0 40.2 ;
      RECT  17.0 31.0 17.6 30.0 ;
      RECT  15.2 31.6 17.6 31.0 ;
      RECT  4.0 31.8 4.8 23.4 ;
      RECT  16.8 39.6 18.2 39.0 ;
      RECT  13.2 30.2 15.4 29.6 ;
      RECT  8.4 26.8 9.2 23.4 ;
      RECT  6.2 33.6 11.2 33.0 ;
      RECT  23.2 24.4 24.0 22.8 ;
      RECT  16.8 34.0 20.6 33.4 ;
      RECT  16.8 39.0 17.6 38.2 ;
      RECT  2.8 42.8 24.6 41.6 ;
      RECT  10.4 33.0 11.2 32.8 ;
      RECT  7.8 34.8 8.6 34.6 ;
      RECT  13.4 28.8 14.2 28.6 ;
      RECT  21.6 41.0 22.4 36.6 ;
      RECT  4.8 35.6 6.4 35.4 ;
      RECT  7.2 28.2 8.0 27.4 ;
      RECT  12.8 41.0 13.6 39.0 ;
      RECT  6.2 33.8 7.0 33.6 ;
      RECT  7.2 30.2 8.0 30.0 ;
      RECT  18.6 36.8 19.4 36.6 ;
      RECT  8.8 38.4 9.6 37.6 ;
      RECT  20.0 41.6 20.8 37.2 ;
      RECT  14.6 30.4 15.4 30.2 ;
      RECT  11.0 41.6 12.0 39.0 ;
      RECT  9.0 37.6 9.6 35.4 ;
      RECT  14.4 27.4 15.2 22.8 ;
      RECT  11.2 27.4 12.0 22.8 ;
      RECT  14.6 35.6 15.4 35.4 ;
      RECT  9.0 31.8 13.8 31.4 ;
      RECT  4.0 32.2 9.8 32.0 ;
      RECT  12.8 27.4 13.6 23.4 ;
      RECT  19.8 33.4 20.6 33.2 ;
      RECT  4.0 32.0 13.8 31.8 ;
      RECT  11.8 30.2 12.6 30.0 ;
      RECT  17.0 41.0 18.2 39.6 ;
      RECT  10.6 37.8 11.4 37.6 ;
      RECT  17.0 30.0 18.4 29.2 ;
      RECT  18.2 32.8 19.0 32.6 ;
      RECT  7.2 39.0 8.0 38.2 ;
      RECT  5.6 41.6 6.4 37.0 ;
      RECT  18.6 36.6 22.4 36.0 ;
      RECT  29.0 23.5 29.8 22.2 ;
      RECT  29.0 42.2 29.8 40.9 ;
      RECT  25.8 40.9 26.6 42.5 ;
      RECT  25.8 25.1 26.6 21.9 ;
      RECT  27.5 40.9 28.1 24.3 ;
      RECT  25.8 25.1 26.6 24.3 ;
      RECT  27.4 25.1 28.2 24.3 ;
      RECT  27.4 25.1 28.2 24.3 ;
      RECT  25.8 25.1 26.6 24.3 ;
      RECT  25.8 40.9 26.6 40.1 ;
      RECT  27.4 40.9 28.2 40.1 ;
      RECT  27.4 40.9 28.2 40.1 ;
      RECT  25.8 40.9 26.6 40.1 ;
      RECT  29.0 23.9 29.8 23.1 ;
      RECT  29.0 41.3 29.8 40.5 ;
      RECT  26.0 33.0 26.8 32.2 ;
      RECT  26.0 33.0 26.8 32.2 ;
      RECT  27.8 32.9 28.4 32.3 ;
      RECT  24.6 22.5 31.0 21.9 ;
      RECT  24.6 42.5 31.0 41.9 ;
      RECT  35.4 23.5 36.2 22.2 ;
      RECT  35.4 42.2 36.2 40.9 ;
      RECT  32.2 40.1 33.0 42.5 ;
      RECT  32.2 26.7 33.0 21.9 ;
      RECT  33.9 40.1 34.5 25.9 ;
      RECT  32.2 26.7 33.0 25.9 ;
      RECT  33.8 26.7 34.6 25.9 ;
      RECT  33.8 26.7 34.6 25.9 ;
      RECT  32.2 26.7 33.0 25.9 ;
      RECT  32.2 40.1 33.0 39.3 ;
      RECT  33.8 40.1 34.6 39.3 ;
      RECT  33.8 40.1 34.6 39.3 ;
      RECT  32.2 40.1 33.0 39.3 ;
      RECT  35.4 23.9 36.2 23.1 ;
      RECT  35.4 41.3 36.2 40.5 ;
      RECT  32.4 33.4 33.2 32.6 ;
      RECT  32.4 33.4 33.2 32.6 ;
      RECT  34.2 33.3 34.8 32.7 ;
      RECT  31.0 22.5 37.4 21.9 ;
      RECT  31.0 42.5 37.4 41.9 ;
      RECT  26.0 33.0 26.8 32.2 ;
      RECT  35.5 34.8 36.3 34.0 ;
      RECT  30.0 31.6 30.8 30.8 ;
      RECT  2.8 22.8 37.4 21.6 ;
      RECT  2.8 42.8 37.4 41.6 ;
      RECT  2.4 21.8 3.2 22.6 ;
      RECT  2.4 1.8 3.2 2.6 ;
      RECT  2.4 21.8 3.2 22.6 ;
      RECT  2.4 41.8 3.2 42.6 ;
      RECT  53.2 11.5 53.8 12.1 ;
      RECT  53.2 11.8 53.8 12.0 ;
      RECT  53.5 11.5 58.2 12.1 ;
      RECT  59.6 10.9 60.2 11.5 ;
      RECT  59.6 11.2 60.2 11.8 ;
      RECT  59.9 10.9 64.6 11.5 ;
      RECT  66.3 10.9 71.0 11.5 ;
      RECT  54.4 20.9 55.2 22.2 ;
      RECT  54.4 2.2 55.2 3.5 ;
      RECT  51.2 3.1 52.0 1.9 ;
      RECT  51.2 20.1 52.0 22.5 ;
      RECT  52.9 3.1 53.5 20.9 ;
      RECT  51.2 20.1 52.0 20.9 ;
      RECT  52.8 20.1 53.6 20.9 ;
      RECT  52.8 20.1 53.6 20.9 ;
      RECT  51.2 20.1 52.0 20.9 ;
      RECT  51.2 3.1 52.0 3.9 ;
      RECT  52.8 3.1 53.6 3.9 ;
      RECT  52.8 3.1 53.6 3.9 ;
      RECT  51.2 3.1 52.0 3.9 ;
      RECT  54.4 20.5 55.2 21.3 ;
      RECT  54.4 3.1 55.2 3.9 ;
      RECT  51.4 11.6 52.2 12.4 ;
      RECT  51.4 11.6 52.2 12.4 ;
      RECT  53.2 11.7 53.8 12.3 ;
      RECT  50.0 21.9 56.4 22.5 ;
      RECT  50.0 1.9 56.4 2.5 ;
      RECT  60.8 20.9 61.6 22.2 ;
      RECT  60.8 2.2 61.6 3.5 ;
      RECT  57.6 3.5 58.4 1.9 ;
      RECT  57.6 19.3 58.4 22.5 ;
      RECT  59.3 3.5 59.9 20.1 ;
      RECT  57.6 19.3 58.4 20.1 ;
      RECT  59.2 19.3 60.0 20.1 ;
      RECT  59.2 19.3 60.0 20.1 ;
      RECT  57.6 19.3 58.4 20.1 ;
      RECT  57.6 3.5 58.4 4.3 ;
      RECT  59.2 3.5 60.0 4.3 ;
      RECT  59.2 3.5 60.0 4.3 ;
      RECT  57.6 3.5 58.4 4.3 ;
      RECT  60.8 20.5 61.6 21.3 ;
      RECT  60.8 3.1 61.6 3.9 ;
      RECT  57.8 11.4 58.6 12.2 ;
      RECT  57.8 11.4 58.6 12.2 ;
      RECT  59.6 11.5 60.2 12.1 ;
      RECT  56.4 21.9 62.8 22.5 ;
      RECT  56.4 1.9 62.8 2.5 ;
      RECT  67.2 20.9 68.0 22.2 ;
      RECT  67.2 2.2 68.0 3.5 ;
      RECT  64.0 4.7 64.8 1.9 ;
      RECT  64.0 16.9 64.8 22.5 ;
      RECT  65.7 4.7 66.3 17.7 ;
      RECT  64.0 16.9 64.8 17.7 ;
      RECT  65.6 16.9 66.4 17.7 ;
      RECT  65.6 16.9 66.4 17.7 ;
      RECT  64.0 16.9 64.8 17.7 ;
      RECT  64.0 4.7 64.8 5.5 ;
      RECT  65.6 4.7 66.4 5.5 ;
      RECT  65.6 4.7 66.4 5.5 ;
      RECT  64.0 4.7 64.8 5.5 ;
      RECT  67.2 20.5 68.0 21.3 ;
      RECT  67.2 3.1 68.0 3.9 ;
      RECT  64.2 10.8 65.0 11.6 ;
      RECT  64.2 10.8 65.0 11.6 ;
      RECT  66.0 10.9 66.6 11.5 ;
      RECT  62.8 21.9 69.2 22.5 ;
      RECT  62.8 1.9 69.2 2.5 ;
      RECT  76.8 20.9 77.6 22.2 ;
      RECT  76.8 2.2 77.6 3.5 ;
      RECT  70.5 3.5 74.3 1.9 ;
      RECT  70.5 18.3 74.3 22.5 ;
      RECT  73.7 6.1 74.3 16.3 ;
      RECT  70.5 17.3 71.1 18.6 ;
      RECT  73.7 17.3 74.3 18.6 ;
      RECT  72.1 16.0 72.7 17.3 ;
      RECT  75.3 16.0 75.9 17.3 ;
      RECT  70.4 16.9 71.2 17.7 ;
      RECT  73.6 16.9 74.4 17.7 ;
      RECT  72.0 16.9 72.8 17.7 ;
      RECT  75.2 16.9 76.0 17.7 ;
      RECT  72.1 15.7 75.9 16.3 ;
      RECT  70.5 18.3 74.3 18.9 ;
      RECT  70.5 3.8 71.1 5.1 ;
      RECT  73.7 3.8 74.3 5.1 ;
      RECT  72.1 5.1 72.7 6.4 ;
      RECT  75.3 5.1 75.9 6.4 ;
      RECT  70.4 4.7 71.2 5.5 ;
      RECT  73.6 4.7 74.4 5.5 ;
      RECT  72.0 4.7 72.8 5.5 ;
      RECT  75.2 4.7 76.0 5.5 ;
      RECT  72.1 6.1 75.9 6.7 ;
      RECT  70.5 3.5 74.3 4.1 ;
      RECT  76.8 20.5 77.6 21.3 ;
      RECT  76.8 3.1 77.6 3.9 ;
      RECT  70.6 10.8 71.4 11.6 ;
      RECT  70.6 10.8 71.4 11.6 ;
      RECT  74.0 10.9 74.6 11.5 ;
      RECT  69.2 21.9 78.8 22.5 ;
      RECT  69.2 1.9 78.8 2.5 ;
      RECT  51.4 11.6 52.2 12.4 ;
      RECT  74.0 10.9 74.6 11.5 ;
      RECT  50.0 21.9 50.6 22.5 ;
      RECT  50.0 1.9 50.6 2.5 ;
      RECT  54.4 23.5 55.2 22.2 ;
      RECT  54.4 42.2 55.2 40.9 ;
      RECT  51.2 41.3 52.0 42.5 ;
      RECT  51.2 24.3 52.0 21.9 ;
      RECT  52.9 41.3 53.5 23.5 ;
      RECT  51.2 24.3 52.0 23.5 ;
      RECT  52.8 24.3 53.6 23.5 ;
      RECT  52.8 24.3 53.6 23.5 ;
      RECT  51.2 24.3 52.0 23.5 ;
      RECT  51.2 41.3 52.0 40.5 ;
      RECT  52.8 41.3 53.6 40.5 ;
      RECT  52.8 41.3 53.6 40.5 ;
      RECT  51.2 41.3 52.0 40.5 ;
      RECT  54.4 23.9 55.2 23.1 ;
      RECT  54.4 41.3 55.2 40.5 ;
      RECT  51.4 32.8 52.2 32.0 ;
      RECT  51.4 32.8 52.2 32.0 ;
      RECT  53.2 32.7 53.8 32.1 ;
      RECT  50.0 22.5 56.4 21.9 ;
      RECT  50.0 42.5 56.4 41.9 ;
      RECT  64.9 37.7 65.5 37.1 ;
      RECT  64.9 32.7 65.5 32.1 ;
      RECT  62.6 37.7 65.2 37.1 ;
      RECT  64.9 37.4 65.5 32.4 ;
      RECT  65.2 32.7 67.8 32.1 ;
      RECT  57.6 40.9 58.4 42.5 ;
      RECT  57.6 24.3 58.4 21.9 ;
      RECT  60.8 24.3 61.6 21.9 ;
      RECT  62.4 23.5 63.2 22.2 ;
      RECT  62.4 42.2 63.2 40.9 ;
      RECT  57.6 24.3 58.4 23.5 ;
      RECT  59.2 24.3 60.0 23.5 ;
      RECT  59.2 24.3 60.0 23.5 ;
      RECT  57.6 24.3 58.4 23.5 ;
      RECT  59.2 24.3 60.0 23.5 ;
      RECT  60.8 24.3 61.6 23.5 ;
      RECT  60.8 24.3 61.6 23.5 ;
      RECT  59.2 24.3 60.0 23.5 ;
      RECT  57.6 40.9 58.4 40.1 ;
      RECT  59.2 40.9 60.0 40.1 ;
      RECT  59.2 40.9 60.0 40.1 ;
      RECT  57.6 40.9 58.4 40.1 ;
      RECT  59.2 40.9 60.0 40.1 ;
      RECT  60.8 40.9 61.6 40.1 ;
      RECT  60.8 40.9 61.6 40.1 ;
      RECT  59.2 40.9 60.0 40.1 ;
      RECT  62.4 23.9 63.2 23.1 ;
      RECT  62.4 41.3 63.2 40.5 ;
      RECT  60.0 39.2 60.8 38.4 ;
      RECT  58.0 37.8 58.8 37.0 ;
      RECT  59.2 24.3 60.0 23.5 ;
      RECT  60.8 40.9 61.6 40.1 ;
      RECT  62.2 37.8 63.0 37.0 ;
      RECT  58.0 37.8 58.8 37.0 ;
      RECT  60.0 39.2 60.8 38.4 ;
      RECT  62.2 37.8 63.0 37.0 ;
      RECT  56.4 22.5 66.0 21.9 ;
      RECT  56.4 42.5 66.0 41.9 ;
      RECT  69.5 32.7 74.2 32.1 ;
      RECT  75.6 33.3 76.2 32.7 ;
      RECT  75.6 33.0 76.2 32.4 ;
      RECT  75.9 33.3 80.6 32.7 ;
      RECT  70.4 23.5 71.2 22.2 ;
      RECT  70.4 42.2 71.2 40.9 ;
      RECT  67.2 41.3 68.0 42.5 ;
      RECT  67.2 24.3 68.0 21.9 ;
      RECT  68.9 41.3 69.5 23.5 ;
      RECT  67.2 24.3 68.0 23.5 ;
      RECT  68.8 24.3 69.6 23.5 ;
      RECT  68.8 24.3 69.6 23.5 ;
      RECT  67.2 24.3 68.0 23.5 ;
      RECT  67.2 41.3 68.0 40.5 ;
      RECT  68.8 41.3 69.6 40.5 ;
      RECT  68.8 41.3 69.6 40.5 ;
      RECT  67.2 41.3 68.0 40.5 ;
      RECT  70.4 23.9 71.2 23.1 ;
      RECT  70.4 41.3 71.2 40.5 ;
      RECT  67.4 32.8 68.2 32.0 ;
      RECT  67.4 32.8 68.2 32.0 ;
      RECT  69.2 32.7 69.8 32.1 ;
      RECT  66.0 22.5 72.4 21.9 ;
      RECT  66.0 42.5 72.4 41.9 ;
      RECT  76.8 23.5 77.6 22.2 ;
      RECT  76.8 42.2 77.6 40.9 ;
      RECT  73.6 41.3 74.4 42.5 ;
      RECT  73.6 24.3 74.4 21.9 ;
      RECT  75.3 41.3 75.9 23.5 ;
      RECT  73.6 24.3 74.4 23.5 ;
      RECT  75.2 24.3 76.0 23.5 ;
      RECT  75.2 24.3 76.0 23.5 ;
      RECT  73.6 24.3 74.4 23.5 ;
      RECT  73.6 41.3 74.4 40.5 ;
      RECT  75.2 41.3 76.0 40.5 ;
      RECT  75.2 41.3 76.0 40.5 ;
      RECT  73.6 41.3 74.4 40.5 ;
      RECT  76.8 23.9 77.6 23.1 ;
      RECT  76.8 41.3 77.6 40.5 ;
      RECT  73.8 32.8 74.6 32.0 ;
      RECT  73.8 32.8 74.6 32.0 ;
      RECT  75.6 32.7 76.2 32.1 ;
      RECT  72.4 22.5 78.8 21.9 ;
      RECT  72.4 42.5 78.8 41.9 ;
      RECT  83.2 23.5 84.0 22.2 ;
      RECT  83.2 42.2 84.0 40.9 ;
      RECT  80.0 40.1 80.8 42.5 ;
      RECT  80.0 26.7 80.8 21.9 ;
      RECT  81.7 40.1 82.3 25.9 ;
      RECT  80.0 26.7 80.8 25.9 ;
      RECT  81.6 26.7 82.4 25.9 ;
      RECT  81.6 26.7 82.4 25.9 ;
      RECT  80.0 26.7 80.8 25.9 ;
      RECT  80.0 40.1 80.8 39.3 ;
      RECT  81.6 40.1 82.4 39.3 ;
      RECT  81.6 40.1 82.4 39.3 ;
      RECT  80.0 40.1 80.8 39.3 ;
      RECT  83.2 23.9 84.0 23.1 ;
      RECT  83.2 41.3 84.0 40.5 ;
      RECT  80.2 33.4 81.0 32.6 ;
      RECT  80.2 33.4 81.0 32.6 ;
      RECT  82.0 33.3 82.6 32.7 ;
      RECT  78.8 22.5 85.2 21.9 ;
      RECT  78.8 42.5 85.2 41.9 ;
      RECT  67.4 32.8 68.2 32.0 ;
      RECT  82.0 33.3 82.6 32.7 ;
      RECT  66.0 22.5 66.6 21.9 ;
      RECT  66.0 42.5 66.6 41.9 ;
      RECT  58.0 37.8 58.8 37.0 ;
      RECT  60.0 39.2 60.8 38.4 ;
      RECT  82.0 33.3 82.6 32.7 ;
      RECT  56.4 22.5 85.2 21.9 ;
      RECT  56.4 42.5 85.2 41.9 ;
      RECT  58.5 46.7 59.1 47.3 ;
      RECT  58.5 51.7 59.1 52.3 ;
      RECT  56.2 46.7 58.8 47.3 ;
      RECT  58.5 47.0 59.1 52.0 ;
      RECT  58.8 51.7 61.4 52.3 ;
      RECT  51.2 43.5 52.0 41.9 ;
      RECT  51.2 60.1 52.0 62.5 ;
      RECT  54.4 60.1 55.2 62.5 ;
      RECT  56.0 60.9 56.8 62.2 ;
      RECT  56.0 42.2 56.8 43.5 ;
      RECT  51.2 60.1 52.0 60.9 ;
      RECT  52.8 60.1 53.6 60.9 ;
      RECT  52.8 60.1 53.6 60.9 ;
      RECT  51.2 60.1 52.0 60.9 ;
      RECT  52.8 60.1 53.6 60.9 ;
      RECT  54.4 60.1 55.2 60.9 ;
      RECT  54.4 60.1 55.2 60.9 ;
      RECT  52.8 60.1 53.6 60.9 ;
      RECT  51.2 43.5 52.0 44.3 ;
      RECT  52.8 43.5 53.6 44.3 ;
      RECT  52.8 43.5 53.6 44.3 ;
      RECT  51.2 43.5 52.0 44.3 ;
      RECT  52.8 43.5 53.6 44.3 ;
      RECT  54.4 43.5 55.2 44.3 ;
      RECT  54.4 43.5 55.2 44.3 ;
      RECT  52.8 43.5 53.6 44.3 ;
      RECT  56.0 60.5 56.8 61.3 ;
      RECT  56.0 43.1 56.8 43.9 ;
      RECT  53.6 45.2 54.4 46.0 ;
      RECT  51.6 46.6 52.4 47.4 ;
      RECT  52.8 60.1 53.6 60.9 ;
      RECT  54.4 43.5 55.2 44.3 ;
      RECT  55.8 46.6 56.6 47.4 ;
      RECT  51.6 46.6 52.4 47.4 ;
      RECT  53.6 45.2 54.4 46.0 ;
      RECT  55.8 46.6 56.6 47.4 ;
      RECT  50.0 61.9 59.6 62.5 ;
      RECT  50.0 41.9 59.6 42.5 ;
      RECT  63.1 51.7 67.8 52.3 ;
      RECT  69.2 51.1 69.8 51.7 ;
      RECT  69.2 51.4 69.8 52.0 ;
      RECT  69.5 51.1 74.2 51.7 ;
      RECT  64.0 60.9 64.8 62.2 ;
      RECT  64.0 42.2 64.8 43.5 ;
      RECT  60.8 43.1 61.6 41.9 ;
      RECT  60.8 60.1 61.6 62.5 ;
      RECT  62.5 43.1 63.1 60.9 ;
      RECT  60.8 60.1 61.6 60.9 ;
      RECT  62.4 60.1 63.2 60.9 ;
      RECT  62.4 60.1 63.2 60.9 ;
      RECT  60.8 60.1 61.6 60.9 ;
      RECT  60.8 43.1 61.6 43.9 ;
      RECT  62.4 43.1 63.2 43.9 ;
      RECT  62.4 43.1 63.2 43.9 ;
      RECT  60.8 43.1 61.6 43.9 ;
      RECT  64.0 60.5 64.8 61.3 ;
      RECT  64.0 43.1 64.8 43.9 ;
      RECT  61.0 51.6 61.8 52.4 ;
      RECT  61.0 51.6 61.8 52.4 ;
      RECT  62.8 51.7 63.4 52.3 ;
      RECT  59.6 61.9 66.0 62.5 ;
      RECT  59.6 41.9 66.0 42.5 ;
      RECT  70.4 60.9 71.2 62.2 ;
      RECT  70.4 42.2 71.2 43.5 ;
      RECT  67.2 43.1 68.0 41.9 ;
      RECT  67.2 60.1 68.0 62.5 ;
      RECT  68.9 43.1 69.5 60.9 ;
      RECT  67.2 60.1 68.0 60.9 ;
      RECT  68.8 60.1 69.6 60.9 ;
      RECT  68.8 60.1 69.6 60.9 ;
      RECT  67.2 60.1 68.0 60.9 ;
      RECT  67.2 43.1 68.0 43.9 ;
      RECT  68.8 43.1 69.6 43.9 ;
      RECT  68.8 43.1 69.6 43.9 ;
      RECT  67.2 43.1 68.0 43.9 ;
      RECT  70.4 60.5 71.2 61.3 ;
      RECT  70.4 43.1 71.2 43.9 ;
      RECT  67.4 51.6 68.2 52.4 ;
      RECT  67.4 51.6 68.2 52.4 ;
      RECT  69.2 51.7 69.8 52.3 ;
      RECT  66.0 61.9 72.4 62.5 ;
      RECT  66.0 41.9 72.4 42.5 ;
      RECT  76.8 60.9 77.6 62.2 ;
      RECT  76.8 42.2 77.6 43.5 ;
      RECT  73.6 44.3 74.4 41.9 ;
      RECT  73.6 57.7 74.4 62.5 ;
      RECT  75.3 44.3 75.9 58.5 ;
      RECT  73.6 57.7 74.4 58.5 ;
      RECT  75.2 57.7 76.0 58.5 ;
      RECT  75.2 57.7 76.0 58.5 ;
      RECT  73.6 57.7 74.4 58.5 ;
      RECT  73.6 44.3 74.4 45.1 ;
      RECT  75.2 44.3 76.0 45.1 ;
      RECT  75.2 44.3 76.0 45.1 ;
      RECT  73.6 44.3 74.4 45.1 ;
      RECT  76.8 60.5 77.6 61.3 ;
      RECT  76.8 43.1 77.6 43.9 ;
      RECT  73.8 51.0 74.6 51.8 ;
      RECT  73.8 51.0 74.6 51.8 ;
      RECT  75.6 51.1 76.2 51.7 ;
      RECT  72.4 61.9 78.8 62.5 ;
      RECT  72.4 41.9 78.8 42.5 ;
      RECT  61.0 51.6 61.8 52.4 ;
      RECT  75.6 51.1 76.2 51.7 ;
      RECT  59.6 61.9 60.2 62.5 ;
      RECT  59.6 41.9 60.2 42.5 ;
      RECT  51.6 46.6 52.4 47.4 ;
      RECT  53.6 45.2 54.4 46.0 ;
      RECT  75.6 51.1 76.2 51.7 ;
      RECT  50.0 61.9 78.8 62.5 ;
      RECT  50.0 41.9 78.8 42.5 ;
      RECT  53.5 72.7 58.2 72.1 ;
      RECT  59.6 72.9 60.2 72.3 ;
      RECT  59.6 72.6 60.2 72.4 ;
      RECT  59.9 72.9 64.6 72.3 ;
      RECT  66.0 73.5 66.6 72.9 ;
      RECT  66.0 73.2 66.6 72.6 ;
      RECT  66.3 73.5 71.0 72.9 ;
      RECT  54.4 63.5 55.2 62.2 ;
      RECT  54.4 82.2 55.2 80.9 ;
      RECT  51.2 81.3 52.0 82.5 ;
      RECT  51.2 64.3 52.0 61.9 ;
      RECT  52.9 81.3 53.5 63.5 ;
      RECT  51.2 64.3 52.0 63.5 ;
      RECT  52.8 64.3 53.6 63.5 ;
      RECT  52.8 64.3 53.6 63.5 ;
      RECT  51.2 64.3 52.0 63.5 ;
      RECT  51.2 81.3 52.0 80.5 ;
      RECT  52.8 81.3 53.6 80.5 ;
      RECT  52.8 81.3 53.6 80.5 ;
      RECT  51.2 81.3 52.0 80.5 ;
      RECT  54.4 63.9 55.2 63.1 ;
      RECT  54.4 81.3 55.2 80.5 ;
      RECT  51.4 72.8 52.2 72.0 ;
      RECT  51.4 72.8 52.2 72.0 ;
      RECT  53.2 72.7 53.8 72.1 ;
      RECT  50.0 62.5 56.4 61.9 ;
      RECT  50.0 82.5 56.4 81.9 ;
      RECT  60.8 63.5 61.6 62.2 ;
      RECT  60.8 82.2 61.6 80.9 ;
      RECT  57.6 81.3 58.4 82.5 ;
      RECT  57.6 64.3 58.4 61.9 ;
      RECT  59.3 81.3 59.9 63.5 ;
      RECT  57.6 64.3 58.4 63.5 ;
      RECT  59.2 64.3 60.0 63.5 ;
      RECT  59.2 64.3 60.0 63.5 ;
      RECT  57.6 64.3 58.4 63.5 ;
      RECT  57.6 81.3 58.4 80.5 ;
      RECT  59.2 81.3 60.0 80.5 ;
      RECT  59.2 81.3 60.0 80.5 ;
      RECT  57.6 81.3 58.4 80.5 ;
      RECT  60.8 63.9 61.6 63.1 ;
      RECT  60.8 81.3 61.6 80.5 ;
      RECT  57.8 72.8 58.6 72.0 ;
      RECT  57.8 72.8 58.6 72.0 ;
      RECT  59.6 72.7 60.2 72.1 ;
      RECT  56.4 62.5 62.8 61.9 ;
      RECT  56.4 82.5 62.8 81.9 ;
      RECT  67.2 63.5 68.0 62.2 ;
      RECT  67.2 82.2 68.0 80.9 ;
      RECT  64.0 80.9 64.8 82.5 ;
      RECT  64.0 65.1 64.8 61.9 ;
      RECT  65.7 80.9 66.3 64.3 ;
      RECT  64.0 65.1 64.8 64.3 ;
      RECT  65.6 65.1 66.4 64.3 ;
      RECT  65.6 65.1 66.4 64.3 ;
      RECT  64.0 65.1 64.8 64.3 ;
      RECT  64.0 80.9 64.8 80.1 ;
      RECT  65.6 80.9 66.4 80.1 ;
      RECT  65.6 80.9 66.4 80.1 ;
      RECT  64.0 80.9 64.8 80.1 ;
      RECT  67.2 63.9 68.0 63.1 ;
      RECT  67.2 81.3 68.0 80.5 ;
      RECT  64.2 73.0 65.0 72.2 ;
      RECT  64.2 73.0 65.0 72.2 ;
      RECT  66.0 72.9 66.6 72.3 ;
      RECT  62.8 62.5 69.2 61.9 ;
      RECT  62.8 82.5 69.2 81.9 ;
      RECT  73.6 63.5 74.4 62.2 ;
      RECT  73.6 82.2 74.4 80.9 ;
      RECT  70.4 79.7 71.2 82.5 ;
      RECT  70.4 67.5 71.2 61.9 ;
      RECT  72.1 79.7 72.7 66.7 ;
      RECT  70.4 67.5 71.2 66.7 ;
      RECT  72.0 67.5 72.8 66.7 ;
      RECT  72.0 67.5 72.8 66.7 ;
      RECT  70.4 67.5 71.2 66.7 ;
      RECT  70.4 79.7 71.2 78.9 ;
      RECT  72.0 79.7 72.8 78.9 ;
      RECT  72.0 79.7 72.8 78.9 ;
      RECT  70.4 79.7 71.2 78.9 ;
      RECT  73.6 63.9 74.4 63.1 ;
      RECT  73.6 81.3 74.4 80.5 ;
      RECT  70.6 73.6 71.4 72.8 ;
      RECT  70.6 73.6 71.4 72.8 ;
      RECT  72.4 73.5 73.0 72.9 ;
      RECT  69.2 62.5 75.6 61.9 ;
      RECT  69.2 82.5 75.6 81.9 ;
      RECT  51.4 72.8 52.2 72.0 ;
      RECT  72.4 73.5 73.0 72.9 ;
      RECT  50.0 62.5 50.6 61.9 ;
      RECT  50.0 82.5 50.6 81.9 ;
      RECT  54.4 140.9 55.2 142.2 ;
      RECT  54.4 122.2 55.2 123.5 ;
      RECT  51.2 123.1 52.0 121.9 ;
      RECT  51.2 140.1 52.0 142.5 ;
      RECT  52.9 123.1 53.5 140.9 ;
      RECT  51.2 140.1 52.0 140.9 ;
      RECT  52.8 140.1 53.6 140.9 ;
      RECT  52.8 140.1 53.6 140.9 ;
      RECT  51.2 140.1 52.0 140.9 ;
      RECT  51.2 123.1 52.0 123.9 ;
      RECT  52.8 123.1 53.6 123.9 ;
      RECT  52.8 123.1 53.6 123.9 ;
      RECT  51.2 123.1 52.0 123.9 ;
      RECT  54.4 140.5 55.2 141.3 ;
      RECT  54.4 123.1 55.2 123.9 ;
      RECT  51.4 131.6 52.2 132.4 ;
      RECT  51.4 131.6 52.2 132.4 ;
      RECT  53.2 131.7 53.8 132.3 ;
      RECT  50.0 141.9 56.4 142.5 ;
      RECT  50.0 121.9 56.4 122.5 ;
      RECT  59.0 87.6 59.6 88.2 ;
      RECT  59.0 90.9 59.6 91.5 ;
      RECT  56.4 87.6 59.3 88.2 ;
      RECT  59.0 87.9 59.6 91.2 ;
      RECT  59.3 90.9 62.2 91.5 ;
      RECT  51.2 83.5 52.0 81.9 ;
      RECT  51.2 100.1 52.0 102.5 ;
      RECT  54.4 100.1 55.2 102.5 ;
      RECT  57.6 100.9 58.4 102.2 ;
      RECT  57.6 82.2 58.4 83.5 ;
      RECT  51.2 100.1 52.0 100.9 ;
      RECT  52.8 100.1 53.6 100.9 ;
      RECT  52.8 100.1 53.6 100.9 ;
      RECT  51.2 100.1 52.0 100.9 ;
      RECT  52.8 100.1 53.6 100.9 ;
      RECT  54.4 100.1 55.2 100.9 ;
      RECT  54.4 100.1 55.2 100.9 ;
      RECT  52.8 100.1 53.6 100.9 ;
      RECT  54.4 100.1 55.2 100.9 ;
      RECT  56.0 100.1 56.8 100.9 ;
      RECT  56.0 100.1 56.8 100.9 ;
      RECT  54.4 100.1 55.2 100.9 ;
      RECT  51.2 83.5 52.0 84.3 ;
      RECT  52.8 83.5 53.6 84.3 ;
      RECT  52.8 83.5 53.6 84.3 ;
      RECT  51.2 83.5 52.0 84.3 ;
      RECT  52.8 83.5 53.6 84.3 ;
      RECT  54.4 83.5 55.2 84.3 ;
      RECT  54.4 83.5 55.2 84.3 ;
      RECT  52.8 83.5 53.6 84.3 ;
      RECT  54.4 83.5 55.2 84.3 ;
      RECT  56.0 83.5 56.8 84.3 ;
      RECT  56.0 83.5 56.8 84.3 ;
      RECT  54.4 83.5 55.2 84.3 ;
      RECT  57.6 100.5 58.4 101.3 ;
      RECT  57.6 83.1 58.4 83.9 ;
      RECT  55.2 84.9 56.0 85.7 ;
      RECT  53.6 86.2 54.4 87.0 ;
      RECT  52.0 87.5 52.8 88.3 ;
      RECT  52.8 100.1 53.6 100.9 ;
      RECT  56.0 100.1 56.8 100.9 ;
      RECT  56.0 83.5 56.8 84.3 ;
      RECT  56.0 87.5 56.8 88.3 ;
      RECT  52.0 87.5 52.8 88.3 ;
      RECT  53.6 86.2 54.4 87.0 ;
      RECT  55.2 84.9 56.0 85.7 ;
      RECT  56.0 87.5 56.8 88.3 ;
      RECT  50.0 101.9 60.4 102.5 ;
      RECT  50.0 81.9 60.4 82.5 ;
      RECT  66.4 100.9 67.2 102.2 ;
      RECT  66.4 82.2 67.2 83.5 ;
      RECT  61.7 83.5 65.5 81.9 ;
      RECT  61.7 98.3 65.5 102.5 ;
      RECT  63.3 84.7 63.9 97.7 ;
      RECT  61.7 97.3 62.3 98.6 ;
      RECT  64.9 97.3 65.5 98.6 ;
      RECT  61.6 96.9 62.4 97.7 ;
      RECT  64.8 96.9 65.6 97.7 ;
      RECT  63.2 96.9 64.0 97.7 ;
      RECT  63.2 96.9 64.0 97.7 ;
      RECT  61.7 98.3 65.5 98.9 ;
      RECT  61.7 83.8 62.3 85.1 ;
      RECT  64.9 83.8 65.5 85.1 ;
      RECT  61.6 84.7 62.4 85.5 ;
      RECT  64.8 84.7 65.6 85.5 ;
      RECT  63.2 84.7 64.0 85.5 ;
      RECT  63.2 84.7 64.0 85.5 ;
      RECT  61.7 83.5 65.5 84.1 ;
      RECT  66.4 100.5 67.2 101.3 ;
      RECT  66.4 83.1 67.2 83.9 ;
      RECT  61.8 90.8 62.6 91.6 ;
      RECT  61.8 90.8 62.6 91.6 ;
      RECT  63.6 90.9 64.2 91.5 ;
      RECT  60.4 101.9 68.4 102.5 ;
      RECT  60.4 81.9 68.4 82.5 ;
      RECT  52.0 87.5 52.8 88.3 ;
      RECT  53.6 86.2 54.4 87.0 ;
      RECT  55.2 84.9 56.0 85.7 ;
      RECT  63.6 90.9 64.2 91.5 ;
      RECT  50.0 101.9 68.4 102.5 ;
      RECT  50.0 81.9 68.4 82.5 ;
      RECT  59.0 156.8 59.6 156.2 ;
      RECT  59.0 152.9 59.6 152.3 ;
      RECT  56.4 156.8 59.3 156.2 ;
      RECT  59.0 156.5 59.6 152.6 ;
      RECT  59.3 152.9 62.2 152.3 ;
      RECT  51.2 160.9 52.0 162.5 ;
      RECT  51.2 144.3 52.0 141.9 ;
      RECT  54.4 144.3 55.2 141.9 ;
      RECT  57.6 143.5 58.4 142.2 ;
      RECT  57.6 162.2 58.4 160.9 ;
      RECT  51.2 144.3 52.0 143.5 ;
      RECT  52.8 144.3 53.6 143.5 ;
      RECT  52.8 144.3 53.6 143.5 ;
      RECT  51.2 144.3 52.0 143.5 ;
      RECT  52.8 144.3 53.6 143.5 ;
      RECT  54.4 144.3 55.2 143.5 ;
      RECT  54.4 144.3 55.2 143.5 ;
      RECT  52.8 144.3 53.6 143.5 ;
      RECT  54.4 144.3 55.2 143.5 ;
      RECT  56.0 144.3 56.8 143.5 ;
      RECT  56.0 144.3 56.8 143.5 ;
      RECT  54.4 144.3 55.2 143.5 ;
      RECT  51.2 160.9 52.0 160.1 ;
      RECT  52.8 160.9 53.6 160.1 ;
      RECT  52.8 160.9 53.6 160.1 ;
      RECT  51.2 160.9 52.0 160.1 ;
      RECT  52.8 160.9 53.6 160.1 ;
      RECT  54.4 160.9 55.2 160.1 ;
      RECT  54.4 160.9 55.2 160.1 ;
      RECT  52.8 160.9 53.6 160.1 ;
      RECT  54.4 160.9 55.2 160.1 ;
      RECT  56.0 160.9 56.8 160.1 ;
      RECT  56.0 160.9 56.8 160.1 ;
      RECT  54.4 160.9 55.2 160.1 ;
      RECT  57.6 143.9 58.4 143.1 ;
      RECT  57.6 161.3 58.4 160.5 ;
      RECT  55.2 159.5 56.0 158.7 ;
      RECT  53.6 158.2 54.4 157.4 ;
      RECT  52.0 156.9 52.8 156.1 ;
      RECT  52.8 144.3 53.6 143.5 ;
      RECT  56.0 144.3 56.8 143.5 ;
      RECT  56.0 160.9 56.8 160.1 ;
      RECT  56.0 156.9 56.8 156.1 ;
      RECT  52.0 156.9 52.8 156.1 ;
      RECT  53.6 158.2 54.4 157.4 ;
      RECT  55.2 159.5 56.0 158.7 ;
      RECT  56.0 156.9 56.8 156.1 ;
      RECT  50.0 142.5 60.4 141.9 ;
      RECT  50.0 162.5 60.4 161.9 ;
      RECT  64.8 143.5 65.6 142.2 ;
      RECT  64.8 162.2 65.6 160.9 ;
      RECT  61.6 160.9 62.4 162.5 ;
      RECT  61.6 145.1 62.4 141.9 ;
      RECT  63.3 160.9 63.9 144.3 ;
      RECT  61.6 145.1 62.4 144.3 ;
      RECT  63.2 145.1 64.0 144.3 ;
      RECT  63.2 145.1 64.0 144.3 ;
      RECT  61.6 145.1 62.4 144.3 ;
      RECT  61.6 160.9 62.4 160.1 ;
      RECT  63.2 160.9 64.0 160.1 ;
      RECT  63.2 160.9 64.0 160.1 ;
      RECT  61.6 160.9 62.4 160.1 ;
      RECT  64.8 143.9 65.6 143.1 ;
      RECT  64.8 161.3 65.6 160.5 ;
      RECT  61.8 153.0 62.6 152.2 ;
      RECT  61.8 153.0 62.6 152.2 ;
      RECT  63.6 152.9 64.2 152.3 ;
      RECT  60.4 142.5 66.8 141.9 ;
      RECT  60.4 162.5 66.8 161.9 ;
      RECT  52.0 156.9 52.8 156.1 ;
      RECT  53.6 158.2 54.4 157.4 ;
      RECT  55.2 159.5 56.0 158.7 ;
      RECT  63.6 152.9 64.2 152.3 ;
      RECT  50.0 142.5 66.8 141.9 ;
      RECT  50.0 162.5 66.8 161.9 ;
      RECT  30.4 174.1 29.6 175.4 ;
      RECT  30.4 165.0 29.6 166.3 ;
      RECT  33.6 165.9 32.8 164.7 ;
      RECT  33.6 173.3 32.8 175.7 ;
      RECT  31.9 165.9 31.3 174.1 ;
      RECT  33.6 173.3 32.8 174.1 ;
      RECT  32.0 173.3 31.2 174.1 ;
      RECT  32.0 173.3 31.2 174.1 ;
      RECT  33.6 173.3 32.8 174.1 ;
      RECT  33.6 165.9 32.8 166.7 ;
      RECT  32.0 165.9 31.2 166.7 ;
      RECT  32.0 165.9 31.2 166.7 ;
      RECT  33.6 165.9 32.8 166.7 ;
      RECT  30.4 173.7 29.6 174.5 ;
      RECT  30.4 165.9 29.6 166.7 ;
      RECT  33.4 169.6 32.6 170.4 ;
      RECT  33.4 169.6 32.6 170.4 ;
      RECT  31.6 169.7 31.0 170.3 ;
      RECT  34.8 175.1 28.4 175.7 ;
      RECT  34.8 164.7 28.4 165.3 ;
      RECT  24.0 174.1 23.2 175.4 ;
      RECT  24.0 165.0 23.2 166.3 ;
      RECT  27.2 165.9 26.4 164.7 ;
      RECT  27.2 173.3 26.4 175.7 ;
      RECT  25.5 165.9 24.9 174.1 ;
      RECT  27.2 173.3 26.4 174.1 ;
      RECT  25.6 173.3 24.8 174.1 ;
      RECT  25.6 173.3 24.8 174.1 ;
      RECT  27.2 173.3 26.4 174.1 ;
      RECT  27.2 165.9 26.4 166.7 ;
      RECT  25.6 165.9 24.8 166.7 ;
      RECT  25.6 165.9 24.8 166.7 ;
      RECT  27.2 165.9 26.4 166.7 ;
      RECT  24.0 173.7 23.2 174.5 ;
      RECT  24.0 165.9 23.2 166.7 ;
      RECT  27.0 169.6 26.2 170.4 ;
      RECT  27.0 169.6 26.2 170.4 ;
      RECT  25.2 169.7 24.6 170.3 ;
      RECT  28.4 175.1 22.0 175.7 ;
      RECT  28.4 164.7 22.0 165.3 ;
      RECT  17.6 174.1 16.8 175.4 ;
      RECT  17.6 165.0 16.8 166.3 ;
      RECT  20.8 165.9 20.0 164.7 ;
      RECT  20.8 173.3 20.0 175.7 ;
      RECT  19.1 165.9 18.5 174.1 ;
      RECT  20.8 173.3 20.0 174.1 ;
      RECT  19.2 173.3 18.4 174.1 ;
      RECT  19.2 173.3 18.4 174.1 ;
      RECT  20.8 173.3 20.0 174.1 ;
      RECT  20.8 165.9 20.0 166.7 ;
      RECT  19.2 165.9 18.4 166.7 ;
      RECT  19.2 165.9 18.4 166.7 ;
      RECT  20.8 165.9 20.0 166.7 ;
      RECT  17.6 173.7 16.8 174.5 ;
      RECT  17.6 165.9 16.8 166.7 ;
      RECT  20.6 169.6 19.8 170.4 ;
      RECT  20.6 169.6 19.8 170.4 ;
      RECT  18.8 169.7 18.2 170.3 ;
      RECT  22.0 175.1 15.6 175.7 ;
      RECT  22.0 164.7 15.6 165.3 ;
      RECT  11.2 174.1 10.4 175.4 ;
      RECT  11.2 165.0 10.4 166.3 ;
      RECT  14.4 165.9 13.6 164.7 ;
      RECT  14.4 173.3 13.6 175.7 ;
      RECT  12.7 165.9 12.1 174.1 ;
      RECT  14.4 173.3 13.6 174.1 ;
      RECT  12.8 173.3 12.0 174.1 ;
      RECT  12.8 173.3 12.0 174.1 ;
      RECT  14.4 173.3 13.6 174.1 ;
      RECT  14.4 165.9 13.6 166.7 ;
      RECT  12.8 165.9 12.0 166.7 ;
      RECT  12.8 165.9 12.0 166.7 ;
      RECT  14.4 165.9 13.6 166.7 ;
      RECT  11.2 173.7 10.4 174.5 ;
      RECT  11.2 165.9 10.4 166.7 ;
      RECT  14.2 169.6 13.4 170.4 ;
      RECT  14.2 169.6 13.4 170.4 ;
      RECT  12.4 169.7 11.8 170.3 ;
      RECT  15.6 175.1 9.2 175.7 ;
      RECT  15.6 164.7 9.2 165.3 ;
      RECT  4.8 174.1 4.0 175.4 ;
      RECT  4.8 165.0 4.0 166.3 ;
      RECT  8.0 165.9 7.2 164.7 ;
      RECT  8.0 173.3 7.2 175.7 ;
      RECT  6.3 165.9 5.7 174.1 ;
      RECT  8.0 173.3 7.2 174.1 ;
      RECT  6.4 173.3 5.6 174.1 ;
      RECT  6.4 173.3 5.6 174.1 ;
      RECT  8.0 173.3 7.2 174.1 ;
      RECT  8.0 165.9 7.2 166.7 ;
      RECT  6.4 165.9 5.6 166.7 ;
      RECT  6.4 165.9 5.6 166.7 ;
      RECT  8.0 165.9 7.2 166.7 ;
      RECT  4.8 173.7 4.0 174.5 ;
      RECT  4.8 165.9 4.0 166.7 ;
      RECT  7.8 169.6 7.0 170.4 ;
      RECT  7.8 169.6 7.0 170.4 ;
      RECT  6.0 169.7 5.4 170.3 ;
      RECT  9.2 175.1 2.8 175.7 ;
      RECT  9.2 164.7 2.8 165.3 ;
      RECT  30.4 176.7 29.6 175.4 ;
      RECT  30.4 185.8 29.6 184.5 ;
      RECT  33.6 184.9 32.8 186.1 ;
      RECT  33.6 177.5 32.8 175.1 ;
      RECT  31.9 184.9 31.3 176.7 ;
      RECT  33.6 177.5 32.8 176.7 ;
      RECT  32.0 177.5 31.2 176.7 ;
      RECT  32.0 177.5 31.2 176.7 ;
      RECT  33.6 177.5 32.8 176.7 ;
      RECT  33.6 184.9 32.8 184.1 ;
      RECT  32.0 184.9 31.2 184.1 ;
      RECT  32.0 184.9 31.2 184.1 ;
      RECT  33.6 184.9 32.8 184.1 ;
      RECT  30.4 177.1 29.6 176.3 ;
      RECT  30.4 184.9 29.6 184.1 ;
      RECT  33.4 181.2 32.6 180.4 ;
      RECT  33.4 181.2 32.6 180.4 ;
      RECT  31.6 181.1 31.0 180.5 ;
      RECT  34.8 175.7 28.4 175.1 ;
      RECT  34.8 186.1 28.4 185.5 ;
      RECT  24.0 176.7 23.2 175.4 ;
      RECT  24.0 185.8 23.2 184.5 ;
      RECT  27.2 184.9 26.4 186.1 ;
      RECT  27.2 177.5 26.4 175.1 ;
      RECT  25.5 184.9 24.9 176.7 ;
      RECT  27.2 177.5 26.4 176.7 ;
      RECT  25.6 177.5 24.8 176.7 ;
      RECT  25.6 177.5 24.8 176.7 ;
      RECT  27.2 177.5 26.4 176.7 ;
      RECT  27.2 184.9 26.4 184.1 ;
      RECT  25.6 184.9 24.8 184.1 ;
      RECT  25.6 184.9 24.8 184.1 ;
      RECT  27.2 184.9 26.4 184.1 ;
      RECT  24.0 177.1 23.2 176.3 ;
      RECT  24.0 184.9 23.2 184.1 ;
      RECT  27.0 181.2 26.2 180.4 ;
      RECT  27.0 181.2 26.2 180.4 ;
      RECT  25.2 181.1 24.6 180.5 ;
      RECT  28.4 175.7 22.0 175.1 ;
      RECT  28.4 186.1 22.0 185.5 ;
      RECT  17.6 176.7 16.8 175.4 ;
      RECT  17.6 185.8 16.8 184.5 ;
      RECT  20.8 184.9 20.0 186.1 ;
      RECT  20.8 177.5 20.0 175.1 ;
      RECT  19.1 184.9 18.5 176.7 ;
      RECT  20.8 177.5 20.0 176.7 ;
      RECT  19.2 177.5 18.4 176.7 ;
      RECT  19.2 177.5 18.4 176.7 ;
      RECT  20.8 177.5 20.0 176.7 ;
      RECT  20.8 184.9 20.0 184.1 ;
      RECT  19.2 184.9 18.4 184.1 ;
      RECT  19.2 184.9 18.4 184.1 ;
      RECT  20.8 184.9 20.0 184.1 ;
      RECT  17.6 177.1 16.8 176.3 ;
      RECT  17.6 184.9 16.8 184.1 ;
      RECT  20.6 181.2 19.8 180.4 ;
      RECT  20.6 181.2 19.8 180.4 ;
      RECT  18.8 181.1 18.2 180.5 ;
      RECT  22.0 175.7 15.6 175.1 ;
      RECT  22.0 186.1 15.6 185.5 ;
      RECT  11.2 176.7 10.4 175.4 ;
      RECT  11.2 185.8 10.4 184.5 ;
      RECT  14.4 184.9 13.6 186.1 ;
      RECT  14.4 177.5 13.6 175.1 ;
      RECT  12.7 184.9 12.1 176.7 ;
      RECT  14.4 177.5 13.6 176.7 ;
      RECT  12.8 177.5 12.0 176.7 ;
      RECT  12.8 177.5 12.0 176.7 ;
      RECT  14.4 177.5 13.6 176.7 ;
      RECT  14.4 184.9 13.6 184.1 ;
      RECT  12.8 184.9 12.0 184.1 ;
      RECT  12.8 184.9 12.0 184.1 ;
      RECT  14.4 184.9 13.6 184.1 ;
      RECT  11.2 177.1 10.4 176.3 ;
      RECT  11.2 184.9 10.4 184.1 ;
      RECT  14.2 181.2 13.4 180.4 ;
      RECT  14.2 181.2 13.4 180.4 ;
      RECT  12.4 181.1 11.8 180.5 ;
      RECT  15.6 175.7 9.2 175.1 ;
      RECT  15.6 186.1 9.2 185.5 ;
      RECT  4.8 176.7 4.0 175.4 ;
      RECT  4.8 185.8 4.0 184.5 ;
      RECT  8.0 184.9 7.2 186.1 ;
      RECT  8.0 177.5 7.2 175.1 ;
      RECT  6.3 184.9 5.7 176.7 ;
      RECT  8.0 177.5 7.2 176.7 ;
      RECT  6.4 177.5 5.6 176.7 ;
      RECT  6.4 177.5 5.6 176.7 ;
      RECT  8.0 177.5 7.2 176.7 ;
      RECT  8.0 184.9 7.2 184.1 ;
      RECT  6.4 184.9 5.6 184.1 ;
      RECT  6.4 184.9 5.6 184.1 ;
      RECT  8.0 184.9 7.2 184.1 ;
      RECT  4.8 177.1 4.0 176.3 ;
      RECT  4.8 184.9 4.0 184.1 ;
      RECT  7.8 181.2 7.0 180.4 ;
      RECT  7.8 181.2 7.0 180.4 ;
      RECT  6.0 181.1 5.4 180.5 ;
      RECT  9.2 175.7 2.8 175.1 ;
      RECT  9.2 186.1 2.8 185.5 ;
      RECT  30.4 194.9 29.6 196.2 ;
      RECT  30.4 185.8 29.6 187.1 ;
      RECT  33.6 186.7 32.8 185.5 ;
      RECT  33.6 194.1 32.8 196.5 ;
      RECT  31.9 186.7 31.3 194.9 ;
      RECT  33.6 194.1 32.8 194.9 ;
      RECT  32.0 194.1 31.2 194.9 ;
      RECT  32.0 194.1 31.2 194.9 ;
      RECT  33.6 194.1 32.8 194.9 ;
      RECT  33.6 186.7 32.8 187.5 ;
      RECT  32.0 186.7 31.2 187.5 ;
      RECT  32.0 186.7 31.2 187.5 ;
      RECT  33.6 186.7 32.8 187.5 ;
      RECT  30.4 194.5 29.6 195.3 ;
      RECT  30.4 186.7 29.6 187.5 ;
      RECT  33.4 190.4 32.6 191.2 ;
      RECT  33.4 190.4 32.6 191.2 ;
      RECT  31.6 190.5 31.0 191.1 ;
      RECT  34.8 195.9 28.4 196.5 ;
      RECT  34.8 185.5 28.4 186.1 ;
      RECT  24.0 194.9 23.2 196.2 ;
      RECT  24.0 185.8 23.2 187.1 ;
      RECT  27.2 186.7 26.4 185.5 ;
      RECT  27.2 194.1 26.4 196.5 ;
      RECT  25.5 186.7 24.9 194.9 ;
      RECT  27.2 194.1 26.4 194.9 ;
      RECT  25.6 194.1 24.8 194.9 ;
      RECT  25.6 194.1 24.8 194.9 ;
      RECT  27.2 194.1 26.4 194.9 ;
      RECT  27.2 186.7 26.4 187.5 ;
      RECT  25.6 186.7 24.8 187.5 ;
      RECT  25.6 186.7 24.8 187.5 ;
      RECT  27.2 186.7 26.4 187.5 ;
      RECT  24.0 194.5 23.2 195.3 ;
      RECT  24.0 186.7 23.2 187.5 ;
      RECT  27.0 190.4 26.2 191.2 ;
      RECT  27.0 190.4 26.2 191.2 ;
      RECT  25.2 190.5 24.6 191.1 ;
      RECT  28.4 195.9 22.0 196.5 ;
      RECT  28.4 185.5 22.0 186.1 ;
      RECT  17.6 194.9 16.8 196.2 ;
      RECT  17.6 185.8 16.8 187.1 ;
      RECT  20.8 186.7 20.0 185.5 ;
      RECT  20.8 194.1 20.0 196.5 ;
      RECT  19.1 186.7 18.5 194.9 ;
      RECT  20.8 194.1 20.0 194.9 ;
      RECT  19.2 194.1 18.4 194.9 ;
      RECT  19.2 194.1 18.4 194.9 ;
      RECT  20.8 194.1 20.0 194.9 ;
      RECT  20.8 186.7 20.0 187.5 ;
      RECT  19.2 186.7 18.4 187.5 ;
      RECT  19.2 186.7 18.4 187.5 ;
      RECT  20.8 186.7 20.0 187.5 ;
      RECT  17.6 194.5 16.8 195.3 ;
      RECT  17.6 186.7 16.8 187.5 ;
      RECT  20.6 190.4 19.8 191.2 ;
      RECT  20.6 190.4 19.8 191.2 ;
      RECT  18.8 190.5 18.2 191.1 ;
      RECT  22.0 195.9 15.6 196.5 ;
      RECT  22.0 185.5 15.6 186.1 ;
      RECT  11.2 194.9 10.4 196.2 ;
      RECT  11.2 185.8 10.4 187.1 ;
      RECT  14.4 186.7 13.6 185.5 ;
      RECT  14.4 194.1 13.6 196.5 ;
      RECT  12.7 186.7 12.1 194.9 ;
      RECT  14.4 194.1 13.6 194.9 ;
      RECT  12.8 194.1 12.0 194.9 ;
      RECT  12.8 194.1 12.0 194.9 ;
      RECT  14.4 194.1 13.6 194.9 ;
      RECT  14.4 186.7 13.6 187.5 ;
      RECT  12.8 186.7 12.0 187.5 ;
      RECT  12.8 186.7 12.0 187.5 ;
      RECT  14.4 186.7 13.6 187.5 ;
      RECT  11.2 194.5 10.4 195.3 ;
      RECT  11.2 186.7 10.4 187.5 ;
      RECT  14.2 190.4 13.4 191.2 ;
      RECT  14.2 190.4 13.4 191.2 ;
      RECT  12.4 190.5 11.8 191.1 ;
      RECT  15.6 195.9 9.2 196.5 ;
      RECT  15.6 185.5 9.2 186.1 ;
      RECT  4.8 194.9 4.0 196.2 ;
      RECT  4.8 185.8 4.0 187.1 ;
      RECT  8.0 186.7 7.2 185.5 ;
      RECT  8.0 194.1 7.2 196.5 ;
      RECT  6.3 186.7 5.7 194.9 ;
      RECT  8.0 194.1 7.2 194.9 ;
      RECT  6.4 194.1 5.6 194.9 ;
      RECT  6.4 194.1 5.6 194.9 ;
      RECT  8.0 194.1 7.2 194.9 ;
      RECT  8.0 186.7 7.2 187.5 ;
      RECT  6.4 186.7 5.6 187.5 ;
      RECT  6.4 186.7 5.6 187.5 ;
      RECT  8.0 186.7 7.2 187.5 ;
      RECT  4.8 194.5 4.0 195.3 ;
      RECT  4.8 186.7 4.0 187.5 ;
      RECT  7.8 190.4 7.0 191.2 ;
      RECT  7.8 190.4 7.0 191.2 ;
      RECT  6.0 190.5 5.4 191.1 ;
      RECT  9.2 195.9 2.8 196.5 ;
      RECT  9.2 185.5 2.8 186.1 ;
      RECT  30.4 197.5 29.6 196.2 ;
      RECT  30.4 206.6 29.6 205.3 ;
      RECT  33.6 205.7 32.8 206.9 ;
      RECT  33.6 198.3 32.8 195.9 ;
      RECT  31.9 205.7 31.3 197.5 ;
      RECT  33.6 198.3 32.8 197.5 ;
      RECT  32.0 198.3 31.2 197.5 ;
      RECT  32.0 198.3 31.2 197.5 ;
      RECT  33.6 198.3 32.8 197.5 ;
      RECT  33.6 205.7 32.8 204.9 ;
      RECT  32.0 205.7 31.2 204.9 ;
      RECT  32.0 205.7 31.2 204.9 ;
      RECT  33.6 205.7 32.8 204.9 ;
      RECT  30.4 197.9 29.6 197.1 ;
      RECT  30.4 205.7 29.6 204.9 ;
      RECT  33.4 202.0 32.6 201.2 ;
      RECT  33.4 202.0 32.6 201.2 ;
      RECT  31.6 201.9 31.0 201.3 ;
      RECT  34.8 196.5 28.4 195.9 ;
      RECT  34.8 206.9 28.4 206.3 ;
      RECT  24.0 197.5 23.2 196.2 ;
      RECT  24.0 206.6 23.2 205.3 ;
      RECT  27.2 205.7 26.4 206.9 ;
      RECT  27.2 198.3 26.4 195.9 ;
      RECT  25.5 205.7 24.9 197.5 ;
      RECT  27.2 198.3 26.4 197.5 ;
      RECT  25.6 198.3 24.8 197.5 ;
      RECT  25.6 198.3 24.8 197.5 ;
      RECT  27.2 198.3 26.4 197.5 ;
      RECT  27.2 205.7 26.4 204.9 ;
      RECT  25.6 205.7 24.8 204.9 ;
      RECT  25.6 205.7 24.8 204.9 ;
      RECT  27.2 205.7 26.4 204.9 ;
      RECT  24.0 197.9 23.2 197.1 ;
      RECT  24.0 205.7 23.2 204.9 ;
      RECT  27.0 202.0 26.2 201.2 ;
      RECT  27.0 202.0 26.2 201.2 ;
      RECT  25.2 201.9 24.6 201.3 ;
      RECT  28.4 196.5 22.0 195.9 ;
      RECT  28.4 206.9 22.0 206.3 ;
      RECT  17.6 197.5 16.8 196.2 ;
      RECT  17.6 206.6 16.8 205.3 ;
      RECT  20.8 205.7 20.0 206.9 ;
      RECT  20.8 198.3 20.0 195.9 ;
      RECT  19.1 205.7 18.5 197.5 ;
      RECT  20.8 198.3 20.0 197.5 ;
      RECT  19.2 198.3 18.4 197.5 ;
      RECT  19.2 198.3 18.4 197.5 ;
      RECT  20.8 198.3 20.0 197.5 ;
      RECT  20.8 205.7 20.0 204.9 ;
      RECT  19.2 205.7 18.4 204.9 ;
      RECT  19.2 205.7 18.4 204.9 ;
      RECT  20.8 205.7 20.0 204.9 ;
      RECT  17.6 197.9 16.8 197.1 ;
      RECT  17.6 205.7 16.8 204.9 ;
      RECT  20.6 202.0 19.8 201.2 ;
      RECT  20.6 202.0 19.8 201.2 ;
      RECT  18.8 201.9 18.2 201.3 ;
      RECT  22.0 196.5 15.6 195.9 ;
      RECT  22.0 206.9 15.6 206.3 ;
      RECT  11.2 197.5 10.4 196.2 ;
      RECT  11.2 206.6 10.4 205.3 ;
      RECT  14.4 205.7 13.6 206.9 ;
      RECT  14.4 198.3 13.6 195.9 ;
      RECT  12.7 205.7 12.1 197.5 ;
      RECT  14.4 198.3 13.6 197.5 ;
      RECT  12.8 198.3 12.0 197.5 ;
      RECT  12.8 198.3 12.0 197.5 ;
      RECT  14.4 198.3 13.6 197.5 ;
      RECT  14.4 205.7 13.6 204.9 ;
      RECT  12.8 205.7 12.0 204.9 ;
      RECT  12.8 205.7 12.0 204.9 ;
      RECT  14.4 205.7 13.6 204.9 ;
      RECT  11.2 197.9 10.4 197.1 ;
      RECT  11.2 205.7 10.4 204.9 ;
      RECT  14.2 202.0 13.4 201.2 ;
      RECT  14.2 202.0 13.4 201.2 ;
      RECT  12.4 201.9 11.8 201.3 ;
      RECT  15.6 196.5 9.2 195.9 ;
      RECT  15.6 206.9 9.2 206.3 ;
      RECT  4.8 197.5 4.0 196.2 ;
      RECT  4.8 206.6 4.0 205.3 ;
      RECT  8.0 205.7 7.2 206.9 ;
      RECT  8.0 198.3 7.2 195.9 ;
      RECT  6.3 205.7 5.7 197.5 ;
      RECT  8.0 198.3 7.2 197.5 ;
      RECT  6.4 198.3 5.6 197.5 ;
      RECT  6.4 198.3 5.6 197.5 ;
      RECT  8.0 198.3 7.2 197.5 ;
      RECT  8.0 205.7 7.2 204.9 ;
      RECT  6.4 205.7 5.6 204.9 ;
      RECT  6.4 205.7 5.6 204.9 ;
      RECT  8.0 205.7 7.2 204.9 ;
      RECT  4.8 197.9 4.0 197.1 ;
      RECT  4.8 205.7 4.0 204.9 ;
      RECT  7.8 202.0 7.0 201.2 ;
      RECT  7.8 202.0 7.0 201.2 ;
      RECT  6.0 201.9 5.4 201.3 ;
      RECT  9.2 196.5 2.8 195.9 ;
      RECT  9.2 206.9 2.8 206.3 ;
      RECT  30.4 215.7 29.6 217.0 ;
      RECT  30.4 206.6 29.6 207.9 ;
      RECT  33.6 207.5 32.8 206.3 ;
      RECT  33.6 214.9 32.8 217.3 ;
      RECT  31.9 207.5 31.3 215.7 ;
      RECT  33.6 214.9 32.8 215.7 ;
      RECT  32.0 214.9 31.2 215.7 ;
      RECT  32.0 214.9 31.2 215.7 ;
      RECT  33.6 214.9 32.8 215.7 ;
      RECT  33.6 207.5 32.8 208.3 ;
      RECT  32.0 207.5 31.2 208.3 ;
      RECT  32.0 207.5 31.2 208.3 ;
      RECT  33.6 207.5 32.8 208.3 ;
      RECT  30.4 215.3 29.6 216.1 ;
      RECT  30.4 207.5 29.6 208.3 ;
      RECT  33.4 211.2 32.6 212.0 ;
      RECT  33.4 211.2 32.6 212.0 ;
      RECT  31.6 211.3 31.0 211.9 ;
      RECT  34.8 216.7 28.4 217.3 ;
      RECT  34.8 206.3 28.4 206.9 ;
      RECT  24.0 215.7 23.2 217.0 ;
      RECT  24.0 206.6 23.2 207.9 ;
      RECT  27.2 207.5 26.4 206.3 ;
      RECT  27.2 214.9 26.4 217.3 ;
      RECT  25.5 207.5 24.9 215.7 ;
      RECT  27.2 214.9 26.4 215.7 ;
      RECT  25.6 214.9 24.8 215.7 ;
      RECT  25.6 214.9 24.8 215.7 ;
      RECT  27.2 214.9 26.4 215.7 ;
      RECT  27.2 207.5 26.4 208.3 ;
      RECT  25.6 207.5 24.8 208.3 ;
      RECT  25.6 207.5 24.8 208.3 ;
      RECT  27.2 207.5 26.4 208.3 ;
      RECT  24.0 215.3 23.2 216.1 ;
      RECT  24.0 207.5 23.2 208.3 ;
      RECT  27.0 211.2 26.2 212.0 ;
      RECT  27.0 211.2 26.2 212.0 ;
      RECT  25.2 211.3 24.6 211.9 ;
      RECT  28.4 216.7 22.0 217.3 ;
      RECT  28.4 206.3 22.0 206.9 ;
      RECT  17.6 215.7 16.8 217.0 ;
      RECT  17.6 206.6 16.8 207.9 ;
      RECT  20.8 207.5 20.0 206.3 ;
      RECT  20.8 214.9 20.0 217.3 ;
      RECT  19.1 207.5 18.5 215.7 ;
      RECT  20.8 214.9 20.0 215.7 ;
      RECT  19.2 214.9 18.4 215.7 ;
      RECT  19.2 214.9 18.4 215.7 ;
      RECT  20.8 214.9 20.0 215.7 ;
      RECT  20.8 207.5 20.0 208.3 ;
      RECT  19.2 207.5 18.4 208.3 ;
      RECT  19.2 207.5 18.4 208.3 ;
      RECT  20.8 207.5 20.0 208.3 ;
      RECT  17.6 215.3 16.8 216.1 ;
      RECT  17.6 207.5 16.8 208.3 ;
      RECT  20.6 211.2 19.8 212.0 ;
      RECT  20.6 211.2 19.8 212.0 ;
      RECT  18.8 211.3 18.2 211.9 ;
      RECT  22.0 216.7 15.6 217.3 ;
      RECT  22.0 206.3 15.6 206.9 ;
      RECT  11.2 215.7 10.4 217.0 ;
      RECT  11.2 206.6 10.4 207.9 ;
      RECT  14.4 207.5 13.6 206.3 ;
      RECT  14.4 214.9 13.6 217.3 ;
      RECT  12.7 207.5 12.1 215.7 ;
      RECT  14.4 214.9 13.6 215.7 ;
      RECT  12.8 214.9 12.0 215.7 ;
      RECT  12.8 214.9 12.0 215.7 ;
      RECT  14.4 214.9 13.6 215.7 ;
      RECT  14.4 207.5 13.6 208.3 ;
      RECT  12.8 207.5 12.0 208.3 ;
      RECT  12.8 207.5 12.0 208.3 ;
      RECT  14.4 207.5 13.6 208.3 ;
      RECT  11.2 215.3 10.4 216.1 ;
      RECT  11.2 207.5 10.4 208.3 ;
      RECT  14.2 211.2 13.4 212.0 ;
      RECT  14.2 211.2 13.4 212.0 ;
      RECT  12.4 211.3 11.8 211.9 ;
      RECT  15.6 216.7 9.2 217.3 ;
      RECT  15.6 206.3 9.2 206.9 ;
      RECT  4.8 215.7 4.0 217.0 ;
      RECT  4.8 206.6 4.0 207.9 ;
      RECT  8.0 207.5 7.2 206.3 ;
      RECT  8.0 214.9 7.2 217.3 ;
      RECT  6.3 207.5 5.7 215.7 ;
      RECT  8.0 214.9 7.2 215.7 ;
      RECT  6.4 214.9 5.6 215.7 ;
      RECT  6.4 214.9 5.6 215.7 ;
      RECT  8.0 214.9 7.2 215.7 ;
      RECT  8.0 207.5 7.2 208.3 ;
      RECT  6.4 207.5 5.6 208.3 ;
      RECT  6.4 207.5 5.6 208.3 ;
      RECT  8.0 207.5 7.2 208.3 ;
      RECT  4.8 215.3 4.0 216.1 ;
      RECT  4.8 207.5 4.0 208.3 ;
      RECT  7.8 211.2 7.0 212.0 ;
      RECT  7.8 211.2 7.0 212.0 ;
      RECT  6.0 211.3 5.4 211.9 ;
      RECT  9.2 216.7 2.8 217.3 ;
      RECT  9.2 206.3 2.8 206.9 ;
      RECT  30.4 218.3 29.6 217.0 ;
      RECT  30.4 227.4 29.6 226.1 ;
      RECT  33.6 226.5 32.8 227.7 ;
      RECT  33.6 219.1 32.8 216.7 ;
      RECT  31.9 226.5 31.3 218.3 ;
      RECT  33.6 219.1 32.8 218.3 ;
      RECT  32.0 219.1 31.2 218.3 ;
      RECT  32.0 219.1 31.2 218.3 ;
      RECT  33.6 219.1 32.8 218.3 ;
      RECT  33.6 226.5 32.8 225.7 ;
      RECT  32.0 226.5 31.2 225.7 ;
      RECT  32.0 226.5 31.2 225.7 ;
      RECT  33.6 226.5 32.8 225.7 ;
      RECT  30.4 218.7 29.6 217.9 ;
      RECT  30.4 226.5 29.6 225.7 ;
      RECT  33.4 222.8 32.6 222.0 ;
      RECT  33.4 222.8 32.6 222.0 ;
      RECT  31.6 222.7 31.0 222.1 ;
      RECT  34.8 217.3 28.4 216.7 ;
      RECT  34.8 227.7 28.4 227.1 ;
      RECT  24.0 218.3 23.2 217.0 ;
      RECT  24.0 227.4 23.2 226.1 ;
      RECT  27.2 226.5 26.4 227.7 ;
      RECT  27.2 219.1 26.4 216.7 ;
      RECT  25.5 226.5 24.9 218.3 ;
      RECT  27.2 219.1 26.4 218.3 ;
      RECT  25.6 219.1 24.8 218.3 ;
      RECT  25.6 219.1 24.8 218.3 ;
      RECT  27.2 219.1 26.4 218.3 ;
      RECT  27.2 226.5 26.4 225.7 ;
      RECT  25.6 226.5 24.8 225.7 ;
      RECT  25.6 226.5 24.8 225.7 ;
      RECT  27.2 226.5 26.4 225.7 ;
      RECT  24.0 218.7 23.2 217.9 ;
      RECT  24.0 226.5 23.2 225.7 ;
      RECT  27.0 222.8 26.2 222.0 ;
      RECT  27.0 222.8 26.2 222.0 ;
      RECT  25.2 222.7 24.6 222.1 ;
      RECT  28.4 217.3 22.0 216.7 ;
      RECT  28.4 227.7 22.0 227.1 ;
      RECT  17.6 218.3 16.8 217.0 ;
      RECT  17.6 227.4 16.8 226.1 ;
      RECT  20.8 226.5 20.0 227.7 ;
      RECT  20.8 219.1 20.0 216.7 ;
      RECT  19.1 226.5 18.5 218.3 ;
      RECT  20.8 219.1 20.0 218.3 ;
      RECT  19.2 219.1 18.4 218.3 ;
      RECT  19.2 219.1 18.4 218.3 ;
      RECT  20.8 219.1 20.0 218.3 ;
      RECT  20.8 226.5 20.0 225.7 ;
      RECT  19.2 226.5 18.4 225.7 ;
      RECT  19.2 226.5 18.4 225.7 ;
      RECT  20.8 226.5 20.0 225.7 ;
      RECT  17.6 218.7 16.8 217.9 ;
      RECT  17.6 226.5 16.8 225.7 ;
      RECT  20.6 222.8 19.8 222.0 ;
      RECT  20.6 222.8 19.8 222.0 ;
      RECT  18.8 222.7 18.2 222.1 ;
      RECT  22.0 217.3 15.6 216.7 ;
      RECT  22.0 227.7 15.6 227.1 ;
      RECT  11.2 218.3 10.4 217.0 ;
      RECT  11.2 227.4 10.4 226.1 ;
      RECT  14.4 226.5 13.6 227.7 ;
      RECT  14.4 219.1 13.6 216.7 ;
      RECT  12.7 226.5 12.1 218.3 ;
      RECT  14.4 219.1 13.6 218.3 ;
      RECT  12.8 219.1 12.0 218.3 ;
      RECT  12.8 219.1 12.0 218.3 ;
      RECT  14.4 219.1 13.6 218.3 ;
      RECT  14.4 226.5 13.6 225.7 ;
      RECT  12.8 226.5 12.0 225.7 ;
      RECT  12.8 226.5 12.0 225.7 ;
      RECT  14.4 226.5 13.6 225.7 ;
      RECT  11.2 218.7 10.4 217.9 ;
      RECT  11.2 226.5 10.4 225.7 ;
      RECT  14.2 222.8 13.4 222.0 ;
      RECT  14.2 222.8 13.4 222.0 ;
      RECT  12.4 222.7 11.8 222.1 ;
      RECT  15.6 217.3 9.2 216.7 ;
      RECT  15.6 227.7 9.2 227.1 ;
      RECT  4.8 218.3 4.0 217.0 ;
      RECT  4.8 227.4 4.0 226.1 ;
      RECT  8.0 226.5 7.2 227.7 ;
      RECT  8.0 219.1 7.2 216.7 ;
      RECT  6.3 226.5 5.7 218.3 ;
      RECT  8.0 219.1 7.2 218.3 ;
      RECT  6.4 219.1 5.6 218.3 ;
      RECT  6.4 219.1 5.6 218.3 ;
      RECT  8.0 219.1 7.2 218.3 ;
      RECT  8.0 226.5 7.2 225.7 ;
      RECT  6.4 226.5 5.6 225.7 ;
      RECT  6.4 226.5 5.6 225.7 ;
      RECT  8.0 226.5 7.2 225.7 ;
      RECT  4.8 218.7 4.0 217.9 ;
      RECT  4.8 226.5 4.0 225.7 ;
      RECT  7.8 222.8 7.0 222.0 ;
      RECT  7.8 222.8 7.0 222.0 ;
      RECT  6.0 222.7 5.4 222.1 ;
      RECT  9.2 217.3 2.8 216.7 ;
      RECT  9.2 227.7 2.8 227.1 ;
      RECT  30.4 236.5 29.6 237.8 ;
      RECT  30.4 227.4 29.6 228.7 ;
      RECT  33.6 228.3 32.8 227.1 ;
      RECT  33.6 235.7 32.8 238.1 ;
      RECT  31.9 228.3 31.3 236.5 ;
      RECT  33.6 235.7 32.8 236.5 ;
      RECT  32.0 235.7 31.2 236.5 ;
      RECT  32.0 235.7 31.2 236.5 ;
      RECT  33.6 235.7 32.8 236.5 ;
      RECT  33.6 228.3 32.8 229.1 ;
      RECT  32.0 228.3 31.2 229.1 ;
      RECT  32.0 228.3 31.2 229.1 ;
      RECT  33.6 228.3 32.8 229.1 ;
      RECT  30.4 236.1 29.6 236.9 ;
      RECT  30.4 228.3 29.6 229.1 ;
      RECT  33.4 232.0 32.6 232.8 ;
      RECT  33.4 232.0 32.6 232.8 ;
      RECT  31.6 232.1 31.0 232.7 ;
      RECT  34.8 237.5 28.4 238.1 ;
      RECT  34.8 227.1 28.4 227.7 ;
      RECT  24.0 236.5 23.2 237.8 ;
      RECT  24.0 227.4 23.2 228.7 ;
      RECT  27.2 228.3 26.4 227.1 ;
      RECT  27.2 235.7 26.4 238.1 ;
      RECT  25.5 228.3 24.9 236.5 ;
      RECT  27.2 235.7 26.4 236.5 ;
      RECT  25.6 235.7 24.8 236.5 ;
      RECT  25.6 235.7 24.8 236.5 ;
      RECT  27.2 235.7 26.4 236.5 ;
      RECT  27.2 228.3 26.4 229.1 ;
      RECT  25.6 228.3 24.8 229.1 ;
      RECT  25.6 228.3 24.8 229.1 ;
      RECT  27.2 228.3 26.4 229.1 ;
      RECT  24.0 236.1 23.2 236.9 ;
      RECT  24.0 228.3 23.2 229.1 ;
      RECT  27.0 232.0 26.2 232.8 ;
      RECT  27.0 232.0 26.2 232.8 ;
      RECT  25.2 232.1 24.6 232.7 ;
      RECT  28.4 237.5 22.0 238.1 ;
      RECT  28.4 227.1 22.0 227.7 ;
      RECT  17.6 236.5 16.8 237.8 ;
      RECT  17.6 227.4 16.8 228.7 ;
      RECT  20.8 228.3 20.0 227.1 ;
      RECT  20.8 235.7 20.0 238.1 ;
      RECT  19.1 228.3 18.5 236.5 ;
      RECT  20.8 235.7 20.0 236.5 ;
      RECT  19.2 235.7 18.4 236.5 ;
      RECT  19.2 235.7 18.4 236.5 ;
      RECT  20.8 235.7 20.0 236.5 ;
      RECT  20.8 228.3 20.0 229.1 ;
      RECT  19.2 228.3 18.4 229.1 ;
      RECT  19.2 228.3 18.4 229.1 ;
      RECT  20.8 228.3 20.0 229.1 ;
      RECT  17.6 236.1 16.8 236.9 ;
      RECT  17.6 228.3 16.8 229.1 ;
      RECT  20.6 232.0 19.8 232.8 ;
      RECT  20.6 232.0 19.8 232.8 ;
      RECT  18.8 232.1 18.2 232.7 ;
      RECT  22.0 237.5 15.6 238.1 ;
      RECT  22.0 227.1 15.6 227.7 ;
      RECT  11.2 236.5 10.4 237.8 ;
      RECT  11.2 227.4 10.4 228.7 ;
      RECT  14.4 228.3 13.6 227.1 ;
      RECT  14.4 235.7 13.6 238.1 ;
      RECT  12.7 228.3 12.1 236.5 ;
      RECT  14.4 235.7 13.6 236.5 ;
      RECT  12.8 235.7 12.0 236.5 ;
      RECT  12.8 235.7 12.0 236.5 ;
      RECT  14.4 235.7 13.6 236.5 ;
      RECT  14.4 228.3 13.6 229.1 ;
      RECT  12.8 228.3 12.0 229.1 ;
      RECT  12.8 228.3 12.0 229.1 ;
      RECT  14.4 228.3 13.6 229.1 ;
      RECT  11.2 236.1 10.4 236.9 ;
      RECT  11.2 228.3 10.4 229.1 ;
      RECT  14.2 232.0 13.4 232.8 ;
      RECT  14.2 232.0 13.4 232.8 ;
      RECT  12.4 232.1 11.8 232.7 ;
      RECT  15.6 237.5 9.2 238.1 ;
      RECT  15.6 227.1 9.2 227.7 ;
      RECT  4.8 236.5 4.0 237.8 ;
      RECT  4.8 227.4 4.0 228.7 ;
      RECT  8.0 228.3 7.2 227.1 ;
      RECT  8.0 235.7 7.2 238.1 ;
      RECT  6.3 228.3 5.7 236.5 ;
      RECT  8.0 235.7 7.2 236.5 ;
      RECT  6.4 235.7 5.6 236.5 ;
      RECT  6.4 235.7 5.6 236.5 ;
      RECT  8.0 235.7 7.2 236.5 ;
      RECT  8.0 228.3 7.2 229.1 ;
      RECT  6.4 228.3 5.6 229.1 ;
      RECT  6.4 228.3 5.6 229.1 ;
      RECT  8.0 228.3 7.2 229.1 ;
      RECT  4.8 236.1 4.0 236.9 ;
      RECT  4.8 228.3 4.0 229.1 ;
      RECT  7.8 232.0 7.0 232.8 ;
      RECT  7.8 232.0 7.0 232.8 ;
      RECT  6.0 232.1 5.4 232.7 ;
      RECT  9.2 237.5 2.8 238.1 ;
      RECT  9.2 227.1 2.8 227.7 ;
      RECT  30.4 239.1 29.6 237.8 ;
      RECT  30.4 248.2 29.6 246.9 ;
      RECT  33.6 247.3 32.8 248.5 ;
      RECT  33.6 239.9 32.8 237.5 ;
      RECT  31.9 247.3 31.3 239.1 ;
      RECT  33.6 239.9 32.8 239.1 ;
      RECT  32.0 239.9 31.2 239.1 ;
      RECT  32.0 239.9 31.2 239.1 ;
      RECT  33.6 239.9 32.8 239.1 ;
      RECT  33.6 247.3 32.8 246.5 ;
      RECT  32.0 247.3 31.2 246.5 ;
      RECT  32.0 247.3 31.2 246.5 ;
      RECT  33.6 247.3 32.8 246.5 ;
      RECT  30.4 239.5 29.6 238.7 ;
      RECT  30.4 247.3 29.6 246.5 ;
      RECT  33.4 243.6 32.6 242.8 ;
      RECT  33.4 243.6 32.6 242.8 ;
      RECT  31.6 243.5 31.0 242.9 ;
      RECT  34.8 238.1 28.4 237.5 ;
      RECT  34.8 248.5 28.4 247.9 ;
      RECT  24.0 239.1 23.2 237.8 ;
      RECT  24.0 248.2 23.2 246.9 ;
      RECT  27.2 247.3 26.4 248.5 ;
      RECT  27.2 239.9 26.4 237.5 ;
      RECT  25.5 247.3 24.9 239.1 ;
      RECT  27.2 239.9 26.4 239.1 ;
      RECT  25.6 239.9 24.8 239.1 ;
      RECT  25.6 239.9 24.8 239.1 ;
      RECT  27.2 239.9 26.4 239.1 ;
      RECT  27.2 247.3 26.4 246.5 ;
      RECT  25.6 247.3 24.8 246.5 ;
      RECT  25.6 247.3 24.8 246.5 ;
      RECT  27.2 247.3 26.4 246.5 ;
      RECT  24.0 239.5 23.2 238.7 ;
      RECT  24.0 247.3 23.2 246.5 ;
      RECT  27.0 243.6 26.2 242.8 ;
      RECT  27.0 243.6 26.2 242.8 ;
      RECT  25.2 243.5 24.6 242.9 ;
      RECT  28.4 238.1 22.0 237.5 ;
      RECT  28.4 248.5 22.0 247.9 ;
      RECT  17.6 239.1 16.8 237.8 ;
      RECT  17.6 248.2 16.8 246.9 ;
      RECT  20.8 247.3 20.0 248.5 ;
      RECT  20.8 239.9 20.0 237.5 ;
      RECT  19.1 247.3 18.5 239.1 ;
      RECT  20.8 239.9 20.0 239.1 ;
      RECT  19.2 239.9 18.4 239.1 ;
      RECT  19.2 239.9 18.4 239.1 ;
      RECT  20.8 239.9 20.0 239.1 ;
      RECT  20.8 247.3 20.0 246.5 ;
      RECT  19.2 247.3 18.4 246.5 ;
      RECT  19.2 247.3 18.4 246.5 ;
      RECT  20.8 247.3 20.0 246.5 ;
      RECT  17.6 239.5 16.8 238.7 ;
      RECT  17.6 247.3 16.8 246.5 ;
      RECT  20.6 243.6 19.8 242.8 ;
      RECT  20.6 243.6 19.8 242.8 ;
      RECT  18.8 243.5 18.2 242.9 ;
      RECT  22.0 238.1 15.6 237.5 ;
      RECT  22.0 248.5 15.6 247.9 ;
      RECT  11.2 239.1 10.4 237.8 ;
      RECT  11.2 248.2 10.4 246.9 ;
      RECT  14.4 247.3 13.6 248.5 ;
      RECT  14.4 239.9 13.6 237.5 ;
      RECT  12.7 247.3 12.1 239.1 ;
      RECT  14.4 239.9 13.6 239.1 ;
      RECT  12.8 239.9 12.0 239.1 ;
      RECT  12.8 239.9 12.0 239.1 ;
      RECT  14.4 239.9 13.6 239.1 ;
      RECT  14.4 247.3 13.6 246.5 ;
      RECT  12.8 247.3 12.0 246.5 ;
      RECT  12.8 247.3 12.0 246.5 ;
      RECT  14.4 247.3 13.6 246.5 ;
      RECT  11.2 239.5 10.4 238.7 ;
      RECT  11.2 247.3 10.4 246.5 ;
      RECT  14.2 243.6 13.4 242.8 ;
      RECT  14.2 243.6 13.4 242.8 ;
      RECT  12.4 243.5 11.8 242.9 ;
      RECT  15.6 238.1 9.2 237.5 ;
      RECT  15.6 248.5 9.2 247.9 ;
      RECT  4.8 239.1 4.0 237.8 ;
      RECT  4.8 248.2 4.0 246.9 ;
      RECT  8.0 247.3 7.2 248.5 ;
      RECT  8.0 239.9 7.2 237.5 ;
      RECT  6.3 247.3 5.7 239.1 ;
      RECT  8.0 239.9 7.2 239.1 ;
      RECT  6.4 239.9 5.6 239.1 ;
      RECT  6.4 239.9 5.6 239.1 ;
      RECT  8.0 239.9 7.2 239.1 ;
      RECT  8.0 247.3 7.2 246.5 ;
      RECT  6.4 247.3 5.6 246.5 ;
      RECT  6.4 247.3 5.6 246.5 ;
      RECT  8.0 247.3 7.2 246.5 ;
      RECT  4.8 239.5 4.0 238.7 ;
      RECT  4.8 247.3 4.0 246.5 ;
      RECT  7.8 243.6 7.0 242.8 ;
      RECT  7.8 243.6 7.0 242.8 ;
      RECT  6.0 243.5 5.4 242.9 ;
      RECT  9.2 238.1 2.8 237.5 ;
      RECT  9.2 248.5 2.8 247.9 ;
      RECT  30.4 257.3 29.6 258.6 ;
      RECT  30.4 248.2 29.6 249.5 ;
      RECT  33.6 249.1 32.8 247.9 ;
      RECT  33.6 256.5 32.8 258.9 ;
      RECT  31.9 249.1 31.3 257.3 ;
      RECT  33.6 256.5 32.8 257.3 ;
      RECT  32.0 256.5 31.2 257.3 ;
      RECT  32.0 256.5 31.2 257.3 ;
      RECT  33.6 256.5 32.8 257.3 ;
      RECT  33.6 249.1 32.8 249.9 ;
      RECT  32.0 249.1 31.2 249.9 ;
      RECT  32.0 249.1 31.2 249.9 ;
      RECT  33.6 249.1 32.8 249.9 ;
      RECT  30.4 256.9 29.6 257.7 ;
      RECT  30.4 249.1 29.6 249.9 ;
      RECT  33.4 252.8 32.6 253.6 ;
      RECT  33.4 252.8 32.6 253.6 ;
      RECT  31.6 252.9 31.0 253.5 ;
      RECT  34.8 258.3 28.4 258.9 ;
      RECT  34.8 247.9 28.4 248.5 ;
      RECT  24.0 257.3 23.2 258.6 ;
      RECT  24.0 248.2 23.2 249.5 ;
      RECT  27.2 249.1 26.4 247.9 ;
      RECT  27.2 256.5 26.4 258.9 ;
      RECT  25.5 249.1 24.9 257.3 ;
      RECT  27.2 256.5 26.4 257.3 ;
      RECT  25.6 256.5 24.8 257.3 ;
      RECT  25.6 256.5 24.8 257.3 ;
      RECT  27.2 256.5 26.4 257.3 ;
      RECT  27.2 249.1 26.4 249.9 ;
      RECT  25.6 249.1 24.8 249.9 ;
      RECT  25.6 249.1 24.8 249.9 ;
      RECT  27.2 249.1 26.4 249.9 ;
      RECT  24.0 256.9 23.2 257.7 ;
      RECT  24.0 249.1 23.2 249.9 ;
      RECT  27.0 252.8 26.2 253.6 ;
      RECT  27.0 252.8 26.2 253.6 ;
      RECT  25.2 252.9 24.6 253.5 ;
      RECT  28.4 258.3 22.0 258.9 ;
      RECT  28.4 247.9 22.0 248.5 ;
      RECT  17.6 257.3 16.8 258.6 ;
      RECT  17.6 248.2 16.8 249.5 ;
      RECT  20.8 249.1 20.0 247.9 ;
      RECT  20.8 256.5 20.0 258.9 ;
      RECT  19.1 249.1 18.5 257.3 ;
      RECT  20.8 256.5 20.0 257.3 ;
      RECT  19.2 256.5 18.4 257.3 ;
      RECT  19.2 256.5 18.4 257.3 ;
      RECT  20.8 256.5 20.0 257.3 ;
      RECT  20.8 249.1 20.0 249.9 ;
      RECT  19.2 249.1 18.4 249.9 ;
      RECT  19.2 249.1 18.4 249.9 ;
      RECT  20.8 249.1 20.0 249.9 ;
      RECT  17.6 256.9 16.8 257.7 ;
      RECT  17.6 249.1 16.8 249.9 ;
      RECT  20.6 252.8 19.8 253.6 ;
      RECT  20.6 252.8 19.8 253.6 ;
      RECT  18.8 252.9 18.2 253.5 ;
      RECT  22.0 258.3 15.6 258.9 ;
      RECT  22.0 247.9 15.6 248.5 ;
      RECT  11.2 257.3 10.4 258.6 ;
      RECT  11.2 248.2 10.4 249.5 ;
      RECT  14.4 249.1 13.6 247.9 ;
      RECT  14.4 256.5 13.6 258.9 ;
      RECT  12.7 249.1 12.1 257.3 ;
      RECT  14.4 256.5 13.6 257.3 ;
      RECT  12.8 256.5 12.0 257.3 ;
      RECT  12.8 256.5 12.0 257.3 ;
      RECT  14.4 256.5 13.6 257.3 ;
      RECT  14.4 249.1 13.6 249.9 ;
      RECT  12.8 249.1 12.0 249.9 ;
      RECT  12.8 249.1 12.0 249.9 ;
      RECT  14.4 249.1 13.6 249.9 ;
      RECT  11.2 256.9 10.4 257.7 ;
      RECT  11.2 249.1 10.4 249.9 ;
      RECT  14.2 252.8 13.4 253.6 ;
      RECT  14.2 252.8 13.4 253.6 ;
      RECT  12.4 252.9 11.8 253.5 ;
      RECT  15.6 258.3 9.2 258.9 ;
      RECT  15.6 247.9 9.2 248.5 ;
      RECT  4.8 257.3 4.0 258.6 ;
      RECT  4.8 248.2 4.0 249.5 ;
      RECT  8.0 249.1 7.2 247.9 ;
      RECT  8.0 256.5 7.2 258.9 ;
      RECT  6.3 249.1 5.7 257.3 ;
      RECT  8.0 256.5 7.2 257.3 ;
      RECT  6.4 256.5 5.6 257.3 ;
      RECT  6.4 256.5 5.6 257.3 ;
      RECT  8.0 256.5 7.2 257.3 ;
      RECT  8.0 249.1 7.2 249.9 ;
      RECT  6.4 249.1 5.6 249.9 ;
      RECT  6.4 249.1 5.6 249.9 ;
      RECT  8.0 249.1 7.2 249.9 ;
      RECT  4.8 256.9 4.0 257.7 ;
      RECT  4.8 249.1 4.0 249.9 ;
      RECT  7.8 252.8 7.0 253.6 ;
      RECT  7.8 252.8 7.0 253.6 ;
      RECT  6.0 252.9 5.4 253.5 ;
      RECT  9.2 258.3 2.8 258.9 ;
      RECT  9.2 247.9 2.8 248.5 ;
      RECT  27.0 169.6 26.2 170.4 ;
      RECT  20.6 169.6 19.8 170.4 ;
      RECT  14.2 169.6 13.4 170.4 ;
      RECT  7.8 169.6 7.0 170.4 ;
      RECT  33.4 169.6 32.6 170.4 ;
      RECT  31.7 169.6 30.9 170.4 ;
      RECT  27.0 180.4 26.2 181.2 ;
      RECT  20.6 180.4 19.8 181.2 ;
      RECT  14.2 180.4 13.4 181.2 ;
      RECT  7.8 180.4 7.0 181.2 ;
      RECT  33.4 180.4 32.6 181.2 ;
      RECT  31.7 180.4 30.9 181.2 ;
      RECT  27.0 190.4 26.2 191.2 ;
      RECT  20.6 190.4 19.8 191.2 ;
      RECT  14.2 190.4 13.4 191.2 ;
      RECT  7.8 190.4 7.0 191.2 ;
      RECT  33.4 190.4 32.6 191.2 ;
      RECT  31.7 190.4 30.9 191.2 ;
      RECT  27.0 201.2 26.2 202.0 ;
      RECT  20.6 201.2 19.8 202.0 ;
      RECT  14.2 201.2 13.4 202.0 ;
      RECT  7.8 201.2 7.0 202.0 ;
      RECT  33.4 201.2 32.6 202.0 ;
      RECT  31.7 201.2 30.9 202.0 ;
      RECT  27.0 211.2 26.2 212.0 ;
      RECT  20.6 211.2 19.8 212.0 ;
      RECT  14.2 211.2 13.4 212.0 ;
      RECT  7.8 211.2 7.0 212.0 ;
      RECT  33.4 211.2 32.6 212.0 ;
      RECT  31.7 211.2 30.9 212.0 ;
      RECT  27.0 222.0 26.2 222.8 ;
      RECT  20.6 222.0 19.8 222.8 ;
      RECT  14.2 222.0 13.4 222.8 ;
      RECT  7.8 222.0 7.0 222.8 ;
      RECT  33.4 222.0 32.6 222.8 ;
      RECT  31.7 222.0 30.9 222.8 ;
      RECT  27.0 232.0 26.2 232.8 ;
      RECT  20.6 232.0 19.8 232.8 ;
      RECT  14.2 232.0 13.4 232.8 ;
      RECT  7.8 232.0 7.0 232.8 ;
      RECT  33.4 232.0 32.6 232.8 ;
      RECT  31.7 232.0 30.9 232.8 ;
      RECT  27.0 242.8 26.2 243.6 ;
      RECT  20.6 242.8 19.8 243.6 ;
      RECT  14.2 242.8 13.4 243.6 ;
      RECT  7.8 242.8 7.0 243.6 ;
      RECT  33.4 242.8 32.6 243.6 ;
      RECT  31.7 242.8 30.9 243.6 ;
      RECT  27.0 252.8 26.2 253.6 ;
      RECT  20.6 252.8 19.8 253.6 ;
      RECT  14.2 252.8 13.4 253.6 ;
      RECT  7.8 252.8 7.0 253.6 ;
      RECT  33.4 252.8 32.6 253.6 ;
      RECT  31.7 252.8 30.9 253.6 ;
      RECT  22.4 175.0 21.6 175.8 ;
      RECT  22.4 164.6 21.6 165.4 ;
      RECT  16.0 175.0 15.2 175.8 ;
      RECT  16.0 164.6 15.2 165.4 ;
      RECT  9.6 175.0 8.8 175.8 ;
      RECT  9.6 164.6 8.8 165.4 ;
      RECT  22.4 195.8 21.6 196.6 ;
      RECT  22.4 185.4 21.6 186.2 ;
      RECT  16.0 195.8 15.2 196.6 ;
      RECT  16.0 185.4 15.2 186.2 ;
      RECT  9.6 195.8 8.8 196.6 ;
      RECT  9.6 185.4 8.8 186.2 ;
      RECT  22.4 216.6 21.6 217.4 ;
      RECT  22.4 206.2 21.6 207.0 ;
      RECT  16.0 216.6 15.2 217.4 ;
      RECT  16.0 206.2 15.2 207.0 ;
      RECT  9.6 216.6 8.8 217.4 ;
      RECT  9.6 206.2 8.8 207.0 ;
      RECT  22.4 237.4 21.6 238.2 ;
      RECT  22.4 227.0 21.6 227.8 ;
      RECT  16.0 237.4 15.2 238.2 ;
      RECT  16.0 227.0 15.2 227.8 ;
      RECT  9.6 237.4 8.8 238.2 ;
      RECT  9.6 227.0 8.8 227.8 ;
      RECT  22.4 258.2 21.6 259.0 ;
      RECT  22.4 247.8 21.6 248.6 ;
      RECT  16.0 258.2 15.2 259.0 ;
      RECT  16.0 247.8 15.2 248.6 ;
      RECT  9.6 258.2 8.8 259.0 ;
      RECT  9.6 247.8 8.8 248.6 ;
      RECT  22.4 247.8 21.6 248.6 ;
      RECT  16.0 247.8 15.2 248.6 ;
      RECT  9.6 247.8 8.8 248.6 ;
      RECT  33.4 169.6 32.6 170.4 ;
      RECT  7.8 252.8 7.0 253.6 ;
      RECT  51.2 120.9 52.0 122.5 ;
      RECT  51.2 104.3 52.0 101.9 ;
      RECT  54.4 104.3 55.2 101.9 ;
      RECT  56.0 103.5 56.8 102.2 ;
      RECT  56.0 122.2 56.8 120.9 ;
      RECT  51.2 104.3 52.0 103.5 ;
      RECT  52.8 104.3 53.6 103.5 ;
      RECT  52.8 104.3 53.6 103.5 ;
      RECT  51.2 104.3 52.0 103.5 ;
      RECT  52.8 104.3 53.6 103.5 ;
      RECT  54.4 104.3 55.2 103.5 ;
      RECT  54.4 104.3 55.2 103.5 ;
      RECT  52.8 104.3 53.6 103.5 ;
      RECT  51.2 120.9 52.0 120.1 ;
      RECT  52.8 120.9 53.6 120.1 ;
      RECT  52.8 120.9 53.6 120.1 ;
      RECT  51.2 120.9 52.0 120.1 ;
      RECT  52.8 120.9 53.6 120.1 ;
      RECT  54.4 120.9 55.2 120.1 ;
      RECT  54.4 120.9 55.2 120.1 ;
      RECT  52.8 120.9 53.6 120.1 ;
      RECT  56.0 103.9 56.8 103.1 ;
      RECT  56.0 121.3 56.8 120.5 ;
      RECT  53.6 119.2 54.4 118.4 ;
      RECT  51.6 117.8 52.4 117.0 ;
      RECT  52.8 104.3 53.6 103.5 ;
      RECT  54.4 120.9 55.2 120.1 ;
      RECT  55.8 117.8 56.6 117.0 ;
      RECT  51.6 117.8 52.4 117.0 ;
      RECT  53.6 119.2 54.4 118.4 ;
      RECT  55.8 117.8 56.6 117.0 ;
      RECT  50.0 102.5 59.6 101.9 ;
      RECT  50.0 122.5 59.6 121.9 ;
      RECT  63.1 112.7 67.8 112.1 ;
      RECT  64.0 103.5 64.8 102.2 ;
      RECT  64.0 122.2 64.8 120.9 ;
      RECT  60.8 121.3 61.6 122.5 ;
      RECT  60.8 104.3 61.6 101.9 ;
      RECT  62.5 121.3 63.1 103.5 ;
      RECT  60.8 104.3 61.6 103.5 ;
      RECT  62.4 104.3 63.2 103.5 ;
      RECT  62.4 104.3 63.2 103.5 ;
      RECT  60.8 104.3 61.6 103.5 ;
      RECT  60.8 121.3 61.6 120.5 ;
      RECT  62.4 121.3 63.2 120.5 ;
      RECT  62.4 121.3 63.2 120.5 ;
      RECT  60.8 121.3 61.6 120.5 ;
      RECT  64.0 103.9 64.8 103.1 ;
      RECT  64.0 121.3 64.8 120.5 ;
      RECT  61.0 112.8 61.8 112.0 ;
      RECT  61.0 112.8 61.8 112.0 ;
      RECT  62.8 112.7 63.4 112.1 ;
      RECT  59.6 102.5 66.0 101.9 ;
      RECT  59.6 122.5 66.0 121.9 ;
      RECT  70.4 103.5 71.2 102.2 ;
      RECT  70.4 122.2 71.2 120.9 ;
      RECT  67.2 121.3 68.0 122.5 ;
      RECT  67.2 104.3 68.0 101.9 ;
      RECT  68.9 121.3 69.5 103.5 ;
      RECT  67.2 104.3 68.0 103.5 ;
      RECT  68.8 104.3 69.6 103.5 ;
      RECT  68.8 104.3 69.6 103.5 ;
      RECT  67.2 104.3 68.0 103.5 ;
      RECT  67.2 121.3 68.0 120.5 ;
      RECT  68.8 121.3 69.6 120.5 ;
      RECT  68.8 121.3 69.6 120.5 ;
      RECT  67.2 121.3 68.0 120.5 ;
      RECT  70.4 103.9 71.2 103.1 ;
      RECT  70.4 121.3 71.2 120.5 ;
      RECT  67.4 112.8 68.2 112.0 ;
      RECT  67.4 112.8 68.2 112.0 ;
      RECT  69.2 112.7 69.8 112.1 ;
      RECT  66.0 102.5 72.4 101.9 ;
      RECT  66.0 122.5 72.4 121.9 ;
      RECT  61.0 112.8 61.8 112.0 ;
      RECT  69.2 112.7 69.8 112.1 ;
      RECT  59.6 102.5 60.2 101.9 ;
      RECT  59.6 122.5 60.2 121.9 ;
      RECT  5.5 44.6 6.3 45.4 ;
      RECT  44.3 44.6 45.1 45.4 ;
      RECT  40.1 72.0 40.9 72.8 ;
      RECT  53.1 131.6 53.9 132.4 ;
      RECT  38.7 131.6 39.5 132.4 ;
      RECT  42.9 87.5 43.7 88.3 ;
      RECT  37.3 86.2 38.1 87.0 ;
      RECT  40.1 84.9 40.9 85.7 ;
      RECT  38.7 156.1 39.5 156.9 ;
      RECT  40.1 157.4 40.9 158.2 ;
      RECT  45.7 158.7 46.5 159.5 ;
      RECT  5.2 101.5 6.0 102.3 ;
      RECT  38.7 101.5 39.5 102.3 ;
      RECT  41.5 117.0 42.3 117.8 ;
      RECT  38.7 118.4 39.5 119.2 ;
      RECT  56.2 112.0 57.0 112.8 ;
      RECT  51.4 11.6 52.2 12.4 ;
      RECT  73.9 10.8 74.7 11.6 ;
      RECT  44.3 32.0 45.1 32.8 ;
      RECT  58.0 37.0 58.8 37.8 ;
      RECT  81.9 32.6 82.7 33.4 ;
      RECT  44.3 46.6 45.1 47.4 ;
      RECT  47.1 45.2 47.9 46.0 ;
      RECT  75.5 51.0 76.3 51.8 ;
      RECT  84.8 21.8 85.6 22.6 ;
      RECT  84.8 1.8 85.6 2.6 ;
      RECT  84.8 21.8 85.6 22.6 ;
      RECT  84.8 41.8 85.6 42.6 ;
      RECT  84.8 61.8 85.6 62.6 ;
      RECT  84.8 41.8 85.6 42.6 ;
      RECT  84.8 61.8 85.6 62.6 ;
      RECT  84.8 81.8 85.6 82.6 ;
      RECT  84.8 101.8 85.6 102.6 ;
      RECT  84.8 81.8 85.6 82.6 ;
      RECT  84.8 101.8 85.6 102.6 ;
      RECT  84.8 121.8 85.6 122.6 ;
      RECT  84.8 141.8 85.6 142.6 ;
      RECT  84.8 121.8 85.6 122.6 ;
      RECT  84.8 141.8 85.6 142.6 ;
      RECT  84.8 161.8 85.6 162.6 ;
      RECT  63.9 152.3 86.6 152.9 ;
      RECT  63.9 90.9 86.6 91.5 ;
      RECT  69.5 112.1 86.6 112.7 ;
      RECT  72.7 72.9 86.6 73.5 ;
      RECT  74.3 10.9 86.6 11.5 ;
      RECT  78.8 300.8 79.6 301.0 ;
      RECT  66.0 294.0 66.8 298.8 ;
      RECT  74.8 307.0 75.4 307.6 ;
      RECT  72.6 306.4 76.2 307.0 ;
      RECT  66.0 302.6 71.6 302.8 ;
      RECT  66.8 299.6 77.8 300.2 ;
      RECT  83.6 303.0 84.4 311.6 ;
      RECT  74.8 296.0 75.4 296.6 ;
      RECT  70.4 294.0 71.2 295.4 ;
      RECT  72.6 306.2 73.4 306.4 ;
      RECT  78.8 306.8 79.6 307.6 ;
      RECT  75.2 303.6 75.8 304.8 ;
      RECT  69.2 307.6 71.2 308.2 ;
      RECT  76.4 293.4 77.2 296.0 ;
      RECT  72.6 296.6 75.4 297.2 ;
      RECT  69.2 295.4 71.2 296.0 ;
      RECT  83.6 299.0 84.4 302.4 ;
      RECT  79.0 307.6 80.2 311.6 ;
      RECT  67.6 303.8 68.4 312.2 ;
      RECT  69.2 304.2 74.6 304.8 ;
      RECT  77.2 300.2 77.8 303.4 ;
      RECT  64.8 312.2 86.6 313.4 ;
      RECT  80.2 302.4 84.4 303.0 ;
      RECT  82.0 303.6 82.8 312.2 ;
      RECT  85.2 293.4 86.0 294.8 ;
      RECT  79.0 304.0 79.6 305.0 ;
      RECT  77.2 303.4 79.6 304.0 ;
      RECT  66.0 303.2 66.8 311.6 ;
      RECT  78.8 295.4 80.2 296.0 ;
      RECT  75.2 304.8 77.4 305.4 ;
      RECT  70.4 308.2 71.2 311.6 ;
      RECT  68.2 301.4 73.2 302.0 ;
      RECT  85.2 310.6 86.0 312.2 ;
      RECT  78.8 301.0 82.6 301.6 ;
      RECT  78.8 296.0 79.6 296.8 ;
      RECT  64.8 292.2 86.6 293.4 ;
      RECT  72.4 302.0 73.2 302.2 ;
      RECT  69.8 300.2 70.6 300.4 ;
      RECT  75.4 306.2 76.2 306.4 ;
      RECT  83.6 294.0 84.4 298.4 ;
      RECT  66.8 299.4 68.4 299.6 ;
      RECT  69.2 306.8 70.0 307.6 ;
      RECT  74.8 294.0 75.6 296.0 ;
      RECT  68.2 301.2 69.0 301.4 ;
      RECT  69.2 304.8 70.0 305.0 ;
      RECT  80.6 298.2 81.4 298.4 ;
      RECT  70.8 296.6 71.6 297.4 ;
      RECT  82.0 293.4 82.8 297.8 ;
      RECT  76.6 304.6 77.4 304.8 ;
      RECT  73.0 293.4 74.0 296.0 ;
      RECT  71.0 297.4 71.6 299.6 ;
      RECT  76.4 307.6 77.2 312.2 ;
      RECT  73.2 307.6 74.0 312.2 ;
      RECT  76.6 299.4 77.4 299.6 ;
      RECT  71.0 303.2 75.8 303.6 ;
      RECT  66.0 302.8 71.8 303.0 ;
      RECT  74.8 307.6 75.6 311.6 ;
      RECT  81.8 301.6 82.6 301.8 ;
      RECT  66.0 303.0 75.8 303.2 ;
      RECT  73.8 304.8 74.6 305.0 ;
      RECT  79.0 294.0 80.2 295.4 ;
      RECT  72.6 297.2 73.4 297.4 ;
      RECT  79.0 305.0 80.4 305.8 ;
      RECT  80.2 302.2 81.0 302.4 ;
      RECT  69.2 296.0 70.0 296.8 ;
      RECT  67.6 293.4 68.4 298.0 ;
      RECT  80.6 298.4 84.4 299.0 ;
      RECT  78.8 324.8 79.6 324.6 ;
      RECT  66.0 331.6 66.8 326.8 ;
      RECT  74.8 318.6 75.4 318.0 ;
      RECT  72.6 319.2 76.2 318.6 ;
      RECT  66.0 323.0 71.6 322.8 ;
      RECT  66.8 326.0 77.8 325.4 ;
      RECT  83.6 322.6 84.4 314.0 ;
      RECT  74.8 329.6 75.4 329.0 ;
      RECT  70.4 331.6 71.2 330.2 ;
      RECT  72.6 319.4 73.4 319.2 ;
      RECT  78.8 318.8 79.6 318.0 ;
      RECT  75.2 322.0 75.8 320.8 ;
      RECT  69.2 318.0 71.2 317.4 ;
      RECT  76.4 332.2 77.2 329.6 ;
      RECT  72.6 329.0 75.4 328.4 ;
      RECT  69.2 330.2 71.2 329.6 ;
      RECT  83.6 326.6 84.4 323.2 ;
      RECT  79.0 318.0 80.2 314.0 ;
      RECT  67.6 321.8 68.4 313.4 ;
      RECT  69.2 321.4 74.6 320.8 ;
      RECT  77.2 325.4 77.8 322.2 ;
      RECT  64.8 313.4 86.6 312.2 ;
      RECT  80.2 323.2 84.4 322.6 ;
      RECT  82.0 322.0 82.8 313.4 ;
      RECT  85.2 332.2 86.0 330.8 ;
      RECT  79.0 321.6 79.6 320.6 ;
      RECT  77.2 322.2 79.6 321.6 ;
      RECT  66.0 322.4 66.8 314.0 ;
      RECT  78.8 330.2 80.2 329.6 ;
      RECT  75.2 320.8 77.4 320.2 ;
      RECT  70.4 317.4 71.2 314.0 ;
      RECT  68.2 324.2 73.2 323.6 ;
      RECT  85.2 315.0 86.0 313.4 ;
      RECT  78.8 324.6 82.6 324.0 ;
      RECT  78.8 329.6 79.6 328.8 ;
      RECT  64.8 333.4 86.6 332.2 ;
      RECT  72.4 323.6 73.2 323.4 ;
      RECT  69.8 325.4 70.6 325.2 ;
      RECT  75.4 319.4 76.2 319.2 ;
      RECT  83.6 331.6 84.4 327.2 ;
      RECT  66.8 326.2 68.4 326.0 ;
      RECT  69.2 318.8 70.0 318.0 ;
      RECT  74.8 331.6 75.6 329.6 ;
      RECT  68.2 324.4 69.0 324.2 ;
      RECT  69.2 320.8 70.0 320.6 ;
      RECT  80.6 327.4 81.4 327.2 ;
      RECT  70.8 329.0 71.6 328.2 ;
      RECT  82.0 332.2 82.8 327.8 ;
      RECT  76.6 321.0 77.4 320.8 ;
      RECT  73.0 332.2 74.0 329.6 ;
      RECT  71.0 328.2 71.6 326.0 ;
      RECT  76.4 318.0 77.2 313.4 ;
      RECT  73.2 318.0 74.0 313.4 ;
      RECT  76.6 326.2 77.4 326.0 ;
      RECT  71.0 322.4 75.8 322.0 ;
      RECT  66.0 322.8 71.8 322.6 ;
      RECT  74.8 318.0 75.6 314.0 ;
      RECT  81.8 324.0 82.6 323.8 ;
      RECT  66.0 322.6 75.8 322.4 ;
      RECT  73.8 320.8 74.6 320.6 ;
      RECT  79.0 331.6 80.2 330.2 ;
      RECT  72.6 328.4 73.4 328.2 ;
      RECT  79.0 320.6 80.4 319.8 ;
      RECT  80.2 323.4 81.0 323.2 ;
      RECT  69.2 329.6 70.0 328.8 ;
      RECT  67.6 332.2 68.4 327.6 ;
      RECT  80.6 327.2 84.4 326.6 ;
      RECT  78.8 340.8 79.6 341.0 ;
      RECT  66.0 334.0 66.8 338.8 ;
      RECT  74.8 347.0 75.4 347.6 ;
      RECT  72.6 346.4 76.2 347.0 ;
      RECT  66.0 342.6 71.6 342.8 ;
      RECT  66.8 339.6 77.8 340.2 ;
      RECT  83.6 343.0 84.4 351.6 ;
      RECT  74.8 336.0 75.4 336.6 ;
      RECT  70.4 334.0 71.2 335.4 ;
      RECT  72.6 346.2 73.4 346.4 ;
      RECT  78.8 346.8 79.6 347.6 ;
      RECT  75.2 343.6 75.8 344.8 ;
      RECT  69.2 347.6 71.2 348.2 ;
      RECT  76.4 333.4 77.2 336.0 ;
      RECT  72.6 336.6 75.4 337.2 ;
      RECT  69.2 335.4 71.2 336.0 ;
      RECT  83.6 339.0 84.4 342.4 ;
      RECT  79.0 347.6 80.2 351.6 ;
      RECT  67.6 343.8 68.4 352.2 ;
      RECT  69.2 344.2 74.6 344.8 ;
      RECT  77.2 340.2 77.8 343.4 ;
      RECT  64.8 352.2 86.6 353.4 ;
      RECT  80.2 342.4 84.4 343.0 ;
      RECT  82.0 343.6 82.8 352.2 ;
      RECT  85.2 333.4 86.0 334.8 ;
      RECT  79.0 344.0 79.6 345.0 ;
      RECT  77.2 343.4 79.6 344.0 ;
      RECT  66.0 343.2 66.8 351.6 ;
      RECT  78.8 335.4 80.2 336.0 ;
      RECT  75.2 344.8 77.4 345.4 ;
      RECT  70.4 348.2 71.2 351.6 ;
      RECT  68.2 341.4 73.2 342.0 ;
      RECT  85.2 350.6 86.0 352.2 ;
      RECT  78.8 341.0 82.6 341.6 ;
      RECT  78.8 336.0 79.6 336.8 ;
      RECT  64.8 332.2 86.6 333.4 ;
      RECT  72.4 342.0 73.2 342.2 ;
      RECT  69.8 340.2 70.6 340.4 ;
      RECT  75.4 346.2 76.2 346.4 ;
      RECT  83.6 334.0 84.4 338.4 ;
      RECT  66.8 339.4 68.4 339.6 ;
      RECT  69.2 346.8 70.0 347.6 ;
      RECT  74.8 334.0 75.6 336.0 ;
      RECT  68.2 341.2 69.0 341.4 ;
      RECT  69.2 344.8 70.0 345.0 ;
      RECT  80.6 338.2 81.4 338.4 ;
      RECT  70.8 336.6 71.6 337.4 ;
      RECT  82.0 333.4 82.8 337.8 ;
      RECT  76.6 344.6 77.4 344.8 ;
      RECT  73.0 333.4 74.0 336.0 ;
      RECT  71.0 337.4 71.6 339.6 ;
      RECT  76.4 347.6 77.2 352.2 ;
      RECT  73.2 347.6 74.0 352.2 ;
      RECT  76.6 339.4 77.4 339.6 ;
      RECT  71.0 343.2 75.8 343.6 ;
      RECT  66.0 342.8 71.8 343.0 ;
      RECT  74.8 347.6 75.6 351.6 ;
      RECT  81.8 341.6 82.6 341.8 ;
      RECT  66.0 343.0 75.8 343.2 ;
      RECT  73.8 344.8 74.6 345.0 ;
      RECT  79.0 334.0 80.2 335.4 ;
      RECT  72.6 337.2 73.4 337.4 ;
      RECT  79.0 345.0 80.4 345.8 ;
      RECT  80.2 342.2 81.0 342.4 ;
      RECT  69.2 336.0 70.0 336.8 ;
      RECT  67.6 333.4 68.4 338.0 ;
      RECT  80.6 338.4 84.4 339.0 ;
      RECT  78.8 364.8 79.6 364.6 ;
      RECT  66.0 371.6 66.8 366.8 ;
      RECT  74.8 358.6 75.4 358.0 ;
      RECT  72.6 359.2 76.2 358.6 ;
      RECT  66.0 363.0 71.6 362.8 ;
      RECT  66.8 366.0 77.8 365.4 ;
      RECT  83.6 362.6 84.4 354.0 ;
      RECT  74.8 369.6 75.4 369.0 ;
      RECT  70.4 371.6 71.2 370.2 ;
      RECT  72.6 359.4 73.4 359.2 ;
      RECT  78.8 358.8 79.6 358.0 ;
      RECT  75.2 362.0 75.8 360.8 ;
      RECT  69.2 358.0 71.2 357.4 ;
      RECT  76.4 372.2 77.2 369.6 ;
      RECT  72.6 369.0 75.4 368.4 ;
      RECT  69.2 370.2 71.2 369.6 ;
      RECT  83.6 366.6 84.4 363.2 ;
      RECT  79.0 358.0 80.2 354.0 ;
      RECT  67.6 361.8 68.4 353.4 ;
      RECT  69.2 361.4 74.6 360.8 ;
      RECT  77.2 365.4 77.8 362.2 ;
      RECT  64.8 353.4 86.6 352.2 ;
      RECT  80.2 363.2 84.4 362.6 ;
      RECT  82.0 362.0 82.8 353.4 ;
      RECT  85.2 372.2 86.0 370.8 ;
      RECT  79.0 361.6 79.6 360.6 ;
      RECT  77.2 362.2 79.6 361.6 ;
      RECT  66.0 362.4 66.8 354.0 ;
      RECT  78.8 370.2 80.2 369.6 ;
      RECT  75.2 360.8 77.4 360.2 ;
      RECT  70.4 357.4 71.2 354.0 ;
      RECT  68.2 364.2 73.2 363.6 ;
      RECT  85.2 355.0 86.0 353.4 ;
      RECT  78.8 364.6 82.6 364.0 ;
      RECT  78.8 369.6 79.6 368.8 ;
      RECT  64.8 373.4 86.6 372.2 ;
      RECT  72.4 363.6 73.2 363.4 ;
      RECT  69.8 365.4 70.6 365.2 ;
      RECT  75.4 359.4 76.2 359.2 ;
      RECT  83.6 371.6 84.4 367.2 ;
      RECT  66.8 366.2 68.4 366.0 ;
      RECT  69.2 358.8 70.0 358.0 ;
      RECT  74.8 371.6 75.6 369.6 ;
      RECT  68.2 364.4 69.0 364.2 ;
      RECT  69.2 360.8 70.0 360.6 ;
      RECT  80.6 367.4 81.4 367.2 ;
      RECT  70.8 369.0 71.6 368.2 ;
      RECT  82.0 372.2 82.8 367.8 ;
      RECT  76.6 361.0 77.4 360.8 ;
      RECT  73.0 372.2 74.0 369.6 ;
      RECT  71.0 368.2 71.6 366.0 ;
      RECT  76.4 358.0 77.2 353.4 ;
      RECT  73.2 358.0 74.0 353.4 ;
      RECT  76.6 366.2 77.4 366.0 ;
      RECT  71.0 362.4 75.8 362.0 ;
      RECT  66.0 362.8 71.8 362.6 ;
      RECT  74.8 358.0 75.6 354.0 ;
      RECT  81.8 364.0 82.6 363.8 ;
      RECT  66.0 362.6 75.8 362.4 ;
      RECT  73.8 360.8 74.6 360.6 ;
      RECT  79.0 371.6 80.2 370.2 ;
      RECT  72.6 368.4 73.4 368.2 ;
      RECT  79.0 360.6 80.4 359.8 ;
      RECT  80.2 363.4 81.0 363.2 ;
      RECT  69.2 369.6 70.0 368.8 ;
      RECT  67.6 372.2 68.4 367.6 ;
      RECT  80.6 367.2 84.4 366.6 ;
      RECT  75.3 312.4 76.1 313.2 ;
      RECT  75.3 292.4 76.1 293.2 ;
      RECT  75.3 312.4 76.1 313.2 ;
      RECT  75.3 332.4 76.1 333.2 ;
      RECT  75.3 352.4 76.1 353.2 ;
      RECT  75.3 332.4 76.1 333.2 ;
      RECT  75.3 352.4 76.1 353.2 ;
      RECT  75.3 372.4 76.1 373.2 ;
      RECT  199.8 56.0 200.6 56.2 ;
      RECT  187.0 49.2 187.8 54.0 ;
      RECT  195.8 62.2 196.4 62.8 ;
      RECT  193.6 61.6 197.2 62.2 ;
      RECT  187.0 57.8 192.6 58.0 ;
      RECT  187.8 54.8 198.8 55.4 ;
      RECT  204.6 58.2 205.4 66.8 ;
      RECT  195.8 51.2 196.4 51.8 ;
      RECT  191.4 49.2 192.2 50.6 ;
      RECT  193.6 61.4 194.4 61.6 ;
      RECT  199.8 62.0 200.6 62.8 ;
      RECT  196.2 58.8 196.8 60.0 ;
      RECT  190.2 62.8 192.2 63.4 ;
      RECT  197.4 48.6 198.2 51.2 ;
      RECT  193.6 51.8 196.4 52.4 ;
      RECT  190.2 50.6 192.2 51.2 ;
      RECT  204.6 54.2 205.4 57.6 ;
      RECT  200.0 62.8 201.2 66.8 ;
      RECT  188.6 59.0 189.4 67.4 ;
      RECT  190.2 59.4 195.6 60.0 ;
      RECT  198.2 55.4 198.8 58.6 ;
      RECT  185.8 67.4 207.6 68.6 ;
      RECT  201.2 57.6 205.4 58.2 ;
      RECT  203.0 58.8 203.8 67.4 ;
      RECT  206.2 48.6 207.0 50.0 ;
      RECT  200.0 59.2 200.6 60.2 ;
      RECT  198.2 58.6 200.6 59.2 ;
      RECT  187.0 58.4 187.8 66.8 ;
      RECT  199.8 50.6 201.2 51.2 ;
      RECT  196.2 60.0 198.4 60.6 ;
      RECT  191.4 63.4 192.2 66.8 ;
      RECT  189.2 56.6 194.2 57.2 ;
      RECT  206.2 65.8 207.0 67.4 ;
      RECT  199.8 56.2 203.6 56.8 ;
      RECT  199.8 51.2 200.6 52.0 ;
      RECT  185.8 47.4 207.6 48.6 ;
      RECT  193.4 57.2 194.2 57.4 ;
      RECT  190.8 55.4 191.6 55.6 ;
      RECT  196.4 61.4 197.2 61.6 ;
      RECT  204.6 49.2 205.4 53.6 ;
      RECT  187.8 54.6 189.4 54.8 ;
      RECT  190.2 62.0 191.0 62.8 ;
      RECT  195.8 49.2 196.6 51.2 ;
      RECT  189.2 56.4 190.0 56.6 ;
      RECT  190.2 60.0 191.0 60.2 ;
      RECT  201.6 53.4 202.4 53.6 ;
      RECT  191.8 51.8 192.6 52.6 ;
      RECT  203.0 48.6 203.8 53.0 ;
      RECT  197.6 59.8 198.4 60.0 ;
      RECT  194.0 48.6 195.0 51.2 ;
      RECT  192.0 52.6 192.6 54.8 ;
      RECT  197.4 62.8 198.2 67.4 ;
      RECT  194.2 62.8 195.0 67.4 ;
      RECT  197.6 54.6 198.4 54.8 ;
      RECT  192.0 58.4 196.8 58.8 ;
      RECT  187.0 58.0 192.8 58.2 ;
      RECT  195.8 62.8 196.6 66.8 ;
      RECT  202.8 56.8 203.6 57.0 ;
      RECT  187.0 58.2 196.8 58.4 ;
      RECT  194.8 60.0 195.6 60.2 ;
      RECT  200.0 49.2 201.2 50.6 ;
      RECT  193.6 52.4 194.4 52.6 ;
      RECT  200.0 60.2 201.4 61.0 ;
      RECT  201.2 57.4 202.0 57.6 ;
      RECT  190.2 51.2 191.0 52.0 ;
      RECT  188.6 48.6 189.4 53.2 ;
      RECT  201.6 53.6 205.4 54.2 ;
      RECT  221.6 56.0 222.4 56.2 ;
      RECT  208.8 49.2 209.6 54.0 ;
      RECT  217.6 62.2 218.2 62.8 ;
      RECT  215.4 61.6 219.0 62.2 ;
      RECT  208.8 57.8 214.4 58.0 ;
      RECT  209.6 54.8 220.6 55.4 ;
      RECT  226.4 58.2 227.2 66.8 ;
      RECT  217.6 51.2 218.2 51.8 ;
      RECT  213.2 49.2 214.0 50.6 ;
      RECT  215.4 61.4 216.2 61.6 ;
      RECT  221.6 62.0 222.4 62.8 ;
      RECT  218.0 58.8 218.6 60.0 ;
      RECT  212.0 62.8 214.0 63.4 ;
      RECT  219.2 48.6 220.0 51.2 ;
      RECT  215.4 51.8 218.2 52.4 ;
      RECT  212.0 50.6 214.0 51.2 ;
      RECT  226.4 54.2 227.2 57.6 ;
      RECT  221.8 62.8 223.0 66.8 ;
      RECT  210.4 59.0 211.2 67.4 ;
      RECT  212.0 59.4 217.4 60.0 ;
      RECT  220.0 55.4 220.6 58.6 ;
      RECT  207.6 67.4 229.4 68.6 ;
      RECT  223.0 57.6 227.2 58.2 ;
      RECT  224.8 58.8 225.6 67.4 ;
      RECT  228.0 48.6 228.8 50.0 ;
      RECT  221.8 59.2 222.4 60.2 ;
      RECT  220.0 58.6 222.4 59.2 ;
      RECT  208.8 58.4 209.6 66.8 ;
      RECT  221.6 50.6 223.0 51.2 ;
      RECT  218.0 60.0 220.2 60.6 ;
      RECT  213.2 63.4 214.0 66.8 ;
      RECT  211.0 56.6 216.0 57.2 ;
      RECT  228.0 65.8 228.8 67.4 ;
      RECT  221.6 56.2 225.4 56.8 ;
      RECT  221.6 51.2 222.4 52.0 ;
      RECT  207.6 47.4 229.4 48.6 ;
      RECT  215.2 57.2 216.0 57.4 ;
      RECT  212.6 55.4 213.4 55.6 ;
      RECT  218.2 61.4 219.0 61.6 ;
      RECT  226.4 49.2 227.2 53.6 ;
      RECT  209.6 54.6 211.2 54.8 ;
      RECT  212.0 62.0 212.8 62.8 ;
      RECT  217.6 49.2 218.4 51.2 ;
      RECT  211.0 56.4 211.8 56.6 ;
      RECT  212.0 60.0 212.8 60.2 ;
      RECT  223.4 53.4 224.2 53.6 ;
      RECT  213.6 51.8 214.4 52.6 ;
      RECT  224.8 48.6 225.6 53.0 ;
      RECT  219.4 59.8 220.2 60.0 ;
      RECT  215.8 48.6 216.8 51.2 ;
      RECT  213.8 52.6 214.4 54.8 ;
      RECT  219.2 62.8 220.0 67.4 ;
      RECT  216.0 62.8 216.8 67.4 ;
      RECT  219.4 54.6 220.2 54.8 ;
      RECT  213.8 58.4 218.6 58.8 ;
      RECT  208.8 58.0 214.6 58.2 ;
      RECT  217.6 62.8 218.4 66.8 ;
      RECT  224.6 56.8 225.4 57.0 ;
      RECT  208.8 58.2 218.6 58.4 ;
      RECT  216.6 60.0 217.4 60.2 ;
      RECT  221.8 49.2 223.0 50.6 ;
      RECT  215.4 52.4 216.2 52.6 ;
      RECT  221.8 60.2 223.2 61.0 ;
      RECT  223.0 57.4 223.8 57.6 ;
      RECT  212.0 51.2 212.8 52.0 ;
      RECT  210.4 48.6 211.2 53.2 ;
      RECT  223.4 53.6 227.2 54.2 ;
      RECT  196.3 67.6 197.1 68.4 ;
      RECT  196.3 47.6 197.1 48.4 ;
      RECT  218.1 67.6 218.9 68.4 ;
      RECT  218.1 47.6 218.9 48.4 ;
      RECT  87.6 10.8 88.4 11.6 ;
      RECT  86.2 152.2 87.0 153.0 ;
      RECT  86.2 90.8 87.0 91.6 ;
      RECT  86.2 112.0 87.0 112.8 ;
      RECT  86.2 72.8 87.0 73.6 ;
      RECT  202.4 70.4 203.2 71.2 ;
      RECT  204.6 70.4 205.4 71.2 ;
      RECT  209.2 71.8 210.0 72.6 ;
      RECT  226.4 71.8 227.2 72.6 ;
   LAYER  metal2 ;
      RECT  87.7 11.2 88.3 298.2 ;
      RECT  87.6 11.2 88.4 53.4 ;
      RECT  87.7 11.2 88.3 53.4 ;
      RECT  180.2 152.6 180.8 191.4 ;
      RECT  178.8 75.0 179.4 91.2 ;
      RECT  181.6 75.0 182.2 112.4 ;
      RECT  183.0 73.2 183.6 75.0 ;
      RECT  193.9 167.5 194.5 173.4 ;
      RECT  89.5 236.2 90.1 302.6 ;
      RECT  90.9 236.2 91.5 323.0 ;
      RECT  92.3 236.2 92.9 342.6 ;
      RECT  93.7 236.2 94.3 363.0 ;
      RECT  202.5 70.8 203.1 76.0 ;
      RECT  204.7 57.8 205.3 70.8 ;
      RECT  209.3 72.2 209.9 76.0 ;
      RECT  226.5 57.8 227.1 72.2 ;
      RECT  200.7 169.2 201.3 171.3 ;
      RECT  200.7 171.3 201.3 173.4 ;
      RECT  204.3 169.2 204.9 171.3 ;
      RECT  204.3 171.3 204.9 173.4 ;
      RECT  207.5 169.2 208.1 171.3 ;
      RECT  207.5 171.3 208.1 173.4 ;
      RECT  211.1 169.2 211.7 171.3 ;
      RECT  211.1 171.3 211.7 173.4 ;
      RECT  193.9 169.2 194.5 171.3 ;
      RECT  193.9 171.3 194.5 173.4 ;
      RECT  197.5 169.2 198.1 171.3 ;
      RECT  197.5 171.3 198.1 173.4 ;
      RECT  181.6 133.2 182.2 160.1 ;
      RECT  183.0 133.2 183.6 191.6 ;
      RECT  178.8 80.1 179.4 133.2 ;
      RECT  180.2 133.2 180.8 149.9 ;
      RECT  161.5 186.2 162.1 194.6 ;
      RECT  202.4 204.2 203.2 205.0 ;
      RECT  199.0 194.2 199.8 205.0 ;
      RECT  204.2 195.8 205.0 205.0 ;
      RECT  200.6 194.2 201.4 205.0 ;
      RECT  203.4 195.0 205.0 195.8 ;
      RECT  205.8 194.2 206.6 205.0 ;
      RECT  204.2 194.2 205.0 195.0 ;
      RECT  202.4 205.0 203.2 204.2 ;
      RECT  199.0 215.0 199.8 204.2 ;
      RECT  204.2 213.4 205.0 204.2 ;
      RECT  200.6 215.0 201.4 204.2 ;
      RECT  203.4 214.2 205.0 213.4 ;
      RECT  205.8 215.0 206.6 204.2 ;
      RECT  204.2 215.0 205.0 214.2 ;
      RECT  202.4 225.0 203.2 225.8 ;
      RECT  199.0 215.0 199.8 225.8 ;
      RECT  204.2 216.6 205.0 225.8 ;
      RECT  200.6 215.0 201.4 225.8 ;
      RECT  203.4 215.8 205.0 216.6 ;
      RECT  205.8 215.0 206.6 225.8 ;
      RECT  204.2 215.0 205.0 215.8 ;
      RECT  202.4 225.8 203.2 225.0 ;
      RECT  199.0 235.8 199.8 225.0 ;
      RECT  204.2 234.2 205.0 225.0 ;
      RECT  200.6 235.8 201.4 225.0 ;
      RECT  203.4 235.0 205.0 234.2 ;
      RECT  205.8 235.8 206.6 225.0 ;
      RECT  204.2 235.8 205.0 235.0 ;
      RECT  202.4 245.8 203.2 246.6 ;
      RECT  199.0 235.8 199.8 246.6 ;
      RECT  204.2 237.4 205.0 246.6 ;
      RECT  200.6 235.8 201.4 246.6 ;
      RECT  203.4 236.6 205.0 237.4 ;
      RECT  205.8 235.8 206.6 246.6 ;
      RECT  204.2 235.8 205.0 236.6 ;
      RECT  202.4 246.6 203.2 245.8 ;
      RECT  199.0 256.6 199.8 245.8 ;
      RECT  204.2 255.0 205.0 245.8 ;
      RECT  200.6 256.6 201.4 245.8 ;
      RECT  203.4 255.8 205.0 255.0 ;
      RECT  205.8 256.6 206.6 245.8 ;
      RECT  204.2 256.6 205.0 255.8 ;
      RECT  202.4 266.6 203.2 267.4 ;
      RECT  199.0 256.6 199.8 267.4 ;
      RECT  204.2 258.2 205.0 267.4 ;
      RECT  200.6 256.6 201.4 267.4 ;
      RECT  203.4 257.4 205.0 258.2 ;
      RECT  205.8 256.6 206.6 267.4 ;
      RECT  204.2 256.6 205.0 257.4 ;
      RECT  202.4 267.4 203.2 266.6 ;
      RECT  199.0 277.4 199.8 266.6 ;
      RECT  204.2 275.8 205.0 266.6 ;
      RECT  200.6 277.4 201.4 266.6 ;
      RECT  203.4 276.6 205.0 275.8 ;
      RECT  205.8 277.4 206.6 266.6 ;
      RECT  204.2 277.4 205.0 276.6 ;
      RECT  202.4 287.4 203.2 288.2 ;
      RECT  199.0 277.4 199.8 288.2 ;
      RECT  204.2 279.0 205.0 288.2 ;
      RECT  200.6 277.4 201.4 288.2 ;
      RECT  203.4 278.2 205.0 279.0 ;
      RECT  205.8 277.4 206.6 288.2 ;
      RECT  204.2 277.4 205.0 278.2 ;
      RECT  202.4 288.2 203.2 287.4 ;
      RECT  199.0 298.2 199.8 287.4 ;
      RECT  204.2 296.6 205.0 287.4 ;
      RECT  200.6 298.2 201.4 287.4 ;
      RECT  203.4 297.4 205.0 296.6 ;
      RECT  205.8 298.2 206.6 287.4 ;
      RECT  204.2 298.2 205.0 297.4 ;
      RECT  202.4 308.2 203.2 309.0 ;
      RECT  199.0 298.2 199.8 309.0 ;
      RECT  204.2 299.8 205.0 309.0 ;
      RECT  200.6 298.2 201.4 309.0 ;
      RECT  203.4 299.0 205.0 299.8 ;
      RECT  205.8 298.2 206.6 309.0 ;
      RECT  204.2 298.2 205.0 299.0 ;
      RECT  202.4 309.0 203.2 308.2 ;
      RECT  199.0 319.0 199.8 308.2 ;
      RECT  204.2 317.4 205.0 308.2 ;
      RECT  200.6 319.0 201.4 308.2 ;
      RECT  203.4 318.2 205.0 317.4 ;
      RECT  205.8 319.0 206.6 308.2 ;
      RECT  204.2 319.0 205.0 318.2 ;
      RECT  202.4 329.0 203.2 329.8 ;
      RECT  199.0 319.0 199.8 329.8 ;
      RECT  204.2 320.6 205.0 329.8 ;
      RECT  200.6 319.0 201.4 329.8 ;
      RECT  203.4 319.8 205.0 320.6 ;
      RECT  205.8 319.0 206.6 329.8 ;
      RECT  204.2 319.0 205.0 319.8 ;
      RECT  202.4 329.8 203.2 329.0 ;
      RECT  199.0 339.8 199.8 329.0 ;
      RECT  204.2 338.2 205.0 329.0 ;
      RECT  200.6 339.8 201.4 329.0 ;
      RECT  203.4 339.0 205.0 338.2 ;
      RECT  205.8 339.8 206.6 329.0 ;
      RECT  204.2 339.8 205.0 339.0 ;
      RECT  202.4 349.8 203.2 350.6 ;
      RECT  199.0 339.8 199.8 350.6 ;
      RECT  204.2 341.4 205.0 350.6 ;
      RECT  200.6 339.8 201.4 350.6 ;
      RECT  203.4 340.6 205.0 341.4 ;
      RECT  205.8 339.8 206.6 350.6 ;
      RECT  204.2 339.8 205.0 340.6 ;
      RECT  202.4 350.6 203.2 349.8 ;
      RECT  199.0 360.6 199.8 349.8 ;
      RECT  204.2 359.0 205.0 349.8 ;
      RECT  200.6 360.6 201.4 349.8 ;
      RECT  203.4 359.8 205.0 359.0 ;
      RECT  205.8 360.6 206.6 349.8 ;
      RECT  204.2 360.6 205.0 359.8 ;
      RECT  209.2 204.2 210.0 205.0 ;
      RECT  205.8 194.2 206.6 205.0 ;
      RECT  211.0 195.8 211.8 205.0 ;
      RECT  207.4 194.2 208.2 205.0 ;
      RECT  210.2 195.0 211.8 195.8 ;
      RECT  212.6 194.2 213.4 205.0 ;
      RECT  211.0 194.2 211.8 195.0 ;
      RECT  209.2 205.0 210.0 204.2 ;
      RECT  205.8 215.0 206.6 204.2 ;
      RECT  211.0 213.4 211.8 204.2 ;
      RECT  207.4 215.0 208.2 204.2 ;
      RECT  210.2 214.2 211.8 213.4 ;
      RECT  212.6 215.0 213.4 204.2 ;
      RECT  211.0 215.0 211.8 214.2 ;
      RECT  209.2 225.0 210.0 225.8 ;
      RECT  205.8 215.0 206.6 225.8 ;
      RECT  211.0 216.6 211.8 225.8 ;
      RECT  207.4 215.0 208.2 225.8 ;
      RECT  210.2 215.8 211.8 216.6 ;
      RECT  212.6 215.0 213.4 225.8 ;
      RECT  211.0 215.0 211.8 215.8 ;
      RECT  209.2 225.8 210.0 225.0 ;
      RECT  205.8 235.8 206.6 225.0 ;
      RECT  211.0 234.2 211.8 225.0 ;
      RECT  207.4 235.8 208.2 225.0 ;
      RECT  210.2 235.0 211.8 234.2 ;
      RECT  212.6 235.8 213.4 225.0 ;
      RECT  211.0 235.8 211.8 235.0 ;
      RECT  209.2 245.8 210.0 246.6 ;
      RECT  205.8 235.8 206.6 246.6 ;
      RECT  211.0 237.4 211.8 246.6 ;
      RECT  207.4 235.8 208.2 246.6 ;
      RECT  210.2 236.6 211.8 237.4 ;
      RECT  212.6 235.8 213.4 246.6 ;
      RECT  211.0 235.8 211.8 236.6 ;
      RECT  209.2 246.6 210.0 245.8 ;
      RECT  205.8 256.6 206.6 245.8 ;
      RECT  211.0 255.0 211.8 245.8 ;
      RECT  207.4 256.6 208.2 245.8 ;
      RECT  210.2 255.8 211.8 255.0 ;
      RECT  212.6 256.6 213.4 245.8 ;
      RECT  211.0 256.6 211.8 255.8 ;
      RECT  209.2 266.6 210.0 267.4 ;
      RECT  205.8 256.6 206.6 267.4 ;
      RECT  211.0 258.2 211.8 267.4 ;
      RECT  207.4 256.6 208.2 267.4 ;
      RECT  210.2 257.4 211.8 258.2 ;
      RECT  212.6 256.6 213.4 267.4 ;
      RECT  211.0 256.6 211.8 257.4 ;
      RECT  209.2 267.4 210.0 266.6 ;
      RECT  205.8 277.4 206.6 266.6 ;
      RECT  211.0 275.8 211.8 266.6 ;
      RECT  207.4 277.4 208.2 266.6 ;
      RECT  210.2 276.6 211.8 275.8 ;
      RECT  212.6 277.4 213.4 266.6 ;
      RECT  211.0 277.4 211.8 276.6 ;
      RECT  209.2 287.4 210.0 288.2 ;
      RECT  205.8 277.4 206.6 288.2 ;
      RECT  211.0 279.0 211.8 288.2 ;
      RECT  207.4 277.4 208.2 288.2 ;
      RECT  210.2 278.2 211.8 279.0 ;
      RECT  212.6 277.4 213.4 288.2 ;
      RECT  211.0 277.4 211.8 278.2 ;
      RECT  209.2 288.2 210.0 287.4 ;
      RECT  205.8 298.2 206.6 287.4 ;
      RECT  211.0 296.6 211.8 287.4 ;
      RECT  207.4 298.2 208.2 287.4 ;
      RECT  210.2 297.4 211.8 296.6 ;
      RECT  212.6 298.2 213.4 287.4 ;
      RECT  211.0 298.2 211.8 297.4 ;
      RECT  209.2 308.2 210.0 309.0 ;
      RECT  205.8 298.2 206.6 309.0 ;
      RECT  211.0 299.8 211.8 309.0 ;
      RECT  207.4 298.2 208.2 309.0 ;
      RECT  210.2 299.0 211.8 299.8 ;
      RECT  212.6 298.2 213.4 309.0 ;
      RECT  211.0 298.2 211.8 299.0 ;
      RECT  209.2 309.0 210.0 308.2 ;
      RECT  205.8 319.0 206.6 308.2 ;
      RECT  211.0 317.4 211.8 308.2 ;
      RECT  207.4 319.0 208.2 308.2 ;
      RECT  210.2 318.2 211.8 317.4 ;
      RECT  212.6 319.0 213.4 308.2 ;
      RECT  211.0 319.0 211.8 318.2 ;
      RECT  209.2 329.0 210.0 329.8 ;
      RECT  205.8 319.0 206.6 329.8 ;
      RECT  211.0 320.6 211.8 329.8 ;
      RECT  207.4 319.0 208.2 329.8 ;
      RECT  210.2 319.8 211.8 320.6 ;
      RECT  212.6 319.0 213.4 329.8 ;
      RECT  211.0 319.0 211.8 319.8 ;
      RECT  209.2 329.8 210.0 329.0 ;
      RECT  205.8 339.8 206.6 329.0 ;
      RECT  211.0 338.2 211.8 329.0 ;
      RECT  207.4 339.8 208.2 329.0 ;
      RECT  210.2 339.0 211.8 338.2 ;
      RECT  212.6 339.8 213.4 329.0 ;
      RECT  211.0 339.8 211.8 339.0 ;
      RECT  209.2 349.8 210.0 350.6 ;
      RECT  205.8 339.8 206.6 350.6 ;
      RECT  211.0 341.4 211.8 350.6 ;
      RECT  207.4 339.8 208.2 350.6 ;
      RECT  210.2 340.6 211.8 341.4 ;
      RECT  212.6 339.8 213.4 350.6 ;
      RECT  211.0 339.8 211.8 340.6 ;
      RECT  209.2 350.6 210.0 349.8 ;
      RECT  205.8 360.6 206.6 349.8 ;
      RECT  211.0 359.0 211.8 349.8 ;
      RECT  207.4 360.6 208.2 349.8 ;
      RECT  210.2 359.8 211.8 359.0 ;
      RECT  212.6 360.6 213.4 349.8 ;
      RECT  211.0 360.6 211.8 359.8 ;
      RECT  202.4 204.2 203.2 205.0 ;
      RECT  199.0 199.2 199.8 200.0 ;
      RECT  205.8 199.2 206.6 200.0 ;
      RECT  209.2 204.2 210.0 205.0 ;
      RECT  205.8 199.2 206.6 200.0 ;
      RECT  212.6 199.2 213.4 200.0 ;
      RECT  202.4 204.2 203.2 205.0 ;
      RECT  199.0 209.2 199.8 210.0 ;
      RECT  205.8 209.2 206.6 210.0 ;
      RECT  209.2 204.2 210.0 205.0 ;
      RECT  205.8 209.2 206.6 210.0 ;
      RECT  212.6 209.2 213.4 210.0 ;
      RECT  202.4 225.0 203.2 225.8 ;
      RECT  199.0 220.0 199.8 220.8 ;
      RECT  205.8 220.0 206.6 220.8 ;
      RECT  209.2 225.0 210.0 225.8 ;
      RECT  205.8 220.0 206.6 220.8 ;
      RECT  212.6 220.0 213.4 220.8 ;
      RECT  202.4 225.0 203.2 225.8 ;
      RECT  199.0 230.0 199.8 230.8 ;
      RECT  205.8 230.0 206.6 230.8 ;
      RECT  209.2 225.0 210.0 225.8 ;
      RECT  205.8 230.0 206.6 230.8 ;
      RECT  212.6 230.0 213.4 230.8 ;
      RECT  202.4 245.8 203.2 246.6 ;
      RECT  199.0 240.8 199.8 241.6 ;
      RECT  205.8 240.8 206.6 241.6 ;
      RECT  209.2 245.8 210.0 246.6 ;
      RECT  205.8 240.8 206.6 241.6 ;
      RECT  212.6 240.8 213.4 241.6 ;
      RECT  202.4 245.8 203.2 246.6 ;
      RECT  199.0 250.8 199.8 251.6 ;
      RECT  205.8 250.8 206.6 251.6 ;
      RECT  209.2 245.8 210.0 246.6 ;
      RECT  205.8 250.8 206.6 251.6 ;
      RECT  212.6 250.8 213.4 251.6 ;
      RECT  202.4 266.6 203.2 267.4 ;
      RECT  199.0 261.6 199.8 262.4 ;
      RECT  205.8 261.6 206.6 262.4 ;
      RECT  209.2 266.6 210.0 267.4 ;
      RECT  205.8 261.6 206.6 262.4 ;
      RECT  212.6 261.6 213.4 262.4 ;
      RECT  202.4 266.6 203.2 267.4 ;
      RECT  199.0 271.6 199.8 272.4 ;
      RECT  205.8 271.6 206.6 272.4 ;
      RECT  209.2 266.6 210.0 267.4 ;
      RECT  205.8 271.6 206.6 272.4 ;
      RECT  212.6 271.6 213.4 272.4 ;
      RECT  202.4 287.4 203.2 288.2 ;
      RECT  199.0 282.4 199.8 283.2 ;
      RECT  205.8 282.4 206.6 283.2 ;
      RECT  209.2 287.4 210.0 288.2 ;
      RECT  205.8 282.4 206.6 283.2 ;
      RECT  212.6 282.4 213.4 283.2 ;
      RECT  202.4 287.4 203.2 288.2 ;
      RECT  199.0 292.4 199.8 293.2 ;
      RECT  205.8 292.4 206.6 293.2 ;
      RECT  209.2 287.4 210.0 288.2 ;
      RECT  205.8 292.4 206.6 293.2 ;
      RECT  212.6 292.4 213.4 293.2 ;
      RECT  202.4 308.2 203.2 309.0 ;
      RECT  199.0 303.2 199.8 304.0 ;
      RECT  205.8 303.2 206.6 304.0 ;
      RECT  209.2 308.2 210.0 309.0 ;
      RECT  205.8 303.2 206.6 304.0 ;
      RECT  212.6 303.2 213.4 304.0 ;
      RECT  202.4 308.2 203.2 309.0 ;
      RECT  199.0 313.2 199.8 314.0 ;
      RECT  205.8 313.2 206.6 314.0 ;
      RECT  209.2 308.2 210.0 309.0 ;
      RECT  205.8 313.2 206.6 314.0 ;
      RECT  212.6 313.2 213.4 314.0 ;
      RECT  202.4 329.0 203.2 329.8 ;
      RECT  199.0 324.0 199.8 324.8 ;
      RECT  205.8 324.0 206.6 324.8 ;
      RECT  209.2 329.0 210.0 329.8 ;
      RECT  205.8 324.0 206.6 324.8 ;
      RECT  212.6 324.0 213.4 324.8 ;
      RECT  202.4 329.0 203.2 329.8 ;
      RECT  199.0 334.0 199.8 334.8 ;
      RECT  205.8 334.0 206.6 334.8 ;
      RECT  209.2 329.0 210.0 329.8 ;
      RECT  205.8 334.0 206.6 334.8 ;
      RECT  212.6 334.0 213.4 334.8 ;
      RECT  202.4 349.8 203.2 350.6 ;
      RECT  199.0 344.8 199.8 345.6 ;
      RECT  205.8 344.8 206.6 345.6 ;
      RECT  209.2 349.8 210.0 350.6 ;
      RECT  205.8 344.8 206.6 345.6 ;
      RECT  212.6 344.8 213.4 345.6 ;
      RECT  202.4 349.8 203.2 350.6 ;
      RECT  199.0 354.8 199.8 355.6 ;
      RECT  205.8 354.8 206.6 355.6 ;
      RECT  209.2 349.8 210.0 350.6 ;
      RECT  205.8 354.8 206.6 355.6 ;
      RECT  212.6 354.8 213.4 355.6 ;
      RECT  200.6 194.2 201.4 360.6 ;
      RECT  204.2 194.2 205.0 360.6 ;
      RECT  207.4 194.2 208.2 360.6 ;
      RECT  211.0 194.2 211.8 360.6 ;
      RECT  195.6 183.4 196.4 184.2 ;
      RECT  192.2 173.4 193.0 184.2 ;
      RECT  193.8 173.4 194.6 184.2 ;
      RECT  197.4 173.4 198.2 184.2 ;
      RECT  199.0 173.4 199.8 184.2 ;
      RECT  195.6 184.2 196.4 183.4 ;
      RECT  192.2 194.2 193.0 183.4 ;
      RECT  197.4 192.6 198.2 183.4 ;
      RECT  193.8 194.2 194.6 183.4 ;
      RECT  196.6 193.4 198.2 192.6 ;
      RECT  199.0 194.2 199.8 183.4 ;
      RECT  197.4 194.2 198.2 193.4 ;
      RECT  195.6 204.2 196.4 205.0 ;
      RECT  192.2 194.2 193.0 205.0 ;
      RECT  197.4 195.8 198.2 205.0 ;
      RECT  193.8 194.2 194.6 205.0 ;
      RECT  196.6 195.0 198.2 195.8 ;
      RECT  199.0 194.2 199.8 205.0 ;
      RECT  197.4 194.2 198.2 195.0 ;
      RECT  195.6 205.0 196.4 204.2 ;
      RECT  192.2 215.0 193.0 204.2 ;
      RECT  197.4 213.4 198.2 204.2 ;
      RECT  193.8 215.0 194.6 204.2 ;
      RECT  196.6 214.2 198.2 213.4 ;
      RECT  199.0 215.0 199.8 204.2 ;
      RECT  197.4 215.0 198.2 214.2 ;
      RECT  195.6 225.0 196.4 225.8 ;
      RECT  192.2 215.0 193.0 225.8 ;
      RECT  197.4 216.6 198.2 225.8 ;
      RECT  193.8 215.0 194.6 225.8 ;
      RECT  196.6 215.8 198.2 216.6 ;
      RECT  199.0 215.0 199.8 225.8 ;
      RECT  197.4 215.0 198.2 215.8 ;
      RECT  195.6 225.8 196.4 225.0 ;
      RECT  192.2 235.8 193.0 225.0 ;
      RECT  197.4 234.2 198.2 225.0 ;
      RECT  193.8 235.8 194.6 225.0 ;
      RECT  196.6 235.0 198.2 234.2 ;
      RECT  199.0 235.8 199.8 225.0 ;
      RECT  197.4 235.8 198.2 235.0 ;
      RECT  195.6 245.8 196.4 246.6 ;
      RECT  192.2 235.8 193.0 246.6 ;
      RECT  197.4 237.4 198.2 246.6 ;
      RECT  193.8 235.8 194.6 246.6 ;
      RECT  196.6 236.6 198.2 237.4 ;
      RECT  199.0 235.8 199.8 246.6 ;
      RECT  197.4 235.8 198.2 236.6 ;
      RECT  195.6 246.6 196.4 245.8 ;
      RECT  192.2 256.6 193.0 245.8 ;
      RECT  197.4 255.0 198.2 245.8 ;
      RECT  193.8 256.6 194.6 245.8 ;
      RECT  196.6 255.8 198.2 255.0 ;
      RECT  199.0 256.6 199.8 245.8 ;
      RECT  197.4 256.6 198.2 255.8 ;
      RECT  195.6 266.6 196.4 267.4 ;
      RECT  192.2 256.6 193.0 267.4 ;
      RECT  197.4 258.2 198.2 267.4 ;
      RECT  193.8 256.6 194.6 267.4 ;
      RECT  196.6 257.4 198.2 258.2 ;
      RECT  199.0 256.6 199.8 267.4 ;
      RECT  197.4 256.6 198.2 257.4 ;
      RECT  195.6 267.4 196.4 266.6 ;
      RECT  192.2 277.4 193.0 266.6 ;
      RECT  197.4 275.8 198.2 266.6 ;
      RECT  193.8 277.4 194.6 266.6 ;
      RECT  196.6 276.6 198.2 275.8 ;
      RECT  199.0 277.4 199.8 266.6 ;
      RECT  197.4 277.4 198.2 276.6 ;
      RECT  195.6 287.4 196.4 288.2 ;
      RECT  192.2 277.4 193.0 288.2 ;
      RECT  197.4 279.0 198.2 288.2 ;
      RECT  193.8 277.4 194.6 288.2 ;
      RECT  196.6 278.2 198.2 279.0 ;
      RECT  199.0 277.4 199.8 288.2 ;
      RECT  197.4 277.4 198.2 278.2 ;
      RECT  195.6 288.2 196.4 287.4 ;
      RECT  192.2 298.2 193.0 287.4 ;
      RECT  197.4 296.6 198.2 287.4 ;
      RECT  193.8 298.2 194.6 287.4 ;
      RECT  196.6 297.4 198.2 296.6 ;
      RECT  199.0 298.2 199.8 287.4 ;
      RECT  197.4 298.2 198.2 297.4 ;
      RECT  195.6 308.2 196.4 309.0 ;
      RECT  192.2 298.2 193.0 309.0 ;
      RECT  197.4 299.8 198.2 309.0 ;
      RECT  193.8 298.2 194.6 309.0 ;
      RECT  196.6 299.0 198.2 299.8 ;
      RECT  199.0 298.2 199.8 309.0 ;
      RECT  197.4 298.2 198.2 299.0 ;
      RECT  195.6 309.0 196.4 308.2 ;
      RECT  192.2 319.0 193.0 308.2 ;
      RECT  197.4 317.4 198.2 308.2 ;
      RECT  193.8 319.0 194.6 308.2 ;
      RECT  196.6 318.2 198.2 317.4 ;
      RECT  199.0 319.0 199.8 308.2 ;
      RECT  197.4 319.0 198.2 318.2 ;
      RECT  195.6 329.0 196.4 329.8 ;
      RECT  192.2 319.0 193.0 329.8 ;
      RECT  197.4 320.6 198.2 329.8 ;
      RECT  193.8 319.0 194.6 329.8 ;
      RECT  196.6 319.8 198.2 320.6 ;
      RECT  199.0 319.0 199.8 329.8 ;
      RECT  197.4 319.0 198.2 319.8 ;
      RECT  195.6 329.8 196.4 329.0 ;
      RECT  192.2 339.8 193.0 329.0 ;
      RECT  197.4 338.2 198.2 329.0 ;
      RECT  193.8 339.8 194.6 329.0 ;
      RECT  196.6 339.0 198.2 338.2 ;
      RECT  199.0 339.8 199.8 329.0 ;
      RECT  197.4 339.8 198.2 339.0 ;
      RECT  195.6 349.8 196.4 350.6 ;
      RECT  192.2 339.8 193.0 350.6 ;
      RECT  197.4 341.4 198.2 350.6 ;
      RECT  193.8 339.8 194.6 350.6 ;
      RECT  196.6 340.6 198.2 341.4 ;
      RECT  199.0 339.8 199.8 350.6 ;
      RECT  197.4 339.8 198.2 340.6 ;
      RECT  195.6 350.6 196.4 349.8 ;
      RECT  192.2 360.6 193.0 349.8 ;
      RECT  197.4 359.0 198.2 349.8 ;
      RECT  193.8 360.6 194.6 349.8 ;
      RECT  196.6 359.8 198.2 359.0 ;
      RECT  199.0 360.6 199.8 349.8 ;
      RECT  197.4 360.6 198.2 359.8 ;
      RECT  195.6 370.6 196.4 371.4 ;
      RECT  192.2 360.6 193.0 371.4 ;
      RECT  193.8 360.6 194.6 371.4 ;
      RECT  197.4 360.6 198.2 371.4 ;
      RECT  199.0 360.6 199.8 371.4 ;
      RECT  195.6 266.6 196.4 267.4 ;
      RECT  195.6 183.4 196.4 184.2 ;
      RECT  195.6 287.4 196.4 288.2 ;
      RECT  195.6 225.0 196.4 225.8 ;
      RECT  195.6 370.6 196.4 371.4 ;
      RECT  195.6 245.8 196.4 246.6 ;
      RECT  195.6 349.8 196.4 350.6 ;
      RECT  195.6 204.2 196.4 205.0 ;
      RECT  195.6 329.0 196.4 329.8 ;
      RECT  195.6 308.2 196.4 309.0 ;
      RECT  199.0 256.6 199.8 267.4 ;
      RECT  192.2 245.8 193.0 256.6 ;
      RECT  192.2 225.0 193.0 235.8 ;
      RECT  192.2 256.6 193.0 267.4 ;
      RECT  199.0 277.4 199.8 288.2 ;
      RECT  199.0 360.6 199.8 371.4 ;
      RECT  199.0 183.4 199.8 194.2 ;
      RECT  192.2 204.2 193.0 215.0 ;
      RECT  192.2 360.6 193.0 371.4 ;
      RECT  199.0 266.6 199.8 277.4 ;
      RECT  192.2 308.2 193.0 319.0 ;
      RECT  199.0 287.4 199.8 298.2 ;
      RECT  199.0 339.8 199.8 350.6 ;
      RECT  199.0 194.2 199.8 205.0 ;
      RECT  199.0 245.8 199.8 256.6 ;
      RECT  192.2 266.6 193.0 277.4 ;
      RECT  192.2 235.8 193.0 246.6 ;
      RECT  199.0 308.2 199.8 319.0 ;
      RECT  192.2 173.4 193.0 184.2 ;
      RECT  192.2 298.2 193.0 309.0 ;
      RECT  199.0 349.8 199.8 360.6 ;
      RECT  192.2 215.0 193.0 225.8 ;
      RECT  192.2 277.4 193.0 288.2 ;
      RECT  199.0 298.2 199.8 309.0 ;
      RECT  199.0 173.4 199.8 184.2 ;
      RECT  199.0 235.8 199.8 246.6 ;
      RECT  199.0 215.0 199.8 225.8 ;
      RECT  192.2 329.0 193.0 339.8 ;
      RECT  199.0 225.0 199.8 235.8 ;
      RECT  192.2 183.4 193.0 194.2 ;
      RECT  192.2 287.4 193.0 298.2 ;
      RECT  192.2 319.0 193.0 329.8 ;
      RECT  199.0 329.0 199.8 339.8 ;
      RECT  192.2 194.2 193.0 205.0 ;
      RECT  199.0 319.0 199.8 329.8 ;
      RECT  192.2 339.8 193.0 350.6 ;
      RECT  199.0 204.2 199.8 215.0 ;
      RECT  192.2 349.8 193.0 360.6 ;
      RECT  202.4 184.2 203.2 183.4 ;
      RECT  199.0 194.2 199.8 183.4 ;
      RECT  200.6 194.2 201.4 183.4 ;
      RECT  204.2 194.2 205.0 183.4 ;
      RECT  205.8 194.2 206.6 183.4 ;
      RECT  209.2 184.2 210.0 183.4 ;
      RECT  205.8 194.2 206.6 183.4 ;
      RECT  207.4 194.2 208.2 183.4 ;
      RECT  211.0 194.2 211.8 183.4 ;
      RECT  212.6 194.2 213.4 183.4 ;
      RECT  202.4 184.2 203.2 183.4 ;
      RECT  199.0 189.2 199.8 188.4 ;
      RECT  205.8 189.2 206.6 188.4 ;
      RECT  209.2 184.2 210.0 183.4 ;
      RECT  205.8 189.2 206.6 188.4 ;
      RECT  212.6 189.2 213.4 188.4 ;
      RECT  200.6 194.2 201.4 183.8 ;
      RECT  204.2 194.2 205.0 183.8 ;
      RECT  207.4 194.2 208.2 183.8 ;
      RECT  211.0 194.2 211.8 183.8 ;
      RECT  202.4 183.4 203.2 184.2 ;
      RECT  199.0 173.4 199.8 184.2 ;
      RECT  200.6 173.4 201.4 184.2 ;
      RECT  204.2 173.4 205.0 184.2 ;
      RECT  205.8 173.4 206.6 184.2 ;
      RECT  209.2 183.4 210.0 184.2 ;
      RECT  205.8 173.4 206.6 184.2 ;
      RECT  207.4 173.4 208.2 184.2 ;
      RECT  211.0 173.4 211.8 184.2 ;
      RECT  212.6 173.4 213.4 184.2 ;
      RECT  202.4 183.4 203.2 184.2 ;
      RECT  199.0 178.4 199.8 179.2 ;
      RECT  205.8 178.4 206.6 179.2 ;
      RECT  209.2 183.4 210.0 184.2 ;
      RECT  205.8 178.4 206.6 179.2 ;
      RECT  212.6 178.4 213.4 179.2 ;
      RECT  200.6 173.4 201.4 183.8 ;
      RECT  204.2 173.4 205.0 183.8 ;
      RECT  207.4 173.4 208.2 183.8 ;
      RECT  211.0 173.4 211.8 183.8 ;
      RECT  202.4 370.6 203.2 371.4 ;
      RECT  199.0 360.6 199.8 371.4 ;
      RECT  200.6 360.6 201.4 371.4 ;
      RECT  204.2 360.6 205.0 371.4 ;
      RECT  205.8 360.6 206.6 371.4 ;
      RECT  209.2 370.6 210.0 371.4 ;
      RECT  205.8 360.6 206.6 371.4 ;
      RECT  207.4 360.6 208.2 371.4 ;
      RECT  211.0 360.6 211.8 371.4 ;
      RECT  212.6 360.6 213.4 371.4 ;
      RECT  202.4 370.6 203.2 371.4 ;
      RECT  199.0 365.6 199.8 366.4 ;
      RECT  205.8 365.6 206.6 366.4 ;
      RECT  209.2 370.6 210.0 371.4 ;
      RECT  205.8 365.6 206.6 366.4 ;
      RECT  212.6 365.6 213.4 366.4 ;
      RECT  200.6 360.6 201.4 371.0 ;
      RECT  204.2 360.6 205.0 371.0 ;
      RECT  207.4 360.6 208.2 371.0 ;
      RECT  211.0 360.6 211.8 371.0 ;
      RECT  188.8 183.4 189.6 184.2 ;
      RECT  185.4 173.4 186.2 184.2 ;
      RECT  187.0 173.4 187.8 184.2 ;
      RECT  190.6 173.4 191.4 184.2 ;
      RECT  192.2 173.4 193.0 184.2 ;
      RECT  188.8 184.2 189.6 183.4 ;
      RECT  185.4 194.2 186.2 183.4 ;
      RECT  187.0 194.2 187.8 183.4 ;
      RECT  190.6 194.2 191.4 183.4 ;
      RECT  192.2 194.2 193.0 183.4 ;
      RECT  188.8 204.2 189.6 205.0 ;
      RECT  185.4 194.2 186.2 205.0 ;
      RECT  187.0 194.2 187.8 205.0 ;
      RECT  190.6 194.2 191.4 205.0 ;
      RECT  192.2 194.2 193.0 205.0 ;
      RECT  188.8 205.0 189.6 204.2 ;
      RECT  185.4 215.0 186.2 204.2 ;
      RECT  187.0 215.0 187.8 204.2 ;
      RECT  190.6 215.0 191.4 204.2 ;
      RECT  192.2 215.0 193.0 204.2 ;
      RECT  188.8 225.0 189.6 225.8 ;
      RECT  185.4 215.0 186.2 225.8 ;
      RECT  187.0 215.0 187.8 225.8 ;
      RECT  190.6 215.0 191.4 225.8 ;
      RECT  192.2 215.0 193.0 225.8 ;
      RECT  188.8 225.8 189.6 225.0 ;
      RECT  185.4 235.8 186.2 225.0 ;
      RECT  187.0 235.8 187.8 225.0 ;
      RECT  190.6 235.8 191.4 225.0 ;
      RECT  192.2 235.8 193.0 225.0 ;
      RECT  188.8 245.8 189.6 246.6 ;
      RECT  185.4 235.8 186.2 246.6 ;
      RECT  187.0 235.8 187.8 246.6 ;
      RECT  190.6 235.8 191.4 246.6 ;
      RECT  192.2 235.8 193.0 246.6 ;
      RECT  188.8 246.6 189.6 245.8 ;
      RECT  185.4 256.6 186.2 245.8 ;
      RECT  187.0 256.6 187.8 245.8 ;
      RECT  190.6 256.6 191.4 245.8 ;
      RECT  192.2 256.6 193.0 245.8 ;
      RECT  188.8 266.6 189.6 267.4 ;
      RECT  185.4 256.6 186.2 267.4 ;
      RECT  187.0 256.6 187.8 267.4 ;
      RECT  190.6 256.6 191.4 267.4 ;
      RECT  192.2 256.6 193.0 267.4 ;
      RECT  188.8 267.4 189.6 266.6 ;
      RECT  185.4 277.4 186.2 266.6 ;
      RECT  187.0 277.4 187.8 266.6 ;
      RECT  190.6 277.4 191.4 266.6 ;
      RECT  192.2 277.4 193.0 266.6 ;
      RECT  188.8 287.4 189.6 288.2 ;
      RECT  185.4 277.4 186.2 288.2 ;
      RECT  187.0 277.4 187.8 288.2 ;
      RECT  190.6 277.4 191.4 288.2 ;
      RECT  192.2 277.4 193.0 288.2 ;
      RECT  188.8 288.2 189.6 287.4 ;
      RECT  185.4 298.2 186.2 287.4 ;
      RECT  187.0 298.2 187.8 287.4 ;
      RECT  190.6 298.2 191.4 287.4 ;
      RECT  192.2 298.2 193.0 287.4 ;
      RECT  188.8 308.2 189.6 309.0 ;
      RECT  185.4 298.2 186.2 309.0 ;
      RECT  187.0 298.2 187.8 309.0 ;
      RECT  190.6 298.2 191.4 309.0 ;
      RECT  192.2 298.2 193.0 309.0 ;
      RECT  188.8 309.0 189.6 308.2 ;
      RECT  185.4 319.0 186.2 308.2 ;
      RECT  187.0 319.0 187.8 308.2 ;
      RECT  190.6 319.0 191.4 308.2 ;
      RECT  192.2 319.0 193.0 308.2 ;
      RECT  188.8 329.0 189.6 329.8 ;
      RECT  185.4 319.0 186.2 329.8 ;
      RECT  187.0 319.0 187.8 329.8 ;
      RECT  190.6 319.0 191.4 329.8 ;
      RECT  192.2 319.0 193.0 329.8 ;
      RECT  188.8 329.8 189.6 329.0 ;
      RECT  185.4 339.8 186.2 329.0 ;
      RECT  187.0 339.8 187.8 329.0 ;
      RECT  190.6 339.8 191.4 329.0 ;
      RECT  192.2 339.8 193.0 329.0 ;
      RECT  188.8 349.8 189.6 350.6 ;
      RECT  185.4 339.8 186.2 350.6 ;
      RECT  187.0 339.8 187.8 350.6 ;
      RECT  190.6 339.8 191.4 350.6 ;
      RECT  192.2 339.8 193.0 350.6 ;
      RECT  188.8 350.6 189.6 349.8 ;
      RECT  185.4 360.6 186.2 349.8 ;
      RECT  187.0 360.6 187.8 349.8 ;
      RECT  190.6 360.6 191.4 349.8 ;
      RECT  192.2 360.6 193.0 349.8 ;
      RECT  188.8 370.6 189.6 371.4 ;
      RECT  185.4 360.6 186.2 371.4 ;
      RECT  187.0 360.6 187.8 371.4 ;
      RECT  190.6 360.6 191.4 371.4 ;
      RECT  192.2 360.6 193.0 371.4 ;
      RECT  188.8 183.4 189.6 184.2 ;
      RECT  185.4 178.4 186.2 179.2 ;
      RECT  192.2 178.4 193.0 179.2 ;
      RECT  188.8 183.4 189.6 184.2 ;
      RECT  185.4 188.4 186.2 189.2 ;
      RECT  192.2 188.4 193.0 189.2 ;
      RECT  188.8 204.2 189.6 205.0 ;
      RECT  185.4 199.2 186.2 200.0 ;
      RECT  192.2 199.2 193.0 200.0 ;
      RECT  188.8 204.2 189.6 205.0 ;
      RECT  185.4 209.2 186.2 210.0 ;
      RECT  192.2 209.2 193.0 210.0 ;
      RECT  188.8 225.0 189.6 225.8 ;
      RECT  185.4 220.0 186.2 220.8 ;
      RECT  192.2 220.0 193.0 220.8 ;
      RECT  188.8 225.0 189.6 225.8 ;
      RECT  185.4 230.0 186.2 230.8 ;
      RECT  192.2 230.0 193.0 230.8 ;
      RECT  188.8 245.8 189.6 246.6 ;
      RECT  185.4 240.8 186.2 241.6 ;
      RECT  192.2 240.8 193.0 241.6 ;
      RECT  188.8 245.8 189.6 246.6 ;
      RECT  185.4 250.8 186.2 251.6 ;
      RECT  192.2 250.8 193.0 251.6 ;
      RECT  188.8 266.6 189.6 267.4 ;
      RECT  185.4 261.6 186.2 262.4 ;
      RECT  192.2 261.6 193.0 262.4 ;
      RECT  188.8 266.6 189.6 267.4 ;
      RECT  185.4 271.6 186.2 272.4 ;
      RECT  192.2 271.6 193.0 272.4 ;
      RECT  188.8 287.4 189.6 288.2 ;
      RECT  185.4 282.4 186.2 283.2 ;
      RECT  192.2 282.4 193.0 283.2 ;
      RECT  188.8 287.4 189.6 288.2 ;
      RECT  185.4 292.4 186.2 293.2 ;
      RECT  192.2 292.4 193.0 293.2 ;
      RECT  188.8 308.2 189.6 309.0 ;
      RECT  185.4 303.2 186.2 304.0 ;
      RECT  192.2 303.2 193.0 304.0 ;
      RECT  188.8 308.2 189.6 309.0 ;
      RECT  185.4 313.2 186.2 314.0 ;
      RECT  192.2 313.2 193.0 314.0 ;
      RECT  188.8 329.0 189.6 329.8 ;
      RECT  185.4 324.0 186.2 324.8 ;
      RECT  192.2 324.0 193.0 324.8 ;
      RECT  188.8 329.0 189.6 329.8 ;
      RECT  185.4 334.0 186.2 334.8 ;
      RECT  192.2 334.0 193.0 334.8 ;
      RECT  188.8 349.8 189.6 350.6 ;
      RECT  185.4 344.8 186.2 345.6 ;
      RECT  192.2 344.8 193.0 345.6 ;
      RECT  188.8 349.8 189.6 350.6 ;
      RECT  185.4 354.8 186.2 355.6 ;
      RECT  192.2 354.8 193.0 355.6 ;
      RECT  188.8 370.6 189.6 371.4 ;
      RECT  185.4 365.6 186.2 366.4 ;
      RECT  192.2 365.6 193.0 366.4 ;
      RECT  187.0 173.4 187.8 371.0 ;
      RECT  190.6 173.4 191.4 371.0 ;
      RECT  216.0 183.4 216.8 184.2 ;
      RECT  212.6 173.4 213.4 184.2 ;
      RECT  214.2 173.4 215.0 184.2 ;
      RECT  217.8 173.4 218.6 184.2 ;
      RECT  219.4 173.4 220.2 184.2 ;
      RECT  216.0 184.2 216.8 183.4 ;
      RECT  212.6 194.2 213.4 183.4 ;
      RECT  214.2 194.2 215.0 183.4 ;
      RECT  217.8 194.2 218.6 183.4 ;
      RECT  219.4 194.2 220.2 183.4 ;
      RECT  216.0 204.2 216.8 205.0 ;
      RECT  212.6 194.2 213.4 205.0 ;
      RECT  214.2 194.2 215.0 205.0 ;
      RECT  217.8 194.2 218.6 205.0 ;
      RECT  219.4 194.2 220.2 205.0 ;
      RECT  216.0 205.0 216.8 204.2 ;
      RECT  212.6 215.0 213.4 204.2 ;
      RECT  214.2 215.0 215.0 204.2 ;
      RECT  217.8 215.0 218.6 204.2 ;
      RECT  219.4 215.0 220.2 204.2 ;
      RECT  216.0 225.0 216.8 225.8 ;
      RECT  212.6 215.0 213.4 225.8 ;
      RECT  214.2 215.0 215.0 225.8 ;
      RECT  217.8 215.0 218.6 225.8 ;
      RECT  219.4 215.0 220.2 225.8 ;
      RECT  216.0 225.8 216.8 225.0 ;
      RECT  212.6 235.8 213.4 225.0 ;
      RECT  214.2 235.8 215.0 225.0 ;
      RECT  217.8 235.8 218.6 225.0 ;
      RECT  219.4 235.8 220.2 225.0 ;
      RECT  216.0 245.8 216.8 246.6 ;
      RECT  212.6 235.8 213.4 246.6 ;
      RECT  214.2 235.8 215.0 246.6 ;
      RECT  217.8 235.8 218.6 246.6 ;
      RECT  219.4 235.8 220.2 246.6 ;
      RECT  216.0 246.6 216.8 245.8 ;
      RECT  212.6 256.6 213.4 245.8 ;
      RECT  214.2 256.6 215.0 245.8 ;
      RECT  217.8 256.6 218.6 245.8 ;
      RECT  219.4 256.6 220.2 245.8 ;
      RECT  216.0 266.6 216.8 267.4 ;
      RECT  212.6 256.6 213.4 267.4 ;
      RECT  214.2 256.6 215.0 267.4 ;
      RECT  217.8 256.6 218.6 267.4 ;
      RECT  219.4 256.6 220.2 267.4 ;
      RECT  216.0 267.4 216.8 266.6 ;
      RECT  212.6 277.4 213.4 266.6 ;
      RECT  214.2 277.4 215.0 266.6 ;
      RECT  217.8 277.4 218.6 266.6 ;
      RECT  219.4 277.4 220.2 266.6 ;
      RECT  216.0 287.4 216.8 288.2 ;
      RECT  212.6 277.4 213.4 288.2 ;
      RECT  214.2 277.4 215.0 288.2 ;
      RECT  217.8 277.4 218.6 288.2 ;
      RECT  219.4 277.4 220.2 288.2 ;
      RECT  216.0 288.2 216.8 287.4 ;
      RECT  212.6 298.2 213.4 287.4 ;
      RECT  214.2 298.2 215.0 287.4 ;
      RECT  217.8 298.2 218.6 287.4 ;
      RECT  219.4 298.2 220.2 287.4 ;
      RECT  216.0 308.2 216.8 309.0 ;
      RECT  212.6 298.2 213.4 309.0 ;
      RECT  214.2 298.2 215.0 309.0 ;
      RECT  217.8 298.2 218.6 309.0 ;
      RECT  219.4 298.2 220.2 309.0 ;
      RECT  216.0 309.0 216.8 308.2 ;
      RECT  212.6 319.0 213.4 308.2 ;
      RECT  214.2 319.0 215.0 308.2 ;
      RECT  217.8 319.0 218.6 308.2 ;
      RECT  219.4 319.0 220.2 308.2 ;
      RECT  216.0 329.0 216.8 329.8 ;
      RECT  212.6 319.0 213.4 329.8 ;
      RECT  214.2 319.0 215.0 329.8 ;
      RECT  217.8 319.0 218.6 329.8 ;
      RECT  219.4 319.0 220.2 329.8 ;
      RECT  216.0 329.8 216.8 329.0 ;
      RECT  212.6 339.8 213.4 329.0 ;
      RECT  214.2 339.8 215.0 329.0 ;
      RECT  217.8 339.8 218.6 329.0 ;
      RECT  219.4 339.8 220.2 329.0 ;
      RECT  216.0 349.8 216.8 350.6 ;
      RECT  212.6 339.8 213.4 350.6 ;
      RECT  214.2 339.8 215.0 350.6 ;
      RECT  217.8 339.8 218.6 350.6 ;
      RECT  219.4 339.8 220.2 350.6 ;
      RECT  216.0 350.6 216.8 349.8 ;
      RECT  212.6 360.6 213.4 349.8 ;
      RECT  214.2 360.6 215.0 349.8 ;
      RECT  217.8 360.6 218.6 349.8 ;
      RECT  219.4 360.6 220.2 349.8 ;
      RECT  216.0 370.6 216.8 371.4 ;
      RECT  212.6 360.6 213.4 371.4 ;
      RECT  214.2 360.6 215.0 371.4 ;
      RECT  217.8 360.6 218.6 371.4 ;
      RECT  219.4 360.6 220.2 371.4 ;
      RECT  216.0 183.4 216.8 184.2 ;
      RECT  212.6 178.4 213.4 179.2 ;
      RECT  219.4 178.4 220.2 179.2 ;
      RECT  216.0 183.4 216.8 184.2 ;
      RECT  212.6 188.4 213.4 189.2 ;
      RECT  219.4 188.4 220.2 189.2 ;
      RECT  216.0 204.2 216.8 205.0 ;
      RECT  212.6 199.2 213.4 200.0 ;
      RECT  219.4 199.2 220.2 200.0 ;
      RECT  216.0 204.2 216.8 205.0 ;
      RECT  212.6 209.2 213.4 210.0 ;
      RECT  219.4 209.2 220.2 210.0 ;
      RECT  216.0 225.0 216.8 225.8 ;
      RECT  212.6 220.0 213.4 220.8 ;
      RECT  219.4 220.0 220.2 220.8 ;
      RECT  216.0 225.0 216.8 225.8 ;
      RECT  212.6 230.0 213.4 230.8 ;
      RECT  219.4 230.0 220.2 230.8 ;
      RECT  216.0 245.8 216.8 246.6 ;
      RECT  212.6 240.8 213.4 241.6 ;
      RECT  219.4 240.8 220.2 241.6 ;
      RECT  216.0 245.8 216.8 246.6 ;
      RECT  212.6 250.8 213.4 251.6 ;
      RECT  219.4 250.8 220.2 251.6 ;
      RECT  216.0 266.6 216.8 267.4 ;
      RECT  212.6 261.6 213.4 262.4 ;
      RECT  219.4 261.6 220.2 262.4 ;
      RECT  216.0 266.6 216.8 267.4 ;
      RECT  212.6 271.6 213.4 272.4 ;
      RECT  219.4 271.6 220.2 272.4 ;
      RECT  216.0 287.4 216.8 288.2 ;
      RECT  212.6 282.4 213.4 283.2 ;
      RECT  219.4 282.4 220.2 283.2 ;
      RECT  216.0 287.4 216.8 288.2 ;
      RECT  212.6 292.4 213.4 293.2 ;
      RECT  219.4 292.4 220.2 293.2 ;
      RECT  216.0 308.2 216.8 309.0 ;
      RECT  212.6 303.2 213.4 304.0 ;
      RECT  219.4 303.2 220.2 304.0 ;
      RECT  216.0 308.2 216.8 309.0 ;
      RECT  212.6 313.2 213.4 314.0 ;
      RECT  219.4 313.2 220.2 314.0 ;
      RECT  216.0 329.0 216.8 329.8 ;
      RECT  212.6 324.0 213.4 324.8 ;
      RECT  219.4 324.0 220.2 324.8 ;
      RECT  216.0 329.0 216.8 329.8 ;
      RECT  212.6 334.0 213.4 334.8 ;
      RECT  219.4 334.0 220.2 334.8 ;
      RECT  216.0 349.8 216.8 350.6 ;
      RECT  212.6 344.8 213.4 345.6 ;
      RECT  219.4 344.8 220.2 345.6 ;
      RECT  216.0 349.8 216.8 350.6 ;
      RECT  212.6 354.8 213.4 355.6 ;
      RECT  219.4 354.8 220.2 355.6 ;
      RECT  216.0 370.6 216.8 371.4 ;
      RECT  212.6 365.6 213.4 366.4 ;
      RECT  219.4 365.6 220.2 366.4 ;
      RECT  214.2 173.4 215.0 371.0 ;
      RECT  217.8 173.4 218.6 371.0 ;
      RECT  195.6 266.6 196.4 267.4 ;
      RECT  195.6 183.4 196.4 184.2 ;
      RECT  195.6 287.4 196.4 288.2 ;
      RECT  195.6 225.0 196.4 225.8 ;
      RECT  195.6 370.6 196.4 371.4 ;
      RECT  195.6 245.8 196.4 246.6 ;
      RECT  195.6 349.8 196.4 350.6 ;
      RECT  195.6 204.2 196.4 205.0 ;
      RECT  195.6 329.0 196.4 329.8 ;
      RECT  195.6 308.2 196.4 309.0 ;
      RECT  199.0 261.6 199.8 262.4 ;
      RECT  192.2 250.8 193.0 251.6 ;
      RECT  192.2 261.6 193.0 262.4 ;
      RECT  192.2 230.0 193.0 230.8 ;
      RECT  199.0 282.4 199.8 283.2 ;
      RECT  199.0 365.6 199.8 366.4 ;
      RECT  199.0 188.4 199.8 189.2 ;
      RECT  192.2 209.2 193.0 210.0 ;
      RECT  192.2 365.6 193.0 366.4 ;
      RECT  192.2 313.2 193.0 314.0 ;
      RECT  199.0 271.6 199.8 272.4 ;
      RECT  199.0 292.4 199.8 293.2 ;
      RECT  199.0 344.8 199.8 345.6 ;
      RECT  199.0 199.2 199.8 200.0 ;
      RECT  199.0 250.8 199.8 251.6 ;
      RECT  192.2 271.6 193.0 272.4 ;
      RECT  199.0 313.2 199.8 314.0 ;
      RECT  192.2 240.8 193.0 241.6 ;
      RECT  192.2 178.4 193.0 179.2 ;
      RECT  192.2 303.2 193.0 304.0 ;
      RECT  199.0 354.8 199.8 355.6 ;
      RECT  192.2 220.0 193.0 220.8 ;
      RECT  192.2 282.4 193.0 283.2 ;
      RECT  199.0 303.2 199.8 304.0 ;
      RECT  199.0 178.4 199.8 179.2 ;
      RECT  199.0 240.8 199.8 241.6 ;
      RECT  199.0 220.0 199.8 220.8 ;
      RECT  192.2 334.0 193.0 334.8 ;
      RECT  199.0 230.0 199.8 230.8 ;
      RECT  192.2 188.4 193.0 189.2 ;
      RECT  192.2 292.4 193.0 293.2 ;
      RECT  192.2 324.0 193.0 324.8 ;
      RECT  199.0 334.0 199.8 334.8 ;
      RECT  192.2 199.2 193.0 200.0 ;
      RECT  199.0 324.0 199.8 324.8 ;
      RECT  192.2 344.8 193.0 345.6 ;
      RECT  199.0 209.2 199.8 210.0 ;
      RECT  192.2 354.8 193.0 355.6 ;
      RECT  200.6 173.4 201.4 371.0 ;
      RECT  204.2 173.4 205.0 371.0 ;
      RECT  207.4 173.4 208.2 371.0 ;
      RECT  211.0 173.4 211.8 371.0 ;
      RECT  193.8 173.4 194.6 371.0 ;
      RECT  197.4 173.4 198.2 371.0 ;
      RECT  201.5 118.7 202.1 118.1 ;
      RECT  201.5 140.9 202.1 118.4 ;
      RECT  201.5 118.4 202.1 114.6 ;
      RECT  203.5 117.3 204.1 116.7 ;
      RECT  203.5 140.9 204.1 117.0 ;
      RECT  203.5 117.0 204.1 113.1 ;
      RECT  208.3 118.7 208.9 118.1 ;
      RECT  208.3 140.9 208.9 118.4 ;
      RECT  208.3 118.4 208.9 114.6 ;
      RECT  210.3 117.3 210.9 116.7 ;
      RECT  210.3 140.9 210.9 117.0 ;
      RECT  210.3 117.0 210.9 113.1 ;
      RECT  200.7 155.5 202.1 154.9 ;
      RECT  200.7 162.9 201.3 155.2 ;
      RECT  201.5 155.2 202.1 140.9 ;
      RECT  203.5 154.1 204.9 153.5 ;
      RECT  204.3 162.9 204.9 153.8 ;
      RECT  203.5 153.8 204.1 140.9 ;
      RECT  207.5 155.5 208.9 154.9 ;
      RECT  207.5 162.9 208.1 155.2 ;
      RECT  208.3 155.2 208.9 140.9 ;
      RECT  210.3 154.1 211.7 153.5 ;
      RECT  211.1 162.9 211.7 153.8 ;
      RECT  210.3 153.8 210.9 140.9 ;
      RECT  195.4 163.0 196.2 163.8 ;
      RECT  195.4 163.0 196.2 163.8 ;
      RECT  193.8 163.0 194.6 163.8 ;
      RECT  193.8 158.2 194.6 159.0 ;
      RECT  197.4 163.0 198.2 163.8 ;
      RECT  197.4 158.2 198.2 159.0 ;
      RECT  193.9 156.6 194.5 169.2 ;
      RECT  197.5 156.6 198.1 169.2 ;
      RECT  202.2 163.0 203.0 163.8 ;
      RECT  202.2 163.0 203.0 163.8 ;
      RECT  200.6 163.0 201.4 163.8 ;
      RECT  200.6 158.2 201.4 159.0 ;
      RECT  204.2 163.0 205.0 163.8 ;
      RECT  204.2 158.2 205.0 159.0 ;
      RECT  200.7 156.6 201.3 169.2 ;
      RECT  204.3 156.6 204.9 169.2 ;
      RECT  209.0 163.0 209.8 163.8 ;
      RECT  209.0 163.0 209.8 163.8 ;
      RECT  207.4 163.0 208.2 163.8 ;
      RECT  207.4 158.2 208.2 159.0 ;
      RECT  211.0 163.0 211.8 163.8 ;
      RECT  211.0 158.2 211.8 159.0 ;
      RECT  207.5 156.6 208.1 169.2 ;
      RECT  211.1 156.6 211.7 169.2 ;
      RECT  193.9 156.6 194.5 169.2 ;
      RECT  197.5 156.6 198.1 169.2 ;
      RECT  200.7 156.6 201.3 169.2 ;
      RECT  204.3 156.6 204.9 169.2 ;
      RECT  207.5 156.6 208.1 169.2 ;
      RECT  211.1 156.6 211.7 169.2 ;
      RECT  201.4 129.4 202.2 152.4 ;
      RECT  203.4 129.4 204.2 152.4 ;
      RECT  203.4 119.8 204.2 128.6 ;
      RECT  200.0 119.8 200.8 122.8 ;
      RECT  205.8 145.6 206.6 147.2 ;
      RECT  203.4 128.6 204.6 129.4 ;
      RECT  201.4 119.8 202.2 128.6 ;
      RECT  204.8 132.2 205.6 133.8 ;
      RECT  201.4 128.6 202.8 129.4 ;
      RECT  208.2 129.4 209.0 152.4 ;
      RECT  210.2 129.4 211.0 152.4 ;
      RECT  210.2 119.8 211.0 128.6 ;
      RECT  206.8 119.8 207.6 122.8 ;
      RECT  212.6 145.6 213.4 147.2 ;
      RECT  210.2 128.6 211.4 129.4 ;
      RECT  208.2 119.8 209.0 128.6 ;
      RECT  211.6 132.2 212.4 133.8 ;
      RECT  208.2 128.6 209.6 129.4 ;
      RECT  205.8 146.0 206.6 146.8 ;
      RECT  204.8 132.6 205.6 133.4 ;
      RECT  212.6 146.0 213.4 146.8 ;
      RECT  211.6 132.6 212.4 133.4 ;
      RECT  200.0 119.8 200.8 122.8 ;
      RECT  201.4 129.4 202.2 152.4 ;
      RECT  203.4 129.4 204.2 152.4 ;
      RECT  206.8 119.8 207.6 122.8 ;
      RECT  208.2 129.4 209.0 152.4 ;
      RECT  210.2 129.4 211.0 152.4 ;
      RECT  203.4 110.6 204.2 115.6 ;
      RECT  204.6 92.2 205.4 93.0 ;
      RECT  203.2 87.8 204.0 88.6 ;
      RECT  201.4 113.6 202.2 115.6 ;
      RECT  201.8 106.8 202.6 107.6 ;
      RECT  202.6 98.6 203.4 99.4 ;
      RECT  202.4 75.0 203.2 77.0 ;
      RECT  203.2 81.2 204.0 82.0 ;
      RECT  210.2 110.6 211.0 115.6 ;
      RECT  211.4 92.2 212.2 93.0 ;
      RECT  210.0 87.8 210.8 88.6 ;
      RECT  208.2 113.6 209.0 115.6 ;
      RECT  208.6 106.8 209.4 107.6 ;
      RECT  209.4 98.6 210.2 99.4 ;
      RECT  209.2 75.0 210.0 77.0 ;
      RECT  210.0 81.2 210.8 82.0 ;
      RECT  203.2 81.2 204.0 82.0 ;
      RECT  202.6 98.6 203.4 99.4 ;
      RECT  203.2 87.8 204.0 88.6 ;
      RECT  204.6 92.2 205.4 93.0 ;
      RECT  201.8 106.8 202.6 107.6 ;
      RECT  210.0 81.2 210.8 82.0 ;
      RECT  209.4 98.6 210.2 99.4 ;
      RECT  210.0 87.8 210.8 88.6 ;
      RECT  211.4 92.2 212.2 93.0 ;
      RECT  208.6 106.8 209.4 107.6 ;
      RECT  202.4 75.0 203.2 77.0 ;
      RECT  209.2 75.0 210.0 77.0 ;
      RECT  201.4 113.6 202.2 115.6 ;
      RECT  203.4 110.6 204.2 115.6 ;
      RECT  208.2 113.6 209.0 115.6 ;
      RECT  210.2 110.6 211.0 115.6 ;
      RECT  193.9 169.2 194.5 156.6 ;
      RECT  197.5 169.2 198.1 156.6 ;
      RECT  200.7 169.2 201.3 156.6 ;
      RECT  204.3 169.2 204.9 156.6 ;
      RECT  207.5 169.2 208.1 156.6 ;
      RECT  211.1 169.2 211.7 156.6 ;
      RECT  200.0 122.8 200.8 119.8 ;
      RECT  206.8 122.8 207.6 119.8 ;
      RECT  202.4 77.0 203.2 75.0 ;
      RECT  209.2 77.0 210.0 75.0 ;
      RECT  126.9 199.9 127.5 204.8 ;
      RECT  126.9 210.7 127.5 215.6 ;
      RECT  126.9 220.7 127.5 225.6 ;
      RECT  126.9 231.5 127.5 236.4 ;
      RECT  126.9 241.5 127.5 246.4 ;
      RECT  126.9 252.3 127.5 257.2 ;
      RECT  126.9 262.3 127.5 267.2 ;
      RECT  126.9 273.1 127.5 278.0 ;
      RECT  108.5 195.8 109.1 236.2 ;
      RECT  109.9 195.8 110.5 236.2 ;
      RECT  111.3 195.8 111.9 236.2 ;
      RECT  112.7 195.8 113.3 236.2 ;
      RECT  120.0 203.0 120.6 203.6 ;
      RECT  120.0 196.0 120.6 196.6 ;
      RECT  117.3 203.0 120.3 203.6 ;
      RECT  120.0 199.4 120.6 203.3 ;
      RECT  120.0 196.3 120.6 199.4 ;
      RECT  118.9 196.0 120.3 196.6 ;
      RECT  116.9 202.9 117.7 203.7 ;
      RECT  118.5 195.9 119.3 196.7 ;
      RECT  119.9 199.0 120.7 199.8 ;
      RECT  120.0 207.0 120.6 206.4 ;
      RECT  120.0 214.0 120.6 213.4 ;
      RECT  117.3 207.0 120.3 206.4 ;
      RECT  120.0 210.6 120.6 206.7 ;
      RECT  120.0 213.7 120.6 210.6 ;
      RECT  118.9 214.0 120.3 213.4 ;
      RECT  116.9 207.1 117.7 206.3 ;
      RECT  118.5 214.1 119.3 213.3 ;
      RECT  119.9 211.0 120.7 210.2 ;
      RECT  120.0 223.8 120.6 224.4 ;
      RECT  120.0 216.8 120.6 217.4 ;
      RECT  117.3 223.8 120.3 224.4 ;
      RECT  120.0 220.2 120.6 224.1 ;
      RECT  120.0 217.1 120.6 220.2 ;
      RECT  118.9 216.8 120.3 217.4 ;
      RECT  116.9 223.7 117.7 224.5 ;
      RECT  118.5 216.7 119.3 217.5 ;
      RECT  119.9 219.8 120.7 220.6 ;
      RECT  120.0 227.8 120.6 227.2 ;
      RECT  120.0 234.8 120.6 234.2 ;
      RECT  117.3 227.8 120.3 227.2 ;
      RECT  120.0 231.4 120.6 227.5 ;
      RECT  120.0 234.5 120.6 231.4 ;
      RECT  118.9 234.8 120.3 234.2 ;
      RECT  116.9 227.9 117.7 227.1 ;
      RECT  118.5 234.9 119.3 234.1 ;
      RECT  119.9 231.8 120.7 231.0 ;
      RECT  108.4 202.8 109.2 203.6 ;
      RECT  96.7 199.2 97.5 200.0 ;
      RECT  109.8 213.2 110.6 214.0 ;
      RECT  98.1 210.0 98.9 210.8 ;
      RECT  96.7 216.4 97.5 217.2 ;
      RECT  111.2 216.4 112.0 217.2 ;
      RECT  98.1 226.8 98.9 227.6 ;
      RECT  112.6 226.8 113.4 227.6 ;
      RECT  108.4 199.0 109.2 199.8 ;
      RECT  109.8 197.6 110.6 198.4 ;
      RECT  111.2 210.2 112.0 211.0 ;
      RECT  109.8 211.6 110.6 212.4 ;
      RECT  108.4 219.8 109.2 220.6 ;
      RECT  112.6 218.4 113.4 219.2 ;
      RECT  111.2 231.0 112.0 231.8 ;
      RECT  112.6 232.4 113.4 233.2 ;
      RECT  105.3 204.6 106.1 205.4 ;
      RECT  105.3 204.6 106.1 205.4 ;
      RECT  122.7 204.6 123.5 205.4 ;
      RECT  122.7 204.6 123.5 205.4 ;
      RECT  105.3 194.2 106.1 195.0 ;
      RECT  105.3 194.2 106.1 195.0 ;
      RECT  122.7 194.2 123.5 195.0 ;
      RECT  122.7 194.2 123.5 195.0 ;
      RECT  105.3 204.6 106.1 205.4 ;
      RECT  105.3 204.6 106.1 205.4 ;
      RECT  122.7 204.6 123.5 205.4 ;
      RECT  122.7 204.6 123.5 205.4 ;
      RECT  105.3 215.0 106.1 215.8 ;
      RECT  105.3 215.0 106.1 215.8 ;
      RECT  122.7 215.0 123.5 215.8 ;
      RECT  122.7 215.0 123.5 215.8 ;
      RECT  105.3 225.4 106.1 226.2 ;
      RECT  105.3 225.4 106.1 226.2 ;
      RECT  122.7 225.4 123.5 226.2 ;
      RECT  122.7 225.4 123.5 226.2 ;
      RECT  105.3 215.0 106.1 215.8 ;
      RECT  105.3 215.0 106.1 215.8 ;
      RECT  122.7 215.0 123.5 215.8 ;
      RECT  122.7 215.0 123.5 215.8 ;
      RECT  105.3 225.4 106.1 226.2 ;
      RECT  105.3 225.4 106.1 226.2 ;
      RECT  122.7 225.4 123.5 226.2 ;
      RECT  122.7 225.4 123.5 226.2 ;
      RECT  105.3 235.8 106.1 236.6 ;
      RECT  105.3 235.8 106.1 236.6 ;
      RECT  122.7 235.8 123.5 236.6 ;
      RECT  122.7 235.8 123.5 236.6 ;
      RECT  96.8 195.8 97.4 236.2 ;
      RECT  98.2 195.8 98.8 236.2 ;
      RECT  108.5 237.4 109.1 277.8 ;
      RECT  109.9 237.4 110.5 277.8 ;
      RECT  111.3 237.4 111.9 277.8 ;
      RECT  112.7 237.4 113.3 277.8 ;
      RECT  120.0 244.6 120.6 245.2 ;
      RECT  120.0 237.6 120.6 238.2 ;
      RECT  117.3 244.6 120.3 245.2 ;
      RECT  120.0 241.0 120.6 244.9 ;
      RECT  120.0 237.9 120.6 241.0 ;
      RECT  118.9 237.6 120.3 238.2 ;
      RECT  116.9 244.5 117.7 245.3 ;
      RECT  118.5 237.5 119.3 238.3 ;
      RECT  119.9 240.6 120.7 241.4 ;
      RECT  120.0 248.6 120.6 248.0 ;
      RECT  120.0 255.6 120.6 255.0 ;
      RECT  117.3 248.6 120.3 248.0 ;
      RECT  120.0 252.2 120.6 248.3 ;
      RECT  120.0 255.3 120.6 252.2 ;
      RECT  118.9 255.6 120.3 255.0 ;
      RECT  116.9 248.7 117.7 247.9 ;
      RECT  118.5 255.7 119.3 254.9 ;
      RECT  119.9 252.6 120.7 251.8 ;
      RECT  120.0 265.4 120.6 266.0 ;
      RECT  120.0 258.4 120.6 259.0 ;
      RECT  117.3 265.4 120.3 266.0 ;
      RECT  120.0 261.8 120.6 265.7 ;
      RECT  120.0 258.7 120.6 261.8 ;
      RECT  118.9 258.4 120.3 259.0 ;
      RECT  116.9 265.3 117.7 266.1 ;
      RECT  118.5 258.3 119.3 259.1 ;
      RECT  119.9 261.4 120.7 262.2 ;
      RECT  120.0 269.4 120.6 268.8 ;
      RECT  120.0 276.4 120.6 275.8 ;
      RECT  117.3 269.4 120.3 268.8 ;
      RECT  120.0 273.0 120.6 269.1 ;
      RECT  120.0 276.1 120.6 273.0 ;
      RECT  118.9 276.4 120.3 275.8 ;
      RECT  116.9 269.5 117.7 268.7 ;
      RECT  118.5 276.5 119.3 275.7 ;
      RECT  119.9 273.4 120.7 272.6 ;
      RECT  108.4 244.4 109.2 245.2 ;
      RECT  96.7 240.8 97.5 241.6 ;
      RECT  109.8 254.8 110.6 255.6 ;
      RECT  98.1 251.6 98.9 252.4 ;
      RECT  96.7 258.0 97.5 258.8 ;
      RECT  111.2 258.0 112.0 258.8 ;
      RECT  98.1 268.4 98.9 269.2 ;
      RECT  112.6 268.4 113.4 269.2 ;
      RECT  108.4 240.6 109.2 241.4 ;
      RECT  109.8 239.2 110.6 240.0 ;
      RECT  111.2 251.8 112.0 252.6 ;
      RECT  109.8 253.2 110.6 254.0 ;
      RECT  108.4 261.4 109.2 262.2 ;
      RECT  112.6 260.0 113.4 260.8 ;
      RECT  111.2 272.6 112.0 273.4 ;
      RECT  112.6 274.0 113.4 274.8 ;
      RECT  105.3 246.2 106.1 247.0 ;
      RECT  105.3 246.2 106.1 247.0 ;
      RECT  122.7 246.2 123.5 247.0 ;
      RECT  122.7 246.2 123.5 247.0 ;
      RECT  105.3 235.8 106.1 236.6 ;
      RECT  105.3 235.8 106.1 236.6 ;
      RECT  122.7 235.8 123.5 236.6 ;
      RECT  122.7 235.8 123.5 236.6 ;
      RECT  105.3 246.2 106.1 247.0 ;
      RECT  105.3 246.2 106.1 247.0 ;
      RECT  122.7 246.2 123.5 247.0 ;
      RECT  122.7 246.2 123.5 247.0 ;
      RECT  105.3 256.6 106.1 257.4 ;
      RECT  105.3 256.6 106.1 257.4 ;
      RECT  122.7 256.6 123.5 257.4 ;
      RECT  122.7 256.6 123.5 257.4 ;
      RECT  105.3 267.0 106.1 267.8 ;
      RECT  105.3 267.0 106.1 267.8 ;
      RECT  122.7 267.0 123.5 267.8 ;
      RECT  122.7 267.0 123.5 267.8 ;
      RECT  105.3 256.6 106.1 257.4 ;
      RECT  105.3 256.6 106.1 257.4 ;
      RECT  122.7 256.6 123.5 257.4 ;
      RECT  122.7 256.6 123.5 257.4 ;
      RECT  105.3 267.0 106.1 267.8 ;
      RECT  105.3 267.0 106.1 267.8 ;
      RECT  122.7 267.0 123.5 267.8 ;
      RECT  122.7 267.0 123.5 267.8 ;
      RECT  105.3 277.4 106.1 278.2 ;
      RECT  105.3 277.4 106.1 278.2 ;
      RECT  122.7 277.4 123.5 278.2 ;
      RECT  122.7 277.4 123.5 278.2 ;
      RECT  96.8 237.4 97.4 277.8 ;
      RECT  98.2 237.4 98.8 277.8 ;
      RECT  147.2 203.0 147.8 203.6 ;
      RECT  147.2 196.0 147.8 196.6 ;
      RECT  144.5 203.0 147.5 203.6 ;
      RECT  147.2 199.4 147.8 203.3 ;
      RECT  147.2 196.3 147.8 199.4 ;
      RECT  146.1 196.0 147.5 196.6 ;
      RECT  144.1 202.9 144.9 203.7 ;
      RECT  145.7 195.9 146.5 196.7 ;
      RECT  147.1 199.0 147.9 199.8 ;
      RECT  147.2 207.0 147.8 206.4 ;
      RECT  147.2 214.0 147.8 213.4 ;
      RECT  144.5 207.0 147.5 206.4 ;
      RECT  147.2 210.6 147.8 206.7 ;
      RECT  147.2 213.7 147.8 210.6 ;
      RECT  146.1 214.0 147.5 213.4 ;
      RECT  144.1 207.1 144.9 206.3 ;
      RECT  145.7 214.1 146.5 213.3 ;
      RECT  147.1 211.0 147.9 210.2 ;
      RECT  147.2 223.8 147.8 224.4 ;
      RECT  147.2 216.8 147.8 217.4 ;
      RECT  144.5 223.8 147.5 224.4 ;
      RECT  147.2 220.2 147.8 224.1 ;
      RECT  147.2 217.1 147.8 220.2 ;
      RECT  146.1 216.8 147.5 217.4 ;
      RECT  144.1 223.7 144.9 224.5 ;
      RECT  145.7 216.7 146.5 217.5 ;
      RECT  147.1 219.8 147.9 220.6 ;
      RECT  147.2 227.8 147.8 227.2 ;
      RECT  147.2 234.8 147.8 234.2 ;
      RECT  144.5 227.8 147.5 227.2 ;
      RECT  147.2 231.4 147.8 227.5 ;
      RECT  147.2 234.5 147.8 231.4 ;
      RECT  146.1 234.8 147.5 234.2 ;
      RECT  144.1 227.9 144.9 227.1 ;
      RECT  145.7 234.9 146.5 234.1 ;
      RECT  147.1 231.8 147.9 231.0 ;
      RECT  147.2 244.6 147.8 245.2 ;
      RECT  147.2 237.6 147.8 238.2 ;
      RECT  144.5 244.6 147.5 245.2 ;
      RECT  147.2 241.0 147.8 244.9 ;
      RECT  147.2 237.9 147.8 241.0 ;
      RECT  146.1 237.6 147.5 238.2 ;
      RECT  144.1 244.5 144.9 245.3 ;
      RECT  145.7 237.5 146.5 238.3 ;
      RECT  147.1 240.6 147.9 241.4 ;
      RECT  147.2 248.6 147.8 248.0 ;
      RECT  147.2 255.6 147.8 255.0 ;
      RECT  144.5 248.6 147.5 248.0 ;
      RECT  147.2 252.2 147.8 248.3 ;
      RECT  147.2 255.3 147.8 252.2 ;
      RECT  146.1 255.6 147.5 255.0 ;
      RECT  144.1 248.7 144.9 247.9 ;
      RECT  145.7 255.7 146.5 254.9 ;
      RECT  147.1 252.6 147.9 251.8 ;
      RECT  147.2 265.4 147.8 266.0 ;
      RECT  147.2 258.4 147.8 259.0 ;
      RECT  144.5 265.4 147.5 266.0 ;
      RECT  147.2 261.8 147.8 265.7 ;
      RECT  147.2 258.7 147.8 261.8 ;
      RECT  146.1 258.4 147.5 259.0 ;
      RECT  144.1 265.3 144.9 266.1 ;
      RECT  145.7 258.3 146.5 259.1 ;
      RECT  147.1 261.4 147.9 262.2 ;
      RECT  147.2 269.4 147.8 268.8 ;
      RECT  147.2 276.4 147.8 275.8 ;
      RECT  144.5 269.4 147.5 268.8 ;
      RECT  147.2 273.0 147.8 269.1 ;
      RECT  147.2 276.1 147.8 273.0 ;
      RECT  146.1 276.4 147.5 275.8 ;
      RECT  144.1 269.5 144.9 268.7 ;
      RECT  145.7 276.5 146.5 275.7 ;
      RECT  147.1 273.4 147.9 272.6 ;
      RECT  147.2 286.2 147.8 286.8 ;
      RECT  147.2 279.2 147.8 279.8 ;
      RECT  144.5 286.2 147.5 286.8 ;
      RECT  147.2 282.6 147.8 286.5 ;
      RECT  147.2 279.5 147.8 282.6 ;
      RECT  146.1 279.2 147.5 279.8 ;
      RECT  144.1 286.1 144.9 286.9 ;
      RECT  145.7 279.1 146.5 279.9 ;
      RECT  147.1 282.2 147.9 283.0 ;
      RECT  147.2 290.2 147.8 289.6 ;
      RECT  147.2 297.2 147.8 296.6 ;
      RECT  144.5 290.2 147.5 289.6 ;
      RECT  147.2 293.8 147.8 289.9 ;
      RECT  147.2 296.9 147.8 293.8 ;
      RECT  146.1 297.2 147.5 296.6 ;
      RECT  144.1 290.3 144.9 289.5 ;
      RECT  145.7 297.3 146.5 296.5 ;
      RECT  147.1 294.2 147.9 293.4 ;
      RECT  147.2 307.0 147.8 307.6 ;
      RECT  147.2 300.0 147.8 300.6 ;
      RECT  144.5 307.0 147.5 307.6 ;
      RECT  147.2 303.4 147.8 307.3 ;
      RECT  147.2 300.3 147.8 303.4 ;
      RECT  146.1 300.0 147.5 300.6 ;
      RECT  144.1 306.9 144.9 307.7 ;
      RECT  145.7 299.9 146.5 300.7 ;
      RECT  147.1 303.0 147.9 303.8 ;
      RECT  147.2 311.0 147.8 310.4 ;
      RECT  147.2 318.0 147.8 317.4 ;
      RECT  144.5 311.0 147.5 310.4 ;
      RECT  147.2 314.6 147.8 310.7 ;
      RECT  147.2 317.7 147.8 314.6 ;
      RECT  146.1 318.0 147.5 317.4 ;
      RECT  144.1 311.1 144.9 310.3 ;
      RECT  145.7 318.1 146.5 317.3 ;
      RECT  147.1 315.0 147.9 314.2 ;
      RECT  147.2 327.8 147.8 328.4 ;
      RECT  147.2 320.8 147.8 321.4 ;
      RECT  144.5 327.8 147.5 328.4 ;
      RECT  147.2 324.2 147.8 328.1 ;
      RECT  147.2 321.1 147.8 324.2 ;
      RECT  146.1 320.8 147.5 321.4 ;
      RECT  144.1 327.7 144.9 328.5 ;
      RECT  145.7 320.7 146.5 321.5 ;
      RECT  147.1 323.8 147.9 324.6 ;
      RECT  147.2 331.8 147.8 331.2 ;
      RECT  147.2 338.8 147.8 338.2 ;
      RECT  144.5 331.8 147.5 331.2 ;
      RECT  147.2 335.4 147.8 331.5 ;
      RECT  147.2 338.5 147.8 335.4 ;
      RECT  146.1 338.8 147.5 338.2 ;
      RECT  144.1 331.9 144.9 331.1 ;
      RECT  145.7 338.9 146.5 338.1 ;
      RECT  147.1 335.8 147.9 335.0 ;
      RECT  147.2 348.6 147.8 349.2 ;
      RECT  147.2 341.6 147.8 342.2 ;
      RECT  144.5 348.6 147.5 349.2 ;
      RECT  147.2 345.0 147.8 348.9 ;
      RECT  147.2 341.9 147.8 345.0 ;
      RECT  146.1 341.6 147.5 342.2 ;
      RECT  144.1 348.5 144.9 349.3 ;
      RECT  145.7 341.5 146.5 342.3 ;
      RECT  147.1 344.6 147.9 345.4 ;
      RECT  147.2 352.6 147.8 352.0 ;
      RECT  147.2 359.6 147.8 359.0 ;
      RECT  144.5 352.6 147.5 352.0 ;
      RECT  147.2 356.2 147.8 352.3 ;
      RECT  147.2 359.3 147.8 356.2 ;
      RECT  146.1 359.6 147.5 359.0 ;
      RECT  144.1 352.7 144.9 351.9 ;
      RECT  145.7 359.7 146.5 358.9 ;
      RECT  147.1 356.6 147.9 355.8 ;
      RECT  96.7 205.8 97.5 206.6 ;
      RECT  89.4 205.8 90.2 206.6 ;
      RECT  98.1 216.2 98.9 217.0 ;
      RECT  90.8 216.2 91.6 217.0 ;
      RECT  96.7 247.4 97.5 248.2 ;
      RECT  92.2 247.4 93.0 248.2 ;
      RECT  98.1 257.8 98.9 258.6 ;
      RECT  93.6 257.8 94.4 258.6 ;
      RECT  126.8 199.2 127.6 200.0 ;
      RECT  126.8 204.4 127.6 205.2 ;
      RECT  130.3 204.4 131.1 205.2 ;
      RECT  126.8 210.0 127.6 210.8 ;
      RECT  126.8 215.2 127.6 216.0 ;
      RECT  131.7 215.2 132.5 216.0 ;
      RECT  126.8 220.0 127.6 220.8 ;
      RECT  126.8 225.2 127.6 226.0 ;
      RECT  133.1 225.2 133.9 226.0 ;
      RECT  126.8 230.8 127.6 231.6 ;
      RECT  126.8 236.0 127.6 236.8 ;
      RECT  134.5 236.0 135.3 236.8 ;
      RECT  126.8 240.8 127.6 241.6 ;
      RECT  126.8 246.0 127.6 246.8 ;
      RECT  135.9 246.0 136.7 246.8 ;
      RECT  126.8 251.6 127.6 252.4 ;
      RECT  126.8 256.8 127.6 257.6 ;
      RECT  137.3 256.8 138.1 257.6 ;
      RECT  126.8 261.6 127.6 262.4 ;
      RECT  126.8 266.8 127.6 267.6 ;
      RECT  138.7 266.8 139.5 267.6 ;
      RECT  126.8 272.4 127.6 273.2 ;
      RECT  126.8 277.6 127.6 278.4 ;
      RECT  140.1 277.6 140.9 278.4 ;
      RECT  130.3 199.0 131.1 199.8 ;
      RECT  135.9 197.6 136.7 198.4 ;
      RECT  131.7 210.2 132.5 211.0 ;
      RECT  135.9 211.6 136.7 212.4 ;
      RECT  133.1 219.8 133.9 220.6 ;
      RECT  135.9 218.4 136.7 219.2 ;
      RECT  134.5 231.0 135.3 231.8 ;
      RECT  135.9 232.4 136.7 233.2 ;
      RECT  130.3 240.6 131.1 241.4 ;
      RECT  137.3 239.2 138.1 240.0 ;
      RECT  131.7 251.8 132.5 252.6 ;
      RECT  137.3 253.2 138.1 254.0 ;
      RECT  133.1 261.4 133.9 262.2 ;
      RECT  137.3 260.0 138.1 260.8 ;
      RECT  134.5 272.6 135.3 273.4 ;
      RECT  137.3 274.0 138.1 274.8 ;
      RECT  130.3 282.2 131.1 283.0 ;
      RECT  138.7 280.8 139.5 281.6 ;
      RECT  131.7 293.4 132.5 294.2 ;
      RECT  138.7 294.8 139.5 295.6 ;
      RECT  133.1 303.0 133.9 303.8 ;
      RECT  138.7 301.6 139.5 302.4 ;
      RECT  134.5 314.2 135.3 315.0 ;
      RECT  138.7 315.6 139.5 316.4 ;
      RECT  130.3 323.8 131.1 324.6 ;
      RECT  140.1 322.4 140.9 323.2 ;
      RECT  131.7 335.0 132.5 335.8 ;
      RECT  140.1 336.4 140.9 337.2 ;
      RECT  133.1 344.6 133.9 345.4 ;
      RECT  140.1 343.2 140.9 344.0 ;
      RECT  134.5 355.8 135.3 356.6 ;
      RECT  140.1 357.2 140.9 358.0 ;
      RECT  145.7 204.6 146.5 205.4 ;
      RECT  145.7 204.6 146.5 205.4 ;
      RECT  145.7 194.2 146.5 195.0 ;
      RECT  145.7 194.2 146.5 195.0 ;
      RECT  145.7 204.6 146.5 205.4 ;
      RECT  145.7 204.6 146.5 205.4 ;
      RECT  145.7 215.0 146.5 215.8 ;
      RECT  145.7 215.0 146.5 215.8 ;
      RECT  145.7 225.4 146.5 226.2 ;
      RECT  145.7 225.4 146.5 226.2 ;
      RECT  145.7 215.0 146.5 215.8 ;
      RECT  145.7 215.0 146.5 215.8 ;
      RECT  145.7 225.4 146.5 226.2 ;
      RECT  145.7 225.4 146.5 226.2 ;
      RECT  145.7 235.8 146.5 236.6 ;
      RECT  145.7 235.8 146.5 236.6 ;
      RECT  145.7 246.2 146.5 247.0 ;
      RECT  145.7 246.2 146.5 247.0 ;
      RECT  145.7 235.8 146.5 236.6 ;
      RECT  145.7 235.8 146.5 236.6 ;
      RECT  145.7 246.2 146.5 247.0 ;
      RECT  145.7 246.2 146.5 247.0 ;
      RECT  145.7 256.6 146.5 257.4 ;
      RECT  145.7 256.6 146.5 257.4 ;
      RECT  145.7 267.0 146.5 267.8 ;
      RECT  145.7 267.0 146.5 267.8 ;
      RECT  145.7 256.6 146.5 257.4 ;
      RECT  145.7 256.6 146.5 257.4 ;
      RECT  145.7 267.0 146.5 267.8 ;
      RECT  145.7 267.0 146.5 267.8 ;
      RECT  145.7 277.4 146.5 278.2 ;
      RECT  145.7 277.4 146.5 278.2 ;
      RECT  145.7 287.8 146.5 288.6 ;
      RECT  145.7 287.8 146.5 288.6 ;
      RECT  145.7 277.4 146.5 278.2 ;
      RECT  145.7 277.4 146.5 278.2 ;
      RECT  145.7 287.8 146.5 288.6 ;
      RECT  145.7 287.8 146.5 288.6 ;
      RECT  145.7 298.2 146.5 299.0 ;
      RECT  145.7 298.2 146.5 299.0 ;
      RECT  145.7 308.6 146.5 309.4 ;
      RECT  145.7 308.6 146.5 309.4 ;
      RECT  145.7 298.2 146.5 299.0 ;
      RECT  145.7 298.2 146.5 299.0 ;
      RECT  145.7 308.6 146.5 309.4 ;
      RECT  145.7 308.6 146.5 309.4 ;
      RECT  145.7 319.0 146.5 319.8 ;
      RECT  145.7 319.0 146.5 319.8 ;
      RECT  145.7 329.4 146.5 330.2 ;
      RECT  145.7 329.4 146.5 330.2 ;
      RECT  145.7 319.0 146.5 319.8 ;
      RECT  145.7 319.0 146.5 319.8 ;
      RECT  145.7 329.4 146.5 330.2 ;
      RECT  145.7 329.4 146.5 330.2 ;
      RECT  145.7 339.8 146.5 340.6 ;
      RECT  145.7 339.8 146.5 340.6 ;
      RECT  145.7 350.2 146.5 351.0 ;
      RECT  145.7 350.2 146.5 351.0 ;
      RECT  145.7 339.8 146.5 340.6 ;
      RECT  145.7 339.8 146.5 340.6 ;
      RECT  145.7 350.2 146.5 351.0 ;
      RECT  145.7 350.2 146.5 351.0 ;
      RECT  145.7 360.6 146.5 361.4 ;
      RECT  145.7 360.6 146.5 361.4 ;
      RECT  89.5 194.6 90.1 277.8 ;
      RECT  90.9 194.6 91.5 277.8 ;
      RECT  92.3 194.6 92.9 277.8 ;
      RECT  93.7 194.6 94.3 277.8 ;
      RECT  162.8 197.7 163.4 198.3 ;
      RECT  162.8 197.4 163.4 198.0 ;
      RECT  163.1 197.7 167.5 198.3 ;
      RECT  162.8 211.7 163.4 212.3 ;
      RECT  162.8 212.0 163.4 212.6 ;
      RECT  163.1 211.7 167.5 212.3 ;
      RECT  162.8 218.5 163.4 219.1 ;
      RECT  162.8 218.2 163.4 218.8 ;
      RECT  163.1 218.5 167.5 219.1 ;
      RECT  162.8 232.5 163.4 233.1 ;
      RECT  162.8 232.8 163.4 233.4 ;
      RECT  163.1 232.5 167.5 233.1 ;
      RECT  162.8 239.3 163.4 239.9 ;
      RECT  162.8 239.0 163.4 239.6 ;
      RECT  163.1 239.3 167.5 239.9 ;
      RECT  162.8 253.3 163.4 253.9 ;
      RECT  162.8 253.6 163.4 254.2 ;
      RECT  163.1 253.3 167.5 253.9 ;
      RECT  162.8 260.1 163.4 260.7 ;
      RECT  162.8 259.8 163.4 260.4 ;
      RECT  163.1 260.1 167.5 260.7 ;
      RECT  162.8 274.1 163.4 274.7 ;
      RECT  162.8 274.4 163.4 275.0 ;
      RECT  163.1 274.1 167.5 274.7 ;
      RECT  162.8 280.9 163.4 281.5 ;
      RECT  162.8 280.6 163.4 281.2 ;
      RECT  163.1 280.9 167.5 281.5 ;
      RECT  162.8 294.9 163.4 295.5 ;
      RECT  162.8 295.2 163.4 295.8 ;
      RECT  163.1 294.9 167.5 295.5 ;
      RECT  162.8 301.7 163.4 302.3 ;
      RECT  162.8 301.4 163.4 302.0 ;
      RECT  163.1 301.7 167.5 302.3 ;
      RECT  162.8 315.7 163.4 316.3 ;
      RECT  162.8 316.0 163.4 316.6 ;
      RECT  163.1 315.7 167.5 316.3 ;
      RECT  162.8 322.5 163.4 323.1 ;
      RECT  162.8 322.2 163.4 322.8 ;
      RECT  163.1 322.5 167.5 323.1 ;
      RECT  162.8 336.5 163.4 337.1 ;
      RECT  162.8 336.8 163.4 337.4 ;
      RECT  163.1 336.5 167.5 337.1 ;
      RECT  162.8 343.3 163.4 343.9 ;
      RECT  162.8 343.0 163.4 343.6 ;
      RECT  163.1 343.3 167.5 343.9 ;
      RECT  162.8 357.3 163.4 357.9 ;
      RECT  162.8 357.6 163.4 358.2 ;
      RECT  163.1 357.3 167.5 357.9 ;
      RECT  169.8 203.0 170.4 203.6 ;
      RECT  169.8 196.0 170.4 196.6 ;
      RECT  167.1 203.0 170.1 203.6 ;
      RECT  169.8 199.4 170.4 203.3 ;
      RECT  169.8 196.3 170.4 199.4 ;
      RECT  168.7 196.0 170.1 196.6 ;
      RECT  166.7 202.9 167.5 203.7 ;
      RECT  168.3 195.9 169.1 196.7 ;
      RECT  169.7 199.0 170.5 199.8 ;
      RECT  169.8 207.0 170.4 206.4 ;
      RECT  169.8 214.0 170.4 213.4 ;
      RECT  167.1 207.0 170.1 206.4 ;
      RECT  169.8 210.6 170.4 206.7 ;
      RECT  169.8 213.7 170.4 210.6 ;
      RECT  168.7 214.0 170.1 213.4 ;
      RECT  166.7 207.1 167.5 206.3 ;
      RECT  168.3 214.1 169.1 213.3 ;
      RECT  169.7 211.0 170.5 210.2 ;
      RECT  169.8 223.8 170.4 224.4 ;
      RECT  169.8 216.8 170.4 217.4 ;
      RECT  167.1 223.8 170.1 224.4 ;
      RECT  169.8 220.2 170.4 224.1 ;
      RECT  169.8 217.1 170.4 220.2 ;
      RECT  168.7 216.8 170.1 217.4 ;
      RECT  166.7 223.7 167.5 224.5 ;
      RECT  168.3 216.7 169.1 217.5 ;
      RECT  169.7 219.8 170.5 220.6 ;
      RECT  169.8 227.8 170.4 227.2 ;
      RECT  169.8 234.8 170.4 234.2 ;
      RECT  167.1 227.8 170.1 227.2 ;
      RECT  169.8 231.4 170.4 227.5 ;
      RECT  169.8 234.5 170.4 231.4 ;
      RECT  168.7 234.8 170.1 234.2 ;
      RECT  166.7 227.9 167.5 227.1 ;
      RECT  168.3 234.9 169.1 234.1 ;
      RECT  169.7 231.8 170.5 231.0 ;
      RECT  169.8 244.6 170.4 245.2 ;
      RECT  169.8 237.6 170.4 238.2 ;
      RECT  167.1 244.6 170.1 245.2 ;
      RECT  169.8 241.0 170.4 244.9 ;
      RECT  169.8 237.9 170.4 241.0 ;
      RECT  168.7 237.6 170.1 238.2 ;
      RECT  166.7 244.5 167.5 245.3 ;
      RECT  168.3 237.5 169.1 238.3 ;
      RECT  169.7 240.6 170.5 241.4 ;
      RECT  169.8 248.6 170.4 248.0 ;
      RECT  169.8 255.6 170.4 255.0 ;
      RECT  167.1 248.6 170.1 248.0 ;
      RECT  169.8 252.2 170.4 248.3 ;
      RECT  169.8 255.3 170.4 252.2 ;
      RECT  168.7 255.6 170.1 255.0 ;
      RECT  166.7 248.7 167.5 247.9 ;
      RECT  168.3 255.7 169.1 254.9 ;
      RECT  169.7 252.6 170.5 251.8 ;
      RECT  169.8 265.4 170.4 266.0 ;
      RECT  169.8 258.4 170.4 259.0 ;
      RECT  167.1 265.4 170.1 266.0 ;
      RECT  169.8 261.8 170.4 265.7 ;
      RECT  169.8 258.7 170.4 261.8 ;
      RECT  168.7 258.4 170.1 259.0 ;
      RECT  166.7 265.3 167.5 266.1 ;
      RECT  168.3 258.3 169.1 259.1 ;
      RECT  169.7 261.4 170.5 262.2 ;
      RECT  169.8 269.4 170.4 268.8 ;
      RECT  169.8 276.4 170.4 275.8 ;
      RECT  167.1 269.4 170.1 268.8 ;
      RECT  169.8 273.0 170.4 269.1 ;
      RECT  169.8 276.1 170.4 273.0 ;
      RECT  168.7 276.4 170.1 275.8 ;
      RECT  166.7 269.5 167.5 268.7 ;
      RECT  168.3 276.5 169.1 275.7 ;
      RECT  169.7 273.4 170.5 272.6 ;
      RECT  169.8 286.2 170.4 286.8 ;
      RECT  169.8 279.2 170.4 279.8 ;
      RECT  167.1 286.2 170.1 286.8 ;
      RECT  169.8 282.6 170.4 286.5 ;
      RECT  169.8 279.5 170.4 282.6 ;
      RECT  168.7 279.2 170.1 279.8 ;
      RECT  166.7 286.1 167.5 286.9 ;
      RECT  168.3 279.1 169.1 279.9 ;
      RECT  169.7 282.2 170.5 283.0 ;
      RECT  169.8 290.2 170.4 289.6 ;
      RECT  169.8 297.2 170.4 296.6 ;
      RECT  167.1 290.2 170.1 289.6 ;
      RECT  169.8 293.8 170.4 289.9 ;
      RECT  169.8 296.9 170.4 293.8 ;
      RECT  168.7 297.2 170.1 296.6 ;
      RECT  166.7 290.3 167.5 289.5 ;
      RECT  168.3 297.3 169.1 296.5 ;
      RECT  169.7 294.2 170.5 293.4 ;
      RECT  169.8 307.0 170.4 307.6 ;
      RECT  169.8 300.0 170.4 300.6 ;
      RECT  167.1 307.0 170.1 307.6 ;
      RECT  169.8 303.4 170.4 307.3 ;
      RECT  169.8 300.3 170.4 303.4 ;
      RECT  168.7 300.0 170.1 300.6 ;
      RECT  166.7 306.9 167.5 307.7 ;
      RECT  168.3 299.9 169.1 300.7 ;
      RECT  169.7 303.0 170.5 303.8 ;
      RECT  169.8 311.0 170.4 310.4 ;
      RECT  169.8 318.0 170.4 317.4 ;
      RECT  167.1 311.0 170.1 310.4 ;
      RECT  169.8 314.6 170.4 310.7 ;
      RECT  169.8 317.7 170.4 314.6 ;
      RECT  168.7 318.0 170.1 317.4 ;
      RECT  166.7 311.1 167.5 310.3 ;
      RECT  168.3 318.1 169.1 317.3 ;
      RECT  169.7 315.0 170.5 314.2 ;
      RECT  169.8 327.8 170.4 328.4 ;
      RECT  169.8 320.8 170.4 321.4 ;
      RECT  167.1 327.8 170.1 328.4 ;
      RECT  169.8 324.2 170.4 328.1 ;
      RECT  169.8 321.1 170.4 324.2 ;
      RECT  168.7 320.8 170.1 321.4 ;
      RECT  166.7 327.7 167.5 328.5 ;
      RECT  168.3 320.7 169.1 321.5 ;
      RECT  169.7 323.8 170.5 324.6 ;
      RECT  169.8 331.8 170.4 331.2 ;
      RECT  169.8 338.8 170.4 338.2 ;
      RECT  167.1 331.8 170.1 331.2 ;
      RECT  169.8 335.4 170.4 331.5 ;
      RECT  169.8 338.5 170.4 335.4 ;
      RECT  168.7 338.8 170.1 338.2 ;
      RECT  166.7 331.9 167.5 331.1 ;
      RECT  168.3 338.9 169.1 338.1 ;
      RECT  169.7 335.8 170.5 335.0 ;
      RECT  169.8 348.6 170.4 349.2 ;
      RECT  169.8 341.6 170.4 342.2 ;
      RECT  167.1 348.6 170.1 349.2 ;
      RECT  169.8 345.0 170.4 348.9 ;
      RECT  169.8 341.9 170.4 345.0 ;
      RECT  168.7 341.6 170.1 342.2 ;
      RECT  166.7 348.5 167.5 349.3 ;
      RECT  168.3 341.5 169.1 342.3 ;
      RECT  169.7 344.6 170.5 345.4 ;
      RECT  169.8 352.6 170.4 352.0 ;
      RECT  169.8 359.6 170.4 359.0 ;
      RECT  167.1 352.6 170.1 352.0 ;
      RECT  169.8 356.2 170.4 352.3 ;
      RECT  169.8 359.3 170.4 356.2 ;
      RECT  168.7 359.6 170.1 359.0 ;
      RECT  166.7 352.7 167.5 351.9 ;
      RECT  168.3 359.7 169.1 358.9 ;
      RECT  169.7 356.6 170.5 355.8 ;
      RECT  161.4 199.0 162.2 199.8 ;
      RECT  162.7 197.0 163.5 197.8 ;
      RECT  166.7 197.6 167.5 198.4 ;
      RECT  161.4 210.2 162.2 211.0 ;
      RECT  162.7 212.2 163.5 213.0 ;
      RECT  166.7 211.6 167.5 212.4 ;
      RECT  161.4 219.8 162.2 220.6 ;
      RECT  162.7 217.8 163.5 218.6 ;
      RECT  166.7 218.4 167.5 219.2 ;
      RECT  161.4 231.0 162.2 231.8 ;
      RECT  162.7 233.0 163.5 233.8 ;
      RECT  166.7 232.4 167.5 233.2 ;
      RECT  161.4 240.6 162.2 241.4 ;
      RECT  162.7 238.6 163.5 239.4 ;
      RECT  166.7 239.2 167.5 240.0 ;
      RECT  161.4 251.8 162.2 252.6 ;
      RECT  162.7 253.8 163.5 254.6 ;
      RECT  166.7 253.2 167.5 254.0 ;
      RECT  161.4 261.4 162.2 262.2 ;
      RECT  162.7 259.4 163.5 260.2 ;
      RECT  166.7 260.0 167.5 260.8 ;
      RECT  161.4 272.6 162.2 273.4 ;
      RECT  162.7 274.6 163.5 275.4 ;
      RECT  166.7 274.0 167.5 274.8 ;
      RECT  161.4 282.2 162.2 283.0 ;
      RECT  162.7 280.2 163.5 281.0 ;
      RECT  166.7 280.8 167.5 281.6 ;
      RECT  161.4 293.4 162.2 294.2 ;
      RECT  162.7 295.4 163.5 296.2 ;
      RECT  166.7 294.8 167.5 295.6 ;
      RECT  161.4 303.0 162.2 303.8 ;
      RECT  162.7 301.0 163.5 301.8 ;
      RECT  166.7 301.6 167.5 302.4 ;
      RECT  161.4 314.2 162.2 315.0 ;
      RECT  162.7 316.2 163.5 317.0 ;
      RECT  166.7 315.6 167.5 316.4 ;
      RECT  161.4 323.8 162.2 324.6 ;
      RECT  162.7 321.8 163.5 322.6 ;
      RECT  166.7 322.4 167.5 323.2 ;
      RECT  161.4 335.0 162.2 335.8 ;
      RECT  162.7 337.0 163.5 337.8 ;
      RECT  166.7 336.4 167.5 337.2 ;
      RECT  161.4 344.6 162.2 345.4 ;
      RECT  162.7 342.6 163.5 343.4 ;
      RECT  166.7 343.2 167.5 344.0 ;
      RECT  161.4 355.8 162.2 356.6 ;
      RECT  162.7 357.8 163.5 358.6 ;
      RECT  166.7 357.2 167.5 358.0 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 194.2 173.9 195.0 ;
      RECT  173.1 194.2 173.9 195.0 ;
      RECT  173.1 194.2 173.9 195.0 ;
      RECT  173.1 194.2 173.9 195.0 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 360.6 173.9 361.4 ;
      RECT  173.1 360.6 173.9 361.4 ;
      RECT  173.1 360.6 173.9 361.4 ;
      RECT  173.1 360.6 173.9 361.4 ;
      RECT  161.5 194.6 162.1 361.0 ;
      RECT  89.5 194.6 90.1 277.8 ;
      RECT  90.9 194.6 91.5 277.8 ;
      RECT  92.3 194.6 92.9 277.8 ;
      RECT  93.7 194.6 94.3 277.8 ;
      RECT  161.5 194.6 162.1 361.0 ;
      RECT  181.5 159.7 182.3 160.5 ;
      RECT  181.5 159.7 182.3 160.5 ;
      RECT  182.9 191.2 183.7 192.0 ;
      RECT  182.9 191.2 183.7 192.0 ;
      RECT  178.7 79.7 179.5 80.5 ;
      RECT  178.7 79.7 179.5 80.5 ;
      RECT  180.1 149.5 180.9 150.3 ;
      RECT  180.1 149.5 180.9 150.3 ;
      RECT  161.4 185.8 162.2 186.6 ;
      RECT  182.9 185.8 183.7 186.6 ;
      RECT  200.0 119.8 200.8 122.8 ;
      RECT  206.8 119.8 207.6 122.8 ;
      RECT  202.4 75.0 203.2 77.0 ;
      RECT  209.2 75.0 210.0 77.0 ;
      RECT  89.5 194.6 90.1 277.8 ;
      RECT  90.9 194.6 91.5 277.8 ;
      RECT  92.3 194.6 92.9 277.8 ;
      RECT  93.7 194.6 94.3 277.8 ;
      RECT  180.2 75.0 180.8 191.4 ;
      RECT  181.6 75.0 182.2 191.4 ;
      RECT  178.8 75.0 179.4 191.4 ;
      RECT  183.0 75.0 183.6 191.4 ;
      RECT  37.4 2.2 38.0 163.6 ;
      RECT  38.8 2.2 39.4 163.6 ;
      RECT  40.2 2.2 40.8 163.6 ;
      RECT  41.6 2.2 42.2 163.6 ;
      RECT  43.0 2.2 43.6 163.6 ;
      RECT  44.4 2.2 45.0 163.6 ;
      RECT  45.8 2.2 46.4 163.6 ;
      RECT  47.2 2.2 47.8 163.6 ;
      RECT  47.2 13.2 47.8 82.9 ;
      RECT  43.0 31.2 43.6 82.9 ;
      RECT  45.8 34.4 46.4 82.9 ;
      RECT  5.6 42.2 6.2 45.0 ;
      RECT  40.2 72.4 40.8 82.9 ;
      RECT  37.4 82.9 38.0 132.0 ;
      RECT  38.8 82.9 39.4 132.0 ;
      RECT  43.0 82.9 43.6 87.9 ;
      RECT  37.4 82.9 38.0 86.6 ;
      RECT  40.2 82.9 40.8 85.3 ;
      RECT  38.8 82.9 39.4 156.5 ;
      RECT  40.2 82.9 40.8 157.8 ;
      RECT  45.8 82.9 46.4 159.1 ;
      RECT  5.3 101.9 5.9 165.0 ;
      RECT  41.6 82.9 42.2 117.4 ;
      RECT  38.8 82.9 39.4 118.8 ;
      RECT  56.3 112.4 56.9 117.4 ;
      RECT  74.0 5.0 74.6 11.2 ;
      RECT  44.4 5.0 45.0 82.9 ;
      RECT  44.4 32.4 45.0 82.9 ;
      RECT  47.2 37.4 47.8 82.9 ;
      RECT  40.2 33.0 40.8 82.9 ;
      RECT  44.4 47.0 45.0 82.9 ;
      RECT  47.2 45.6 47.8 82.9 ;
      RECT  41.6 51.4 42.2 82.9 ;
      RECT  10.4 10.8 11.2 11.6 ;
      RECT  21.6 11.6 22.4 12.4 ;
      RECT  5.6 8.8 6.4 9.6 ;
      RECT  4.0 7.4 4.8 13.0 ;
      RECT  7.2 5.4 8.0 17.0 ;
      RECT  16.8 5.4 17.6 17.0 ;
      RECT  21.6 11.6 22.4 12.4 ;
      RECT  26.0 11.4 26.8 12.2 ;
      RECT  26.0 11.4 26.8 12.2 ;
      RECT  35.5 9.6 36.3 10.4 ;
      RECT  30.0 12.8 30.8 13.6 ;
      RECT  10.4 10.8 11.2 11.6 ;
      RECT  35.6 9.7 36.2 10.3 ;
      RECT  30.2 12.9 30.8 13.5 ;
      RECT  5.6 8.8 6.4 9.6 ;
      RECT  10.4 33.6 11.2 32.8 ;
      RECT  21.6 32.8 22.4 32.0 ;
      RECT  5.6 35.6 6.4 34.8 ;
      RECT  4.0 37.0 4.8 31.4 ;
      RECT  7.2 39.0 8.0 27.4 ;
      RECT  16.8 39.0 17.6 27.4 ;
      RECT  21.6 32.8 22.4 32.0 ;
      RECT  26.0 33.0 26.8 32.2 ;
      RECT  26.0 33.0 26.8 32.2 ;
      RECT  35.5 34.8 36.3 34.0 ;
      RECT  30.0 31.6 30.8 30.8 ;
      RECT  10.4 33.6 11.2 32.8 ;
      RECT  35.6 34.7 36.2 34.1 ;
      RECT  30.2 31.5 30.8 30.9 ;
      RECT  5.6 35.6 6.4 34.8 ;
      RECT  2.4 21.8 3.2 22.6 ;
      RECT  2.4 21.8 3.2 22.6 ;
      RECT  2.4 1.8 3.2 2.6 ;
      RECT  2.4 1.8 3.2 2.6 ;
      RECT  2.4 21.8 3.2 22.6 ;
      RECT  2.4 21.8 3.2 22.6 ;
      RECT  2.4 41.8 3.2 42.6 ;
      RECT  2.4 41.8 3.2 42.6 ;
      RECT  10.4 10.8 11.2 11.6 ;
      RECT  10.4 32.8 11.2 33.6 ;
      RECT  35.6 9.7 36.2 10.3 ;
      RECT  30.2 12.9 30.8 13.5 ;
      RECT  35.6 34.1 36.2 34.7 ;
      RECT  30.2 30.9 30.8 31.5 ;
      RECT  5.6 2.2 6.2 42.2 ;
      RECT  62.3 24.2 62.9 23.6 ;
      RECT  62.3 40.8 62.9 40.2 ;
      RECT  59.6 24.2 62.6 23.6 ;
      RECT  62.3 37.4 62.9 23.9 ;
      RECT  62.3 40.5 62.9 37.4 ;
      RECT  61.2 40.8 62.6 40.2 ;
      RECT  59.2 24.3 60.0 23.5 ;
      RECT  60.8 40.9 61.6 40.1 ;
      RECT  62.2 37.8 63.0 37.0 ;
      RECT  55.9 60.2 56.5 60.8 ;
      RECT  55.9 43.6 56.5 44.2 ;
      RECT  53.2 60.2 56.2 60.8 ;
      RECT  55.9 47.0 56.5 60.5 ;
      RECT  55.9 43.9 56.5 47.0 ;
      RECT  54.8 43.6 56.2 44.2 ;
      RECT  52.8 60.1 53.6 60.9 ;
      RECT  54.4 43.5 55.2 44.3 ;
      RECT  55.8 46.6 56.6 47.4 ;
      RECT  56.1 84.3 56.7 100.1 ;
      RECT  52.9 87.6 53.5 88.2 ;
      RECT  56.1 87.6 56.7 88.2 ;
      RECT  52.9 87.9 53.5 100.1 ;
      RECT  53.2 87.6 56.4 88.2 ;
      RECT  56.1 84.3 56.7 87.9 ;
      RECT  52.8 100.1 53.6 100.9 ;
      RECT  56.0 100.1 56.8 100.9 ;
      RECT  56.0 83.5 56.8 84.3 ;
      RECT  56.0 87.5 56.8 88.3 ;
      RECT  56.1 160.1 56.7 144.3 ;
      RECT  52.9 156.8 53.5 156.2 ;
      RECT  56.1 156.8 56.7 156.2 ;
      RECT  52.9 156.5 53.5 144.3 ;
      RECT  53.2 156.8 56.4 156.2 ;
      RECT  56.1 160.1 56.7 156.5 ;
      RECT  52.8 144.3 53.6 143.5 ;
      RECT  56.0 144.3 56.8 143.5 ;
      RECT  56.0 160.9 56.8 160.1 ;
      RECT  56.0 156.9 56.8 156.1 ;
      RECT  31.6 175.1 31.0 175.7 ;
      RECT  33.3 175.1 32.7 175.7 ;
      RECT  31.6 170.0 31.0 175.4 ;
      RECT  33.0 175.1 31.3 175.7 ;
      RECT  33.3 175.4 32.7 180.8 ;
      RECT  31.6 185.5 31.0 186.1 ;
      RECT  33.3 185.5 32.7 186.1 ;
      RECT  31.6 180.8 31.0 185.8 ;
      RECT  33.0 185.5 31.3 186.1 ;
      RECT  33.3 185.8 32.7 190.8 ;
      RECT  31.6 195.9 31.0 196.5 ;
      RECT  33.3 195.9 32.7 196.5 ;
      RECT  31.6 190.8 31.0 196.2 ;
      RECT  33.0 195.9 31.3 196.5 ;
      RECT  33.3 196.2 32.7 201.6 ;
      RECT  31.6 206.3 31.0 206.9 ;
      RECT  33.3 206.3 32.7 206.9 ;
      RECT  31.6 201.6 31.0 206.6 ;
      RECT  33.0 206.3 31.3 206.9 ;
      RECT  33.3 206.6 32.7 211.6 ;
      RECT  31.6 216.7 31.0 217.3 ;
      RECT  33.3 216.7 32.7 217.3 ;
      RECT  31.6 211.6 31.0 217.0 ;
      RECT  33.0 216.7 31.3 217.3 ;
      RECT  33.3 217.0 32.7 222.4 ;
      RECT  31.6 227.1 31.0 227.7 ;
      RECT  33.3 227.1 32.7 227.7 ;
      RECT  31.6 222.4 31.0 227.4 ;
      RECT  33.0 227.1 31.3 227.7 ;
      RECT  33.3 227.4 32.7 232.4 ;
      RECT  31.6 237.5 31.0 238.1 ;
      RECT  33.3 237.5 32.7 238.1 ;
      RECT  31.6 232.4 31.0 237.8 ;
      RECT  33.0 237.5 31.3 238.1 ;
      RECT  33.3 237.8 32.7 243.2 ;
      RECT  31.6 247.9 31.0 248.5 ;
      RECT  33.3 247.9 32.7 248.5 ;
      RECT  31.6 243.2 31.0 248.2 ;
      RECT  33.0 247.9 31.3 248.5 ;
      RECT  33.3 248.2 32.7 253.2 ;
      RECT  5.9 252.9 5.3 253.5 ;
      RECT  7.4 252.9 5.6 253.5 ;
      RECT  5.9 165.0 5.3 253.2 ;
      RECT  27.0 169.6 26.2 170.4 ;
      RECT  27.0 169.6 26.2 170.4 ;
      RECT  20.6 169.6 19.8 170.4 ;
      RECT  20.6 169.6 19.8 170.4 ;
      RECT  14.2 169.6 13.4 170.4 ;
      RECT  14.2 169.6 13.4 170.4 ;
      RECT  7.8 169.6 7.0 170.4 ;
      RECT  7.8 169.6 7.0 170.4 ;
      RECT  33.4 169.6 32.6 170.4 ;
      RECT  31.7 169.6 30.9 170.4 ;
      RECT  31.7 169.6 30.9 170.4 ;
      RECT  27.0 180.4 26.2 181.2 ;
      RECT  27.0 180.4 26.2 181.2 ;
      RECT  20.6 180.4 19.8 181.2 ;
      RECT  20.6 180.4 19.8 181.2 ;
      RECT  14.2 180.4 13.4 181.2 ;
      RECT  14.2 180.4 13.4 181.2 ;
      RECT  7.8 180.4 7.0 181.2 ;
      RECT  7.8 180.4 7.0 181.2 ;
      RECT  33.4 180.4 32.6 181.2 ;
      RECT  31.7 180.4 30.9 181.2 ;
      RECT  31.7 180.4 30.9 181.2 ;
      RECT  27.0 190.4 26.2 191.2 ;
      RECT  27.0 190.4 26.2 191.2 ;
      RECT  20.6 190.4 19.8 191.2 ;
      RECT  20.6 190.4 19.8 191.2 ;
      RECT  14.2 190.4 13.4 191.2 ;
      RECT  14.2 190.4 13.4 191.2 ;
      RECT  7.8 190.4 7.0 191.2 ;
      RECT  7.8 190.4 7.0 191.2 ;
      RECT  33.4 190.4 32.6 191.2 ;
      RECT  31.7 190.4 30.9 191.2 ;
      RECT  31.7 190.4 30.9 191.2 ;
      RECT  27.0 201.2 26.2 202.0 ;
      RECT  27.0 201.2 26.2 202.0 ;
      RECT  20.6 201.2 19.8 202.0 ;
      RECT  20.6 201.2 19.8 202.0 ;
      RECT  14.2 201.2 13.4 202.0 ;
      RECT  14.2 201.2 13.4 202.0 ;
      RECT  7.8 201.2 7.0 202.0 ;
      RECT  7.8 201.2 7.0 202.0 ;
      RECT  33.4 201.2 32.6 202.0 ;
      RECT  31.7 201.2 30.9 202.0 ;
      RECT  31.7 201.2 30.9 202.0 ;
      RECT  27.0 211.2 26.2 212.0 ;
      RECT  27.0 211.2 26.2 212.0 ;
      RECT  20.6 211.2 19.8 212.0 ;
      RECT  20.6 211.2 19.8 212.0 ;
      RECT  14.2 211.2 13.4 212.0 ;
      RECT  14.2 211.2 13.4 212.0 ;
      RECT  7.8 211.2 7.0 212.0 ;
      RECT  7.8 211.2 7.0 212.0 ;
      RECT  33.4 211.2 32.6 212.0 ;
      RECT  31.7 211.2 30.9 212.0 ;
      RECT  31.7 211.2 30.9 212.0 ;
      RECT  27.0 222.0 26.2 222.8 ;
      RECT  27.0 222.0 26.2 222.8 ;
      RECT  20.6 222.0 19.8 222.8 ;
      RECT  20.6 222.0 19.8 222.8 ;
      RECT  14.2 222.0 13.4 222.8 ;
      RECT  14.2 222.0 13.4 222.8 ;
      RECT  7.8 222.0 7.0 222.8 ;
      RECT  7.8 222.0 7.0 222.8 ;
      RECT  33.4 222.0 32.6 222.8 ;
      RECT  31.7 222.0 30.9 222.8 ;
      RECT  31.7 222.0 30.9 222.8 ;
      RECT  27.0 232.0 26.2 232.8 ;
      RECT  27.0 232.0 26.2 232.8 ;
      RECT  20.6 232.0 19.8 232.8 ;
      RECT  20.6 232.0 19.8 232.8 ;
      RECT  14.2 232.0 13.4 232.8 ;
      RECT  14.2 232.0 13.4 232.8 ;
      RECT  7.8 232.0 7.0 232.8 ;
      RECT  7.8 232.0 7.0 232.8 ;
      RECT  33.4 232.0 32.6 232.8 ;
      RECT  31.7 232.0 30.9 232.8 ;
      RECT  31.7 232.0 30.9 232.8 ;
      RECT  27.0 242.8 26.2 243.6 ;
      RECT  27.0 242.8 26.2 243.6 ;
      RECT  20.6 242.8 19.8 243.6 ;
      RECT  20.6 242.8 19.8 243.6 ;
      RECT  14.2 242.8 13.4 243.6 ;
      RECT  14.2 242.8 13.4 243.6 ;
      RECT  7.8 242.8 7.0 243.6 ;
      RECT  7.8 242.8 7.0 243.6 ;
      RECT  33.4 242.8 32.6 243.6 ;
      RECT  31.7 242.8 30.9 243.6 ;
      RECT  31.7 242.8 30.9 243.6 ;
      RECT  27.0 252.8 26.2 253.6 ;
      RECT  27.0 252.8 26.2 253.6 ;
      RECT  20.6 252.8 19.8 253.6 ;
      RECT  20.6 252.8 19.8 253.6 ;
      RECT  14.2 252.8 13.4 253.6 ;
      RECT  14.2 252.8 13.4 253.6 ;
      RECT  7.8 252.8 7.0 253.6 ;
      RECT  7.8 252.8 7.0 253.6 ;
      RECT  33.4 252.8 32.6 253.6 ;
      RECT  31.7 252.8 30.9 253.6 ;
      RECT  31.7 252.8 30.9 253.6 ;
      RECT  22.4 175.0 21.6 175.8 ;
      RECT  22.4 175.0 21.6 175.8 ;
      RECT  22.4 164.6 21.6 165.4 ;
      RECT  22.4 164.6 21.6 165.4 ;
      RECT  16.0 175.0 15.2 175.8 ;
      RECT  16.0 175.0 15.2 175.8 ;
      RECT  16.0 164.6 15.2 165.4 ;
      RECT  16.0 164.6 15.2 165.4 ;
      RECT  9.6 175.0 8.8 175.8 ;
      RECT  9.6 175.0 8.8 175.8 ;
      RECT  9.6 164.6 8.8 165.4 ;
      RECT  9.6 164.6 8.8 165.4 ;
      RECT  22.4 195.8 21.6 196.6 ;
      RECT  22.4 195.8 21.6 196.6 ;
      RECT  22.4 185.4 21.6 186.2 ;
      RECT  22.4 185.4 21.6 186.2 ;
      RECT  16.0 195.8 15.2 196.6 ;
      RECT  16.0 195.8 15.2 196.6 ;
      RECT  16.0 185.4 15.2 186.2 ;
      RECT  16.0 185.4 15.2 186.2 ;
      RECT  9.6 195.8 8.8 196.6 ;
      RECT  9.6 195.8 8.8 196.6 ;
      RECT  9.6 185.4 8.8 186.2 ;
      RECT  9.6 185.4 8.8 186.2 ;
      RECT  22.4 216.6 21.6 217.4 ;
      RECT  22.4 216.6 21.6 217.4 ;
      RECT  22.4 206.2 21.6 207.0 ;
      RECT  22.4 206.2 21.6 207.0 ;
      RECT  16.0 216.6 15.2 217.4 ;
      RECT  16.0 216.6 15.2 217.4 ;
      RECT  16.0 206.2 15.2 207.0 ;
      RECT  16.0 206.2 15.2 207.0 ;
      RECT  9.6 216.6 8.8 217.4 ;
      RECT  9.6 216.6 8.8 217.4 ;
      RECT  9.6 206.2 8.8 207.0 ;
      RECT  9.6 206.2 8.8 207.0 ;
      RECT  22.4 237.4 21.6 238.2 ;
      RECT  22.4 237.4 21.6 238.2 ;
      RECT  22.4 227.0 21.6 227.8 ;
      RECT  22.4 227.0 21.6 227.8 ;
      RECT  16.0 237.4 15.2 238.2 ;
      RECT  16.0 237.4 15.2 238.2 ;
      RECT  16.0 227.0 15.2 227.8 ;
      RECT  16.0 227.0 15.2 227.8 ;
      RECT  9.6 237.4 8.8 238.2 ;
      RECT  9.6 237.4 8.8 238.2 ;
      RECT  9.6 227.0 8.8 227.8 ;
      RECT  9.6 227.0 8.8 227.8 ;
      RECT  22.4 258.2 21.6 259.0 ;
      RECT  22.4 258.2 21.6 259.0 ;
      RECT  22.4 247.8 21.6 248.6 ;
      RECT  22.4 247.8 21.6 248.6 ;
      RECT  16.0 258.2 15.2 259.0 ;
      RECT  16.0 258.2 15.2 259.0 ;
      RECT  16.0 247.8 15.2 248.6 ;
      RECT  16.0 247.8 15.2 248.6 ;
      RECT  9.6 258.2 8.8 259.0 ;
      RECT  9.6 258.2 8.8 259.0 ;
      RECT  9.6 247.8 8.8 248.6 ;
      RECT  9.6 247.8 8.8 248.6 ;
      RECT  22.4 247.8 21.6 248.6 ;
      RECT  22.4 247.8 21.6 248.6 ;
      RECT  16.0 247.8 15.2 248.6 ;
      RECT  16.0 247.8 15.2 248.6 ;
      RECT  9.6 247.8 8.8 248.6 ;
      RECT  9.6 247.8 8.8 248.6 ;
      RECT  33.4 169.6 32.6 170.4 ;
      RECT  7.8 252.8 7.0 253.6 ;
      RECT  33.4 165.0 32.8 170.0 ;
      RECT  5.9 165.0 5.3 253.2 ;
      RECT  55.9 104.2 56.5 103.6 ;
      RECT  55.9 120.8 56.5 120.2 ;
      RECT  53.2 104.2 56.2 103.6 ;
      RECT  55.9 117.4 56.5 103.9 ;
      RECT  55.9 120.5 56.5 117.4 ;
      RECT  54.8 120.8 56.2 120.2 ;
      RECT  52.8 104.3 53.6 103.5 ;
      RECT  54.4 120.9 55.2 120.1 ;
      RECT  55.8 117.8 56.6 117.0 ;
      RECT  47.1 12.8 47.9 13.6 ;
      RECT  30.1 12.8 30.9 13.6 ;
      RECT  42.9 30.8 43.7 31.6 ;
      RECT  30.1 30.8 30.9 31.6 ;
      RECT  45.7 34.0 46.5 34.8 ;
      RECT  35.5 34.0 36.3 34.8 ;
      RECT  5.5 44.6 6.3 45.4 ;
      RECT  44.3 44.6 45.1 45.4 ;
      RECT  40.1 72.0 40.9 72.8 ;
      RECT  37.3 131.6 38.1 132.4 ;
      RECT  53.1 131.6 53.9 132.4 ;
      RECT  53.1 131.6 53.9 132.4 ;
      RECT  38.7 131.6 39.5 132.4 ;
      RECT  42.9 87.5 43.7 88.3 ;
      RECT  37.3 86.2 38.1 87.0 ;
      RECT  40.1 84.9 40.9 85.7 ;
      RECT  38.7 156.1 39.5 156.9 ;
      RECT  40.1 157.4 40.9 158.2 ;
      RECT  45.7 158.7 46.5 159.5 ;
      RECT  5.2 101.5 6.0 102.3 ;
      RECT  38.7 101.5 39.5 102.3 ;
      RECT  41.5 117.0 42.3 117.8 ;
      RECT  38.7 118.4 39.5 119.2 ;
      RECT  56.2 112.0 57.0 112.8 ;
      RECT  51.4 11.6 52.2 12.4 ;
      RECT  73.9 4.6 74.7 5.4 ;
      RECT  44.3 4.6 45.1 5.4 ;
      RECT  73.9 10.8 74.7 11.6 ;
      RECT  44.3 32.0 45.1 32.8 ;
      RECT  47.1 37.0 47.9 37.8 ;
      RECT  58.0 37.0 58.8 37.8 ;
      RECT  58.0 37.0 58.8 37.8 ;
      RECT  40.1 32.6 40.9 33.4 ;
      RECT  81.9 32.6 82.7 33.4 ;
      RECT  81.9 32.6 82.7 33.4 ;
      RECT  44.3 46.6 45.1 47.4 ;
      RECT  47.1 45.2 47.9 46.0 ;
      RECT  41.5 51.0 42.3 51.8 ;
      RECT  75.5 51.0 76.3 51.8 ;
      RECT  75.5 51.0 76.3 51.8 ;
      RECT  84.8 21.8 85.6 22.6 ;
      RECT  84.8 21.8 85.6 22.6 ;
      RECT  84.8 1.8 85.6 2.6 ;
      RECT  84.8 1.8 85.6 2.6 ;
      RECT  84.8 21.8 85.6 22.6 ;
      RECT  84.8 21.8 85.6 22.6 ;
      RECT  84.8 41.8 85.6 42.6 ;
      RECT  84.8 41.8 85.6 42.6 ;
      RECT  84.8 61.8 85.6 62.6 ;
      RECT  84.8 61.8 85.6 62.6 ;
      RECT  84.8 41.8 85.6 42.6 ;
      RECT  84.8 41.8 85.6 42.6 ;
      RECT  84.8 61.8 85.6 62.6 ;
      RECT  84.8 61.8 85.6 62.6 ;
      RECT  84.8 81.8 85.6 82.6 ;
      RECT  84.8 81.8 85.6 82.6 ;
      RECT  84.8 101.8 85.6 102.6 ;
      RECT  84.8 101.8 85.6 102.6 ;
      RECT  84.8 81.8 85.6 82.6 ;
      RECT  84.8 81.8 85.6 82.6 ;
      RECT  84.8 101.8 85.6 102.6 ;
      RECT  84.8 101.8 85.6 102.6 ;
      RECT  84.8 121.8 85.6 122.6 ;
      RECT  84.8 121.8 85.6 122.6 ;
      RECT  84.8 141.8 85.6 142.6 ;
      RECT  84.8 141.8 85.6 142.6 ;
      RECT  84.8 121.8 85.6 122.6 ;
      RECT  84.8 121.8 85.6 122.6 ;
      RECT  84.8 141.8 85.6 142.6 ;
      RECT  84.8 141.8 85.6 142.6 ;
      RECT  84.8 161.8 85.6 162.6 ;
      RECT  84.8 161.8 85.6 162.6 ;
      RECT  10.4 10.8 11.2 11.6 ;
      RECT  10.4 32.8 11.2 33.6 ;
      RECT  51.5 2.2 52.1 12.0 ;
      RECT  32.8 165.0 33.4 170.0 ;
      RECT  67.6 292.8 68.2 372.8 ;
      RECT  72.4 301.4 73.2 302.2 ;
      RECT  83.6 302.2 84.4 303.0 ;
      RECT  67.6 299.4 68.4 300.2 ;
      RECT  66.0 298.0 66.8 303.6 ;
      RECT  69.2 296.0 70.0 307.6 ;
      RECT  78.8 296.0 79.6 307.6 ;
      RECT  72.4 324.2 73.2 323.4 ;
      RECT  83.6 323.4 84.4 322.6 ;
      RECT  67.6 326.2 68.4 325.4 ;
      RECT  66.0 327.6 66.8 322.0 ;
      RECT  69.2 329.6 70.0 318.0 ;
      RECT  78.8 329.6 79.6 318.0 ;
      RECT  72.4 341.4 73.2 342.2 ;
      RECT  83.6 342.2 84.4 343.0 ;
      RECT  67.6 339.4 68.4 340.2 ;
      RECT  66.0 338.0 66.8 343.6 ;
      RECT  69.2 336.0 70.0 347.6 ;
      RECT  78.8 336.0 79.6 347.6 ;
      RECT  72.4 364.2 73.2 363.4 ;
      RECT  83.6 363.4 84.4 362.6 ;
      RECT  67.6 366.2 68.4 365.4 ;
      RECT  66.0 367.6 66.8 362.0 ;
      RECT  69.2 369.6 70.0 358.0 ;
      RECT  78.8 369.6 79.6 358.0 ;
      RECT  75.3 312.4 76.1 313.2 ;
      RECT  75.3 312.4 76.1 313.2 ;
      RECT  75.3 292.4 76.1 293.2 ;
      RECT  75.3 292.4 76.1 293.2 ;
      RECT  75.3 312.4 76.1 313.2 ;
      RECT  75.3 312.4 76.1 313.2 ;
      RECT  75.3 332.4 76.1 333.2 ;
      RECT  75.3 332.4 76.1 333.2 ;
      RECT  75.3 352.4 76.1 353.2 ;
      RECT  75.3 352.4 76.1 353.2 ;
      RECT  75.3 332.4 76.1 333.2 ;
      RECT  75.3 332.4 76.1 333.2 ;
      RECT  75.3 352.4 76.1 353.2 ;
      RECT  75.3 352.4 76.1 353.2 ;
      RECT  75.3 372.4 76.1 373.2 ;
      RECT  75.3 372.4 76.1 373.2 ;
      RECT  67.6 297.8 68.4 298.6 ;
      RECT  72.4 301.4 73.2 302.2 ;
      RECT  72.4 323.4 73.2 324.2 ;
      RECT  72.4 341.4 73.2 342.2 ;
      RECT  72.4 363.4 73.2 364.2 ;
      RECT  83.6 302.2 84.4 303.0 ;
      RECT  83.6 322.6 84.4 323.4 ;
      RECT  83.6 342.2 84.4 343.0 ;
      RECT  83.6 362.6 84.4 363.4 ;
      RECT  188.6 48.0 189.2 68.0 ;
      RECT  210.4 48.0 211.0 68.0 ;
      RECT  193.4 56.6 194.2 57.4 ;
      RECT  204.6 57.4 205.4 58.2 ;
      RECT  188.6 54.6 189.4 55.4 ;
      RECT  187.0 53.2 187.8 58.8 ;
      RECT  190.2 51.2 191.0 62.8 ;
      RECT  199.8 51.2 200.6 62.8 ;
      RECT  215.2 56.6 216.0 57.4 ;
      RECT  226.4 57.4 227.2 58.2 ;
      RECT  210.4 54.6 211.2 55.4 ;
      RECT  208.8 53.2 209.6 58.8 ;
      RECT  212.0 51.2 212.8 62.8 ;
      RECT  221.6 51.2 222.4 62.8 ;
      RECT  196.3 67.6 197.1 68.4 ;
      RECT  196.3 67.6 197.1 68.4 ;
      RECT  196.3 47.6 197.1 48.4 ;
      RECT  196.3 47.6 197.1 48.4 ;
      RECT  218.1 67.6 218.9 68.4 ;
      RECT  218.1 67.6 218.9 68.4 ;
      RECT  218.1 47.6 218.9 48.4 ;
      RECT  218.1 47.6 218.9 48.4 ;
      RECT  188.6 53.0 189.4 53.8 ;
      RECT  210.4 53.0 211.2 53.8 ;
      RECT  193.4 56.6 194.2 57.4 ;
      RECT  215.2 56.6 216.0 57.4 ;
      RECT  204.6 57.4 205.4 58.2 ;
      RECT  226.4 57.4 227.2 58.2 ;
      RECT  87.6 10.8 88.4 11.6 ;
      RECT  87.6 297.8 88.4 298.6 ;
      RECT  87.6 53.0 88.4 53.8 ;
      RECT  180.1 152.2 180.9 153.0 ;
      RECT  86.2 152.2 87.0 153.0 ;
      RECT  86.2 152.2 87.0 153.0 ;
      RECT  178.7 90.8 179.5 91.6 ;
      RECT  86.2 90.8 87.0 91.6 ;
      RECT  86.2 90.8 87.0 91.6 ;
      RECT  181.5 112.0 182.3 112.8 ;
      RECT  86.2 112.0 87.0 112.8 ;
      RECT  86.2 112.0 87.0 112.8 ;
      RECT  182.9 72.8 183.7 73.6 ;
      RECT  86.2 72.8 87.0 73.6 ;
      RECT  86.2 72.8 87.0 73.6 ;
      RECT  193.8 167.1 194.6 167.9 ;
      RECT  33.0 167.1 33.8 167.9 ;
      RECT  89.4 302.2 90.2 303.0 ;
      RECT  83.6 302.2 84.4 303.0 ;
      RECT  90.8 322.6 91.6 323.4 ;
      RECT  83.6 322.6 84.4 323.4 ;
      RECT  92.2 342.2 93.0 343.0 ;
      RECT  83.6 342.2 84.4 343.0 ;
      RECT  93.6 362.6 94.4 363.4 ;
      RECT  83.6 362.6 84.4 363.4 ;
      RECT  202.4 70.4 203.2 71.2 ;
      RECT  204.6 70.4 205.4 71.2 ;
      RECT  209.2 71.8 210.0 72.6 ;
      RECT  226.4 71.8 227.2 72.6 ;
   LAYER  metal3 ;
      RECT  86.6 297.9 88.0 298.5 ;
      RECT  88.0 53.1 207.6 53.7 ;
      RECT  86.6 152.3 180.5 152.9 ;
      RECT  86.6 90.9 179.1 91.5 ;
      RECT  86.6 112.1 181.9 112.7 ;
      RECT  86.6 72.9 183.3 73.5 ;
      RECT  33.4 167.2 194.2 167.8 ;
      RECT  84.0 302.3 89.8 302.9 ;
      RECT  84.0 322.7 91.2 323.3 ;
      RECT  84.0 342.3 92.6 342.9 ;
      RECT  84.0 362.7 94.0 363.3 ;
      RECT  0.0 21.6 3.6 22.8 ;
      RECT  7.2 216.0 10.8 219.6 ;
      RECT  7.2 235.2 10.8 238.8 ;
      RECT  7.2 194.4 10.8 198.0 ;
      RECT  7.2 256.8 10.8 260.4 ;
      RECT  7.2 172.8 10.8 176.4 ;
      RECT  14.4 235.2 18.0 238.8 ;
      RECT  14.4 256.8 18.0 260.4 ;
      RECT  14.4 194.4 18.0 198.0 ;
      RECT  14.4 172.8 18.0 176.4 ;
      RECT  14.4 216.0 18.0 219.6 ;
      RECT  19.2 194.4 22.8 198.0 ;
      RECT  19.2 256.8 22.8 260.4 ;
      RECT  19.2 172.8 20.4 176.4 ;
      RECT  19.2 175.2 22.8 176.4 ;
      RECT  19.8 175.0 22.4 175.8 ;
      RECT  19.2 235.2 20.4 238.8 ;
      RECT  19.2 237.6 22.8 238.8 ;
      RECT  19.8 237.4 22.4 238.2 ;
      RECT  19.2 216.0 20.4 219.6 ;
      RECT  19.2 216.0 22.8 217.2 ;
      RECT  19.8 216.6 22.4 217.4 ;
      RECT  74.4 350.4 78.0 354.0 ;
      RECT  74.4 312.0 75.6 315.6 ;
      RECT  74.4 314.4 78.0 315.6 ;
      RECT  75.3 312.4 76.1 315.0 ;
      RECT  84.0 100.8 87.6 104.4 ;
      RECT  84.0 21.6 87.6 22.8 ;
      RECT  84.0 60.0 87.6 63.6 ;
      RECT  84.0 141.6 87.6 142.8 ;
      RECT  103.2 266.4 106.8 270.0 ;
      RECT  103.2 244.8 106.8 248.4 ;
      RECT  103.2 204.0 106.8 207.6 ;
      RECT  103.2 223.2 106.8 226.8 ;
      RECT  122.4 223.2 123.6 226.8 ;
      RECT  122.4 204.0 123.6 207.6 ;
      RECT  122.4 266.4 123.6 270.0 ;
      RECT  122.4 244.8 123.6 248.4 ;
      RECT  144.0 244.8 147.6 248.4 ;
      RECT  144.0 348.0 147.6 351.6 ;
      RECT  144.0 307.2 147.6 310.8 ;
      RECT  144.0 285.6 147.6 289.2 ;
      RECT  144.0 223.2 147.6 226.8 ;
      RECT  144.0 328.8 147.6 332.4 ;
      RECT  144.0 204.0 147.6 207.6 ;
      RECT  144.0 266.4 147.6 270.0 ;
      RECT  172.8 244.8 174.0 248.4 ;
      RECT  172.8 204.0 174.0 207.6 ;
      RECT  172.8 328.8 174.0 332.4 ;
      RECT  172.8 348.0 174.0 351.6 ;
      RECT  172.8 223.2 174.0 226.8 ;
      RECT  172.8 285.6 174.0 289.2 ;
      RECT  172.8 266.4 174.0 270.0 ;
      RECT  172.8 307.2 174.0 310.8 ;
      RECT  187.2 204.0 190.8 205.2 ;
      RECT  187.2 285.6 190.8 289.2 ;
      RECT  187.2 328.8 190.8 330.0 ;
      RECT  187.2 348.0 190.8 351.6 ;
      RECT  187.2 369.6 190.8 373.2 ;
      RECT  187.2 182.4 190.8 186.0 ;
      RECT  187.2 244.8 190.8 248.4 ;
      RECT  187.2 223.2 190.8 226.8 ;
      RECT  187.2 307.2 190.8 310.8 ;
      RECT  187.2 266.4 190.8 267.6 ;
      RECT  194.4 160.8 198.0 164.4 ;
      RECT  194.4 307.2 198.0 310.8 ;
      RECT  194.4 244.8 198.0 248.4 ;
      RECT  194.4 204.0 198.0 205.2 ;
      RECT  194.4 266.4 198.0 267.6 ;
      RECT  194.4 223.2 198.0 226.8 ;
      RECT  194.4 328.8 198.0 330.0 ;
      RECT  194.4 182.4 198.0 186.0 ;
      RECT  194.4 348.0 198.0 351.6 ;
      RECT  194.4 369.6 198.0 373.2 ;
      RECT  194.4 285.6 198.0 289.2 ;
      RECT  194.4 69.6 198.0 70.8 ;
      RECT  196.8 67.2 198.0 70.8 ;
      RECT  196.3 67.6 197.1 70.2 ;
      RECT  201.6 160.8 205.2 164.4 ;
      RECT  201.6 244.8 205.2 248.4 ;
      RECT  201.6 369.6 205.2 373.2 ;
      RECT  201.6 348.0 205.2 351.6 ;
      RECT  201.6 204.0 205.2 205.2 ;
      RECT  201.6 266.4 205.2 267.6 ;
      RECT  201.6 307.2 205.2 310.8 ;
      RECT  201.6 182.4 205.2 186.0 ;
      RECT  201.6 223.2 205.2 226.8 ;
      RECT  201.6 285.6 205.2 289.2 ;
      RECT  201.6 328.8 205.2 330.0 ;
      RECT  201.6 98.4 205.2 99.6 ;
      RECT  201.6 79.2 205.2 82.8 ;
      RECT  204.0 132.0 207.6 135.6 ;
      RECT  208.8 160.8 210.0 164.4 ;
      RECT  208.8 307.2 212.4 310.8 ;
      RECT  208.8 204.0 212.4 205.2 ;
      RECT  208.8 328.8 212.4 330.0 ;
      RECT  208.8 244.8 212.4 248.4 ;
      RECT  208.8 223.2 212.4 226.8 ;
      RECT  208.8 369.6 212.4 373.2 ;
      RECT  208.8 348.0 212.4 351.6 ;
      RECT  208.8 182.4 212.4 186.0 ;
      RECT  208.8 266.4 212.4 267.6 ;
      RECT  208.8 285.6 212.4 289.2 ;
      RECT  208.8 98.4 212.4 99.6 ;
      RECT  208.8 79.2 212.4 82.8 ;
      RECT  211.2 132.0 214.8 135.6 ;
      RECT  213.6 328.8 217.2 330.0 ;
      RECT  213.6 285.6 217.2 289.2 ;
      RECT  213.6 204.0 217.2 205.2 ;
      RECT  213.6 244.8 217.2 248.4 ;
      RECT  213.6 223.2 217.2 226.8 ;
      RECT  213.6 307.2 217.2 310.8 ;
      RECT  213.6 348.0 217.2 351.6 ;
      RECT  213.6 369.6 217.2 373.2 ;
      RECT  213.6 266.4 217.2 267.6 ;
      RECT  213.6 182.4 217.2 186.0 ;
      RECT  218.4 67.2 219.6 70.8 ;
      RECT  216.0 69.6 219.6 70.8 ;
      RECT  218.1 67.6 218.9 70.2 ;
      RECT  0.0 40.8 3.6 44.4 ;
      RECT  0.0 0.0 3.6 3.6 ;
      RECT  7.2 163.2 10.8 166.8 ;
      RECT  7.2 184.8 10.8 188.4 ;
      RECT  7.2 225.6 10.8 229.2 ;
      RECT  7.2 247.2 10.8 250.8 ;
      RECT  7.2 204.0 10.8 207.6 ;
      RECT  14.4 225.6 18.0 229.2 ;
      RECT  14.4 247.2 18.0 250.8 ;
      RECT  14.4 163.2 18.0 166.8 ;
      RECT  14.4 184.8 18.0 188.4 ;
      RECT  14.4 204.0 18.0 207.6 ;
      RECT  19.2 204.0 20.4 207.6 ;
      RECT  19.2 206.4 22.8 207.6 ;
      RECT  19.8 206.2 22.4 207.0 ;
      RECT  19.2 163.2 22.8 166.8 ;
      RECT  19.2 184.8 20.4 188.4 ;
      RECT  19.2 184.8 22.8 186.0 ;
      RECT  19.8 185.4 22.4 186.2 ;
      RECT  19.2 225.6 22.8 229.2 ;
      RECT  19.2 247.2 20.4 250.8 ;
      RECT  19.2 247.2 22.8 248.4 ;
      RECT  19.8 247.8 22.4 248.6 ;
      RECT  74.4 290.4 78.0 294.0 ;
      RECT  74.4 372.0 75.6 375.6 ;
      RECT  74.4 374.4 78.0 375.6 ;
      RECT  75.3 372.4 76.1 375.0 ;
      RECT  74.4 331.2 78.0 334.8 ;
      RECT  84.0 0.0 87.6 3.6 ;
      RECT  84.0 160.8 87.6 164.4 ;
      RECT  84.0 40.8 87.6 44.4 ;
      RECT  84.0 81.6 87.6 82.8 ;
      RECT  84.0 120.0 87.6 123.6 ;
      RECT  103.2 254.4 106.8 258.0 ;
      RECT  103.2 235.2 106.8 238.8 ;
      RECT  103.2 192.0 106.8 195.6 ;
      RECT  103.2 213.6 106.8 217.2 ;
      RECT  103.2 276.0 106.8 279.6 ;
      RECT  122.4 192.0 123.6 195.6 ;
      RECT  122.4 235.2 123.6 238.8 ;
      RECT  122.4 254.4 123.6 258.0 ;
      RECT  122.4 213.6 123.6 217.2 ;
      RECT  122.4 276.0 123.6 279.6 ;
      RECT  144.0 254.4 147.6 258.0 ;
      RECT  144.0 297.6 147.6 301.2 ;
      RECT  144.0 338.4 147.6 342.0 ;
      RECT  144.0 235.2 147.6 238.8 ;
      RECT  144.0 192.0 147.6 195.6 ;
      RECT  144.0 316.8 147.6 320.4 ;
      RECT  144.0 276.0 147.6 279.6 ;
      RECT  144.0 360.0 147.6 363.6 ;
      RECT  144.0 213.6 147.6 217.2 ;
      RECT  172.8 235.2 174.0 238.8 ;
      RECT  172.8 192.0 174.0 195.6 ;
      RECT  172.8 360.0 174.0 363.6 ;
      RECT  172.8 276.0 174.0 279.6 ;
      RECT  172.8 297.6 174.0 301.2 ;
      RECT  172.8 254.4 174.0 258.0 ;
      RECT  172.8 316.8 174.0 320.4 ;
      RECT  172.8 338.4 174.0 342.0 ;
      RECT  172.8 213.6 174.0 217.2 ;
      RECT  184.8 177.6 188.4 181.2 ;
      RECT  184.8 218.4 188.4 222.0 ;
      RECT  184.8 228.0 188.4 231.6 ;
      RECT  184.8 352.8 188.4 356.4 ;
      RECT  184.8 333.6 188.4 337.2 ;
      RECT  184.8 196.8 188.4 200.4 ;
      RECT  184.8 280.8 188.4 284.4 ;
      RECT  184.8 187.2 188.4 190.8 ;
      RECT  184.8 364.8 188.4 368.4 ;
      RECT  184.8 249.6 188.4 253.2 ;
      RECT  184.8 271.2 188.4 274.8 ;
      RECT  184.8 321.6 188.4 325.2 ;
      RECT  184.8 290.4 188.4 294.0 ;
      RECT  184.8 259.2 188.4 262.8 ;
      RECT  184.8 302.4 188.4 306.0 ;
      RECT  184.8 312.0 188.4 315.6 ;
      RECT  184.8 208.8 188.4 212.4 ;
      RECT  184.8 343.2 188.4 346.8 ;
      RECT  184.8 240.0 188.4 243.6 ;
      RECT  192.0 259.2 193.2 262.8 ;
      RECT  192.0 240.0 193.2 243.6 ;
      RECT  192.0 333.6 193.2 337.2 ;
      RECT  192.0 302.4 193.2 306.0 ;
      RECT  192.0 208.8 193.2 212.4 ;
      RECT  192.0 196.8 193.2 200.4 ;
      RECT  192.0 343.2 193.2 346.8 ;
      RECT  192.0 290.4 193.2 294.0 ;
      RECT  192.0 271.2 193.2 274.8 ;
      RECT  192.0 352.8 193.2 356.4 ;
      RECT  192.0 364.8 193.2 368.4 ;
      RECT  192.0 321.6 193.2 325.2 ;
      RECT  192.0 177.6 193.2 181.2 ;
      RECT  192.0 228.0 193.2 231.6 ;
      RECT  192.0 249.6 193.2 253.2 ;
      RECT  192.0 187.2 193.2 190.8 ;
      RECT  192.0 312.0 193.2 315.6 ;
      RECT  192.0 280.8 193.2 284.4 ;
      RECT  192.0 218.4 193.2 222.0 ;
      RECT  194.4 45.6 198.0 49.2 ;
      RECT  196.8 177.6 200.4 181.2 ;
      RECT  196.8 259.2 200.4 262.8 ;
      RECT  196.8 271.2 200.4 274.8 ;
      RECT  196.8 249.6 200.4 253.2 ;
      RECT  196.8 187.2 200.4 190.8 ;
      RECT  196.8 196.8 200.4 200.4 ;
      RECT  196.8 321.6 200.4 325.2 ;
      RECT  196.8 290.4 200.4 294.0 ;
      RECT  196.8 228.0 200.4 231.6 ;
      RECT  196.8 240.0 200.4 243.6 ;
      RECT  196.8 343.2 200.4 346.8 ;
      RECT  196.8 302.4 200.4 306.0 ;
      RECT  196.8 364.8 200.4 368.4 ;
      RECT  196.8 352.8 200.4 356.4 ;
      RECT  196.8 208.8 200.4 212.4 ;
      RECT  196.8 218.4 200.4 222.0 ;
      RECT  196.8 333.6 200.4 337.2 ;
      RECT  196.8 312.0 200.4 315.6 ;
      RECT  196.8 280.8 200.4 284.4 ;
      RECT  201.6 105.6 202.8 109.2 ;
      RECT  201.6 86.4 205.2 90.0 ;
      RECT  204.0 91.2 207.6 94.8 ;
      RECT  204.0 343.2 207.6 346.8 ;
      RECT  204.0 302.4 207.6 306.0 ;
      RECT  204.0 177.6 207.6 181.2 ;
      RECT  204.0 228.0 207.6 231.6 ;
      RECT  204.0 280.8 207.6 284.4 ;
      RECT  204.0 196.8 207.6 200.4 ;
      RECT  204.0 271.2 207.6 274.8 ;
      RECT  204.0 290.4 207.6 294.0 ;
      RECT  204.0 333.6 207.6 337.2 ;
      RECT  204.0 321.6 207.6 325.2 ;
      RECT  204.0 259.2 207.6 262.8 ;
      RECT  204.0 312.0 207.6 315.6 ;
      RECT  204.0 240.0 207.6 243.6 ;
      RECT  204.0 187.2 207.6 190.8 ;
      RECT  204.0 218.4 207.6 222.0 ;
      RECT  204.0 144.0 207.6 147.6 ;
      RECT  204.0 249.6 207.6 253.2 ;
      RECT  204.0 352.8 207.6 356.4 ;
      RECT  204.0 364.8 207.6 368.4 ;
      RECT  204.0 208.8 207.6 212.4 ;
      RECT  206.4 105.6 210.0 109.2 ;
      RECT  208.8 86.4 212.4 90.0 ;
      RECT  211.2 91.2 212.4 94.8 ;
      RECT  211.2 290.4 214.8 294.0 ;
      RECT  211.2 352.8 214.8 356.4 ;
      RECT  211.2 144.0 214.8 147.6 ;
      RECT  211.2 321.6 214.8 325.2 ;
      RECT  211.2 228.0 214.8 231.6 ;
      RECT  211.2 240.0 214.8 243.6 ;
      RECT  211.2 218.4 214.8 222.0 ;
      RECT  211.2 196.8 214.8 200.4 ;
      RECT  211.2 364.8 214.8 368.4 ;
      RECT  211.2 280.8 214.8 284.4 ;
      RECT  211.2 271.2 214.8 274.8 ;
      RECT  211.2 302.4 214.8 306.0 ;
      RECT  211.2 177.6 214.8 181.2 ;
      RECT  211.2 312.0 214.8 315.6 ;
      RECT  211.2 208.8 214.8 212.4 ;
      RECT  211.2 249.6 214.8 253.2 ;
      RECT  211.2 259.2 214.8 262.8 ;
      RECT  211.2 187.2 214.8 190.8 ;
      RECT  211.2 333.6 214.8 337.2 ;
      RECT  211.2 343.2 214.8 346.8 ;
      RECT  216.0 45.6 219.6 49.2 ;
      RECT  218.4 259.2 222.0 262.8 ;
      RECT  218.4 280.8 222.0 284.4 ;
      RECT  218.4 321.6 222.0 325.2 ;
      RECT  218.4 312.0 222.0 315.6 ;
      RECT  218.4 302.4 222.0 306.0 ;
      RECT  218.4 271.2 222.0 274.8 ;
      RECT  218.4 352.8 222.0 356.4 ;
      RECT  218.4 187.2 222.0 190.8 ;
      RECT  218.4 333.6 222.0 337.2 ;
      RECT  218.4 196.8 222.0 200.4 ;
      RECT  218.4 240.0 222.0 243.6 ;
      RECT  218.4 218.4 222.0 222.0 ;
      RECT  218.4 249.6 222.0 253.2 ;
      RECT  218.4 343.2 222.0 346.8 ;
      RECT  218.4 177.6 222.0 181.2 ;
      RECT  218.4 290.4 222.0 294.0 ;
      RECT  218.4 208.8 222.0 212.4 ;
      RECT  218.4 364.8 222.0 368.4 ;
      RECT  218.4 228.0 222.0 231.6 ;
      RECT  105.6 247.2 106.8 248.4 ;
      RECT  105.6 204.0 106.8 205.2 ;
      RECT  122.4 228.0 123.6 229.2 ;
      RECT  122.4 226.2 123.6 228.6 ;
      RECT  122.4 225.6 123.6 226.8 ;
      RECT  122.4 228.0 123.6 229.2 ;
      RECT  122.4 208.8 123.6 210.0 ;
      RECT  122.4 207.0 123.6 209.4 ;
      RECT  122.4 206.4 123.6 207.6 ;
      RECT  122.4 208.8 123.6 210.0 ;
      RECT  120.0 266.4 121.2 267.6 ;
      RECT  120.6 266.4 123.0 267.6 ;
      RECT  122.4 266.4 123.6 267.6 ;
      RECT  120.0 266.4 121.2 267.6 ;
      RECT  122.4 242.4 123.6 243.6 ;
      RECT  122.4 243.0 123.6 245.4 ;
      RECT  122.4 244.8 123.6 246.0 ;
      RECT  122.4 242.4 123.6 243.6 ;
      RECT  187.2 369.6 188.4 370.8 ;
      RECT  196.8 369.6 198.0 370.8 ;
      RECT  201.6 369.6 202.8 370.8 ;
      RECT  211.2 369.6 212.4 370.8 ;
      RECT  216.0 369.6 217.2 370.8 ;
      RECT  74.4 369.6 75.6 370.8 ;
      RECT  74.4 370.2 75.6 372.6 ;
      RECT  74.4 372.0 75.6 373.2 ;
      RECT  74.4 369.6 75.6 370.8 ;
      RECT  103.2 211.2 104.4 212.4 ;
      RECT  103.2 211.8 104.4 214.2 ;
      RECT  103.2 213.6 104.4 214.8 ;
      RECT  103.2 211.2 104.4 212.4 ;
      RECT  122.4 240.0 123.6 241.2 ;
      RECT  122.4 238.2 123.6 240.6 ;
      RECT  122.4 237.6 123.6 238.8 ;
      RECT  122.4 240.0 123.6 241.2 ;
      RECT  122.4 211.2 123.6 212.4 ;
      RECT  122.4 211.8 123.6 214.2 ;
      RECT  122.4 213.6 123.6 214.8 ;
      RECT  122.4 211.2 123.6 212.4 ;
      RECT  120.0 278.4 121.2 279.6 ;
      RECT  120.6 278.4 123.0 279.6 ;
      RECT  122.4 278.4 123.6 279.6 ;
      RECT  120.0 278.4 121.2 279.6 ;
      RECT  202.4 204.2 203.2 205.0 ;
      RECT  199.0 199.2 199.8 200.0 ;
      RECT  205.8 199.2 206.6 200.0 ;
      RECT  209.2 204.2 210.0 205.0 ;
      RECT  205.8 199.2 206.6 200.0 ;
      RECT  212.6 199.2 213.4 200.0 ;
      RECT  202.4 204.2 203.2 205.0 ;
      RECT  199.0 209.2 199.8 210.0 ;
      RECT  205.8 209.2 206.6 210.0 ;
      RECT  209.2 204.2 210.0 205.0 ;
      RECT  205.8 209.2 206.6 210.0 ;
      RECT  212.6 209.2 213.4 210.0 ;
      RECT  202.4 225.0 203.2 225.8 ;
      RECT  199.0 220.0 199.8 220.8 ;
      RECT  205.8 220.0 206.6 220.8 ;
      RECT  209.2 225.0 210.0 225.8 ;
      RECT  205.8 220.0 206.6 220.8 ;
      RECT  212.6 220.0 213.4 220.8 ;
      RECT  202.4 225.0 203.2 225.8 ;
      RECT  199.0 230.0 199.8 230.8 ;
      RECT  205.8 230.0 206.6 230.8 ;
      RECT  209.2 225.0 210.0 225.8 ;
      RECT  205.8 230.0 206.6 230.8 ;
      RECT  212.6 230.0 213.4 230.8 ;
      RECT  202.4 245.8 203.2 246.6 ;
      RECT  199.0 240.8 199.8 241.6 ;
      RECT  205.8 240.8 206.6 241.6 ;
      RECT  209.2 245.8 210.0 246.6 ;
      RECT  205.8 240.8 206.6 241.6 ;
      RECT  212.6 240.8 213.4 241.6 ;
      RECT  202.4 245.8 203.2 246.6 ;
      RECT  199.0 250.8 199.8 251.6 ;
      RECT  205.8 250.8 206.6 251.6 ;
      RECT  209.2 245.8 210.0 246.6 ;
      RECT  205.8 250.8 206.6 251.6 ;
      RECT  212.6 250.8 213.4 251.6 ;
      RECT  202.4 266.6 203.2 267.4 ;
      RECT  199.0 261.6 199.8 262.4 ;
      RECT  205.8 261.6 206.6 262.4 ;
      RECT  209.2 266.6 210.0 267.4 ;
      RECT  205.8 261.6 206.6 262.4 ;
      RECT  212.6 261.6 213.4 262.4 ;
      RECT  202.4 266.6 203.2 267.4 ;
      RECT  199.0 271.6 199.8 272.4 ;
      RECT  205.8 271.6 206.6 272.4 ;
      RECT  209.2 266.6 210.0 267.4 ;
      RECT  205.8 271.6 206.6 272.4 ;
      RECT  212.6 271.6 213.4 272.4 ;
      RECT  202.4 287.4 203.2 288.2 ;
      RECT  199.0 282.4 199.8 283.2 ;
      RECT  205.8 282.4 206.6 283.2 ;
      RECT  209.2 287.4 210.0 288.2 ;
      RECT  205.8 282.4 206.6 283.2 ;
      RECT  212.6 282.4 213.4 283.2 ;
      RECT  202.4 287.4 203.2 288.2 ;
      RECT  199.0 292.4 199.8 293.2 ;
      RECT  205.8 292.4 206.6 293.2 ;
      RECT  209.2 287.4 210.0 288.2 ;
      RECT  205.8 292.4 206.6 293.2 ;
      RECT  212.6 292.4 213.4 293.2 ;
      RECT  202.4 308.2 203.2 309.0 ;
      RECT  199.0 303.2 199.8 304.0 ;
      RECT  205.8 303.2 206.6 304.0 ;
      RECT  209.2 308.2 210.0 309.0 ;
      RECT  205.8 303.2 206.6 304.0 ;
      RECT  212.6 303.2 213.4 304.0 ;
      RECT  202.4 308.2 203.2 309.0 ;
      RECT  199.0 313.2 199.8 314.0 ;
      RECT  205.8 313.2 206.6 314.0 ;
      RECT  209.2 308.2 210.0 309.0 ;
      RECT  205.8 313.2 206.6 314.0 ;
      RECT  212.6 313.2 213.4 314.0 ;
      RECT  202.4 329.0 203.2 329.8 ;
      RECT  199.0 324.0 199.8 324.8 ;
      RECT  205.8 324.0 206.6 324.8 ;
      RECT  209.2 329.0 210.0 329.8 ;
      RECT  205.8 324.0 206.6 324.8 ;
      RECT  212.6 324.0 213.4 324.8 ;
      RECT  202.4 329.0 203.2 329.8 ;
      RECT  199.0 334.0 199.8 334.8 ;
      RECT  205.8 334.0 206.6 334.8 ;
      RECT  209.2 329.0 210.0 329.8 ;
      RECT  205.8 334.0 206.6 334.8 ;
      RECT  212.6 334.0 213.4 334.8 ;
      RECT  202.4 349.8 203.2 350.6 ;
      RECT  199.0 344.8 199.8 345.6 ;
      RECT  205.8 344.8 206.6 345.6 ;
      RECT  209.2 349.8 210.0 350.6 ;
      RECT  205.8 344.8 206.6 345.6 ;
      RECT  212.6 344.8 213.4 345.6 ;
      RECT  202.4 349.8 203.2 350.6 ;
      RECT  199.0 354.8 199.8 355.6 ;
      RECT  205.8 354.8 206.6 355.6 ;
      RECT  209.2 349.8 210.0 350.6 ;
      RECT  205.8 354.8 206.6 355.6 ;
      RECT  212.6 354.8 213.4 355.6 ;
      RECT  209.2 349.8 210.0 350.6 ;
      RECT  209.2 204.2 210.0 205.0 ;
      RECT  202.4 308.2 203.2 309.0 ;
      RECT  202.4 204.2 203.2 205.0 ;
      RECT  209.2 245.8 210.0 246.6 ;
      RECT  202.4 225.0 203.2 225.8 ;
      RECT  209.2 225.0 210.0 225.8 ;
      RECT  209.2 287.4 210.0 288.2 ;
      RECT  202.4 349.8 203.2 350.6 ;
      RECT  202.4 245.8 203.2 246.6 ;
      RECT  209.2 308.2 210.0 309.0 ;
      RECT  202.4 266.6 203.2 267.4 ;
      RECT  202.4 329.0 203.2 329.8 ;
      RECT  202.4 287.4 203.2 288.2 ;
      RECT  209.2 266.6 210.0 267.4 ;
      RECT  209.2 329.0 210.0 329.8 ;
      RECT  205.8 292.4 206.6 293.2 ;
      RECT  205.8 313.2 206.6 314.0 ;
      RECT  199.0 220.0 199.8 220.8 ;
      RECT  205.8 250.8 206.6 251.6 ;
      RECT  199.0 303.2 199.8 304.0 ;
      RECT  205.8 209.2 206.6 210.0 ;
      RECT  205.8 261.6 206.6 262.4 ;
      RECT  205.8 271.6 206.6 272.4 ;
      RECT  212.6 344.8 213.4 345.6 ;
      RECT  199.0 334.0 199.8 334.8 ;
      RECT  212.6 230.0 213.4 230.8 ;
      RECT  212.6 209.2 213.4 210.0 ;
      RECT  199.0 292.4 199.8 293.2 ;
      RECT  212.6 313.2 213.4 314.0 ;
      RECT  205.8 240.8 206.6 241.6 ;
      RECT  205.8 334.0 206.6 334.8 ;
      RECT  199.0 199.2 199.8 200.0 ;
      RECT  212.6 261.6 213.4 262.4 ;
      RECT  212.6 303.2 213.4 304.0 ;
      RECT  199.0 240.8 199.8 241.6 ;
      RECT  205.8 220.0 206.6 220.8 ;
      RECT  199.0 230.0 199.8 230.8 ;
      RECT  199.0 344.8 199.8 345.6 ;
      RECT  205.8 344.8 206.6 345.6 ;
      RECT  205.8 324.0 206.6 324.8 ;
      RECT  212.6 250.8 213.4 251.6 ;
      RECT  205.8 303.2 206.6 304.0 ;
      RECT  212.6 199.2 213.4 200.0 ;
      RECT  199.0 271.6 199.8 272.4 ;
      RECT  199.0 324.0 199.8 324.8 ;
      RECT  199.0 354.8 199.8 355.6 ;
      RECT  205.8 354.8 206.6 355.6 ;
      RECT  205.8 230.0 206.6 230.8 ;
      RECT  212.6 271.6 213.4 272.4 ;
      RECT  199.0 261.6 199.8 262.4 ;
      RECT  212.6 334.0 213.4 334.8 ;
      RECT  205.8 282.4 206.6 283.2 ;
      RECT  199.0 282.4 199.8 283.2 ;
      RECT  205.8 199.2 206.6 200.0 ;
      RECT  212.6 240.8 213.4 241.6 ;
      RECT  212.6 354.8 213.4 355.6 ;
      RECT  199.0 209.2 199.8 210.0 ;
      RECT  212.6 292.4 213.4 293.2 ;
      RECT  212.6 220.0 213.4 220.8 ;
      RECT  212.6 324.0 213.4 324.8 ;
      RECT  199.0 250.8 199.8 251.6 ;
      RECT  199.0 313.2 199.8 314.0 ;
      RECT  212.6 282.4 213.4 283.2 ;
      RECT  202.4 184.2 203.2 183.4 ;
      RECT  199.0 189.2 199.8 188.4 ;
      RECT  205.8 189.2 206.6 188.4 ;
      RECT  209.2 184.2 210.0 183.4 ;
      RECT  205.8 189.2 206.6 188.4 ;
      RECT  212.6 189.2 213.4 188.4 ;
      RECT  209.2 184.2 210.0 183.4 ;
      RECT  202.4 184.2 203.2 183.4 ;
      RECT  212.6 189.2 213.4 188.4 ;
      RECT  205.8 189.2 206.6 188.4 ;
      RECT  199.0 189.2 199.8 188.4 ;
      RECT  202.4 183.4 203.2 184.2 ;
      RECT  199.0 178.4 199.8 179.2 ;
      RECT  205.8 178.4 206.6 179.2 ;
      RECT  209.2 183.4 210.0 184.2 ;
      RECT  205.8 178.4 206.6 179.2 ;
      RECT  212.6 178.4 213.4 179.2 ;
      RECT  209.2 183.4 210.0 184.2 ;
      RECT  202.4 183.4 203.2 184.2 ;
      RECT  212.6 178.4 213.4 179.2 ;
      RECT  205.8 178.4 206.6 179.2 ;
      RECT  199.0 178.4 199.8 179.2 ;
      RECT  202.4 370.6 203.2 371.4 ;
      RECT  199.0 365.6 199.8 366.4 ;
      RECT  205.8 365.6 206.6 366.4 ;
      RECT  209.2 370.6 210.0 371.4 ;
      RECT  205.8 365.6 206.6 366.4 ;
      RECT  212.6 365.6 213.4 366.4 ;
      RECT  209.2 370.6 210.0 371.4 ;
      RECT  202.4 370.6 203.2 371.4 ;
      RECT  212.6 365.6 213.4 366.4 ;
      RECT  205.8 365.6 206.6 366.4 ;
      RECT  199.0 365.6 199.8 366.4 ;
      RECT  188.8 183.4 189.6 184.2 ;
      RECT  185.4 178.4 186.2 179.2 ;
      RECT  192.2 178.4 193.0 179.2 ;
      RECT  188.8 183.4 189.6 184.2 ;
      RECT  185.4 188.4 186.2 189.2 ;
      RECT  192.2 188.4 193.0 189.2 ;
      RECT  188.8 204.2 189.6 205.0 ;
      RECT  185.4 199.2 186.2 200.0 ;
      RECT  192.2 199.2 193.0 200.0 ;
      RECT  188.8 204.2 189.6 205.0 ;
      RECT  185.4 209.2 186.2 210.0 ;
      RECT  192.2 209.2 193.0 210.0 ;
      RECT  188.8 225.0 189.6 225.8 ;
      RECT  185.4 220.0 186.2 220.8 ;
      RECT  192.2 220.0 193.0 220.8 ;
      RECT  188.8 225.0 189.6 225.8 ;
      RECT  185.4 230.0 186.2 230.8 ;
      RECT  192.2 230.0 193.0 230.8 ;
      RECT  188.8 245.8 189.6 246.6 ;
      RECT  185.4 240.8 186.2 241.6 ;
      RECT  192.2 240.8 193.0 241.6 ;
      RECT  188.8 245.8 189.6 246.6 ;
      RECT  185.4 250.8 186.2 251.6 ;
      RECT  192.2 250.8 193.0 251.6 ;
      RECT  188.8 266.6 189.6 267.4 ;
      RECT  185.4 261.6 186.2 262.4 ;
      RECT  192.2 261.6 193.0 262.4 ;
      RECT  188.8 266.6 189.6 267.4 ;
      RECT  185.4 271.6 186.2 272.4 ;
      RECT  192.2 271.6 193.0 272.4 ;
      RECT  188.8 287.4 189.6 288.2 ;
      RECT  185.4 282.4 186.2 283.2 ;
      RECT  192.2 282.4 193.0 283.2 ;
      RECT  188.8 287.4 189.6 288.2 ;
      RECT  185.4 292.4 186.2 293.2 ;
      RECT  192.2 292.4 193.0 293.2 ;
      RECT  188.8 308.2 189.6 309.0 ;
      RECT  185.4 303.2 186.2 304.0 ;
      RECT  192.2 303.2 193.0 304.0 ;
      RECT  188.8 308.2 189.6 309.0 ;
      RECT  185.4 313.2 186.2 314.0 ;
      RECT  192.2 313.2 193.0 314.0 ;
      RECT  188.8 329.0 189.6 329.8 ;
      RECT  185.4 324.0 186.2 324.8 ;
      RECT  192.2 324.0 193.0 324.8 ;
      RECT  188.8 329.0 189.6 329.8 ;
      RECT  185.4 334.0 186.2 334.8 ;
      RECT  192.2 334.0 193.0 334.8 ;
      RECT  188.8 349.8 189.6 350.6 ;
      RECT  185.4 344.8 186.2 345.6 ;
      RECT  192.2 344.8 193.0 345.6 ;
      RECT  188.8 349.8 189.6 350.6 ;
      RECT  185.4 354.8 186.2 355.6 ;
      RECT  192.2 354.8 193.0 355.6 ;
      RECT  188.8 370.6 189.6 371.4 ;
      RECT  185.4 365.6 186.2 366.4 ;
      RECT  192.2 365.6 193.0 366.4 ;
      RECT  188.8 287.4 189.6 288.2 ;
      RECT  188.8 183.4 189.6 184.2 ;
      RECT  188.8 204.2 189.6 205.0 ;
      RECT  188.8 329.0 189.6 329.8 ;
      RECT  188.8 349.8 189.6 350.6 ;
      RECT  188.8 225.0 189.6 225.8 ;
      RECT  188.8 370.6 189.6 371.4 ;
      RECT  188.8 245.8 189.6 246.6 ;
      RECT  188.8 308.2 189.6 309.0 ;
      RECT  188.8 266.6 189.6 267.4 ;
      RECT  192.2 271.6 193.0 272.4 ;
      RECT  192.2 292.4 193.0 293.2 ;
      RECT  185.4 199.2 186.2 200.0 ;
      RECT  192.2 230.0 193.0 230.8 ;
      RECT  185.4 282.4 186.2 283.2 ;
      RECT  192.2 188.4 193.0 189.2 ;
      RECT  192.2 344.8 193.0 345.6 ;
      RECT  192.2 240.8 193.0 241.6 ;
      RECT  192.2 250.8 193.0 251.6 ;
      RECT  192.2 365.6 193.0 366.4 ;
      RECT  185.4 271.6 186.2 272.4 ;
      RECT  192.2 220.0 193.0 220.8 ;
      RECT  192.2 313.2 193.0 314.0 ;
      RECT  192.2 354.8 193.0 355.6 ;
      RECT  185.4 178.4 186.2 179.2 ;
      RECT  185.4 220.0 186.2 220.8 ;
      RECT  192.2 199.2 193.0 200.0 ;
      RECT  185.4 209.2 186.2 210.0 ;
      RECT  185.4 324.0 186.2 324.8 ;
      RECT  192.2 324.0 193.0 324.8 ;
      RECT  192.2 303.2 193.0 304.0 ;
      RECT  185.4 365.6 186.2 366.4 ;
      RECT  192.2 282.4 193.0 283.2 ;
      RECT  185.4 344.8 186.2 345.6 ;
      RECT  185.4 303.2 186.2 304.0 ;
      RECT  185.4 250.8 186.2 251.6 ;
      RECT  185.4 334.0 186.2 334.8 ;
      RECT  192.2 334.0 193.0 334.8 ;
      RECT  192.2 209.2 193.0 210.0 ;
      RECT  185.4 240.8 186.2 241.6 ;
      RECT  192.2 261.6 193.0 262.4 ;
      RECT  185.4 261.6 186.2 262.4 ;
      RECT  192.2 178.4 193.0 179.2 ;
      RECT  185.4 188.4 186.2 189.2 ;
      RECT  185.4 354.8 186.2 355.6 ;
      RECT  185.4 230.0 186.2 230.8 ;
      RECT  185.4 292.4 186.2 293.2 ;
      RECT  185.4 313.2 186.2 314.0 ;
      RECT  216.0 183.4 216.8 184.2 ;
      RECT  212.6 178.4 213.4 179.2 ;
      RECT  219.4 178.4 220.2 179.2 ;
      RECT  216.0 183.4 216.8 184.2 ;
      RECT  212.6 188.4 213.4 189.2 ;
      RECT  219.4 188.4 220.2 189.2 ;
      RECT  216.0 204.2 216.8 205.0 ;
      RECT  212.6 199.2 213.4 200.0 ;
      RECT  219.4 199.2 220.2 200.0 ;
      RECT  216.0 204.2 216.8 205.0 ;
      RECT  212.6 209.2 213.4 210.0 ;
      RECT  219.4 209.2 220.2 210.0 ;
      RECT  216.0 225.0 216.8 225.8 ;
      RECT  212.6 220.0 213.4 220.8 ;
      RECT  219.4 220.0 220.2 220.8 ;
      RECT  216.0 225.0 216.8 225.8 ;
      RECT  212.6 230.0 213.4 230.8 ;
      RECT  219.4 230.0 220.2 230.8 ;
      RECT  216.0 245.8 216.8 246.6 ;
      RECT  212.6 240.8 213.4 241.6 ;
      RECT  219.4 240.8 220.2 241.6 ;
      RECT  216.0 245.8 216.8 246.6 ;
      RECT  212.6 250.8 213.4 251.6 ;
      RECT  219.4 250.8 220.2 251.6 ;
      RECT  216.0 266.6 216.8 267.4 ;
      RECT  212.6 261.6 213.4 262.4 ;
      RECT  219.4 261.6 220.2 262.4 ;
      RECT  216.0 266.6 216.8 267.4 ;
      RECT  212.6 271.6 213.4 272.4 ;
      RECT  219.4 271.6 220.2 272.4 ;
      RECT  216.0 287.4 216.8 288.2 ;
      RECT  212.6 282.4 213.4 283.2 ;
      RECT  219.4 282.4 220.2 283.2 ;
      RECT  216.0 287.4 216.8 288.2 ;
      RECT  212.6 292.4 213.4 293.2 ;
      RECT  219.4 292.4 220.2 293.2 ;
      RECT  216.0 308.2 216.8 309.0 ;
      RECT  212.6 303.2 213.4 304.0 ;
      RECT  219.4 303.2 220.2 304.0 ;
      RECT  216.0 308.2 216.8 309.0 ;
      RECT  212.6 313.2 213.4 314.0 ;
      RECT  219.4 313.2 220.2 314.0 ;
      RECT  216.0 329.0 216.8 329.8 ;
      RECT  212.6 324.0 213.4 324.8 ;
      RECT  219.4 324.0 220.2 324.8 ;
      RECT  216.0 329.0 216.8 329.8 ;
      RECT  212.6 334.0 213.4 334.8 ;
      RECT  219.4 334.0 220.2 334.8 ;
      RECT  216.0 349.8 216.8 350.6 ;
      RECT  212.6 344.8 213.4 345.6 ;
      RECT  219.4 344.8 220.2 345.6 ;
      RECT  216.0 349.8 216.8 350.6 ;
      RECT  212.6 354.8 213.4 355.6 ;
      RECT  219.4 354.8 220.2 355.6 ;
      RECT  216.0 370.6 216.8 371.4 ;
      RECT  212.6 365.6 213.4 366.4 ;
      RECT  219.4 365.6 220.2 366.4 ;
      RECT  216.0 287.4 216.8 288.2 ;
      RECT  216.0 183.4 216.8 184.2 ;
      RECT  216.0 204.2 216.8 205.0 ;
      RECT  216.0 329.0 216.8 329.8 ;
      RECT  216.0 349.8 216.8 350.6 ;
      RECT  216.0 225.0 216.8 225.8 ;
      RECT  216.0 370.6 216.8 371.4 ;
      RECT  216.0 245.8 216.8 246.6 ;
      RECT  216.0 308.2 216.8 309.0 ;
      RECT  216.0 266.6 216.8 267.4 ;
      RECT  219.4 271.6 220.2 272.4 ;
      RECT  219.4 292.4 220.2 293.2 ;
      RECT  212.6 199.2 213.4 200.0 ;
      RECT  219.4 230.0 220.2 230.8 ;
      RECT  212.6 282.4 213.4 283.2 ;
      RECT  219.4 188.4 220.2 189.2 ;
      RECT  219.4 344.8 220.2 345.6 ;
      RECT  219.4 240.8 220.2 241.6 ;
      RECT  219.4 250.8 220.2 251.6 ;
      RECT  219.4 365.6 220.2 366.4 ;
      RECT  212.6 271.6 213.4 272.4 ;
      RECT  219.4 220.0 220.2 220.8 ;
      RECT  219.4 313.2 220.2 314.0 ;
      RECT  219.4 354.8 220.2 355.6 ;
      RECT  212.6 178.4 213.4 179.2 ;
      RECT  212.6 220.0 213.4 220.8 ;
      RECT  219.4 199.2 220.2 200.0 ;
      RECT  212.6 209.2 213.4 210.0 ;
      RECT  212.6 324.0 213.4 324.8 ;
      RECT  219.4 324.0 220.2 324.8 ;
      RECT  219.4 303.2 220.2 304.0 ;
      RECT  212.6 365.6 213.4 366.4 ;
      RECT  219.4 282.4 220.2 283.2 ;
      RECT  212.6 344.8 213.4 345.6 ;
      RECT  212.6 303.2 213.4 304.0 ;
      RECT  212.6 250.8 213.4 251.6 ;
      RECT  212.6 334.0 213.4 334.8 ;
      RECT  219.4 334.0 220.2 334.8 ;
      RECT  219.4 209.2 220.2 210.0 ;
      RECT  212.6 240.8 213.4 241.6 ;
      RECT  219.4 261.6 220.2 262.4 ;
      RECT  212.6 261.6 213.4 262.4 ;
      RECT  219.4 178.4 220.2 179.2 ;
      RECT  212.6 188.4 213.4 189.2 ;
      RECT  212.6 354.8 213.4 355.6 ;
      RECT  212.6 230.0 213.4 230.8 ;
      RECT  212.6 292.4 213.4 293.2 ;
      RECT  212.6 313.2 213.4 314.0 ;
      RECT  195.6 266.6 196.4 267.4 ;
      RECT  195.6 183.4 196.4 184.2 ;
      RECT  195.6 287.4 196.4 288.2 ;
      RECT  195.6 225.0 196.4 225.8 ;
      RECT  195.6 370.6 196.4 371.4 ;
      RECT  195.6 245.8 196.4 246.6 ;
      RECT  195.6 349.8 196.4 350.6 ;
      RECT  195.6 204.2 196.4 205.0 ;
      RECT  195.6 329.0 196.4 329.8 ;
      RECT  195.6 308.2 196.4 309.0 ;
      RECT  199.0 261.6 199.8 262.4 ;
      RECT  192.2 250.8 193.0 251.6 ;
      RECT  192.2 261.6 193.0 262.4 ;
      RECT  192.2 230.0 193.0 230.8 ;
      RECT  199.0 282.4 199.8 283.2 ;
      RECT  199.0 365.6 199.8 366.4 ;
      RECT  199.0 188.4 199.8 189.2 ;
      RECT  192.2 209.2 193.0 210.0 ;
      RECT  192.2 365.6 193.0 366.4 ;
      RECT  192.2 313.2 193.0 314.0 ;
      RECT  199.0 271.6 199.8 272.4 ;
      RECT  199.0 292.4 199.8 293.2 ;
      RECT  199.0 344.8 199.8 345.6 ;
      RECT  199.0 199.2 199.8 200.0 ;
      RECT  199.0 250.8 199.8 251.6 ;
      RECT  192.2 271.6 193.0 272.4 ;
      RECT  199.0 313.2 199.8 314.0 ;
      RECT  192.2 240.8 193.0 241.6 ;
      RECT  192.2 178.4 193.0 179.2 ;
      RECT  192.2 303.2 193.0 304.0 ;
      RECT  199.0 354.8 199.8 355.6 ;
      RECT  192.2 220.0 193.0 220.8 ;
      RECT  192.2 282.4 193.0 283.2 ;
      RECT  199.0 303.2 199.8 304.0 ;
      RECT  199.0 178.4 199.8 179.2 ;
      RECT  199.0 240.8 199.8 241.6 ;
      RECT  199.0 220.0 199.8 220.8 ;
      RECT  192.2 334.0 193.0 334.8 ;
      RECT  199.0 230.0 199.8 230.8 ;
      RECT  192.2 188.4 193.0 189.2 ;
      RECT  192.2 292.4 193.0 293.2 ;
      RECT  192.2 324.0 193.0 324.8 ;
      RECT  199.0 334.0 199.8 334.8 ;
      RECT  192.2 199.2 193.0 200.0 ;
      RECT  199.0 324.0 199.8 324.8 ;
      RECT  192.2 344.8 193.0 345.6 ;
      RECT  199.0 209.2 199.8 210.0 ;
      RECT  192.2 354.8 193.0 355.6 ;
      RECT  188.9 204.3 189.5 204.9 ;
      RECT  209.3 370.7 209.9 371.3 ;
      RECT  188.9 225.1 189.5 225.7 ;
      RECT  216.1 266.7 216.7 267.3 ;
      RECT  216.1 329.1 216.7 329.7 ;
      RECT  216.1 349.9 216.7 350.5 ;
      RECT  216.1 225.1 216.7 225.7 ;
      RECT  195.6 370.6 196.4 371.4 ;
      RECT  202.5 370.7 203.1 371.3 ;
      RECT  209.3 183.5 209.9 184.1 ;
      RECT  195.6 204.2 196.4 205.0 ;
      RECT  216.1 370.7 216.7 371.3 ;
      RECT  202.5 266.7 203.1 267.3 ;
      RECT  209.3 266.7 209.9 267.3 ;
      RECT  202.5 245.9 203.1 246.5 ;
      RECT  216.1 183.5 216.7 184.1 ;
      RECT  209.3 225.1 209.9 225.7 ;
      RECT  202.5 329.1 203.1 329.7 ;
      RECT  202.5 204.3 203.1 204.9 ;
      RECT  209.3 308.3 209.9 308.9 ;
      RECT  188.9 370.7 189.5 371.3 ;
      RECT  216.1 308.3 216.7 308.9 ;
      RECT  188.9 266.7 189.5 267.3 ;
      RECT  209.3 349.9 209.9 350.5 ;
      RECT  195.6 308.2 196.4 309.0 ;
      RECT  202.5 287.5 203.1 288.1 ;
      RECT  216.1 287.5 216.7 288.1 ;
      RECT  195.6 349.8 196.4 350.6 ;
      RECT  188.9 245.9 189.5 246.5 ;
      RECT  216.1 245.9 216.7 246.5 ;
      RECT  195.6 266.6 196.4 267.4 ;
      RECT  209.3 329.1 209.9 329.7 ;
      RECT  188.9 183.5 189.5 184.1 ;
      RECT  195.6 287.4 196.4 288.2 ;
      RECT  188.9 287.5 189.5 288.1 ;
      RECT  202.5 308.3 203.1 308.9 ;
      RECT  195.6 329.0 196.4 329.8 ;
      RECT  195.6 183.4 196.4 184.2 ;
      RECT  216.1 204.3 216.7 204.9 ;
      RECT  209.3 245.9 209.9 246.5 ;
      RECT  188.9 329.1 189.5 329.7 ;
      RECT  202.5 225.1 203.1 225.7 ;
      RECT  195.6 225.0 196.4 225.8 ;
      RECT  202.5 183.5 203.1 184.1 ;
      RECT  188.9 349.9 189.5 350.5 ;
      RECT  202.5 349.9 203.1 350.5 ;
      RECT  209.3 204.3 209.9 204.9 ;
      RECT  209.3 287.5 209.9 288.1 ;
      RECT  195.6 245.8 196.4 246.6 ;
      RECT  188.9 308.3 189.5 308.9 ;
      RECT  192.2 292.4 193.0 293.2 ;
      RECT  192.2 344.8 193.0 345.6 ;
      RECT  219.5 354.9 220.1 355.5 ;
      RECT  192.2 230.0 193.0 230.8 ;
      RECT  192.2 188.4 193.0 189.2 ;
      RECT  192.3 199.3 192.9 199.9 ;
      RECT  192.3 324.1 192.9 324.7 ;
      RECT  219.5 178.5 220.1 179.1 ;
      RECT  205.9 324.1 206.5 324.7 ;
      RECT  205.9 282.5 206.5 283.1 ;
      RECT  199.1 209.3 199.7 209.9 ;
      RECT  205.9 344.9 206.5 345.5 ;
      RECT  205.9 209.3 206.5 209.9 ;
      RECT  192.2 199.2 193.0 200.0 ;
      RECT  212.7 199.3 213.3 199.9 ;
      RECT  199.1 188.5 199.7 189.1 ;
      RECT  192.2 303.2 193.0 304.0 ;
      RECT  219.5 313.3 220.1 313.9 ;
      RECT  199.0 230.0 199.8 230.8 ;
      RECT  212.7 188.5 213.3 189.1 ;
      RECT  192.3 334.1 192.9 334.7 ;
      RECT  192.3 209.3 192.9 209.9 ;
      RECT  205.9 313.3 206.5 313.9 ;
      RECT  185.5 282.5 186.1 283.1 ;
      RECT  205.9 354.9 206.5 355.5 ;
      RECT  199.1 199.3 199.7 199.9 ;
      RECT  219.5 324.1 220.1 324.7 ;
      RECT  185.5 334.1 186.1 334.7 ;
      RECT  199.0 334.0 199.8 334.8 ;
      RECT  199.1 303.3 199.7 303.9 ;
      RECT  219.5 240.9 220.1 241.5 ;
      RECT  219.5 344.9 220.1 345.5 ;
      RECT  192.3 292.5 192.9 293.1 ;
      RECT  199.0 271.6 199.8 272.4 ;
      RECT  212.7 209.3 213.3 209.9 ;
      RECT  212.7 313.3 213.3 313.9 ;
      RECT  185.5 324.1 186.1 324.7 ;
      RECT  212.7 292.5 213.3 293.1 ;
      RECT  219.5 282.5 220.1 283.1 ;
      RECT  219.5 365.7 220.1 366.3 ;
      RECT  212.7 178.5 213.3 179.1 ;
      RECT  192.3 250.9 192.9 251.5 ;
      RECT  199.0 209.2 199.8 210.0 ;
      RECT  205.9 240.9 206.5 241.5 ;
      RECT  185.5 354.9 186.1 355.5 ;
      RECT  199.0 292.4 199.8 293.2 ;
      RECT  185.5 199.3 186.1 199.9 ;
      RECT  199.0 240.8 199.8 241.6 ;
      RECT  192.3 282.5 192.9 283.1 ;
      RECT  185.5 344.9 186.1 345.5 ;
      RECT  192.2 209.2 193.0 210.0 ;
      RECT  205.9 178.5 206.5 179.1 ;
      RECT  199.1 313.3 199.7 313.9 ;
      RECT  205.9 220.1 206.5 220.7 ;
      RECT  219.5 334.1 220.1 334.7 ;
      RECT  185.5 271.7 186.1 272.3 ;
      RECT  192.2 178.4 193.0 179.2 ;
      RECT  199.1 354.9 199.7 355.5 ;
      RECT  185.5 313.3 186.1 313.9 ;
      RECT  199.1 365.7 199.7 366.3 ;
      RECT  205.9 199.3 206.5 199.9 ;
      RECT  212.7 354.9 213.3 355.5 ;
      RECT  185.5 292.5 186.1 293.1 ;
      RECT  199.0 344.8 199.8 345.6 ;
      RECT  192.2 271.6 193.0 272.4 ;
      RECT  199.0 324.0 199.8 324.8 ;
      RECT  212.7 303.3 213.3 303.9 ;
      RECT  199.1 261.7 199.7 262.3 ;
      RECT  212.7 271.7 213.3 272.3 ;
      RECT  192.3 365.7 192.9 366.3 ;
      RECT  185.5 230.1 186.1 230.7 ;
      RECT  192.2 313.2 193.0 314.0 ;
      RECT  192.2 354.8 193.0 355.6 ;
      RECT  185.5 209.3 186.1 209.9 ;
      RECT  199.0 282.4 199.8 283.2 ;
      RECT  205.9 188.5 206.5 189.1 ;
      RECT  192.3 220.1 192.9 220.7 ;
      RECT  192.3 344.9 192.9 345.5 ;
      RECT  192.2 324.0 193.0 324.8 ;
      RECT  199.1 292.5 199.7 293.1 ;
      RECT  192.2 282.4 193.0 283.2 ;
      RECT  192.3 230.1 192.9 230.7 ;
      RECT  192.3 271.7 192.9 272.3 ;
      RECT  185.5 188.5 186.1 189.1 ;
      RECT  199.0 354.8 199.8 355.6 ;
      RECT  205.9 365.7 206.5 366.3 ;
      RECT  205.9 230.1 206.5 230.7 ;
      RECT  192.3 178.5 192.9 179.1 ;
      RECT  199.0 250.8 199.8 251.6 ;
      RECT  205.9 334.1 206.5 334.7 ;
      RECT  199.1 178.5 199.7 179.1 ;
      RECT  212.7 324.1 213.3 324.7 ;
      RECT  192.2 261.6 193.0 262.4 ;
      RECT  185.5 365.7 186.1 366.3 ;
      RECT  185.5 178.5 186.1 179.1 ;
      RECT  205.9 250.9 206.5 251.5 ;
      RECT  199.0 220.0 199.8 220.8 ;
      RECT  212.7 365.7 213.3 366.3 ;
      RECT  219.5 271.7 220.1 272.3 ;
      RECT  199.1 282.5 199.7 283.1 ;
      RECT  192.3 313.3 192.9 313.9 ;
      RECT  212.7 334.1 213.3 334.7 ;
      RECT  199.0 303.2 199.8 304.0 ;
      RECT  219.5 261.7 220.1 262.3 ;
      RECT  219.5 250.9 220.1 251.5 ;
      RECT  219.5 220.1 220.1 220.7 ;
      RECT  185.5 303.3 186.1 303.9 ;
      RECT  205.9 271.7 206.5 272.3 ;
      RECT  192.2 240.8 193.0 241.6 ;
      RECT  199.1 271.7 199.7 272.3 ;
      RECT  192.2 250.8 193.0 251.6 ;
      RECT  212.7 344.9 213.3 345.5 ;
      RECT  192.3 354.9 192.9 355.5 ;
      RECT  192.2 365.6 193.0 366.4 ;
      RECT  212.7 230.1 213.3 230.7 ;
      RECT  199.1 334.1 199.7 334.7 ;
      RECT  219.5 303.3 220.1 303.9 ;
      RECT  192.3 261.7 192.9 262.3 ;
      RECT  199.0 188.4 199.8 189.2 ;
      RECT  192.2 220.0 193.0 220.8 ;
      RECT  185.5 240.9 186.1 241.5 ;
      RECT  212.7 250.9 213.3 251.5 ;
      RECT  219.5 188.5 220.1 189.1 ;
      RECT  219.5 199.3 220.1 199.9 ;
      RECT  199.1 344.9 199.7 345.5 ;
      RECT  192.3 303.3 192.9 303.9 ;
      RECT  212.7 282.5 213.3 283.1 ;
      RECT  199.1 250.9 199.7 251.5 ;
      RECT  192.3 240.9 192.9 241.5 ;
      RECT  185.5 250.9 186.1 251.5 ;
      RECT  199.1 240.9 199.7 241.5 ;
      RECT  199.1 220.1 199.7 220.7 ;
      RECT  219.5 209.3 220.1 209.9 ;
      RECT  199.0 178.4 199.8 179.2 ;
      RECT  185.5 220.1 186.1 220.7 ;
      RECT  192.2 334.0 193.0 334.8 ;
      RECT  212.7 240.9 213.3 241.5 ;
      RECT  205.9 292.5 206.5 293.1 ;
      RECT  199.1 324.1 199.7 324.7 ;
      RECT  199.1 230.1 199.7 230.7 ;
      RECT  199.0 313.2 199.8 314.0 ;
      RECT  185.5 261.7 186.1 262.3 ;
      RECT  205.9 303.3 206.5 303.9 ;
      RECT  219.5 292.5 220.1 293.1 ;
      RECT  199.0 365.6 199.8 366.4 ;
      RECT  199.0 199.2 199.8 200.0 ;
      RECT  212.7 261.7 213.3 262.3 ;
      RECT  212.7 220.1 213.3 220.7 ;
      RECT  192.3 188.5 192.9 189.1 ;
      RECT  219.5 230.1 220.1 230.7 ;
      RECT  205.9 261.7 206.5 262.3 ;
      RECT  199.0 261.6 199.8 262.4 ;
      RECT  195.4 163.0 196.2 163.8 ;
      RECT  195.4 163.0 196.2 163.8 ;
      RECT  202.2 163.0 203.0 163.8 ;
      RECT  202.2 163.0 203.0 163.8 ;
      RECT  209.0 163.0 209.8 163.8 ;
      RECT  209.0 163.0 209.8 163.8 ;
      RECT  202.2 163.0 203.0 163.8 ;
      RECT  195.4 163.0 196.2 163.8 ;
      RECT  209.0 163.0 209.8 163.8 ;
      RECT  205.8 146.0 206.6 146.8 ;
      RECT  204.8 132.6 205.6 133.4 ;
      RECT  212.6 146.0 213.4 146.8 ;
      RECT  211.6 132.6 212.4 133.4 ;
      RECT  211.7 132.7 212.3 133.3 ;
      RECT  204.9 132.7 205.5 133.3 ;
      RECT  212.7 146.1 213.3 146.7 ;
      RECT  205.9 146.1 206.5 146.7 ;
      RECT  203.2 81.2 204.0 82.0 ;
      RECT  202.6 98.6 203.4 99.4 ;
      RECT  203.2 87.8 204.0 88.6 ;
      RECT  204.6 92.2 205.4 93.0 ;
      RECT  201.8 106.8 202.6 107.6 ;
      RECT  210.0 81.2 210.8 82.0 ;
      RECT  209.4 98.6 210.2 99.4 ;
      RECT  210.0 87.8 210.8 88.6 ;
      RECT  211.4 92.2 212.2 93.0 ;
      RECT  208.6 106.8 209.4 107.6 ;
      RECT  210.1 81.3 210.7 81.9 ;
      RECT  209.5 98.7 210.1 99.3 ;
      RECT  202.7 98.7 203.3 99.3 ;
      RECT  203.3 81.3 203.9 81.9 ;
      RECT  208.7 106.9 209.3 107.5 ;
      RECT  201.9 106.9 202.5 107.5 ;
      RECT  204.7 92.3 205.3 92.9 ;
      RECT  210.1 87.9 210.7 88.5 ;
      RECT  203.3 87.9 203.9 88.5 ;
      RECT  211.5 92.3 212.1 92.9 ;
      RECT  204.9 133.3 205.5 132.7 ;
      RECT  202.2 163.8 203.0 163.0 ;
      RECT  203.3 81.9 203.9 81.3 ;
      RECT  210.1 81.9 210.7 81.3 ;
      RECT  195.4 163.8 196.2 163.0 ;
      RECT  209.0 163.8 209.8 163.0 ;
      RECT  211.7 133.3 212.3 132.7 ;
      RECT  209.5 99.3 210.1 98.7 ;
      RECT  202.7 99.3 203.3 98.7 ;
      RECT  201.9 107.5 202.5 106.9 ;
      RECT  205.9 146.7 206.5 146.1 ;
      RECT  208.7 107.5 209.3 106.9 ;
      RECT  212.7 146.7 213.3 146.1 ;
      RECT  204.7 92.9 205.3 92.3 ;
      RECT  211.5 92.9 212.1 92.3 ;
      RECT  210.1 88.5 210.7 87.9 ;
      RECT  203.3 88.5 203.9 87.9 ;
      RECT  89.8 205.9 97.1 206.5 ;
      RECT  91.2 216.3 98.5 216.9 ;
      RECT  92.6 247.5 97.1 248.1 ;
      RECT  94.0 257.9 98.5 258.5 ;
      RECT  127.2 204.5 130.7 205.1 ;
      RECT  127.2 215.3 132.1 215.9 ;
      RECT  127.2 225.3 133.5 225.9 ;
      RECT  127.2 236.1 134.9 236.7 ;
      RECT  127.2 246.1 136.3 246.7 ;
      RECT  127.2 256.9 137.7 257.5 ;
      RECT  127.2 266.9 139.1 267.5 ;
      RECT  127.2 277.7 140.5 278.3 ;
      RECT  105.3 204.6 106.1 205.4 ;
      RECT  122.7 204.6 123.5 205.4 ;
      RECT  105.3 194.2 106.1 195.0 ;
      RECT  122.7 194.2 123.5 195.0 ;
      RECT  105.3 204.6 106.1 205.4 ;
      RECT  122.7 204.6 123.5 205.4 ;
      RECT  105.3 215.0 106.1 215.8 ;
      RECT  122.7 215.0 123.5 215.8 ;
      RECT  105.3 225.4 106.1 226.2 ;
      RECT  122.7 225.4 123.5 226.2 ;
      RECT  105.3 215.0 106.1 215.8 ;
      RECT  122.7 215.0 123.5 215.8 ;
      RECT  105.3 225.4 106.1 226.2 ;
      RECT  122.7 225.4 123.5 226.2 ;
      RECT  105.3 235.8 106.1 236.6 ;
      RECT  122.7 235.8 123.5 236.6 ;
      RECT  105.3 204.6 106.1 205.4 ;
      RECT  105.3 225.4 106.1 226.2 ;
      RECT  122.7 225.4 123.5 226.2 ;
      RECT  122.7 204.6 123.5 205.4 ;
      RECT  105.3 215.0 106.1 215.8 ;
      RECT  105.3 194.2 106.1 195.0 ;
      RECT  105.3 235.8 106.1 236.6 ;
      RECT  122.7 194.2 123.5 195.0 ;
      RECT  122.7 215.0 123.5 215.8 ;
      RECT  122.7 235.8 123.5 236.6 ;
      RECT  105.3 246.2 106.1 247.0 ;
      RECT  122.7 246.2 123.5 247.0 ;
      RECT  105.3 235.8 106.1 236.6 ;
      RECT  122.7 235.8 123.5 236.6 ;
      RECT  105.3 246.2 106.1 247.0 ;
      RECT  122.7 246.2 123.5 247.0 ;
      RECT  105.3 256.6 106.1 257.4 ;
      RECT  122.7 256.6 123.5 257.4 ;
      RECT  105.3 267.0 106.1 267.8 ;
      RECT  122.7 267.0 123.5 267.8 ;
      RECT  105.3 256.6 106.1 257.4 ;
      RECT  122.7 256.6 123.5 257.4 ;
      RECT  105.3 267.0 106.1 267.8 ;
      RECT  122.7 267.0 123.5 267.8 ;
      RECT  105.3 277.4 106.1 278.2 ;
      RECT  122.7 277.4 123.5 278.2 ;
      RECT  105.3 246.2 106.1 247.0 ;
      RECT  105.3 267.0 106.1 267.8 ;
      RECT  122.7 267.0 123.5 267.8 ;
      RECT  122.7 246.2 123.5 247.0 ;
      RECT  105.3 256.6 106.1 257.4 ;
      RECT  105.3 235.8 106.1 236.6 ;
      RECT  105.3 277.4 106.1 278.2 ;
      RECT  122.7 235.8 123.5 236.6 ;
      RECT  122.7 256.6 123.5 257.4 ;
      RECT  122.7 277.4 123.5 278.2 ;
      RECT  96.7 205.8 97.5 206.6 ;
      RECT  89.4 205.8 90.2 206.6 ;
      RECT  98.1 216.2 98.9 217.0 ;
      RECT  90.8 216.2 91.6 217.0 ;
      RECT  96.7 247.4 97.5 248.2 ;
      RECT  92.2 247.4 93.0 248.2 ;
      RECT  98.1 257.8 98.9 258.6 ;
      RECT  93.6 257.8 94.4 258.6 ;
      RECT  126.8 204.4 127.6 205.2 ;
      RECT  130.3 204.4 131.1 205.2 ;
      RECT  126.8 215.2 127.6 216.0 ;
      RECT  131.7 215.2 132.5 216.0 ;
      RECT  126.8 225.2 127.6 226.0 ;
      RECT  133.1 225.2 133.9 226.0 ;
      RECT  126.8 236.0 127.6 236.8 ;
      RECT  134.5 236.0 135.3 236.8 ;
      RECT  126.8 246.0 127.6 246.8 ;
      RECT  135.9 246.0 136.7 246.8 ;
      RECT  126.8 256.8 127.6 257.6 ;
      RECT  137.3 256.8 138.1 257.6 ;
      RECT  126.8 266.8 127.6 267.6 ;
      RECT  138.7 266.8 139.5 267.6 ;
      RECT  126.8 277.6 127.6 278.4 ;
      RECT  140.1 277.6 140.9 278.4 ;
      RECT  145.7 204.6 146.5 205.4 ;
      RECT  145.7 194.2 146.5 195.0 ;
      RECT  145.7 204.6 146.5 205.4 ;
      RECT  145.7 215.0 146.5 215.8 ;
      RECT  145.7 225.4 146.5 226.2 ;
      RECT  145.7 215.0 146.5 215.8 ;
      RECT  145.7 225.4 146.5 226.2 ;
      RECT  145.7 235.8 146.5 236.6 ;
      RECT  145.7 246.2 146.5 247.0 ;
      RECT  145.7 235.8 146.5 236.6 ;
      RECT  145.7 246.2 146.5 247.0 ;
      RECT  145.7 256.6 146.5 257.4 ;
      RECT  145.7 267.0 146.5 267.8 ;
      RECT  145.7 256.6 146.5 257.4 ;
      RECT  145.7 267.0 146.5 267.8 ;
      RECT  145.7 277.4 146.5 278.2 ;
      RECT  145.7 287.8 146.5 288.6 ;
      RECT  145.7 277.4 146.5 278.2 ;
      RECT  145.7 287.8 146.5 288.6 ;
      RECT  145.7 298.2 146.5 299.0 ;
      RECT  145.7 308.6 146.5 309.4 ;
      RECT  145.7 298.2 146.5 299.0 ;
      RECT  145.7 308.6 146.5 309.4 ;
      RECT  145.7 319.0 146.5 319.8 ;
      RECT  145.7 329.4 146.5 330.2 ;
      RECT  145.7 319.0 146.5 319.8 ;
      RECT  145.7 329.4 146.5 330.2 ;
      RECT  145.7 339.8 146.5 340.6 ;
      RECT  145.7 350.2 146.5 351.0 ;
      RECT  145.7 339.8 146.5 340.6 ;
      RECT  145.7 350.2 146.5 351.0 ;
      RECT  145.7 360.6 146.5 361.4 ;
      RECT  145.7 225.4 146.5 226.2 ;
      RECT  145.7 350.2 146.5 351.0 ;
      RECT  145.7 246.2 146.5 247.0 ;
      RECT  145.7 204.6 146.5 205.4 ;
      RECT  145.7 287.8 146.5 288.6 ;
      RECT  122.7 204.6 123.5 205.4 ;
      RECT  145.7 329.4 146.5 330.2 ;
      RECT  105.3 225.4 106.1 226.2 ;
      RECT  122.7 225.4 123.5 226.2 ;
      RECT  105.3 267.0 106.1 267.8 ;
      RECT  105.3 246.2 106.1 247.0 ;
      RECT  122.7 246.2 123.5 247.0 ;
      RECT  122.7 267.0 123.5 267.8 ;
      RECT  105.3 204.6 106.1 205.4 ;
      RECT  145.7 308.6 146.5 309.4 ;
      RECT  145.7 267.0 146.5 267.8 ;
      RECT  145.7 360.6 146.5 361.4 ;
      RECT  122.7 277.4 123.5 278.2 ;
      RECT  105.3 256.6 106.1 257.4 ;
      RECT  145.7 298.2 146.5 299.0 ;
      RECT  105.3 277.4 106.1 278.2 ;
      RECT  145.7 277.4 146.5 278.2 ;
      RECT  105.3 215.0 106.1 215.8 ;
      RECT  145.7 319.0 146.5 319.8 ;
      RECT  122.7 235.8 123.5 236.6 ;
      RECT  145.7 235.8 146.5 236.6 ;
      RECT  145.7 215.0 146.5 215.8 ;
      RECT  105.3 235.8 106.1 236.6 ;
      RECT  122.7 256.6 123.5 257.4 ;
      RECT  145.7 256.6 146.5 257.4 ;
      RECT  122.7 194.2 123.5 195.0 ;
      RECT  122.7 215.0 123.5 215.8 ;
      RECT  105.3 194.2 106.1 195.0 ;
      RECT  145.7 339.8 146.5 340.6 ;
      RECT  145.7 194.2 146.5 195.0 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 194.2 173.9 195.0 ;
      RECT  173.1 194.2 173.9 195.0 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 360.6 173.9 361.4 ;
      RECT  173.1 360.6 173.9 361.4 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 194.2 173.9 195.0 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  173.1 360.6 173.9 361.4 ;
      RECT  145.7 329.4 146.5 330.2 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  122.7 246.2 123.5 247.0 ;
      RECT  122.7 225.4 123.5 226.2 ;
      RECT  122.7 267.0 123.5 267.8 ;
      RECT  105.3 267.0 106.1 267.8 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  145.7 350.2 146.5 351.0 ;
      RECT  145.7 246.2 146.5 247.0 ;
      RECT  105.3 246.2 106.1 247.0 ;
      RECT  145.7 225.4 146.5 226.2 ;
      RECT  145.7 204.6 146.5 205.4 ;
      RECT  105.3 225.4 106.1 226.2 ;
      RECT  122.7 204.6 123.5 205.4 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  145.7 287.8 146.5 288.6 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  105.3 204.6 106.1 205.4 ;
      RECT  145.7 267.0 146.5 267.8 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  145.7 308.6 146.5 309.4 ;
      RECT  145.7 256.6 146.5 257.4 ;
      RECT  145.7 235.8 146.5 236.6 ;
      RECT  173.1 194.2 173.9 195.0 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  145.7 339.8 146.5 340.6 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  122.7 215.0 123.5 215.8 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  122.7 277.4 123.5 278.2 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  145.7 277.4 146.5 278.2 ;
      RECT  122.7 235.8 123.5 236.6 ;
      RECT  145.7 215.0 146.5 215.8 ;
      RECT  105.3 194.2 106.1 195.0 ;
      RECT  105.3 235.8 106.1 236.6 ;
      RECT  145.7 360.6 146.5 361.4 ;
      RECT  122.7 194.2 123.5 195.0 ;
      RECT  105.3 215.0 106.1 215.8 ;
      RECT  145.7 298.2 146.5 299.0 ;
      RECT  145.7 319.0 146.5 319.8 ;
      RECT  122.7 256.6 123.5 257.4 ;
      RECT  105.3 277.4 106.1 278.2 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  105.3 256.6 106.1 257.4 ;
      RECT  145.7 194.2 146.5 195.0 ;
      RECT  173.1 360.6 173.9 361.4 ;
      RECT  209.3 370.7 209.9 371.3 ;
      RECT  188.9 225.1 189.5 225.7 ;
      RECT  209.3 183.5 209.9 184.1 ;
      RECT  173.1 267.0 173.9 267.8 ;
      RECT  209.3 225.1 209.9 225.7 ;
      RECT  209.3 308.3 209.9 308.9 ;
      RECT  209.3 349.9 209.9 350.5 ;
      RECT  204.9 132.7 205.5 133.3 ;
      RECT  202.5 287.5 203.1 288.1 ;
      RECT  122.7 225.4 123.5 226.2 ;
      RECT  188.9 183.5 189.5 184.1 ;
      RECT  173.1 350.2 173.9 351.0 ;
      RECT  188.9 287.5 189.5 288.1 ;
      RECT  195.6 183.4 196.4 184.2 ;
      RECT  209.3 245.9 209.9 246.5 ;
      RECT  188.9 329.1 189.5 329.7 ;
      RECT  195.6 225.0 196.4 225.8 ;
      RECT  188.9 204.3 189.5 204.9 ;
      RECT  216.1 266.7 216.7 267.3 ;
      RECT  216.1 329.1 216.7 329.7 ;
      RECT  216.1 349.9 216.7 350.5 ;
      RECT  173.1 225.4 173.9 226.2 ;
      RECT  216.1 370.7 216.7 371.3 ;
      RECT  122.7 246.2 123.5 247.0 ;
      RECT  145.7 287.8 146.5 288.6 ;
      RECT  173.1 329.4 173.9 330.2 ;
      RECT  202.5 245.9 203.1 246.5 ;
      RECT  105.3 225.4 106.1 226.2 ;
      RECT  202.7 98.7 203.3 99.3 ;
      RECT  202.5 329.1 203.1 329.7 ;
      RECT  145.7 267.0 146.5 267.8 ;
      RECT  216.1 287.5 216.7 288.1 ;
      RECT  195.6 349.8 196.4 350.6 ;
      RECT  188.9 245.9 189.5 246.5 ;
      RECT  216.1 245.9 216.7 246.5 ;
      RECT  195.6 266.6 196.4 267.4 ;
      RECT  145.7 329.4 146.5 330.2 ;
      RECT  195.6 287.4 196.4 288.2 ;
      RECT  122.7 204.6 123.5 205.4 ;
      RECT  202.5 308.3 203.1 308.9 ;
      RECT  145.7 246.2 146.5 247.0 ;
      RECT  145.7 204.6 146.5 205.4 ;
      RECT  173.1 246.2 173.9 247.0 ;
      RECT  188.9 349.9 189.5 350.5 ;
      RECT  145.7 225.4 146.5 226.2 ;
      RECT  209.3 204.3 209.9 204.9 ;
      RECT  122.7 267.0 123.5 267.8 ;
      RECT  188.9 308.3 189.5 308.9 ;
      RECT  105.3 246.2 106.1 247.0 ;
      RECT  216.1 225.1 216.7 225.7 ;
      RECT  195.6 370.6 196.4 371.4 ;
      RECT  202.5 370.7 203.1 371.3 ;
      RECT  195.6 204.2 196.4 205.0 ;
      RECT  209.3 266.7 209.9 267.3 ;
      RECT  216.1 183.5 216.7 184.1 ;
      RECT  202.5 204.3 203.1 204.9 ;
      RECT  145.7 308.6 146.5 309.4 ;
      RECT  216.1 308.3 216.7 308.9 ;
      RECT  210.1 81.3 210.7 81.9 ;
      RECT  195.6 308.2 196.4 309.0 ;
      RECT  173.1 308.6 173.9 309.4 ;
      RECT  105.3 267.0 106.1 267.8 ;
      RECT  195.6 329.0 196.4 329.8 ;
      RECT  209.0 163.0 209.8 163.8 ;
      RECT  216.1 204.3 216.7 204.9 ;
      RECT  202.5 225.1 203.1 225.7 ;
      RECT  173.1 287.8 173.9 288.6 ;
      RECT  202.5 349.9 203.1 350.5 ;
      RECT  202.5 183.5 203.1 184.1 ;
      RECT  209.3 287.5 209.9 288.1 ;
      RECT  188.9 266.7 189.5 267.3 ;
      RECT  195.6 245.8 196.4 246.6 ;
      RECT  145.7 350.2 146.5 351.0 ;
      RECT  195.4 163.0 196.2 163.8 ;
      RECT  211.7 132.7 212.3 133.3 ;
      RECT  202.5 266.7 203.1 267.3 ;
      RECT  203.3 81.3 203.9 81.9 ;
      RECT  105.3 204.6 106.1 205.4 ;
      RECT  188.9 370.7 189.5 371.3 ;
      RECT  209.5 98.7 210.1 99.3 ;
      RECT  173.1 204.6 173.9 205.4 ;
      RECT  209.3 329.1 209.9 329.7 ;
      RECT  202.2 163.0 203.0 163.8 ;
      RECT  192.2 292.4 193.0 293.2 ;
      RECT  192.2 344.8 193.0 345.6 ;
      RECT  219.5 354.9 220.1 355.5 ;
      RECT  192.2 230.0 193.0 230.8 ;
      RECT  192.2 188.4 193.0 189.2 ;
      RECT  192.3 199.3 192.9 199.9 ;
      RECT  122.7 235.8 123.5 236.6 ;
      RECT  192.3 324.1 192.9 324.7 ;
      RECT  173.1 339.8 173.9 340.6 ;
      RECT  219.5 178.5 220.1 179.1 ;
      RECT  205.9 324.1 206.5 324.7 ;
      RECT  145.7 194.2 146.5 195.0 ;
      RECT  173.1 319.0 173.9 319.8 ;
      RECT  205.9 282.5 206.5 283.1 ;
      RECT  199.1 209.3 199.7 209.9 ;
      RECT  212.7 146.1 213.3 146.7 ;
      RECT  122.7 215.0 123.5 215.8 ;
      RECT  145.7 298.2 146.5 299.0 ;
      RECT  205.9 344.9 206.5 345.5 ;
      RECT  205.9 209.3 206.5 209.9 ;
      RECT  192.2 199.2 193.0 200.0 ;
      RECT  212.7 199.3 213.3 199.9 ;
      RECT  199.1 188.5 199.7 189.1 ;
      RECT  192.2 303.2 193.0 304.0 ;
      RECT  203.3 87.9 203.9 88.5 ;
      RECT  219.5 313.3 220.1 313.9 ;
      RECT  199.0 230.0 199.8 230.8 ;
      RECT  212.7 188.5 213.3 189.1 ;
      RECT  192.3 334.1 192.9 334.7 ;
      RECT  192.3 209.3 192.9 209.9 ;
      RECT  205.9 313.3 206.5 313.9 ;
      RECT  185.5 282.5 186.1 283.1 ;
      RECT  205.9 354.9 206.5 355.5 ;
      RECT  199.1 199.3 199.7 199.9 ;
      RECT  219.5 324.1 220.1 324.7 ;
      RECT  145.7 339.8 146.5 340.6 ;
      RECT  185.5 334.1 186.1 334.7 ;
      RECT  199.0 334.0 199.8 334.8 ;
      RECT  199.1 303.3 199.7 303.9 ;
      RECT  219.5 240.9 220.1 241.5 ;
      RECT  219.5 344.9 220.1 345.5 ;
      RECT  192.3 292.5 192.9 293.1 ;
      RECT  199.0 271.6 199.8 272.4 ;
      RECT  173.1 277.4 173.9 278.2 ;
      RECT  122.7 277.4 123.5 278.2 ;
      RECT  212.7 209.3 213.3 209.9 ;
      RECT  212.7 313.3 213.3 313.9 ;
      RECT  185.5 324.1 186.1 324.7 ;
      RECT  204.7 92.3 205.3 92.9 ;
      RECT  212.7 292.5 213.3 293.1 ;
      RECT  219.5 282.5 220.1 283.1 ;
      RECT  219.5 365.7 220.1 366.3 ;
      RECT  211.5 92.3 212.1 92.9 ;
      RECT  212.7 178.5 213.3 179.1 ;
      RECT  192.3 250.9 192.9 251.5 ;
      RECT  199.0 209.2 199.8 210.0 ;
      RECT  205.9 240.9 206.5 241.5 ;
      RECT  173.1 298.2 173.9 299.0 ;
      RECT  185.5 354.9 186.1 355.5 ;
      RECT  199.0 292.4 199.8 293.2 ;
      RECT  185.5 199.3 186.1 199.9 ;
      RECT  199.0 240.8 199.8 241.6 ;
      RECT  105.3 194.2 106.1 195.0 ;
      RECT  192.3 282.5 192.9 283.1 ;
      RECT  185.5 344.9 186.1 345.5 ;
      RECT  145.7 215.0 146.5 215.8 ;
      RECT  201.9 106.9 202.5 107.5 ;
      RECT  192.2 209.2 193.0 210.0 ;
      RECT  205.9 178.5 206.5 179.1 ;
      RECT  199.1 313.3 199.7 313.9 ;
      RECT  205.9 220.1 206.5 220.7 ;
      RECT  219.5 334.1 220.1 334.7 ;
      RECT  185.5 271.7 186.1 272.3 ;
      RECT  145.7 277.4 146.5 278.2 ;
      RECT  192.2 178.4 193.0 179.2 ;
      RECT  199.1 354.9 199.7 355.5 ;
      RECT  185.5 313.3 186.1 313.9 ;
      RECT  199.1 365.7 199.7 366.3 ;
      RECT  205.9 199.3 206.5 199.9 ;
      RECT  105.3 215.0 106.1 215.8 ;
      RECT  212.7 354.9 213.3 355.5 ;
      RECT  208.7 106.9 209.3 107.5 ;
      RECT  185.5 292.5 186.1 293.1 ;
      RECT  199.0 344.8 199.8 345.6 ;
      RECT  192.2 271.6 193.0 272.4 ;
      RECT  173.1 235.8 173.9 236.6 ;
      RECT  199.0 324.0 199.8 324.8 ;
      RECT  212.7 303.3 213.3 303.9 ;
      RECT  199.1 261.7 199.7 262.3 ;
      RECT  212.7 271.7 213.3 272.3 ;
      RECT  192.3 365.7 192.9 366.3 ;
      RECT  185.5 230.1 186.1 230.7 ;
      RECT  192.2 313.2 193.0 314.0 ;
      RECT  192.2 354.8 193.0 355.6 ;
      RECT  185.5 209.3 186.1 209.9 ;
      RECT  173.1 360.6 173.9 361.4 ;
      RECT  199.0 282.4 199.8 283.2 ;
      RECT  205.9 188.5 206.5 189.1 ;
      RECT  192.3 220.1 192.9 220.7 ;
      RECT  173.1 215.0 173.9 215.8 ;
      RECT  192.3 344.9 192.9 345.5 ;
      RECT  192.2 324.0 193.0 324.8 ;
      RECT  199.1 292.5 199.7 293.1 ;
      RECT  192.2 282.4 193.0 283.2 ;
      RECT  192.3 230.1 192.9 230.7 ;
      RECT  192.3 271.7 192.9 272.3 ;
      RECT  185.5 188.5 186.1 189.1 ;
      RECT  199.0 354.8 199.8 355.6 ;
      RECT  205.9 365.7 206.5 366.3 ;
      RECT  205.9 230.1 206.5 230.7 ;
      RECT  122.7 194.2 123.5 195.0 ;
      RECT  192.3 178.5 192.9 179.1 ;
      RECT  199.0 250.8 199.8 251.6 ;
      RECT  173.1 194.2 173.9 195.0 ;
      RECT  145.7 360.6 146.5 361.4 ;
      RECT  205.9 334.1 206.5 334.7 ;
      RECT  199.1 178.5 199.7 179.1 ;
      RECT  212.7 324.1 213.3 324.7 ;
      RECT  192.2 261.6 193.0 262.4 ;
      RECT  185.5 365.7 186.1 366.3 ;
      RECT  185.5 178.5 186.1 179.1 ;
      RECT  173.1 256.6 173.9 257.4 ;
      RECT  205.9 250.9 206.5 251.5 ;
      RECT  199.0 220.0 199.8 220.8 ;
      RECT  212.7 365.7 213.3 366.3 ;
      RECT  219.5 271.7 220.1 272.3 ;
      RECT  145.7 256.6 146.5 257.4 ;
      RECT  105.3 235.8 106.1 236.6 ;
      RECT  199.1 282.5 199.7 283.1 ;
      RECT  192.3 313.3 192.9 313.9 ;
      RECT  212.7 334.1 213.3 334.7 ;
      RECT  199.0 303.2 199.8 304.0 ;
      RECT  219.5 261.7 220.1 262.3 ;
      RECT  219.5 250.9 220.1 251.5 ;
      RECT  219.5 220.1 220.1 220.7 ;
      RECT  105.3 256.6 106.1 257.4 ;
      RECT  185.5 303.3 186.1 303.9 ;
      RECT  205.9 271.7 206.5 272.3 ;
      RECT  192.2 240.8 193.0 241.6 ;
      RECT  199.1 271.7 199.7 272.3 ;
      RECT  192.2 250.8 193.0 251.6 ;
      RECT  212.7 344.9 213.3 345.5 ;
      RECT  192.3 354.9 192.9 355.5 ;
      RECT  192.2 365.6 193.0 366.4 ;
      RECT  212.7 230.1 213.3 230.7 ;
      RECT  199.1 334.1 199.7 334.7 ;
      RECT  219.5 303.3 220.1 303.9 ;
      RECT  192.3 261.7 192.9 262.3 ;
      RECT  199.0 188.4 199.8 189.2 ;
      RECT  192.2 220.0 193.0 220.8 ;
      RECT  185.5 240.9 186.1 241.5 ;
      RECT  212.7 250.9 213.3 251.5 ;
      RECT  145.7 235.8 146.5 236.6 ;
      RECT  219.5 188.5 220.1 189.1 ;
      RECT  219.5 199.3 220.1 199.9 ;
      RECT  199.1 344.9 199.7 345.5 ;
      RECT  205.9 146.1 206.5 146.7 ;
      RECT  192.3 303.3 192.9 303.9 ;
      RECT  210.1 87.9 210.7 88.5 ;
      RECT  212.7 282.5 213.3 283.1 ;
      RECT  199.1 250.9 199.7 251.5 ;
      RECT  192.3 240.9 192.9 241.5 ;
      RECT  185.5 250.9 186.1 251.5 ;
      RECT  199.1 240.9 199.7 241.5 ;
      RECT  122.7 256.6 123.5 257.4 ;
      RECT  199.1 220.1 199.7 220.7 ;
      RECT  219.5 209.3 220.1 209.9 ;
      RECT  105.3 277.4 106.1 278.2 ;
      RECT  199.0 178.4 199.8 179.2 ;
      RECT  185.5 220.1 186.1 220.7 ;
      RECT  145.7 319.0 146.5 319.8 ;
      RECT  192.2 334.0 193.0 334.8 ;
      RECT  212.7 240.9 213.3 241.5 ;
      RECT  205.9 292.5 206.5 293.1 ;
      RECT  199.1 324.1 199.7 324.7 ;
      RECT  199.1 230.1 199.7 230.7 ;
      RECT  199.0 313.2 199.8 314.0 ;
      RECT  185.5 261.7 186.1 262.3 ;
      RECT  205.9 303.3 206.5 303.9 ;
      RECT  219.5 292.5 220.1 293.1 ;
      RECT  199.0 365.6 199.8 366.4 ;
      RECT  199.0 199.2 199.8 200.0 ;
      RECT  212.7 261.7 213.3 262.3 ;
      RECT  212.7 220.1 213.3 220.7 ;
      RECT  192.3 188.5 192.9 189.1 ;
      RECT  219.5 230.1 220.1 230.7 ;
      RECT  205.9 261.7 206.5 262.3 ;
      RECT  199.0 261.6 199.8 262.4 ;
      RECT  30.5 12.9 47.5 13.5 ;
      RECT  30.5 30.9 43.3 31.5 ;
      RECT  35.9 34.1 46.1 34.7 ;
      RECT  37.7 131.7 53.5 132.3 ;
      RECT  44.7 4.7 74.3 5.3 ;
      RECT  47.5 37.1 58.4 37.7 ;
      RECT  40.5 32.7 82.3 33.3 ;
      RECT  41.9 51.1 75.9 51.7 ;
      RECT  23.9 11.7 24.5 12.3 ;
      RECT  23.9 11.5 24.5 12.1 ;
      RECT  22.0 11.7 24.2 12.3 ;
      RECT  23.9 11.8 24.5 12.0 ;
      RECT  24.2 11.5 26.4 12.1 ;
      RECT  21.6 11.6 22.4 12.4 ;
      RECT  26.0 11.4 26.8 12.2 ;
      RECT  23.9 32.7 24.5 32.1 ;
      RECT  23.9 32.9 24.5 32.3 ;
      RECT  22.0 32.7 24.2 32.1 ;
      RECT  23.9 32.6 24.5 32.4 ;
      RECT  24.2 32.9 26.4 32.3 ;
      RECT  21.6 32.8 22.4 32.0 ;
      RECT  26.0 33.0 26.8 32.2 ;
      RECT  2.4 21.8 3.2 22.6 ;
      RECT  2.4 1.8 3.2 2.6 ;
      RECT  2.4 21.8 3.2 22.6 ;
      RECT  2.4 41.8 3.2 42.6 ;
      RECT  2.4 21.8 3.2 22.6 ;
      RECT  2.4 1.8 3.2 2.6 ;
      RECT  2.4 41.8 3.2 42.6 ;
      RECT  31.3 169.7 7.4 170.3 ;
      RECT  31.3 180.5 7.4 181.1 ;
      RECT  31.3 190.5 7.4 191.1 ;
      RECT  31.3 201.3 7.4 201.9 ;
      RECT  31.3 211.3 7.4 211.9 ;
      RECT  31.3 222.1 7.4 222.7 ;
      RECT  31.3 232.1 7.4 232.7 ;
      RECT  31.3 242.9 7.4 243.5 ;
      RECT  31.3 252.9 7.4 253.5 ;
      RECT  27.0 169.6 26.2 170.4 ;
      RECT  20.6 169.6 19.8 170.4 ;
      RECT  14.2 169.6 13.4 170.4 ;
      RECT  7.8 169.6 7.0 170.4 ;
      RECT  31.7 169.6 30.9 170.4 ;
      RECT  27.0 180.4 26.2 181.2 ;
      RECT  20.6 180.4 19.8 181.2 ;
      RECT  14.2 180.4 13.4 181.2 ;
      RECT  7.8 180.4 7.0 181.2 ;
      RECT  31.7 180.4 30.9 181.2 ;
      RECT  27.0 190.4 26.2 191.2 ;
      RECT  20.6 190.4 19.8 191.2 ;
      RECT  14.2 190.4 13.4 191.2 ;
      RECT  7.8 190.4 7.0 191.2 ;
      RECT  31.7 190.4 30.9 191.2 ;
      RECT  27.0 201.2 26.2 202.0 ;
      RECT  20.6 201.2 19.8 202.0 ;
      RECT  14.2 201.2 13.4 202.0 ;
      RECT  7.8 201.2 7.0 202.0 ;
      RECT  31.7 201.2 30.9 202.0 ;
      RECT  27.0 211.2 26.2 212.0 ;
      RECT  20.6 211.2 19.8 212.0 ;
      RECT  14.2 211.2 13.4 212.0 ;
      RECT  7.8 211.2 7.0 212.0 ;
      RECT  31.7 211.2 30.9 212.0 ;
      RECT  27.0 222.0 26.2 222.8 ;
      RECT  20.6 222.0 19.8 222.8 ;
      RECT  14.2 222.0 13.4 222.8 ;
      RECT  7.8 222.0 7.0 222.8 ;
      RECT  31.7 222.0 30.9 222.8 ;
      RECT  27.0 232.0 26.2 232.8 ;
      RECT  20.6 232.0 19.8 232.8 ;
      RECT  14.2 232.0 13.4 232.8 ;
      RECT  7.8 232.0 7.0 232.8 ;
      RECT  31.7 232.0 30.9 232.8 ;
      RECT  27.0 242.8 26.2 243.6 ;
      RECT  20.6 242.8 19.8 243.6 ;
      RECT  14.2 242.8 13.4 243.6 ;
      RECT  7.8 242.8 7.0 243.6 ;
      RECT  31.7 242.8 30.9 243.6 ;
      RECT  27.0 252.8 26.2 253.6 ;
      RECT  20.6 252.8 19.8 253.6 ;
      RECT  14.2 252.8 13.4 253.6 ;
      RECT  7.8 252.8 7.0 253.6 ;
      RECT  31.7 252.8 30.9 253.6 ;
      RECT  22.4 175.0 21.6 175.8 ;
      RECT  22.4 164.6 21.6 165.4 ;
      RECT  16.0 175.0 15.2 175.8 ;
      RECT  16.0 164.6 15.2 165.4 ;
      RECT  9.6 175.0 8.8 175.8 ;
      RECT  9.6 164.6 8.8 165.4 ;
      RECT  22.4 195.8 21.6 196.6 ;
      RECT  22.4 185.4 21.6 186.2 ;
      RECT  16.0 195.8 15.2 196.6 ;
      RECT  16.0 185.4 15.2 186.2 ;
      RECT  9.6 195.8 8.8 196.6 ;
      RECT  9.6 185.4 8.8 186.2 ;
      RECT  22.4 216.6 21.6 217.4 ;
      RECT  22.4 206.2 21.6 207.0 ;
      RECT  16.0 216.6 15.2 217.4 ;
      RECT  16.0 206.2 15.2 207.0 ;
      RECT  9.6 216.6 8.8 217.4 ;
      RECT  9.6 206.2 8.8 207.0 ;
      RECT  22.4 237.4 21.6 238.2 ;
      RECT  22.4 227.0 21.6 227.8 ;
      RECT  16.0 237.4 15.2 238.2 ;
      RECT  16.0 227.0 15.2 227.8 ;
      RECT  9.6 237.4 8.8 238.2 ;
      RECT  9.6 227.0 8.8 227.8 ;
      RECT  22.4 258.2 21.6 259.0 ;
      RECT  22.4 247.8 21.6 248.6 ;
      RECT  16.0 258.2 15.2 259.0 ;
      RECT  16.0 247.8 15.2 248.6 ;
      RECT  9.6 258.2 8.8 259.0 ;
      RECT  9.6 247.8 8.8 248.6 ;
      RECT  22.4 247.8 21.6 248.6 ;
      RECT  16.0 247.8 15.2 248.6 ;
      RECT  9.6 247.8 8.8 248.6 ;
      RECT  22.4 237.4 21.6 238.2 ;
      RECT  9.6 258.2 8.8 259.0 ;
      RECT  22.4 258.2 21.6 259.0 ;
      RECT  16.0 175.0 15.2 175.8 ;
      RECT  16.0 258.2 15.2 259.0 ;
      RECT  9.6 195.8 8.8 196.6 ;
      RECT  22.4 216.6 21.6 217.4 ;
      RECT  9.6 237.4 8.8 238.2 ;
      RECT  22.4 195.8 21.6 196.6 ;
      RECT  16.0 195.8 15.2 196.6 ;
      RECT  22.4 175.0 21.6 175.8 ;
      RECT  16.0 216.6 15.2 217.4 ;
      RECT  9.6 216.6 8.8 217.4 ;
      RECT  16.0 237.4 15.2 238.2 ;
      RECT  9.6 175.0 8.8 175.8 ;
      RECT  9.6 185.4 8.8 186.2 ;
      RECT  9.6 164.6 8.8 165.4 ;
      RECT  22.4 227.0 21.6 227.8 ;
      RECT  16.0 227.0 15.2 227.8 ;
      RECT  9.6 227.0 8.8 227.8 ;
      RECT  22.4 185.4 21.6 186.2 ;
      RECT  22.4 247.8 21.6 248.6 ;
      RECT  22.4 206.2 21.6 207.0 ;
      RECT  9.6 206.2 8.8 207.0 ;
      RECT  16.0 206.2 15.2 207.0 ;
      RECT  9.6 247.8 8.8 248.6 ;
      RECT  16.0 164.6 15.2 165.4 ;
      RECT  22.4 164.6 21.6 165.4 ;
      RECT  16.0 185.4 15.2 186.2 ;
      RECT  16.0 247.8 15.2 248.6 ;
      RECT  47.1 12.8 47.9 13.6 ;
      RECT  30.1 12.8 30.9 13.6 ;
      RECT  42.9 30.8 43.7 31.6 ;
      RECT  30.1 30.8 30.9 31.6 ;
      RECT  45.7 34.0 46.5 34.8 ;
      RECT  35.5 34.0 36.3 34.8 ;
      RECT  37.3 131.6 38.1 132.4 ;
      RECT  53.1 131.6 53.9 132.4 ;
      RECT  73.9 4.6 74.7 5.4 ;
      RECT  44.3 4.6 45.1 5.4 ;
      RECT  47.1 37.0 47.9 37.8 ;
      RECT  58.0 37.0 58.8 37.8 ;
      RECT  40.1 32.6 40.9 33.4 ;
      RECT  81.9 32.6 82.7 33.4 ;
      RECT  41.5 51.0 42.3 51.8 ;
      RECT  75.5 51.0 76.3 51.8 ;
      RECT  84.8 21.8 85.6 22.6 ;
      RECT  84.8 1.8 85.6 2.6 ;
      RECT  84.8 21.8 85.6 22.6 ;
      RECT  84.8 41.8 85.6 42.6 ;
      RECT  84.8 61.8 85.6 62.6 ;
      RECT  84.8 41.8 85.6 42.6 ;
      RECT  84.8 61.8 85.6 62.6 ;
      RECT  84.8 81.8 85.6 82.6 ;
      RECT  84.8 101.8 85.6 102.6 ;
      RECT  84.8 81.8 85.6 82.6 ;
      RECT  84.8 101.8 85.6 102.6 ;
      RECT  84.8 121.8 85.6 122.6 ;
      RECT  84.8 141.8 85.6 142.6 ;
      RECT  84.8 121.8 85.6 122.6 ;
      RECT  84.8 141.8 85.6 142.6 ;
      RECT  84.8 161.8 85.6 162.6 ;
      RECT  21.6 195.8 22.4 196.6 ;
      RECT  84.8 101.8 85.6 102.6 ;
      RECT  21.6 258.2 22.4 259.0 ;
      RECT  8.8 175.0 9.6 175.8 ;
      RECT  15.2 258.2 16.0 259.0 ;
      RECT  21.6 216.6 22.4 217.4 ;
      RECT  21.6 175.0 22.4 175.8 ;
      RECT  8.8 195.8 9.6 196.6 ;
      RECT  2.4 21.8 3.2 22.6 ;
      RECT  8.8 258.2 9.6 259.0 ;
      RECT  21.6 237.4 22.4 238.2 ;
      RECT  8.8 216.6 9.6 217.4 ;
      RECT  15.2 216.6 16.0 217.4 ;
      RECT  8.8 237.4 9.6 238.2 ;
      RECT  84.8 21.8 85.6 22.6 ;
      RECT  84.8 61.8 85.6 62.6 ;
      RECT  15.2 175.0 16.0 175.8 ;
      RECT  15.2 237.4 16.0 238.2 ;
      RECT  15.2 195.8 16.0 196.6 ;
      RECT  84.8 141.8 85.6 142.6 ;
      RECT  21.6 227.0 22.4 227.8 ;
      RECT  21.6 206.2 22.4 207.0 ;
      RECT  15.2 185.4 16.0 186.2 ;
      RECT  15.2 247.8 16.0 248.6 ;
      RECT  84.8 161.8 85.6 162.6 ;
      RECT  2.4 41.8 3.2 42.6 ;
      RECT  21.6 247.8 22.4 248.6 ;
      RECT  84.8 1.8 85.6 2.6 ;
      RECT  15.2 227.0 16.0 227.8 ;
      RECT  84.8 41.8 85.6 42.6 ;
      RECT  15.2 164.6 16.0 165.4 ;
      RECT  2.4 1.8 3.2 2.6 ;
      RECT  15.2 206.2 16.0 207.0 ;
      RECT  21.6 185.4 22.4 186.2 ;
      RECT  8.8 185.4 9.6 186.2 ;
      RECT  8.8 227.0 9.6 227.8 ;
      RECT  84.8 121.8 85.6 122.6 ;
      RECT  8.8 164.6 9.6 165.4 ;
      RECT  8.8 206.2 9.6 207.0 ;
      RECT  8.8 247.8 9.6 248.6 ;
      RECT  84.8 81.8 85.6 82.6 ;
      RECT  21.6 164.6 22.4 165.4 ;
      RECT  75.3 312.4 76.1 313.2 ;
      RECT  75.3 292.4 76.1 293.2 ;
      RECT  75.3 312.4 76.1 313.2 ;
      RECT  75.3 332.4 76.1 333.2 ;
      RECT  75.3 352.4 76.1 353.2 ;
      RECT  75.3 332.4 76.1 333.2 ;
      RECT  75.3 352.4 76.1 353.2 ;
      RECT  75.3 372.4 76.1 373.2 ;
      RECT  67.6 297.8 68.4 298.6 ;
      RECT  64.8 297.9 86.6 298.5 ;
      RECT  75.3 352.4 76.1 353.2 ;
      RECT  75.3 312.4 76.1 313.2 ;
      RECT  75.3 372.4 76.1 373.2 ;
      RECT  75.3 332.4 76.1 333.2 ;
      RECT  75.3 292.4 76.1 293.2 ;
      RECT  196.3 67.6 197.1 68.4 ;
      RECT  196.3 47.6 197.1 48.4 ;
      RECT  218.1 67.6 218.9 68.4 ;
      RECT  218.1 47.6 218.9 48.4 ;
      RECT  188.6 53.0 189.4 53.8 ;
      RECT  210.4 53.0 211.2 53.8 ;
      RECT  185.8 53.1 229.4 53.7 ;
      RECT  218.1 67.6 218.9 68.4 ;
      RECT  196.3 67.6 197.1 68.4 ;
      RECT  218.1 47.6 218.9 48.4 ;
      RECT  196.3 47.6 197.1 48.4 ;
      RECT  87.6 297.8 88.4 298.6 ;
      RECT  87.6 53.0 88.4 53.8 ;
      RECT  180.1 152.2 180.9 153.0 ;
      RECT  86.2 152.2 87.0 153.0 ;
      RECT  178.7 90.8 179.5 91.6 ;
      RECT  86.2 90.8 87.0 91.6 ;
      RECT  181.5 112.0 182.3 112.8 ;
      RECT  86.2 112.0 87.0 112.8 ;
      RECT  182.9 72.8 183.7 73.6 ;
      RECT  86.2 72.8 87.0 73.6 ;
      RECT  193.8 167.1 194.6 167.9 ;
      RECT  33.0 167.1 33.8 167.9 ;
      RECT  89.4 302.2 90.2 303.0 ;
      RECT  83.6 302.2 84.4 303.0 ;
      RECT  90.8 322.6 91.6 323.4 ;
      RECT  83.6 322.6 84.4 323.4 ;
      RECT  92.2 342.2 93.0 343.0 ;
      RECT  83.6 342.2 84.4 343.0 ;
      RECT  93.6 362.6 94.4 363.4 ;
      RECT  83.6 362.6 84.4 363.4 ;
      RECT  2.6 0.2 3.4 1.0 ;
      RECT  7.4 0.2 8.2 1.0 ;
      RECT  12.2 0.2 13.0 1.0 ;
      RECT  17.0 0.2 17.8 1.0 ;
      RECT  21.8 0.2 22.6 1.0 ;
      RECT  26.6 0.2 27.4 1.0 ;
      RECT  31.4 0.2 32.2 1.0 ;
      RECT  36.2 0.2 37.0 1.0 ;
      RECT  41.0 0.2 41.8 1.0 ;
      RECT  45.8 0.2 46.6 1.0 ;
      RECT  50.6 0.2 51.4 1.0 ;
      RECT  55.4 0.2 56.2 1.0 ;
      RECT  60.2 0.2 61.0 1.0 ;
      RECT  65.0 0.2 65.8 1.0 ;
      RECT  69.8 0.2 70.6 1.0 ;
      RECT  74.6 0.2 75.4 1.0 ;
      RECT  79.4 0.2 80.2 1.0 ;
      RECT  84.2 0.2 85.0 1.0 ;
      RECT  89.0 0.2 89.8 1.0 ;
      RECT  93.8 0.2 94.6 1.0 ;
      RECT  98.6 0.2 99.4 1.0 ;
      RECT  103.4 0.2 104.2 1.0 ;
      RECT  108.2 0.2 109.0 1.0 ;
      RECT  113.0 0.2 113.8 1.0 ;
      RECT  117.8 0.2 118.6 1.0 ;
      RECT  122.6 0.2 123.4 1.0 ;
      RECT  127.4 0.2 128.2 1.0 ;
      RECT  132.2 0.2 133.0 1.0 ;
      RECT  137.0 0.2 137.8 1.0 ;
      RECT  141.8 0.2 142.6 1.0 ;
      RECT  146.6 0.2 147.4 1.0 ;
      RECT  151.4 0.2 152.2 1.0 ;
      RECT  156.2 0.2 157.0 1.0 ;
      RECT  161.0 0.2 161.8 1.0 ;
      RECT  165.8 0.2 166.6 1.0 ;
      RECT  170.6 0.2 171.4 1.0 ;
      RECT  175.4 0.2 176.2 1.0 ;
      RECT  180.2 0.2 181.0 1.0 ;
      RECT  185.0 0.2 185.8 1.0 ;
      RECT  189.8 0.2 190.6 1.0 ;
      RECT  194.6 0.2 195.4 1.0 ;
      RECT  199.4 0.2 200.2 1.0 ;
      RECT  204.2 0.2 205.0 1.0 ;
      RECT  209.0 0.2 209.8 1.0 ;
      RECT  213.8 0.2 214.6 1.0 ;
      RECT  218.6 0.2 219.4 1.0 ;
      RECT  223.4 0.2 224.2 1.0 ;
      RECT  2.6 5.0 3.4 5.8 ;
      RECT  7.4 5.0 8.2 5.8 ;
      RECT  12.2 5.0 13.0 5.8 ;
      RECT  17.0 5.0 17.8 5.8 ;
      RECT  21.8 5.0 22.6 5.8 ;
      RECT  26.6 5.0 27.4 5.8 ;
      RECT  31.4 5.0 32.2 5.8 ;
      RECT  36.2 5.0 37.0 5.8 ;
      RECT  79.4 5.0 80.2 5.8 ;
      RECT  84.2 5.0 85.0 5.8 ;
      RECT  89.0 5.0 89.8 5.8 ;
      RECT  93.8 5.0 94.6 5.8 ;
      RECT  98.6 5.0 99.4 5.8 ;
      RECT  103.4 5.0 104.2 5.8 ;
      RECT  108.2 5.0 109.0 5.8 ;
      RECT  113.0 5.0 113.8 5.8 ;
      RECT  117.8 5.0 118.6 5.8 ;
      RECT  122.6 5.0 123.4 5.8 ;
      RECT  127.4 5.0 128.2 5.8 ;
      RECT  132.2 5.0 133.0 5.8 ;
      RECT  137.0 5.0 137.8 5.8 ;
      RECT  141.8 5.0 142.6 5.8 ;
      RECT  146.6 5.0 147.4 5.8 ;
      RECT  151.4 5.0 152.2 5.8 ;
      RECT  156.2 5.0 157.0 5.8 ;
      RECT  161.0 5.0 161.8 5.8 ;
      RECT  165.8 5.0 166.6 5.8 ;
      RECT  170.6 5.0 171.4 5.8 ;
      RECT  175.4 5.0 176.2 5.8 ;
      RECT  180.2 5.0 181.0 5.8 ;
      RECT  185.0 5.0 185.8 5.8 ;
      RECT  189.8 5.0 190.6 5.8 ;
      RECT  194.6 5.0 195.4 5.8 ;
      RECT  199.4 5.0 200.2 5.8 ;
      RECT  204.2 5.0 205.0 5.8 ;
      RECT  209.0 5.0 209.8 5.8 ;
      RECT  213.8 5.0 214.6 5.8 ;
      RECT  218.6 5.0 219.4 5.8 ;
      RECT  223.4 5.0 224.2 5.8 ;
      RECT  31.4 9.8 32.2 10.6 ;
      RECT  36.2 9.8 37.0 10.6 ;
      RECT  41.0 9.8 41.8 10.6 ;
      RECT  45.8 9.8 46.6 10.6 ;
      RECT  50.6 9.8 51.4 10.6 ;
      RECT  55.4 9.8 56.2 10.6 ;
      RECT  60.2 9.8 61.0 10.6 ;
      RECT  65.0 9.8 65.8 10.6 ;
      RECT  69.8 9.8 70.6 10.6 ;
      RECT  74.6 9.8 75.4 10.6 ;
      RECT  79.4 9.8 80.2 10.6 ;
      RECT  84.2 9.8 85.0 10.6 ;
      RECT  89.0 9.8 89.8 10.6 ;
      RECT  93.8 9.8 94.6 10.6 ;
      RECT  98.6 9.8 99.4 10.6 ;
      RECT  103.4 9.8 104.2 10.6 ;
      RECT  108.2 9.8 109.0 10.6 ;
      RECT  113.0 9.8 113.8 10.6 ;
      RECT  117.8 9.8 118.6 10.6 ;
      RECT  122.6 9.8 123.4 10.6 ;
      RECT  127.4 9.8 128.2 10.6 ;
      RECT  132.2 9.8 133.0 10.6 ;
      RECT  137.0 9.8 137.8 10.6 ;
      RECT  141.8 9.8 142.6 10.6 ;
      RECT  146.6 9.8 147.4 10.6 ;
      RECT  151.4 9.8 152.2 10.6 ;
      RECT  156.2 9.8 157.0 10.6 ;
      RECT  161.0 9.8 161.8 10.6 ;
      RECT  165.8 9.8 166.6 10.6 ;
      RECT  170.6 9.8 171.4 10.6 ;
      RECT  175.4 9.8 176.2 10.6 ;
      RECT  180.2 9.8 181.0 10.6 ;
      RECT  185.0 9.8 185.8 10.6 ;
      RECT  189.8 9.8 190.6 10.6 ;
      RECT  194.6 9.8 195.4 10.6 ;
      RECT  199.4 9.8 200.2 10.6 ;
      RECT  204.2 9.8 205.0 10.6 ;
      RECT  209.0 9.8 209.8 10.6 ;
      RECT  213.8 9.8 214.6 10.6 ;
      RECT  218.6 9.8 219.4 10.6 ;
      RECT  223.4 9.8 224.2 10.6 ;
      RECT  50.6 14.6 51.4 15.4 ;
      RECT  55.4 14.6 56.2 15.4 ;
      RECT  60.2 14.6 61.0 15.4 ;
      RECT  65.0 14.6 65.8 15.4 ;
      RECT  69.8 14.6 70.6 15.4 ;
      RECT  74.6 14.6 75.4 15.4 ;
      RECT  79.4 14.6 80.2 15.4 ;
      RECT  84.2 14.6 85.0 15.4 ;
      RECT  89.0 14.6 89.8 15.4 ;
      RECT  93.8 14.6 94.6 15.4 ;
      RECT  98.6 14.6 99.4 15.4 ;
      RECT  103.4 14.6 104.2 15.4 ;
      RECT  108.2 14.6 109.0 15.4 ;
      RECT  113.0 14.6 113.8 15.4 ;
      RECT  117.8 14.6 118.6 15.4 ;
      RECT  122.6 14.6 123.4 15.4 ;
      RECT  127.4 14.6 128.2 15.4 ;
      RECT  132.2 14.6 133.0 15.4 ;
      RECT  137.0 14.6 137.8 15.4 ;
      RECT  141.8 14.6 142.6 15.4 ;
      RECT  146.6 14.6 147.4 15.4 ;
      RECT  151.4 14.6 152.2 15.4 ;
      RECT  156.2 14.6 157.0 15.4 ;
      RECT  161.0 14.6 161.8 15.4 ;
      RECT  165.8 14.6 166.6 15.4 ;
      RECT  170.6 14.6 171.4 15.4 ;
      RECT  175.4 14.6 176.2 15.4 ;
      RECT  180.2 14.6 181.0 15.4 ;
      RECT  185.0 14.6 185.8 15.4 ;
      RECT  189.8 14.6 190.6 15.4 ;
      RECT  194.6 14.6 195.4 15.4 ;
      RECT  199.4 14.6 200.2 15.4 ;
      RECT  204.2 14.6 205.0 15.4 ;
      RECT  209.0 14.6 209.8 15.4 ;
      RECT  213.8 14.6 214.6 15.4 ;
      RECT  218.6 14.6 219.4 15.4 ;
      RECT  223.4 14.6 224.2 15.4 ;
      RECT  2.6 19.4 3.4 20.2 ;
      RECT  7.4 19.4 8.2 20.2 ;
      RECT  12.2 19.4 13.0 20.2 ;
      RECT  17.0 19.4 17.8 20.2 ;
      RECT  21.8 19.4 22.6 20.2 ;
      RECT  26.6 19.4 27.4 20.2 ;
      RECT  31.4 19.4 32.2 20.2 ;
      RECT  36.2 19.4 37.0 20.2 ;
      RECT  41.0 19.4 41.8 20.2 ;
      RECT  45.8 19.4 46.6 20.2 ;
      RECT  50.6 19.4 51.4 20.2 ;
      RECT  55.4 19.4 56.2 20.2 ;
      RECT  60.2 19.4 61.0 20.2 ;
      RECT  65.0 19.4 65.8 20.2 ;
      RECT  69.8 19.4 70.6 20.2 ;
      RECT  74.6 19.4 75.4 20.2 ;
      RECT  79.4 19.4 80.2 20.2 ;
      RECT  84.2 19.4 85.0 20.2 ;
      RECT  89.0 19.4 89.8 20.2 ;
      RECT  93.8 19.4 94.6 20.2 ;
      RECT  98.6 19.4 99.4 20.2 ;
      RECT  103.4 19.4 104.2 20.2 ;
      RECT  108.2 19.4 109.0 20.2 ;
      RECT  113.0 19.4 113.8 20.2 ;
      RECT  117.8 19.4 118.6 20.2 ;
      RECT  122.6 19.4 123.4 20.2 ;
      RECT  127.4 19.4 128.2 20.2 ;
      RECT  132.2 19.4 133.0 20.2 ;
      RECT  137.0 19.4 137.8 20.2 ;
      RECT  141.8 19.4 142.6 20.2 ;
      RECT  146.6 19.4 147.4 20.2 ;
      RECT  151.4 19.4 152.2 20.2 ;
      RECT  156.2 19.4 157.0 20.2 ;
      RECT  161.0 19.4 161.8 20.2 ;
      RECT  165.8 19.4 166.6 20.2 ;
      RECT  170.6 19.4 171.4 20.2 ;
      RECT  175.4 19.4 176.2 20.2 ;
      RECT  180.2 19.4 181.0 20.2 ;
      RECT  185.0 19.4 185.8 20.2 ;
      RECT  189.8 19.4 190.6 20.2 ;
      RECT  194.6 19.4 195.4 20.2 ;
      RECT  199.4 19.4 200.2 20.2 ;
      RECT  204.2 19.4 205.0 20.2 ;
      RECT  209.0 19.4 209.8 20.2 ;
      RECT  213.8 19.4 214.6 20.2 ;
      RECT  218.6 19.4 219.4 20.2 ;
      RECT  223.4 19.4 224.2 20.2 ;
      RECT  2.6 24.2 3.4 25.0 ;
      RECT  7.4 24.2 8.2 25.0 ;
      RECT  12.2 24.2 13.0 25.0 ;
      RECT  17.0 24.2 17.8 25.0 ;
      RECT  21.8 24.2 22.6 25.0 ;
      RECT  26.6 24.2 27.4 25.0 ;
      RECT  31.4 24.2 32.2 25.0 ;
      RECT  36.2 24.2 37.0 25.0 ;
      RECT  41.0 24.2 41.8 25.0 ;
      RECT  45.8 24.2 46.6 25.0 ;
      RECT  50.6 24.2 51.4 25.0 ;
      RECT  55.4 24.2 56.2 25.0 ;
      RECT  60.2 24.2 61.0 25.0 ;
      RECT  65.0 24.2 65.8 25.0 ;
      RECT  69.8 24.2 70.6 25.0 ;
      RECT  74.6 24.2 75.4 25.0 ;
      RECT  79.4 24.2 80.2 25.0 ;
      RECT  84.2 24.2 85.0 25.0 ;
      RECT  89.0 24.2 89.8 25.0 ;
      RECT  93.8 24.2 94.6 25.0 ;
      RECT  98.6 24.2 99.4 25.0 ;
      RECT  103.4 24.2 104.2 25.0 ;
      RECT  108.2 24.2 109.0 25.0 ;
      RECT  113.0 24.2 113.8 25.0 ;
      RECT  117.8 24.2 118.6 25.0 ;
      RECT  122.6 24.2 123.4 25.0 ;
      RECT  127.4 24.2 128.2 25.0 ;
      RECT  132.2 24.2 133.0 25.0 ;
      RECT  137.0 24.2 137.8 25.0 ;
      RECT  141.8 24.2 142.6 25.0 ;
      RECT  146.6 24.2 147.4 25.0 ;
      RECT  151.4 24.2 152.2 25.0 ;
      RECT  156.2 24.2 157.0 25.0 ;
      RECT  161.0 24.2 161.8 25.0 ;
      RECT  165.8 24.2 166.6 25.0 ;
      RECT  170.6 24.2 171.4 25.0 ;
      RECT  175.4 24.2 176.2 25.0 ;
      RECT  180.2 24.2 181.0 25.0 ;
      RECT  185.0 24.2 185.8 25.0 ;
      RECT  189.8 24.2 190.6 25.0 ;
      RECT  194.6 24.2 195.4 25.0 ;
      RECT  199.4 24.2 200.2 25.0 ;
      RECT  204.2 24.2 205.0 25.0 ;
      RECT  209.0 24.2 209.8 25.0 ;
      RECT  213.8 24.2 214.6 25.0 ;
      RECT  218.6 24.2 219.4 25.0 ;
      RECT  223.4 24.2 224.2 25.0 ;
      RECT  45.8 29.0 46.6 29.8 ;
      RECT  50.6 29.0 51.4 29.8 ;
      RECT  55.4 29.0 56.2 29.8 ;
      RECT  60.2 29.0 61.0 29.8 ;
      RECT  65.0 29.0 65.8 29.8 ;
      RECT  69.8 29.0 70.6 29.8 ;
      RECT  74.6 29.0 75.4 29.8 ;
      RECT  79.4 29.0 80.2 29.8 ;
      RECT  84.2 29.0 85.0 29.8 ;
      RECT  89.0 29.0 89.8 29.8 ;
      RECT  93.8 29.0 94.6 29.8 ;
      RECT  98.6 29.0 99.4 29.8 ;
      RECT  103.4 29.0 104.2 29.8 ;
      RECT  108.2 29.0 109.0 29.8 ;
      RECT  113.0 29.0 113.8 29.8 ;
      RECT  117.8 29.0 118.6 29.8 ;
      RECT  122.6 29.0 123.4 29.8 ;
      RECT  127.4 29.0 128.2 29.8 ;
      RECT  132.2 29.0 133.0 29.8 ;
      RECT  137.0 29.0 137.8 29.8 ;
      RECT  141.8 29.0 142.6 29.8 ;
      RECT  146.6 29.0 147.4 29.8 ;
      RECT  151.4 29.0 152.2 29.8 ;
      RECT  156.2 29.0 157.0 29.8 ;
      RECT  161.0 29.0 161.8 29.8 ;
      RECT  165.8 29.0 166.6 29.8 ;
      RECT  170.6 29.0 171.4 29.8 ;
      RECT  175.4 29.0 176.2 29.8 ;
      RECT  180.2 29.0 181.0 29.8 ;
      RECT  185.0 29.0 185.8 29.8 ;
      RECT  189.8 29.0 190.6 29.8 ;
      RECT  194.6 29.0 195.4 29.8 ;
      RECT  199.4 29.0 200.2 29.8 ;
      RECT  204.2 29.0 205.0 29.8 ;
      RECT  209.0 29.0 209.8 29.8 ;
      RECT  213.8 29.0 214.6 29.8 ;
      RECT  218.6 29.0 219.4 29.8 ;
      RECT  223.4 29.0 224.2 29.8 ;
      RECT  84.2 33.8 85.0 34.6 ;
      RECT  89.0 33.8 89.8 34.6 ;
      RECT  93.8 33.8 94.6 34.6 ;
      RECT  98.6 33.8 99.4 34.6 ;
      RECT  103.4 33.8 104.2 34.6 ;
      RECT  108.2 33.8 109.0 34.6 ;
      RECT  113.0 33.8 113.8 34.6 ;
      RECT  117.8 33.8 118.6 34.6 ;
      RECT  122.6 33.8 123.4 34.6 ;
      RECT  127.4 33.8 128.2 34.6 ;
      RECT  132.2 33.8 133.0 34.6 ;
      RECT  137.0 33.8 137.8 34.6 ;
      RECT  141.8 33.8 142.6 34.6 ;
      RECT  146.6 33.8 147.4 34.6 ;
      RECT  151.4 33.8 152.2 34.6 ;
      RECT  156.2 33.8 157.0 34.6 ;
      RECT  161.0 33.8 161.8 34.6 ;
      RECT  165.8 33.8 166.6 34.6 ;
      RECT  170.6 33.8 171.4 34.6 ;
      RECT  175.4 33.8 176.2 34.6 ;
      RECT  180.2 33.8 181.0 34.6 ;
      RECT  185.0 33.8 185.8 34.6 ;
      RECT  189.8 33.8 190.6 34.6 ;
      RECT  194.6 33.8 195.4 34.6 ;
      RECT  199.4 33.8 200.2 34.6 ;
      RECT  204.2 33.8 205.0 34.6 ;
      RECT  209.0 33.8 209.8 34.6 ;
      RECT  213.8 33.8 214.6 34.6 ;
      RECT  218.6 33.8 219.4 34.6 ;
      RECT  223.4 33.8 224.2 34.6 ;
      RECT  2.6 38.6 3.4 39.4 ;
      RECT  7.4 38.6 8.2 39.4 ;
      RECT  12.2 38.6 13.0 39.4 ;
      RECT  17.0 38.6 17.8 39.4 ;
      RECT  21.8 38.6 22.6 39.4 ;
      RECT  26.6 38.6 27.4 39.4 ;
      RECT  31.4 38.6 32.2 39.4 ;
      RECT  36.2 38.6 37.0 39.4 ;
      RECT  41.0 38.6 41.8 39.4 ;
      RECT  60.2 38.6 61.0 39.4 ;
      RECT  65.0 38.6 65.8 39.4 ;
      RECT  69.8 38.6 70.6 39.4 ;
      RECT  74.6 38.6 75.4 39.4 ;
      RECT  79.4 38.6 80.2 39.4 ;
      RECT  84.2 38.6 85.0 39.4 ;
      RECT  89.0 38.6 89.8 39.4 ;
      RECT  93.8 38.6 94.6 39.4 ;
      RECT  98.6 38.6 99.4 39.4 ;
      RECT  103.4 38.6 104.2 39.4 ;
      RECT  108.2 38.6 109.0 39.4 ;
      RECT  113.0 38.6 113.8 39.4 ;
      RECT  117.8 38.6 118.6 39.4 ;
      RECT  122.6 38.6 123.4 39.4 ;
      RECT  127.4 38.6 128.2 39.4 ;
      RECT  132.2 38.6 133.0 39.4 ;
      RECT  137.0 38.6 137.8 39.4 ;
      RECT  141.8 38.6 142.6 39.4 ;
      RECT  146.6 38.6 147.4 39.4 ;
      RECT  151.4 38.6 152.2 39.4 ;
      RECT  156.2 38.6 157.0 39.4 ;
      RECT  161.0 38.6 161.8 39.4 ;
      RECT  165.8 38.6 166.6 39.4 ;
      RECT  170.6 38.6 171.4 39.4 ;
      RECT  175.4 38.6 176.2 39.4 ;
      RECT  180.2 38.6 181.0 39.4 ;
      RECT  185.0 38.6 185.8 39.4 ;
      RECT  189.8 38.6 190.6 39.4 ;
      RECT  194.6 38.6 195.4 39.4 ;
      RECT  199.4 38.6 200.2 39.4 ;
      RECT  204.2 38.6 205.0 39.4 ;
      RECT  209.0 38.6 209.8 39.4 ;
      RECT  213.8 38.6 214.6 39.4 ;
      RECT  218.6 38.6 219.4 39.4 ;
      RECT  223.4 38.6 224.2 39.4 ;
      RECT  2.6 43.4 3.4 44.2 ;
      RECT  7.4 43.4 8.2 44.2 ;
      RECT  12.2 43.4 13.0 44.2 ;
      RECT  17.0 43.4 17.8 44.2 ;
      RECT  21.8 43.4 22.6 44.2 ;
      RECT  26.6 43.4 27.4 44.2 ;
      RECT  31.4 43.4 32.2 44.2 ;
      RECT  36.2 43.4 37.0 44.2 ;
      RECT  41.0 43.4 41.8 44.2 ;
      RECT  45.8 43.4 46.6 44.2 ;
      RECT  50.6 43.4 51.4 44.2 ;
      RECT  55.4 43.4 56.2 44.2 ;
      RECT  60.2 43.4 61.0 44.2 ;
      RECT  65.0 43.4 65.8 44.2 ;
      RECT  69.8 43.4 70.6 44.2 ;
      RECT  74.6 43.4 75.4 44.2 ;
      RECT  79.4 43.4 80.2 44.2 ;
      RECT  84.2 43.4 85.0 44.2 ;
      RECT  89.0 43.4 89.8 44.2 ;
      RECT  93.8 43.4 94.6 44.2 ;
      RECT  98.6 43.4 99.4 44.2 ;
      RECT  103.4 43.4 104.2 44.2 ;
      RECT  108.2 43.4 109.0 44.2 ;
      RECT  113.0 43.4 113.8 44.2 ;
      RECT  117.8 43.4 118.6 44.2 ;
      RECT  122.6 43.4 123.4 44.2 ;
      RECT  127.4 43.4 128.2 44.2 ;
      RECT  132.2 43.4 133.0 44.2 ;
      RECT  137.0 43.4 137.8 44.2 ;
      RECT  141.8 43.4 142.6 44.2 ;
      RECT  146.6 43.4 147.4 44.2 ;
      RECT  151.4 43.4 152.2 44.2 ;
      RECT  156.2 43.4 157.0 44.2 ;
      RECT  161.0 43.4 161.8 44.2 ;
      RECT  165.8 43.4 166.6 44.2 ;
      RECT  170.6 43.4 171.4 44.2 ;
      RECT  175.4 43.4 176.2 44.2 ;
      RECT  180.2 43.4 181.0 44.2 ;
      RECT  185.0 43.4 185.8 44.2 ;
      RECT  189.8 43.4 190.6 44.2 ;
      RECT  194.6 43.4 195.4 44.2 ;
      RECT  199.4 43.4 200.2 44.2 ;
      RECT  204.2 43.4 205.0 44.2 ;
      RECT  209.0 43.4 209.8 44.2 ;
      RECT  213.8 43.4 214.6 44.2 ;
      RECT  218.6 43.4 219.4 44.2 ;
      RECT  223.4 43.4 224.2 44.2 ;
      RECT  2.6 48.2 3.4 49.0 ;
      RECT  7.4 48.2 8.2 49.0 ;
      RECT  12.2 48.2 13.0 49.0 ;
      RECT  17.0 48.2 17.8 49.0 ;
      RECT  21.8 48.2 22.6 49.0 ;
      RECT  26.6 48.2 27.4 49.0 ;
      RECT  31.4 48.2 32.2 49.0 ;
      RECT  36.2 48.2 37.0 49.0 ;
      RECT  41.0 48.2 41.8 49.0 ;
      RECT  45.8 48.2 46.6 49.0 ;
      RECT  50.6 48.2 51.4 49.0 ;
      RECT  55.4 48.2 56.2 49.0 ;
      RECT  60.2 48.2 61.0 49.0 ;
      RECT  65.0 48.2 65.8 49.0 ;
      RECT  69.8 48.2 70.6 49.0 ;
      RECT  74.6 48.2 75.4 49.0 ;
      RECT  79.4 48.2 80.2 49.0 ;
      RECT  84.2 48.2 85.0 49.0 ;
      RECT  89.0 48.2 89.8 49.0 ;
      RECT  93.8 48.2 94.6 49.0 ;
      RECT  98.6 48.2 99.4 49.0 ;
      RECT  103.4 48.2 104.2 49.0 ;
      RECT  108.2 48.2 109.0 49.0 ;
      RECT  113.0 48.2 113.8 49.0 ;
      RECT  117.8 48.2 118.6 49.0 ;
      RECT  122.6 48.2 123.4 49.0 ;
      RECT  127.4 48.2 128.2 49.0 ;
      RECT  132.2 48.2 133.0 49.0 ;
      RECT  137.0 48.2 137.8 49.0 ;
      RECT  141.8 48.2 142.6 49.0 ;
      RECT  146.6 48.2 147.4 49.0 ;
      RECT  151.4 48.2 152.2 49.0 ;
      RECT  156.2 48.2 157.0 49.0 ;
      RECT  161.0 48.2 161.8 49.0 ;
      RECT  165.8 48.2 166.6 49.0 ;
      RECT  170.6 48.2 171.4 49.0 ;
      RECT  175.4 48.2 176.2 49.0 ;
      RECT  180.2 48.2 181.0 49.0 ;
      RECT  185.0 48.2 185.8 49.0 ;
      RECT  189.8 48.2 190.6 49.0 ;
      RECT  194.6 48.2 195.4 49.0 ;
      RECT  199.4 48.2 200.2 49.0 ;
      RECT  204.2 48.2 205.0 49.0 ;
      RECT  209.0 48.2 209.8 49.0 ;
      RECT  213.8 48.2 214.6 49.0 ;
      RECT  218.6 48.2 219.4 49.0 ;
      RECT  223.4 48.2 224.2 49.0 ;
      RECT  2.6 53.0 3.4 53.8 ;
      RECT  7.4 53.0 8.2 53.8 ;
      RECT  12.2 53.0 13.0 53.8 ;
      RECT  17.0 53.0 17.8 53.8 ;
      RECT  21.8 53.0 22.6 53.8 ;
      RECT  26.6 53.0 27.4 53.8 ;
      RECT  31.4 53.0 32.2 53.8 ;
      RECT  36.2 53.0 37.0 53.8 ;
      RECT  41.0 53.0 41.8 53.8 ;
      RECT  45.8 53.0 46.6 53.8 ;
      RECT  50.6 53.0 51.4 53.8 ;
      RECT  55.4 53.0 56.2 53.8 ;
      RECT  60.2 53.0 61.0 53.8 ;
      RECT  65.0 53.0 65.8 53.8 ;
      RECT  69.8 53.0 70.6 53.8 ;
      RECT  74.6 53.0 75.4 53.8 ;
      RECT  79.4 53.0 80.2 53.8 ;
      RECT  2.6 57.8 3.4 58.6 ;
      RECT  7.4 57.8 8.2 58.6 ;
      RECT  12.2 57.8 13.0 58.6 ;
      RECT  17.0 57.8 17.8 58.6 ;
      RECT  21.8 57.8 22.6 58.6 ;
      RECT  26.6 57.8 27.4 58.6 ;
      RECT  31.4 57.8 32.2 58.6 ;
      RECT  36.2 57.8 37.0 58.6 ;
      RECT  41.0 57.8 41.8 58.6 ;
      RECT  45.8 57.8 46.6 58.6 ;
      RECT  50.6 57.8 51.4 58.6 ;
      RECT  55.4 57.8 56.2 58.6 ;
      RECT  60.2 57.8 61.0 58.6 ;
      RECT  65.0 57.8 65.8 58.6 ;
      RECT  69.8 57.8 70.6 58.6 ;
      RECT  74.6 57.8 75.4 58.6 ;
      RECT  79.4 57.8 80.2 58.6 ;
      RECT  84.2 57.8 85.0 58.6 ;
      RECT  89.0 57.8 89.8 58.6 ;
      RECT  93.8 57.8 94.6 58.6 ;
      RECT  98.6 57.8 99.4 58.6 ;
      RECT  103.4 57.8 104.2 58.6 ;
      RECT  108.2 57.8 109.0 58.6 ;
      RECT  113.0 57.8 113.8 58.6 ;
      RECT  117.8 57.8 118.6 58.6 ;
      RECT  122.6 57.8 123.4 58.6 ;
      RECT  127.4 57.8 128.2 58.6 ;
      RECT  132.2 57.8 133.0 58.6 ;
      RECT  137.0 57.8 137.8 58.6 ;
      RECT  141.8 57.8 142.6 58.6 ;
      RECT  146.6 57.8 147.4 58.6 ;
      RECT  151.4 57.8 152.2 58.6 ;
      RECT  156.2 57.8 157.0 58.6 ;
      RECT  161.0 57.8 161.8 58.6 ;
      RECT  165.8 57.8 166.6 58.6 ;
      RECT  170.6 57.8 171.4 58.6 ;
      RECT  175.4 57.8 176.2 58.6 ;
      RECT  180.2 57.8 181.0 58.6 ;
      RECT  185.0 57.8 185.8 58.6 ;
      RECT  189.8 57.8 190.6 58.6 ;
      RECT  194.6 57.8 195.4 58.6 ;
      RECT  199.4 57.8 200.2 58.6 ;
      RECT  204.2 57.8 205.0 58.6 ;
      RECT  209.0 57.8 209.8 58.6 ;
      RECT  213.8 57.8 214.6 58.6 ;
      RECT  218.6 57.8 219.4 58.6 ;
      RECT  223.4 57.8 224.2 58.6 ;
      RECT  2.6 62.6 3.4 63.4 ;
      RECT  7.4 62.6 8.2 63.4 ;
      RECT  12.2 62.6 13.0 63.4 ;
      RECT  17.0 62.6 17.8 63.4 ;
      RECT  21.8 62.6 22.6 63.4 ;
      RECT  26.6 62.6 27.4 63.4 ;
      RECT  31.4 62.6 32.2 63.4 ;
      RECT  36.2 62.6 37.0 63.4 ;
      RECT  41.0 62.6 41.8 63.4 ;
      RECT  45.8 62.6 46.6 63.4 ;
      RECT  50.6 62.6 51.4 63.4 ;
      RECT  55.4 62.6 56.2 63.4 ;
      RECT  60.2 62.6 61.0 63.4 ;
      RECT  65.0 62.6 65.8 63.4 ;
      RECT  69.8 62.6 70.6 63.4 ;
      RECT  74.6 62.6 75.4 63.4 ;
      RECT  79.4 62.6 80.2 63.4 ;
      RECT  89.0 62.6 89.8 63.4 ;
      RECT  93.8 62.6 94.6 63.4 ;
      RECT  98.6 62.6 99.4 63.4 ;
      RECT  103.4 62.6 104.2 63.4 ;
      RECT  108.2 62.6 109.0 63.4 ;
      RECT  113.0 62.6 113.8 63.4 ;
      RECT  117.8 62.6 118.6 63.4 ;
      RECT  122.6 62.6 123.4 63.4 ;
      RECT  127.4 62.6 128.2 63.4 ;
      RECT  132.2 62.6 133.0 63.4 ;
      RECT  137.0 62.6 137.8 63.4 ;
      RECT  141.8 62.6 142.6 63.4 ;
      RECT  146.6 62.6 147.4 63.4 ;
      RECT  151.4 62.6 152.2 63.4 ;
      RECT  156.2 62.6 157.0 63.4 ;
      RECT  161.0 62.6 161.8 63.4 ;
      RECT  165.8 62.6 166.6 63.4 ;
      RECT  170.6 62.6 171.4 63.4 ;
      RECT  175.4 62.6 176.2 63.4 ;
      RECT  180.2 62.6 181.0 63.4 ;
      RECT  185.0 62.6 185.8 63.4 ;
      RECT  189.8 62.6 190.6 63.4 ;
      RECT  194.6 62.6 195.4 63.4 ;
      RECT  199.4 62.6 200.2 63.4 ;
      RECT  204.2 62.6 205.0 63.4 ;
      RECT  209.0 62.6 209.8 63.4 ;
      RECT  213.8 62.6 214.6 63.4 ;
      RECT  218.6 62.6 219.4 63.4 ;
      RECT  223.4 62.6 224.2 63.4 ;
      RECT  2.6 67.4 3.4 68.2 ;
      RECT  7.4 67.4 8.2 68.2 ;
      RECT  12.2 67.4 13.0 68.2 ;
      RECT  17.0 67.4 17.8 68.2 ;
      RECT  21.8 67.4 22.6 68.2 ;
      RECT  26.6 67.4 27.4 68.2 ;
      RECT  31.4 67.4 32.2 68.2 ;
      RECT  36.2 67.4 37.0 68.2 ;
      RECT  41.0 67.4 41.8 68.2 ;
      RECT  45.8 67.4 46.6 68.2 ;
      RECT  50.6 67.4 51.4 68.2 ;
      RECT  55.4 67.4 56.2 68.2 ;
      RECT  60.2 67.4 61.0 68.2 ;
      RECT  65.0 67.4 65.8 68.2 ;
      RECT  69.8 67.4 70.6 68.2 ;
      RECT  74.6 67.4 75.4 68.2 ;
      RECT  79.4 67.4 80.2 68.2 ;
      RECT  84.2 67.4 85.0 68.2 ;
      RECT  89.0 67.4 89.8 68.2 ;
      RECT  93.8 67.4 94.6 68.2 ;
      RECT  98.6 67.4 99.4 68.2 ;
      RECT  103.4 67.4 104.2 68.2 ;
      RECT  108.2 67.4 109.0 68.2 ;
      RECT  113.0 67.4 113.8 68.2 ;
      RECT  117.8 67.4 118.6 68.2 ;
      RECT  122.6 67.4 123.4 68.2 ;
      RECT  127.4 67.4 128.2 68.2 ;
      RECT  132.2 67.4 133.0 68.2 ;
      RECT  137.0 67.4 137.8 68.2 ;
      RECT  141.8 67.4 142.6 68.2 ;
      RECT  146.6 67.4 147.4 68.2 ;
      RECT  151.4 67.4 152.2 68.2 ;
      RECT  156.2 67.4 157.0 68.2 ;
      RECT  161.0 67.4 161.8 68.2 ;
      RECT  165.8 67.4 166.6 68.2 ;
      RECT  170.6 67.4 171.4 68.2 ;
      RECT  175.4 67.4 176.2 68.2 ;
      RECT  180.2 67.4 181.0 68.2 ;
      RECT  185.0 67.4 185.8 68.2 ;
      RECT  189.8 67.4 190.6 68.2 ;
      RECT  2.6 72.2 3.4 73.0 ;
      RECT  7.4 72.2 8.2 73.0 ;
      RECT  12.2 72.2 13.0 73.0 ;
      RECT  17.0 72.2 17.8 73.0 ;
      RECT  21.8 72.2 22.6 73.0 ;
      RECT  26.6 72.2 27.4 73.0 ;
      RECT  31.4 72.2 32.2 73.0 ;
      RECT  36.2 72.2 37.0 73.0 ;
      RECT  41.0 72.2 41.8 73.0 ;
      RECT  45.8 72.2 46.6 73.0 ;
      RECT  50.6 72.2 51.4 73.0 ;
      RECT  55.4 72.2 56.2 73.0 ;
      RECT  60.2 72.2 61.0 73.0 ;
      RECT  65.0 72.2 65.8 73.0 ;
      RECT  69.8 72.2 70.6 73.0 ;
      RECT  74.6 72.2 75.4 73.0 ;
      RECT  79.4 72.2 80.2 73.0 ;
      RECT  189.8 72.2 190.6 73.0 ;
      RECT  194.6 72.2 195.4 73.0 ;
      RECT  199.4 72.2 200.2 73.0 ;
      RECT  204.2 72.2 205.0 73.0 ;
      RECT  209.0 72.2 209.8 73.0 ;
      RECT  213.8 72.2 214.6 73.0 ;
      RECT  218.6 72.2 219.4 73.0 ;
      RECT  223.4 72.2 224.2 73.0 ;
      RECT  2.6 77.0 3.4 77.8 ;
      RECT  7.4 77.0 8.2 77.8 ;
      RECT  12.2 77.0 13.0 77.8 ;
      RECT  17.0 77.0 17.8 77.8 ;
      RECT  21.8 77.0 22.6 77.8 ;
      RECT  26.6 77.0 27.4 77.8 ;
      RECT  31.4 77.0 32.2 77.8 ;
      RECT  36.2 77.0 37.0 77.8 ;
      RECT  41.0 77.0 41.8 77.8 ;
      RECT  45.8 77.0 46.6 77.8 ;
      RECT  50.6 77.0 51.4 77.8 ;
      RECT  55.4 77.0 56.2 77.8 ;
      RECT  60.2 77.0 61.0 77.8 ;
      RECT  65.0 77.0 65.8 77.8 ;
      RECT  69.8 77.0 70.6 77.8 ;
      RECT  74.6 77.0 75.4 77.8 ;
      RECT  79.4 77.0 80.2 77.8 ;
      RECT  84.2 77.0 85.0 77.8 ;
      RECT  89.0 77.0 89.8 77.8 ;
      RECT  93.8 77.0 94.6 77.8 ;
      RECT  98.6 77.0 99.4 77.8 ;
      RECT  103.4 77.0 104.2 77.8 ;
      RECT  108.2 77.0 109.0 77.8 ;
      RECT  113.0 77.0 113.8 77.8 ;
      RECT  117.8 77.0 118.6 77.8 ;
      RECT  122.6 77.0 123.4 77.8 ;
      RECT  127.4 77.0 128.2 77.8 ;
      RECT  132.2 77.0 133.0 77.8 ;
      RECT  137.0 77.0 137.8 77.8 ;
      RECT  141.8 77.0 142.6 77.8 ;
      RECT  146.6 77.0 147.4 77.8 ;
      RECT  151.4 77.0 152.2 77.8 ;
      RECT  156.2 77.0 157.0 77.8 ;
      RECT  161.0 77.0 161.8 77.8 ;
      RECT  165.8 77.0 166.6 77.8 ;
      RECT  170.6 77.0 171.4 77.8 ;
      RECT  175.4 77.0 176.2 77.8 ;
      RECT  180.2 77.0 181.0 77.8 ;
      RECT  185.0 77.0 185.8 77.8 ;
      RECT  189.8 77.0 190.6 77.8 ;
      RECT  194.6 77.0 195.4 77.8 ;
      RECT  199.4 77.0 200.2 77.8 ;
      RECT  204.2 77.0 205.0 77.8 ;
      RECT  209.0 77.0 209.8 77.8 ;
      RECT  213.8 77.0 214.6 77.8 ;
      RECT  218.6 77.0 219.4 77.8 ;
      RECT  223.4 77.0 224.2 77.8 ;
      RECT  2.6 81.8 3.4 82.6 ;
      RECT  7.4 81.8 8.2 82.6 ;
      RECT  12.2 81.8 13.0 82.6 ;
      RECT  17.0 81.8 17.8 82.6 ;
      RECT  21.8 81.8 22.6 82.6 ;
      RECT  26.6 81.8 27.4 82.6 ;
      RECT  31.4 81.8 32.2 82.6 ;
      RECT  36.2 81.8 37.0 82.6 ;
      RECT  41.0 81.8 41.8 82.6 ;
      RECT  45.8 81.8 46.6 82.6 ;
      RECT  50.6 81.8 51.4 82.6 ;
      RECT  55.4 81.8 56.2 82.6 ;
      RECT  60.2 81.8 61.0 82.6 ;
      RECT  65.0 81.8 65.8 82.6 ;
      RECT  69.8 81.8 70.6 82.6 ;
      RECT  74.6 81.8 75.4 82.6 ;
      RECT  79.4 81.8 80.2 82.6 ;
      RECT  84.2 81.8 85.0 82.6 ;
      RECT  89.0 81.8 89.8 82.6 ;
      RECT  93.8 81.8 94.6 82.6 ;
      RECT  98.6 81.8 99.4 82.6 ;
      RECT  103.4 81.8 104.2 82.6 ;
      RECT  108.2 81.8 109.0 82.6 ;
      RECT  113.0 81.8 113.8 82.6 ;
      RECT  117.8 81.8 118.6 82.6 ;
      RECT  122.6 81.8 123.4 82.6 ;
      RECT  127.4 81.8 128.2 82.6 ;
      RECT  132.2 81.8 133.0 82.6 ;
      RECT  137.0 81.8 137.8 82.6 ;
      RECT  141.8 81.8 142.6 82.6 ;
      RECT  146.6 81.8 147.4 82.6 ;
      RECT  151.4 81.8 152.2 82.6 ;
      RECT  156.2 81.8 157.0 82.6 ;
      RECT  161.0 81.8 161.8 82.6 ;
      RECT  165.8 81.8 166.6 82.6 ;
      RECT  170.6 81.8 171.4 82.6 ;
      RECT  175.4 81.8 176.2 82.6 ;
      RECT  180.2 81.8 181.0 82.6 ;
      RECT  185.0 81.8 185.8 82.6 ;
      RECT  189.8 81.8 190.6 82.6 ;
      RECT  194.6 81.8 195.4 82.6 ;
      RECT  2.6 86.6 3.4 87.4 ;
      RECT  7.4 86.6 8.2 87.4 ;
      RECT  12.2 86.6 13.0 87.4 ;
      RECT  17.0 86.6 17.8 87.4 ;
      RECT  21.8 86.6 22.6 87.4 ;
      RECT  26.6 86.6 27.4 87.4 ;
      RECT  31.4 86.6 32.2 87.4 ;
      RECT  36.2 86.6 37.0 87.4 ;
      RECT  41.0 86.6 41.8 87.4 ;
      RECT  45.8 86.6 46.6 87.4 ;
      RECT  50.6 86.6 51.4 87.4 ;
      RECT  55.4 86.6 56.2 87.4 ;
      RECT  60.2 86.6 61.0 87.4 ;
      RECT  65.0 86.6 65.8 87.4 ;
      RECT  69.8 86.6 70.6 87.4 ;
      RECT  74.6 86.6 75.4 87.4 ;
      RECT  79.4 86.6 80.2 87.4 ;
      RECT  84.2 86.6 85.0 87.4 ;
      RECT  89.0 86.6 89.8 87.4 ;
      RECT  93.8 86.6 94.6 87.4 ;
      RECT  98.6 86.6 99.4 87.4 ;
      RECT  103.4 86.6 104.2 87.4 ;
      RECT  108.2 86.6 109.0 87.4 ;
      RECT  113.0 86.6 113.8 87.4 ;
      RECT  117.8 86.6 118.6 87.4 ;
      RECT  122.6 86.6 123.4 87.4 ;
      RECT  127.4 86.6 128.2 87.4 ;
      RECT  132.2 86.6 133.0 87.4 ;
      RECT  137.0 86.6 137.8 87.4 ;
      RECT  141.8 86.6 142.6 87.4 ;
      RECT  146.6 86.6 147.4 87.4 ;
      RECT  151.4 86.6 152.2 87.4 ;
      RECT  156.2 86.6 157.0 87.4 ;
      RECT  161.0 86.6 161.8 87.4 ;
      RECT  165.8 86.6 166.6 87.4 ;
      RECT  170.6 86.6 171.4 87.4 ;
      RECT  175.4 86.6 176.2 87.4 ;
      RECT  180.2 86.6 181.0 87.4 ;
      RECT  185.0 86.6 185.8 87.4 ;
      RECT  189.8 86.6 190.6 87.4 ;
      RECT  194.6 86.6 195.4 87.4 ;
      RECT  199.4 86.6 200.2 87.4 ;
      RECT  204.2 86.6 205.0 87.4 ;
      RECT  209.0 86.6 209.8 87.4 ;
      RECT  213.8 86.6 214.6 87.4 ;
      RECT  218.6 86.6 219.4 87.4 ;
      RECT  223.4 86.6 224.2 87.4 ;
      RECT  2.6 91.4 3.4 92.2 ;
      RECT  7.4 91.4 8.2 92.2 ;
      RECT  12.2 91.4 13.0 92.2 ;
      RECT  17.0 91.4 17.8 92.2 ;
      RECT  21.8 91.4 22.6 92.2 ;
      RECT  26.6 91.4 27.4 92.2 ;
      RECT  31.4 91.4 32.2 92.2 ;
      RECT  36.2 91.4 37.0 92.2 ;
      RECT  41.0 91.4 41.8 92.2 ;
      RECT  45.8 91.4 46.6 92.2 ;
      RECT  50.6 91.4 51.4 92.2 ;
      RECT  55.4 91.4 56.2 92.2 ;
      RECT  60.2 91.4 61.0 92.2 ;
      RECT  65.0 91.4 65.8 92.2 ;
      RECT  69.8 91.4 70.6 92.2 ;
      RECT  74.6 91.4 75.4 92.2 ;
      RECT  79.4 91.4 80.2 92.2 ;
      RECT  185.0 91.4 185.8 92.2 ;
      RECT  189.8 91.4 190.6 92.2 ;
      RECT  194.6 91.4 195.4 92.2 ;
      RECT  199.4 91.4 200.2 92.2 ;
      RECT  204.2 91.4 205.0 92.2 ;
      RECT  209.0 91.4 209.8 92.2 ;
      RECT  213.8 91.4 214.6 92.2 ;
      RECT  218.6 91.4 219.4 92.2 ;
      RECT  223.4 91.4 224.2 92.2 ;
      RECT  2.6 96.2 3.4 97.0 ;
      RECT  7.4 96.2 8.2 97.0 ;
      RECT  12.2 96.2 13.0 97.0 ;
      RECT  17.0 96.2 17.8 97.0 ;
      RECT  21.8 96.2 22.6 97.0 ;
      RECT  26.6 96.2 27.4 97.0 ;
      RECT  31.4 96.2 32.2 97.0 ;
      RECT  36.2 96.2 37.0 97.0 ;
      RECT  41.0 96.2 41.8 97.0 ;
      RECT  45.8 96.2 46.6 97.0 ;
      RECT  50.6 96.2 51.4 97.0 ;
      RECT  55.4 96.2 56.2 97.0 ;
      RECT  60.2 96.2 61.0 97.0 ;
      RECT  65.0 96.2 65.8 97.0 ;
      RECT  69.8 96.2 70.6 97.0 ;
      RECT  74.6 96.2 75.4 97.0 ;
      RECT  79.4 96.2 80.2 97.0 ;
      RECT  84.2 96.2 85.0 97.0 ;
      RECT  89.0 96.2 89.8 97.0 ;
      RECT  93.8 96.2 94.6 97.0 ;
      RECT  98.6 96.2 99.4 97.0 ;
      RECT  103.4 96.2 104.2 97.0 ;
      RECT  108.2 96.2 109.0 97.0 ;
      RECT  113.0 96.2 113.8 97.0 ;
      RECT  117.8 96.2 118.6 97.0 ;
      RECT  122.6 96.2 123.4 97.0 ;
      RECT  127.4 96.2 128.2 97.0 ;
      RECT  132.2 96.2 133.0 97.0 ;
      RECT  137.0 96.2 137.8 97.0 ;
      RECT  141.8 96.2 142.6 97.0 ;
      RECT  146.6 96.2 147.4 97.0 ;
      RECT  151.4 96.2 152.2 97.0 ;
      RECT  156.2 96.2 157.0 97.0 ;
      RECT  161.0 96.2 161.8 97.0 ;
      RECT  165.8 96.2 166.6 97.0 ;
      RECT  170.6 96.2 171.4 97.0 ;
      RECT  175.4 96.2 176.2 97.0 ;
      RECT  180.2 96.2 181.0 97.0 ;
      RECT  185.0 96.2 185.8 97.0 ;
      RECT  189.8 96.2 190.6 97.0 ;
      RECT  194.6 96.2 195.4 97.0 ;
      RECT  199.4 96.2 200.2 97.0 ;
      RECT  204.2 96.2 205.0 97.0 ;
      RECT  209.0 96.2 209.8 97.0 ;
      RECT  213.8 96.2 214.6 97.0 ;
      RECT  218.6 96.2 219.4 97.0 ;
      RECT  223.4 96.2 224.2 97.0 ;
      RECT  2.6 101.0 3.4 101.8 ;
      RECT  7.4 101.0 8.2 101.8 ;
      RECT  12.2 101.0 13.0 101.8 ;
      RECT  17.0 101.0 17.8 101.8 ;
      RECT  21.8 101.0 22.6 101.8 ;
      RECT  26.6 101.0 27.4 101.8 ;
      RECT  31.4 101.0 32.2 101.8 ;
      RECT  36.2 101.0 37.0 101.8 ;
      RECT  41.0 101.0 41.8 101.8 ;
      RECT  45.8 101.0 46.6 101.8 ;
      RECT  50.6 101.0 51.4 101.8 ;
      RECT  55.4 101.0 56.2 101.8 ;
      RECT  60.2 101.0 61.0 101.8 ;
      RECT  65.0 101.0 65.8 101.8 ;
      RECT  69.8 101.0 70.6 101.8 ;
      RECT  74.6 101.0 75.4 101.8 ;
      RECT  79.4 101.0 80.2 101.8 ;
      RECT  89.0 101.0 89.8 101.8 ;
      RECT  93.8 101.0 94.6 101.8 ;
      RECT  98.6 101.0 99.4 101.8 ;
      RECT  103.4 101.0 104.2 101.8 ;
      RECT  108.2 101.0 109.0 101.8 ;
      RECT  113.0 101.0 113.8 101.8 ;
      RECT  117.8 101.0 118.6 101.8 ;
      RECT  122.6 101.0 123.4 101.8 ;
      RECT  127.4 101.0 128.2 101.8 ;
      RECT  132.2 101.0 133.0 101.8 ;
      RECT  137.0 101.0 137.8 101.8 ;
      RECT  141.8 101.0 142.6 101.8 ;
      RECT  146.6 101.0 147.4 101.8 ;
      RECT  151.4 101.0 152.2 101.8 ;
      RECT  156.2 101.0 157.0 101.8 ;
      RECT  161.0 101.0 161.8 101.8 ;
      RECT  165.8 101.0 166.6 101.8 ;
      RECT  170.6 101.0 171.4 101.8 ;
      RECT  175.4 101.0 176.2 101.8 ;
      RECT  180.2 101.0 181.0 101.8 ;
      RECT  185.0 101.0 185.8 101.8 ;
      RECT  189.8 101.0 190.6 101.8 ;
      RECT  194.6 101.0 195.4 101.8 ;
      RECT  199.4 101.0 200.2 101.8 ;
      RECT  204.2 101.0 205.0 101.8 ;
      RECT  209.0 101.0 209.8 101.8 ;
      RECT  213.8 101.0 214.6 101.8 ;
      RECT  218.6 101.0 219.4 101.8 ;
      RECT  223.4 101.0 224.2 101.8 ;
      RECT  2.6 105.8 3.4 106.6 ;
      RECT  7.4 105.8 8.2 106.6 ;
      RECT  12.2 105.8 13.0 106.6 ;
      RECT  17.0 105.8 17.8 106.6 ;
      RECT  21.8 105.8 22.6 106.6 ;
      RECT  26.6 105.8 27.4 106.6 ;
      RECT  31.4 105.8 32.2 106.6 ;
      RECT  36.2 105.8 37.0 106.6 ;
      RECT  41.0 105.8 41.8 106.6 ;
      RECT  45.8 105.8 46.6 106.6 ;
      RECT  50.6 105.8 51.4 106.6 ;
      RECT  55.4 105.8 56.2 106.6 ;
      RECT  60.2 105.8 61.0 106.6 ;
      RECT  65.0 105.8 65.8 106.6 ;
      RECT  69.8 105.8 70.6 106.6 ;
      RECT  74.6 105.8 75.4 106.6 ;
      RECT  79.4 105.8 80.2 106.6 ;
      RECT  84.2 105.8 85.0 106.6 ;
      RECT  89.0 105.8 89.8 106.6 ;
      RECT  93.8 105.8 94.6 106.6 ;
      RECT  98.6 105.8 99.4 106.6 ;
      RECT  103.4 105.8 104.2 106.6 ;
      RECT  108.2 105.8 109.0 106.6 ;
      RECT  113.0 105.8 113.8 106.6 ;
      RECT  117.8 105.8 118.6 106.6 ;
      RECT  122.6 105.8 123.4 106.6 ;
      RECT  127.4 105.8 128.2 106.6 ;
      RECT  132.2 105.8 133.0 106.6 ;
      RECT  137.0 105.8 137.8 106.6 ;
      RECT  141.8 105.8 142.6 106.6 ;
      RECT  146.6 105.8 147.4 106.6 ;
      RECT  151.4 105.8 152.2 106.6 ;
      RECT  156.2 105.8 157.0 106.6 ;
      RECT  161.0 105.8 161.8 106.6 ;
      RECT  165.8 105.8 166.6 106.6 ;
      RECT  170.6 105.8 171.4 106.6 ;
      RECT  175.4 105.8 176.2 106.6 ;
      RECT  180.2 105.8 181.0 106.6 ;
      RECT  185.0 105.8 185.8 106.6 ;
      RECT  189.8 105.8 190.6 106.6 ;
      RECT  194.6 105.8 195.4 106.6 ;
      RECT  199.4 105.8 200.2 106.6 ;
      RECT  204.2 105.8 205.0 106.6 ;
      RECT  209.0 105.8 209.8 106.6 ;
      RECT  213.8 105.8 214.6 106.6 ;
      RECT  218.6 105.8 219.4 106.6 ;
      RECT  223.4 105.8 224.2 106.6 ;
      RECT  2.6 110.6 3.4 111.4 ;
      RECT  7.4 110.6 8.2 111.4 ;
      RECT  12.2 110.6 13.0 111.4 ;
      RECT  17.0 110.6 17.8 111.4 ;
      RECT  21.8 110.6 22.6 111.4 ;
      RECT  26.6 110.6 27.4 111.4 ;
      RECT  31.4 110.6 32.2 111.4 ;
      RECT  36.2 110.6 37.0 111.4 ;
      RECT  41.0 110.6 41.8 111.4 ;
      RECT  45.8 110.6 46.6 111.4 ;
      RECT  50.6 110.6 51.4 111.4 ;
      RECT  55.4 110.6 56.2 111.4 ;
      RECT  60.2 110.6 61.0 111.4 ;
      RECT  65.0 110.6 65.8 111.4 ;
      RECT  69.8 110.6 70.6 111.4 ;
      RECT  74.6 110.6 75.4 111.4 ;
      RECT  79.4 110.6 80.2 111.4 ;
      RECT  189.8 110.6 190.6 111.4 ;
      RECT  194.6 110.6 195.4 111.4 ;
      RECT  199.4 110.6 200.2 111.4 ;
      RECT  204.2 110.6 205.0 111.4 ;
      RECT  209.0 110.6 209.8 111.4 ;
      RECT  213.8 110.6 214.6 111.4 ;
      RECT  218.6 110.6 219.4 111.4 ;
      RECT  223.4 110.6 224.2 111.4 ;
      RECT  2.6 115.4 3.4 116.2 ;
      RECT  7.4 115.4 8.2 116.2 ;
      RECT  12.2 115.4 13.0 116.2 ;
      RECT  17.0 115.4 17.8 116.2 ;
      RECT  21.8 115.4 22.6 116.2 ;
      RECT  26.6 115.4 27.4 116.2 ;
      RECT  31.4 115.4 32.2 116.2 ;
      RECT  36.2 115.4 37.0 116.2 ;
      RECT  41.0 115.4 41.8 116.2 ;
      RECT  45.8 115.4 46.6 116.2 ;
      RECT  50.6 115.4 51.4 116.2 ;
      RECT  55.4 115.4 56.2 116.2 ;
      RECT  60.2 115.4 61.0 116.2 ;
      RECT  65.0 115.4 65.8 116.2 ;
      RECT  69.8 115.4 70.6 116.2 ;
      RECT  74.6 115.4 75.4 116.2 ;
      RECT  79.4 115.4 80.2 116.2 ;
      RECT  84.2 115.4 85.0 116.2 ;
      RECT  89.0 115.4 89.8 116.2 ;
      RECT  93.8 115.4 94.6 116.2 ;
      RECT  98.6 115.4 99.4 116.2 ;
      RECT  103.4 115.4 104.2 116.2 ;
      RECT  108.2 115.4 109.0 116.2 ;
      RECT  113.0 115.4 113.8 116.2 ;
      RECT  117.8 115.4 118.6 116.2 ;
      RECT  122.6 115.4 123.4 116.2 ;
      RECT  127.4 115.4 128.2 116.2 ;
      RECT  132.2 115.4 133.0 116.2 ;
      RECT  137.0 115.4 137.8 116.2 ;
      RECT  141.8 115.4 142.6 116.2 ;
      RECT  146.6 115.4 147.4 116.2 ;
      RECT  151.4 115.4 152.2 116.2 ;
      RECT  156.2 115.4 157.0 116.2 ;
      RECT  161.0 115.4 161.8 116.2 ;
      RECT  165.8 115.4 166.6 116.2 ;
      RECT  170.6 115.4 171.4 116.2 ;
      RECT  175.4 115.4 176.2 116.2 ;
      RECT  180.2 115.4 181.0 116.2 ;
      RECT  185.0 115.4 185.8 116.2 ;
      RECT  189.8 115.4 190.6 116.2 ;
      RECT  194.6 115.4 195.4 116.2 ;
      RECT  199.4 115.4 200.2 116.2 ;
      RECT  204.2 115.4 205.0 116.2 ;
      RECT  209.0 115.4 209.8 116.2 ;
      RECT  213.8 115.4 214.6 116.2 ;
      RECT  218.6 115.4 219.4 116.2 ;
      RECT  223.4 115.4 224.2 116.2 ;
      RECT  2.6 120.2 3.4 121.0 ;
      RECT  7.4 120.2 8.2 121.0 ;
      RECT  12.2 120.2 13.0 121.0 ;
      RECT  17.0 120.2 17.8 121.0 ;
      RECT  21.8 120.2 22.6 121.0 ;
      RECT  26.6 120.2 27.4 121.0 ;
      RECT  31.4 120.2 32.2 121.0 ;
      RECT  36.2 120.2 37.0 121.0 ;
      RECT  41.0 120.2 41.8 121.0 ;
      RECT  45.8 120.2 46.6 121.0 ;
      RECT  50.6 120.2 51.4 121.0 ;
      RECT  55.4 120.2 56.2 121.0 ;
      RECT  60.2 120.2 61.0 121.0 ;
      RECT  65.0 120.2 65.8 121.0 ;
      RECT  69.8 120.2 70.6 121.0 ;
      RECT  74.6 120.2 75.4 121.0 ;
      RECT  79.4 120.2 80.2 121.0 ;
      RECT  84.2 120.2 85.0 121.0 ;
      RECT  89.0 120.2 89.8 121.0 ;
      RECT  93.8 120.2 94.6 121.0 ;
      RECT  98.6 120.2 99.4 121.0 ;
      RECT  103.4 120.2 104.2 121.0 ;
      RECT  108.2 120.2 109.0 121.0 ;
      RECT  113.0 120.2 113.8 121.0 ;
      RECT  117.8 120.2 118.6 121.0 ;
      RECT  122.6 120.2 123.4 121.0 ;
      RECT  127.4 120.2 128.2 121.0 ;
      RECT  132.2 120.2 133.0 121.0 ;
      RECT  137.0 120.2 137.8 121.0 ;
      RECT  141.8 120.2 142.6 121.0 ;
      RECT  146.6 120.2 147.4 121.0 ;
      RECT  151.4 120.2 152.2 121.0 ;
      RECT  156.2 120.2 157.0 121.0 ;
      RECT  161.0 120.2 161.8 121.0 ;
      RECT  165.8 120.2 166.6 121.0 ;
      RECT  170.6 120.2 171.4 121.0 ;
      RECT  175.4 120.2 176.2 121.0 ;
      RECT  180.2 120.2 181.0 121.0 ;
      RECT  185.0 120.2 185.8 121.0 ;
      RECT  189.8 120.2 190.6 121.0 ;
      RECT  194.6 120.2 195.4 121.0 ;
      RECT  199.4 120.2 200.2 121.0 ;
      RECT  204.2 120.2 205.0 121.0 ;
      RECT  209.0 120.2 209.8 121.0 ;
      RECT  213.8 120.2 214.6 121.0 ;
      RECT  218.6 120.2 219.4 121.0 ;
      RECT  223.4 120.2 224.2 121.0 ;
      RECT  2.6 125.0 3.4 125.8 ;
      RECT  7.4 125.0 8.2 125.8 ;
      RECT  12.2 125.0 13.0 125.8 ;
      RECT  17.0 125.0 17.8 125.8 ;
      RECT  21.8 125.0 22.6 125.8 ;
      RECT  26.6 125.0 27.4 125.8 ;
      RECT  31.4 125.0 32.2 125.8 ;
      RECT  36.2 125.0 37.0 125.8 ;
      RECT  41.0 125.0 41.8 125.8 ;
      RECT  45.8 125.0 46.6 125.8 ;
      RECT  50.6 125.0 51.4 125.8 ;
      RECT  55.4 125.0 56.2 125.8 ;
      RECT  60.2 125.0 61.0 125.8 ;
      RECT  65.0 125.0 65.8 125.8 ;
      RECT  69.8 125.0 70.6 125.8 ;
      RECT  74.6 125.0 75.4 125.8 ;
      RECT  79.4 125.0 80.2 125.8 ;
      RECT  84.2 125.0 85.0 125.8 ;
      RECT  89.0 125.0 89.8 125.8 ;
      RECT  93.8 125.0 94.6 125.8 ;
      RECT  98.6 125.0 99.4 125.8 ;
      RECT  103.4 125.0 104.2 125.8 ;
      RECT  108.2 125.0 109.0 125.8 ;
      RECT  113.0 125.0 113.8 125.8 ;
      RECT  117.8 125.0 118.6 125.8 ;
      RECT  122.6 125.0 123.4 125.8 ;
      RECT  127.4 125.0 128.2 125.8 ;
      RECT  132.2 125.0 133.0 125.8 ;
      RECT  137.0 125.0 137.8 125.8 ;
      RECT  141.8 125.0 142.6 125.8 ;
      RECT  146.6 125.0 147.4 125.8 ;
      RECT  151.4 125.0 152.2 125.8 ;
      RECT  156.2 125.0 157.0 125.8 ;
      RECT  161.0 125.0 161.8 125.8 ;
      RECT  165.8 125.0 166.6 125.8 ;
      RECT  170.6 125.0 171.4 125.8 ;
      RECT  175.4 125.0 176.2 125.8 ;
      RECT  180.2 125.0 181.0 125.8 ;
      RECT  185.0 125.0 185.8 125.8 ;
      RECT  189.8 125.0 190.6 125.8 ;
      RECT  194.6 125.0 195.4 125.8 ;
      RECT  199.4 125.0 200.2 125.8 ;
      RECT  204.2 125.0 205.0 125.8 ;
      RECT  209.0 125.0 209.8 125.8 ;
      RECT  213.8 125.0 214.6 125.8 ;
      RECT  218.6 125.0 219.4 125.8 ;
      RECT  223.4 125.0 224.2 125.8 ;
      RECT  2.6 129.8 3.4 130.6 ;
      RECT  7.4 129.8 8.2 130.6 ;
      RECT  12.2 129.8 13.0 130.6 ;
      RECT  17.0 129.8 17.8 130.6 ;
      RECT  21.8 129.8 22.6 130.6 ;
      RECT  26.6 129.8 27.4 130.6 ;
      RECT  31.4 129.8 32.2 130.6 ;
      RECT  55.4 129.8 56.2 130.6 ;
      RECT  60.2 129.8 61.0 130.6 ;
      RECT  65.0 129.8 65.8 130.6 ;
      RECT  69.8 129.8 70.6 130.6 ;
      RECT  74.6 129.8 75.4 130.6 ;
      RECT  79.4 129.8 80.2 130.6 ;
      RECT  84.2 129.8 85.0 130.6 ;
      RECT  89.0 129.8 89.8 130.6 ;
      RECT  93.8 129.8 94.6 130.6 ;
      RECT  98.6 129.8 99.4 130.6 ;
      RECT  103.4 129.8 104.2 130.6 ;
      RECT  108.2 129.8 109.0 130.6 ;
      RECT  113.0 129.8 113.8 130.6 ;
      RECT  117.8 129.8 118.6 130.6 ;
      RECT  122.6 129.8 123.4 130.6 ;
      RECT  127.4 129.8 128.2 130.6 ;
      RECT  132.2 129.8 133.0 130.6 ;
      RECT  137.0 129.8 137.8 130.6 ;
      RECT  141.8 129.8 142.6 130.6 ;
      RECT  146.6 129.8 147.4 130.6 ;
      RECT  151.4 129.8 152.2 130.6 ;
      RECT  156.2 129.8 157.0 130.6 ;
      RECT  161.0 129.8 161.8 130.6 ;
      RECT  165.8 129.8 166.6 130.6 ;
      RECT  170.6 129.8 171.4 130.6 ;
      RECT  175.4 129.8 176.2 130.6 ;
      RECT  180.2 129.8 181.0 130.6 ;
      RECT  185.0 129.8 185.8 130.6 ;
      RECT  189.8 129.8 190.6 130.6 ;
      RECT  194.6 129.8 195.4 130.6 ;
      RECT  199.4 129.8 200.2 130.6 ;
      RECT  204.2 129.8 205.0 130.6 ;
      RECT  209.0 129.8 209.8 130.6 ;
      RECT  213.8 129.8 214.6 130.6 ;
      RECT  218.6 129.8 219.4 130.6 ;
      RECT  223.4 129.8 224.2 130.6 ;
      RECT  2.6 134.6 3.4 135.4 ;
      RECT  7.4 134.6 8.2 135.4 ;
      RECT  12.2 134.6 13.0 135.4 ;
      RECT  17.0 134.6 17.8 135.4 ;
      RECT  21.8 134.6 22.6 135.4 ;
      RECT  26.6 134.6 27.4 135.4 ;
      RECT  31.4 134.6 32.2 135.4 ;
      RECT  36.2 134.6 37.0 135.4 ;
      RECT  41.0 134.6 41.8 135.4 ;
      RECT  45.8 134.6 46.6 135.4 ;
      RECT  50.6 134.6 51.4 135.4 ;
      RECT  55.4 134.6 56.2 135.4 ;
      RECT  60.2 134.6 61.0 135.4 ;
      RECT  65.0 134.6 65.8 135.4 ;
      RECT  69.8 134.6 70.6 135.4 ;
      RECT  74.6 134.6 75.4 135.4 ;
      RECT  79.4 134.6 80.2 135.4 ;
      RECT  84.2 134.6 85.0 135.4 ;
      RECT  89.0 134.6 89.8 135.4 ;
      RECT  93.8 134.6 94.6 135.4 ;
      RECT  98.6 134.6 99.4 135.4 ;
      RECT  103.4 134.6 104.2 135.4 ;
      RECT  108.2 134.6 109.0 135.4 ;
      RECT  113.0 134.6 113.8 135.4 ;
      RECT  117.8 134.6 118.6 135.4 ;
      RECT  122.6 134.6 123.4 135.4 ;
      RECT  127.4 134.6 128.2 135.4 ;
      RECT  132.2 134.6 133.0 135.4 ;
      RECT  137.0 134.6 137.8 135.4 ;
      RECT  141.8 134.6 142.6 135.4 ;
      RECT  146.6 134.6 147.4 135.4 ;
      RECT  151.4 134.6 152.2 135.4 ;
      RECT  156.2 134.6 157.0 135.4 ;
      RECT  161.0 134.6 161.8 135.4 ;
      RECT  165.8 134.6 166.6 135.4 ;
      RECT  170.6 134.6 171.4 135.4 ;
      RECT  175.4 134.6 176.2 135.4 ;
      RECT  180.2 134.6 181.0 135.4 ;
      RECT  185.0 134.6 185.8 135.4 ;
      RECT  189.8 134.6 190.6 135.4 ;
      RECT  194.6 134.6 195.4 135.4 ;
      RECT  199.4 134.6 200.2 135.4 ;
      RECT  2.6 139.4 3.4 140.2 ;
      RECT  7.4 139.4 8.2 140.2 ;
      RECT  12.2 139.4 13.0 140.2 ;
      RECT  17.0 139.4 17.8 140.2 ;
      RECT  21.8 139.4 22.6 140.2 ;
      RECT  26.6 139.4 27.4 140.2 ;
      RECT  31.4 139.4 32.2 140.2 ;
      RECT  36.2 139.4 37.0 140.2 ;
      RECT  41.0 139.4 41.8 140.2 ;
      RECT  45.8 139.4 46.6 140.2 ;
      RECT  50.6 139.4 51.4 140.2 ;
      RECT  55.4 139.4 56.2 140.2 ;
      RECT  60.2 139.4 61.0 140.2 ;
      RECT  65.0 139.4 65.8 140.2 ;
      RECT  69.8 139.4 70.6 140.2 ;
      RECT  74.6 139.4 75.4 140.2 ;
      RECT  79.4 139.4 80.2 140.2 ;
      RECT  84.2 139.4 85.0 140.2 ;
      RECT  89.0 139.4 89.8 140.2 ;
      RECT  93.8 139.4 94.6 140.2 ;
      RECT  98.6 139.4 99.4 140.2 ;
      RECT  103.4 139.4 104.2 140.2 ;
      RECT  108.2 139.4 109.0 140.2 ;
      RECT  113.0 139.4 113.8 140.2 ;
      RECT  117.8 139.4 118.6 140.2 ;
      RECT  122.6 139.4 123.4 140.2 ;
      RECT  127.4 139.4 128.2 140.2 ;
      RECT  132.2 139.4 133.0 140.2 ;
      RECT  137.0 139.4 137.8 140.2 ;
      RECT  141.8 139.4 142.6 140.2 ;
      RECT  146.6 139.4 147.4 140.2 ;
      RECT  151.4 139.4 152.2 140.2 ;
      RECT  156.2 139.4 157.0 140.2 ;
      RECT  161.0 139.4 161.8 140.2 ;
      RECT  165.8 139.4 166.6 140.2 ;
      RECT  170.6 139.4 171.4 140.2 ;
      RECT  175.4 139.4 176.2 140.2 ;
      RECT  180.2 139.4 181.0 140.2 ;
      RECT  185.0 139.4 185.8 140.2 ;
      RECT  189.8 139.4 190.6 140.2 ;
      RECT  194.6 139.4 195.4 140.2 ;
      RECT  199.4 139.4 200.2 140.2 ;
      RECT  204.2 139.4 205.0 140.2 ;
      RECT  209.0 139.4 209.8 140.2 ;
      RECT  213.8 139.4 214.6 140.2 ;
      RECT  218.6 139.4 219.4 140.2 ;
      RECT  223.4 139.4 224.2 140.2 ;
      RECT  2.6 144.2 3.4 145.0 ;
      RECT  7.4 144.2 8.2 145.0 ;
      RECT  12.2 144.2 13.0 145.0 ;
      RECT  17.0 144.2 17.8 145.0 ;
      RECT  21.8 144.2 22.6 145.0 ;
      RECT  26.6 144.2 27.4 145.0 ;
      RECT  31.4 144.2 32.2 145.0 ;
      RECT  36.2 144.2 37.0 145.0 ;
      RECT  41.0 144.2 41.8 145.0 ;
      RECT  45.8 144.2 46.6 145.0 ;
      RECT  50.6 144.2 51.4 145.0 ;
      RECT  55.4 144.2 56.2 145.0 ;
      RECT  60.2 144.2 61.0 145.0 ;
      RECT  65.0 144.2 65.8 145.0 ;
      RECT  69.8 144.2 70.6 145.0 ;
      RECT  74.6 144.2 75.4 145.0 ;
      RECT  79.4 144.2 80.2 145.0 ;
      RECT  84.2 144.2 85.0 145.0 ;
      RECT  89.0 144.2 89.8 145.0 ;
      RECT  93.8 144.2 94.6 145.0 ;
      RECT  98.6 144.2 99.4 145.0 ;
      RECT  103.4 144.2 104.2 145.0 ;
      RECT  108.2 144.2 109.0 145.0 ;
      RECT  113.0 144.2 113.8 145.0 ;
      RECT  117.8 144.2 118.6 145.0 ;
      RECT  122.6 144.2 123.4 145.0 ;
      RECT  127.4 144.2 128.2 145.0 ;
      RECT  132.2 144.2 133.0 145.0 ;
      RECT  137.0 144.2 137.8 145.0 ;
      RECT  141.8 144.2 142.6 145.0 ;
      RECT  146.6 144.2 147.4 145.0 ;
      RECT  151.4 144.2 152.2 145.0 ;
      RECT  156.2 144.2 157.0 145.0 ;
      RECT  161.0 144.2 161.8 145.0 ;
      RECT  165.8 144.2 166.6 145.0 ;
      RECT  170.6 144.2 171.4 145.0 ;
      RECT  175.4 144.2 176.2 145.0 ;
      RECT  180.2 144.2 181.0 145.0 ;
      RECT  185.0 144.2 185.8 145.0 ;
      RECT  189.8 144.2 190.6 145.0 ;
      RECT  194.6 144.2 195.4 145.0 ;
      RECT  199.4 144.2 200.2 145.0 ;
      RECT  204.2 144.2 205.0 145.0 ;
      RECT  209.0 144.2 209.8 145.0 ;
      RECT  213.8 144.2 214.6 145.0 ;
      RECT  218.6 144.2 219.4 145.0 ;
      RECT  223.4 144.2 224.2 145.0 ;
      RECT  2.6 149.0 3.4 149.8 ;
      RECT  7.4 149.0 8.2 149.8 ;
      RECT  12.2 149.0 13.0 149.8 ;
      RECT  17.0 149.0 17.8 149.8 ;
      RECT  21.8 149.0 22.6 149.8 ;
      RECT  26.6 149.0 27.4 149.8 ;
      RECT  31.4 149.0 32.2 149.8 ;
      RECT  36.2 149.0 37.0 149.8 ;
      RECT  41.0 149.0 41.8 149.8 ;
      RECT  45.8 149.0 46.6 149.8 ;
      RECT  50.6 149.0 51.4 149.8 ;
      RECT  55.4 149.0 56.2 149.8 ;
      RECT  60.2 149.0 61.0 149.8 ;
      RECT  65.0 149.0 65.8 149.8 ;
      RECT  69.8 149.0 70.6 149.8 ;
      RECT  74.6 149.0 75.4 149.8 ;
      RECT  79.4 149.0 80.2 149.8 ;
      RECT  84.2 149.0 85.0 149.8 ;
      RECT  89.0 149.0 89.8 149.8 ;
      RECT  93.8 149.0 94.6 149.8 ;
      RECT  98.6 149.0 99.4 149.8 ;
      RECT  103.4 149.0 104.2 149.8 ;
      RECT  108.2 149.0 109.0 149.8 ;
      RECT  113.0 149.0 113.8 149.8 ;
      RECT  117.8 149.0 118.6 149.8 ;
      RECT  122.6 149.0 123.4 149.8 ;
      RECT  127.4 149.0 128.2 149.8 ;
      RECT  132.2 149.0 133.0 149.8 ;
      RECT  137.0 149.0 137.8 149.8 ;
      RECT  141.8 149.0 142.6 149.8 ;
      RECT  146.6 149.0 147.4 149.8 ;
      RECT  151.4 149.0 152.2 149.8 ;
      RECT  156.2 149.0 157.0 149.8 ;
      RECT  161.0 149.0 161.8 149.8 ;
      RECT  165.8 149.0 166.6 149.8 ;
      RECT  170.6 149.0 171.4 149.8 ;
      RECT  175.4 149.0 176.2 149.8 ;
      RECT  180.2 149.0 181.0 149.8 ;
      RECT  185.0 149.0 185.8 149.8 ;
      RECT  189.8 149.0 190.6 149.8 ;
      RECT  194.6 149.0 195.4 149.8 ;
      RECT  199.4 149.0 200.2 149.8 ;
      RECT  204.2 149.0 205.0 149.8 ;
      RECT  209.0 149.0 209.8 149.8 ;
      RECT  213.8 149.0 214.6 149.8 ;
      RECT  218.6 149.0 219.4 149.8 ;
      RECT  223.4 149.0 224.2 149.8 ;
      RECT  2.6 153.8 3.4 154.6 ;
      RECT  7.4 153.8 8.2 154.6 ;
      RECT  12.2 153.8 13.0 154.6 ;
      RECT  17.0 153.8 17.8 154.6 ;
      RECT  21.8 153.8 22.6 154.6 ;
      RECT  26.6 153.8 27.4 154.6 ;
      RECT  31.4 153.8 32.2 154.6 ;
      RECT  36.2 153.8 37.0 154.6 ;
      RECT  41.0 153.8 41.8 154.6 ;
      RECT  45.8 153.8 46.6 154.6 ;
      RECT  50.6 153.8 51.4 154.6 ;
      RECT  55.4 153.8 56.2 154.6 ;
      RECT  60.2 153.8 61.0 154.6 ;
      RECT  65.0 153.8 65.8 154.6 ;
      RECT  69.8 153.8 70.6 154.6 ;
      RECT  74.6 153.8 75.4 154.6 ;
      RECT  79.4 153.8 80.2 154.6 ;
      RECT  185.0 153.8 185.8 154.6 ;
      RECT  189.8 153.8 190.6 154.6 ;
      RECT  194.6 153.8 195.4 154.6 ;
      RECT  199.4 153.8 200.2 154.6 ;
      RECT  204.2 153.8 205.0 154.6 ;
      RECT  209.0 153.8 209.8 154.6 ;
      RECT  213.8 153.8 214.6 154.6 ;
      RECT  218.6 153.8 219.4 154.6 ;
      RECT  223.4 153.8 224.2 154.6 ;
      RECT  2.6 158.6 3.4 159.4 ;
      RECT  7.4 158.6 8.2 159.4 ;
      RECT  12.2 158.6 13.0 159.4 ;
      RECT  17.0 158.6 17.8 159.4 ;
      RECT  21.8 158.6 22.6 159.4 ;
      RECT  26.6 158.6 27.4 159.4 ;
      RECT  31.4 158.6 32.2 159.4 ;
      RECT  36.2 158.6 37.0 159.4 ;
      RECT  41.0 158.6 41.8 159.4 ;
      RECT  45.8 158.6 46.6 159.4 ;
      RECT  50.6 158.6 51.4 159.4 ;
      RECT  55.4 158.6 56.2 159.4 ;
      RECT  60.2 158.6 61.0 159.4 ;
      RECT  65.0 158.6 65.8 159.4 ;
      RECT  69.8 158.6 70.6 159.4 ;
      RECT  74.6 158.6 75.4 159.4 ;
      RECT  79.4 158.6 80.2 159.4 ;
      RECT  84.2 158.6 85.0 159.4 ;
      RECT  89.0 158.6 89.8 159.4 ;
      RECT  93.8 158.6 94.6 159.4 ;
      RECT  98.6 158.6 99.4 159.4 ;
      RECT  103.4 158.6 104.2 159.4 ;
      RECT  108.2 158.6 109.0 159.4 ;
      RECT  113.0 158.6 113.8 159.4 ;
      RECT  117.8 158.6 118.6 159.4 ;
      RECT  122.6 158.6 123.4 159.4 ;
      RECT  127.4 158.6 128.2 159.4 ;
      RECT  132.2 158.6 133.0 159.4 ;
      RECT  137.0 158.6 137.8 159.4 ;
      RECT  141.8 158.6 142.6 159.4 ;
      RECT  146.6 158.6 147.4 159.4 ;
      RECT  151.4 158.6 152.2 159.4 ;
      RECT  156.2 158.6 157.0 159.4 ;
      RECT  161.0 158.6 161.8 159.4 ;
      RECT  165.8 158.6 166.6 159.4 ;
      RECT  170.6 158.6 171.4 159.4 ;
      RECT  175.4 158.6 176.2 159.4 ;
      RECT  180.2 158.6 181.0 159.4 ;
      RECT  185.0 158.6 185.8 159.4 ;
      RECT  189.8 158.6 190.6 159.4 ;
      RECT  194.6 158.6 195.4 159.4 ;
      RECT  199.4 158.6 200.2 159.4 ;
      RECT  204.2 158.6 205.0 159.4 ;
      RECT  209.0 158.6 209.8 159.4 ;
      RECT  213.8 158.6 214.6 159.4 ;
      RECT  218.6 158.6 219.4 159.4 ;
      RECT  223.4 158.6 224.2 159.4 ;
      RECT  2.6 163.4 3.4 164.2 ;
      RECT  7.4 163.4 8.2 164.2 ;
      RECT  12.2 163.4 13.0 164.2 ;
      RECT  17.0 163.4 17.8 164.2 ;
      RECT  21.8 163.4 22.6 164.2 ;
      RECT  26.6 163.4 27.4 164.2 ;
      RECT  31.4 163.4 32.2 164.2 ;
      RECT  36.2 163.4 37.0 164.2 ;
      RECT  41.0 163.4 41.8 164.2 ;
      RECT  45.8 163.4 46.6 164.2 ;
      RECT  50.6 163.4 51.4 164.2 ;
      RECT  55.4 163.4 56.2 164.2 ;
      RECT  60.2 163.4 61.0 164.2 ;
      RECT  65.0 163.4 65.8 164.2 ;
      RECT  69.8 163.4 70.6 164.2 ;
      RECT  74.6 163.4 75.4 164.2 ;
      RECT  79.4 163.4 80.2 164.2 ;
      RECT  84.2 163.4 85.0 164.2 ;
      RECT  89.0 163.4 89.8 164.2 ;
      RECT  93.8 163.4 94.6 164.2 ;
      RECT  98.6 163.4 99.4 164.2 ;
      RECT  103.4 163.4 104.2 164.2 ;
      RECT  108.2 163.4 109.0 164.2 ;
      RECT  113.0 163.4 113.8 164.2 ;
      RECT  117.8 163.4 118.6 164.2 ;
      RECT  122.6 163.4 123.4 164.2 ;
      RECT  127.4 163.4 128.2 164.2 ;
      RECT  132.2 163.4 133.0 164.2 ;
      RECT  137.0 163.4 137.8 164.2 ;
      RECT  141.8 163.4 142.6 164.2 ;
      RECT  146.6 163.4 147.4 164.2 ;
      RECT  151.4 163.4 152.2 164.2 ;
      RECT  156.2 163.4 157.0 164.2 ;
      RECT  161.0 163.4 161.8 164.2 ;
      RECT  165.8 163.4 166.6 164.2 ;
      RECT  170.6 163.4 171.4 164.2 ;
      RECT  175.4 163.4 176.2 164.2 ;
      RECT  180.2 163.4 181.0 164.2 ;
      RECT  185.0 163.4 185.8 164.2 ;
      RECT  189.8 163.4 190.6 164.2 ;
      RECT  199.4 168.2 200.2 169.0 ;
      RECT  204.2 168.2 205.0 169.0 ;
      RECT  209.0 168.2 209.8 169.0 ;
      RECT  213.8 168.2 214.6 169.0 ;
      RECT  218.6 168.2 219.4 169.0 ;
      RECT  223.4 168.2 224.2 169.0 ;
      RECT  21.8 173.0 22.6 173.8 ;
      RECT  26.6 173.0 27.4 173.8 ;
      RECT  31.4 173.0 32.2 173.8 ;
      RECT  36.2 173.0 37.0 173.8 ;
      RECT  41.0 173.0 41.8 173.8 ;
      RECT  45.8 173.0 46.6 173.8 ;
      RECT  50.6 173.0 51.4 173.8 ;
      RECT  55.4 173.0 56.2 173.8 ;
      RECT  60.2 173.0 61.0 173.8 ;
      RECT  65.0 173.0 65.8 173.8 ;
      RECT  69.8 173.0 70.6 173.8 ;
      RECT  74.6 173.0 75.4 173.8 ;
      RECT  79.4 173.0 80.2 173.8 ;
      RECT  84.2 173.0 85.0 173.8 ;
      RECT  89.0 173.0 89.8 173.8 ;
      RECT  93.8 173.0 94.6 173.8 ;
      RECT  98.6 173.0 99.4 173.8 ;
      RECT  103.4 173.0 104.2 173.8 ;
      RECT  108.2 173.0 109.0 173.8 ;
      RECT  113.0 173.0 113.8 173.8 ;
      RECT  117.8 173.0 118.6 173.8 ;
      RECT  122.6 173.0 123.4 173.8 ;
      RECT  127.4 173.0 128.2 173.8 ;
      RECT  132.2 173.0 133.0 173.8 ;
      RECT  137.0 173.0 137.8 173.8 ;
      RECT  141.8 173.0 142.6 173.8 ;
      RECT  146.6 173.0 147.4 173.8 ;
      RECT  151.4 173.0 152.2 173.8 ;
      RECT  156.2 173.0 157.0 173.8 ;
      RECT  161.0 173.0 161.8 173.8 ;
      RECT  165.8 173.0 166.6 173.8 ;
      RECT  170.6 173.0 171.4 173.8 ;
      RECT  175.4 173.0 176.2 173.8 ;
      RECT  180.2 173.0 181.0 173.8 ;
      RECT  185.0 173.0 185.8 173.8 ;
      RECT  189.8 173.0 190.6 173.8 ;
      RECT  194.6 173.0 195.4 173.8 ;
      RECT  199.4 173.0 200.2 173.8 ;
      RECT  204.2 173.0 205.0 173.8 ;
      RECT  209.0 173.0 209.8 173.8 ;
      RECT  213.8 173.0 214.6 173.8 ;
      RECT  218.6 173.0 219.4 173.8 ;
      RECT  223.4 173.0 224.2 173.8 ;
      RECT  2.6 177.8 3.4 178.6 ;
      RECT  7.4 177.8 8.2 178.6 ;
      RECT  12.2 177.8 13.0 178.6 ;
      RECT  17.0 177.8 17.8 178.6 ;
      RECT  21.8 177.8 22.6 178.6 ;
      RECT  26.6 177.8 27.4 178.6 ;
      RECT  31.4 177.8 32.2 178.6 ;
      RECT  36.2 177.8 37.0 178.6 ;
      RECT  41.0 177.8 41.8 178.6 ;
      RECT  45.8 177.8 46.6 178.6 ;
      RECT  50.6 177.8 51.4 178.6 ;
      RECT  55.4 177.8 56.2 178.6 ;
      RECT  60.2 177.8 61.0 178.6 ;
      RECT  65.0 177.8 65.8 178.6 ;
      RECT  69.8 177.8 70.6 178.6 ;
      RECT  74.6 177.8 75.4 178.6 ;
      RECT  79.4 177.8 80.2 178.6 ;
      RECT  84.2 177.8 85.0 178.6 ;
      RECT  89.0 177.8 89.8 178.6 ;
      RECT  93.8 177.8 94.6 178.6 ;
      RECT  98.6 177.8 99.4 178.6 ;
      RECT  103.4 177.8 104.2 178.6 ;
      RECT  108.2 177.8 109.0 178.6 ;
      RECT  113.0 177.8 113.8 178.6 ;
      RECT  117.8 177.8 118.6 178.6 ;
      RECT  122.6 177.8 123.4 178.6 ;
      RECT  127.4 177.8 128.2 178.6 ;
      RECT  132.2 177.8 133.0 178.6 ;
      RECT  137.0 177.8 137.8 178.6 ;
      RECT  141.8 177.8 142.6 178.6 ;
      RECT  146.6 177.8 147.4 178.6 ;
      RECT  151.4 177.8 152.2 178.6 ;
      RECT  156.2 177.8 157.0 178.6 ;
      RECT  161.0 177.8 161.8 178.6 ;
      RECT  165.8 177.8 166.6 178.6 ;
      RECT  170.6 177.8 171.4 178.6 ;
      RECT  175.4 177.8 176.2 178.6 ;
      RECT  180.2 177.8 181.0 178.6 ;
      RECT  185.0 177.8 185.8 178.6 ;
      RECT  189.8 177.8 190.6 178.6 ;
      RECT  194.6 177.8 195.4 178.6 ;
      RECT  199.4 177.8 200.2 178.6 ;
      RECT  204.2 177.8 205.0 178.6 ;
      RECT  209.0 177.8 209.8 178.6 ;
      RECT  213.8 177.8 214.6 178.6 ;
      RECT  218.6 177.8 219.4 178.6 ;
      RECT  223.4 177.8 224.2 178.6 ;
      RECT  2.6 182.6 3.4 183.4 ;
      RECT  7.4 182.6 8.2 183.4 ;
      RECT  12.2 182.6 13.0 183.4 ;
      RECT  17.0 182.6 17.8 183.4 ;
      RECT  21.8 182.6 22.6 183.4 ;
      RECT  26.6 182.6 27.4 183.4 ;
      RECT  31.4 182.6 32.2 183.4 ;
      RECT  36.2 182.6 37.0 183.4 ;
      RECT  41.0 182.6 41.8 183.4 ;
      RECT  45.8 182.6 46.6 183.4 ;
      RECT  50.6 182.6 51.4 183.4 ;
      RECT  55.4 182.6 56.2 183.4 ;
      RECT  60.2 182.6 61.0 183.4 ;
      RECT  65.0 182.6 65.8 183.4 ;
      RECT  69.8 182.6 70.6 183.4 ;
      RECT  74.6 182.6 75.4 183.4 ;
      RECT  79.4 182.6 80.2 183.4 ;
      RECT  84.2 182.6 85.0 183.4 ;
      RECT  89.0 182.6 89.8 183.4 ;
      RECT  93.8 182.6 94.6 183.4 ;
      RECT  98.6 182.6 99.4 183.4 ;
      RECT  103.4 182.6 104.2 183.4 ;
      RECT  108.2 182.6 109.0 183.4 ;
      RECT  113.0 182.6 113.8 183.4 ;
      RECT  117.8 182.6 118.6 183.4 ;
      RECT  122.6 182.6 123.4 183.4 ;
      RECT  127.4 182.6 128.2 183.4 ;
      RECT  132.2 182.6 133.0 183.4 ;
      RECT  137.0 182.6 137.8 183.4 ;
      RECT  141.8 182.6 142.6 183.4 ;
      RECT  146.6 182.6 147.4 183.4 ;
      RECT  151.4 182.6 152.2 183.4 ;
      RECT  156.2 182.6 157.0 183.4 ;
      RECT  161.0 182.6 161.8 183.4 ;
      RECT  165.8 182.6 166.6 183.4 ;
      RECT  170.6 182.6 171.4 183.4 ;
      RECT  175.4 182.6 176.2 183.4 ;
      RECT  180.2 182.6 181.0 183.4 ;
      RECT  2.6 187.4 3.4 188.2 ;
      RECT  7.4 187.4 8.2 188.2 ;
      RECT  12.2 187.4 13.0 188.2 ;
      RECT  17.0 187.4 17.8 188.2 ;
      RECT  21.8 187.4 22.6 188.2 ;
      RECT  26.6 187.4 27.4 188.2 ;
      RECT  31.4 187.4 32.2 188.2 ;
      RECT  36.2 187.4 37.0 188.2 ;
      RECT  41.0 187.4 41.8 188.2 ;
      RECT  45.8 187.4 46.6 188.2 ;
      RECT  50.6 187.4 51.4 188.2 ;
      RECT  55.4 187.4 56.2 188.2 ;
      RECT  60.2 187.4 61.0 188.2 ;
      RECT  65.0 187.4 65.8 188.2 ;
      RECT  69.8 187.4 70.6 188.2 ;
      RECT  74.6 187.4 75.4 188.2 ;
      RECT  79.4 187.4 80.2 188.2 ;
      RECT  84.2 187.4 85.0 188.2 ;
      RECT  89.0 187.4 89.8 188.2 ;
      RECT  93.8 187.4 94.6 188.2 ;
      RECT  98.6 187.4 99.4 188.2 ;
      RECT  103.4 187.4 104.2 188.2 ;
      RECT  108.2 187.4 109.0 188.2 ;
      RECT  113.0 187.4 113.8 188.2 ;
      RECT  117.8 187.4 118.6 188.2 ;
      RECT  122.6 187.4 123.4 188.2 ;
      RECT  127.4 187.4 128.2 188.2 ;
      RECT  132.2 187.4 133.0 188.2 ;
      RECT  137.0 187.4 137.8 188.2 ;
      RECT  141.8 187.4 142.6 188.2 ;
      RECT  146.6 187.4 147.4 188.2 ;
      RECT  151.4 187.4 152.2 188.2 ;
      RECT  156.2 187.4 157.0 188.2 ;
      RECT  161.0 187.4 161.8 188.2 ;
      RECT  165.8 187.4 166.6 188.2 ;
      RECT  170.6 187.4 171.4 188.2 ;
      RECT  175.4 187.4 176.2 188.2 ;
      RECT  180.2 187.4 181.0 188.2 ;
      RECT  185.0 187.4 185.8 188.2 ;
      RECT  189.8 187.4 190.6 188.2 ;
      RECT  194.6 187.4 195.4 188.2 ;
      RECT  199.4 187.4 200.2 188.2 ;
      RECT  204.2 187.4 205.0 188.2 ;
      RECT  209.0 187.4 209.8 188.2 ;
      RECT  213.8 187.4 214.6 188.2 ;
      RECT  218.6 187.4 219.4 188.2 ;
      RECT  223.4 187.4 224.2 188.2 ;
      RECT  36.2 192.2 37.0 193.0 ;
      RECT  41.0 192.2 41.8 193.0 ;
      RECT  45.8 192.2 46.6 193.0 ;
      RECT  50.6 192.2 51.4 193.0 ;
      RECT  55.4 192.2 56.2 193.0 ;
      RECT  60.2 192.2 61.0 193.0 ;
      RECT  65.0 192.2 65.8 193.0 ;
      RECT  69.8 192.2 70.6 193.0 ;
      RECT  74.6 192.2 75.4 193.0 ;
      RECT  79.4 192.2 80.2 193.0 ;
      RECT  84.2 192.2 85.0 193.0 ;
      RECT  89.0 192.2 89.8 193.0 ;
      RECT  93.8 192.2 94.6 193.0 ;
      RECT  98.6 192.2 99.4 193.0 ;
      RECT  103.4 192.2 104.2 193.0 ;
      RECT  108.2 192.2 109.0 193.0 ;
      RECT  113.0 192.2 113.8 193.0 ;
      RECT  117.8 192.2 118.6 193.0 ;
      RECT  122.6 192.2 123.4 193.0 ;
      RECT  127.4 192.2 128.2 193.0 ;
      RECT  132.2 192.2 133.0 193.0 ;
      RECT  137.0 192.2 137.8 193.0 ;
      RECT  141.8 192.2 142.6 193.0 ;
      RECT  146.6 192.2 147.4 193.0 ;
      RECT  151.4 192.2 152.2 193.0 ;
      RECT  156.2 192.2 157.0 193.0 ;
      RECT  161.0 192.2 161.8 193.0 ;
      RECT  165.8 192.2 166.6 193.0 ;
      RECT  170.6 192.2 171.4 193.0 ;
      RECT  175.4 192.2 176.2 193.0 ;
      RECT  180.2 192.2 181.0 193.0 ;
      RECT  185.0 192.2 185.8 193.0 ;
      RECT  189.8 192.2 190.6 193.0 ;
      RECT  194.6 192.2 195.4 193.0 ;
      RECT  199.4 192.2 200.2 193.0 ;
      RECT  204.2 192.2 205.0 193.0 ;
      RECT  209.0 192.2 209.8 193.0 ;
      RECT  213.8 192.2 214.6 193.0 ;
      RECT  218.6 192.2 219.4 193.0 ;
      RECT  223.4 192.2 224.2 193.0 ;
      RECT  26.6 197.0 27.4 197.8 ;
      RECT  31.4 197.0 32.2 197.8 ;
      RECT  36.2 197.0 37.0 197.8 ;
      RECT  41.0 197.0 41.8 197.8 ;
      RECT  45.8 197.0 46.6 197.8 ;
      RECT  50.6 197.0 51.4 197.8 ;
      RECT  55.4 197.0 56.2 197.8 ;
      RECT  60.2 197.0 61.0 197.8 ;
      RECT  65.0 197.0 65.8 197.8 ;
      RECT  69.8 197.0 70.6 197.8 ;
      RECT  74.6 197.0 75.4 197.8 ;
      RECT  79.4 197.0 80.2 197.8 ;
      RECT  84.2 197.0 85.0 197.8 ;
      RECT  89.0 197.0 89.8 197.8 ;
      RECT  93.8 197.0 94.6 197.8 ;
      RECT  98.6 197.0 99.4 197.8 ;
      RECT  103.4 197.0 104.2 197.8 ;
      RECT  108.2 197.0 109.0 197.8 ;
      RECT  113.0 197.0 113.8 197.8 ;
      RECT  117.8 197.0 118.6 197.8 ;
      RECT  122.6 197.0 123.4 197.8 ;
      RECT  127.4 197.0 128.2 197.8 ;
      RECT  132.2 197.0 133.0 197.8 ;
      RECT  137.0 197.0 137.8 197.8 ;
      RECT  141.8 197.0 142.6 197.8 ;
      RECT  146.6 197.0 147.4 197.8 ;
      RECT  151.4 197.0 152.2 197.8 ;
      RECT  156.2 197.0 157.0 197.8 ;
      RECT  161.0 197.0 161.8 197.8 ;
      RECT  165.8 197.0 166.6 197.8 ;
      RECT  170.6 197.0 171.4 197.8 ;
      RECT  175.4 197.0 176.2 197.8 ;
      RECT  180.2 197.0 181.0 197.8 ;
      RECT  185.0 197.0 185.8 197.8 ;
      RECT  189.8 197.0 190.6 197.8 ;
      RECT  194.6 197.0 195.4 197.8 ;
      RECT  199.4 197.0 200.2 197.8 ;
      RECT  204.2 197.0 205.0 197.8 ;
      RECT  209.0 197.0 209.8 197.8 ;
      RECT  213.8 197.0 214.6 197.8 ;
      RECT  218.6 197.0 219.4 197.8 ;
      RECT  223.4 197.0 224.2 197.8 ;
      RECT  36.2 201.8 37.0 202.6 ;
      RECT  41.0 201.8 41.8 202.6 ;
      RECT  45.8 201.8 46.6 202.6 ;
      RECT  50.6 201.8 51.4 202.6 ;
      RECT  55.4 201.8 56.2 202.6 ;
      RECT  60.2 201.8 61.0 202.6 ;
      RECT  65.0 201.8 65.8 202.6 ;
      RECT  69.8 201.8 70.6 202.6 ;
      RECT  74.6 201.8 75.4 202.6 ;
      RECT  79.4 201.8 80.2 202.6 ;
      RECT  84.2 201.8 85.0 202.6 ;
      RECT  89.0 201.8 89.8 202.6 ;
      RECT  93.8 201.8 94.6 202.6 ;
      RECT  98.6 201.8 99.4 202.6 ;
      RECT  103.4 201.8 104.2 202.6 ;
      RECT  108.2 201.8 109.0 202.6 ;
      RECT  113.0 201.8 113.8 202.6 ;
      RECT  117.8 201.8 118.6 202.6 ;
      RECT  122.6 201.8 123.4 202.6 ;
      RECT  127.4 201.8 128.2 202.6 ;
      RECT  132.2 201.8 133.0 202.6 ;
      RECT  137.0 201.8 137.8 202.6 ;
      RECT  141.8 201.8 142.6 202.6 ;
      RECT  146.6 201.8 147.4 202.6 ;
      RECT  151.4 201.8 152.2 202.6 ;
      RECT  156.2 201.8 157.0 202.6 ;
      RECT  161.0 201.8 161.8 202.6 ;
      RECT  165.8 201.8 166.6 202.6 ;
      RECT  170.6 201.8 171.4 202.6 ;
      RECT  175.4 201.8 176.2 202.6 ;
      RECT  180.2 201.8 181.0 202.6 ;
      RECT  185.0 201.8 185.8 202.6 ;
      RECT  189.8 201.8 190.6 202.6 ;
      RECT  194.6 201.8 195.4 202.6 ;
      RECT  199.4 201.8 200.2 202.6 ;
      RECT  204.2 201.8 205.0 202.6 ;
      RECT  209.0 201.8 209.8 202.6 ;
      RECT  213.8 201.8 214.6 202.6 ;
      RECT  218.6 201.8 219.4 202.6 ;
      RECT  223.4 201.8 224.2 202.6 ;
      RECT  2.6 206.6 3.4 207.4 ;
      RECT  7.4 206.6 8.2 207.4 ;
      RECT  12.2 206.6 13.0 207.4 ;
      RECT  17.0 206.6 17.8 207.4 ;
      RECT  21.8 206.6 22.6 207.4 ;
      RECT  26.6 206.6 27.4 207.4 ;
      RECT  31.4 206.6 32.2 207.4 ;
      RECT  36.2 206.6 37.0 207.4 ;
      RECT  41.0 206.6 41.8 207.4 ;
      RECT  45.8 206.6 46.6 207.4 ;
      RECT  50.6 206.6 51.4 207.4 ;
      RECT  55.4 206.6 56.2 207.4 ;
      RECT  60.2 206.6 61.0 207.4 ;
      RECT  65.0 206.6 65.8 207.4 ;
      RECT  69.8 206.6 70.6 207.4 ;
      RECT  74.6 206.6 75.4 207.4 ;
      RECT  79.4 206.6 80.2 207.4 ;
      RECT  84.2 206.6 85.0 207.4 ;
      RECT  180.2 206.6 181.0 207.4 ;
      RECT  185.0 206.6 185.8 207.4 ;
      RECT  189.8 206.6 190.6 207.4 ;
      RECT  194.6 206.6 195.4 207.4 ;
      RECT  199.4 206.6 200.2 207.4 ;
      RECT  204.2 206.6 205.0 207.4 ;
      RECT  209.0 206.6 209.8 207.4 ;
      RECT  213.8 206.6 214.6 207.4 ;
      RECT  218.6 206.6 219.4 207.4 ;
      RECT  223.4 206.6 224.2 207.4 ;
      RECT  36.2 211.4 37.0 212.2 ;
      RECT  41.0 211.4 41.8 212.2 ;
      RECT  45.8 211.4 46.6 212.2 ;
      RECT  50.6 211.4 51.4 212.2 ;
      RECT  55.4 211.4 56.2 212.2 ;
      RECT  60.2 211.4 61.0 212.2 ;
      RECT  65.0 211.4 65.8 212.2 ;
      RECT  69.8 211.4 70.6 212.2 ;
      RECT  74.6 211.4 75.4 212.2 ;
      RECT  79.4 211.4 80.2 212.2 ;
      RECT  84.2 211.4 85.0 212.2 ;
      RECT  89.0 211.4 89.8 212.2 ;
      RECT  93.8 211.4 94.6 212.2 ;
      RECT  98.6 211.4 99.4 212.2 ;
      RECT  103.4 211.4 104.2 212.2 ;
      RECT  108.2 211.4 109.0 212.2 ;
      RECT  113.0 211.4 113.8 212.2 ;
      RECT  117.8 211.4 118.6 212.2 ;
      RECT  122.6 211.4 123.4 212.2 ;
      RECT  127.4 211.4 128.2 212.2 ;
      RECT  132.2 211.4 133.0 212.2 ;
      RECT  137.0 211.4 137.8 212.2 ;
      RECT  141.8 211.4 142.6 212.2 ;
      RECT  146.6 211.4 147.4 212.2 ;
      RECT  151.4 211.4 152.2 212.2 ;
      RECT  156.2 211.4 157.0 212.2 ;
      RECT  161.0 211.4 161.8 212.2 ;
      RECT  165.8 211.4 166.6 212.2 ;
      RECT  170.6 211.4 171.4 212.2 ;
      RECT  175.4 211.4 176.2 212.2 ;
      RECT  180.2 211.4 181.0 212.2 ;
      RECT  185.0 211.4 185.8 212.2 ;
      RECT  189.8 211.4 190.6 212.2 ;
      RECT  194.6 211.4 195.4 212.2 ;
      RECT  199.4 211.4 200.2 212.2 ;
      RECT  204.2 211.4 205.0 212.2 ;
      RECT  209.0 211.4 209.8 212.2 ;
      RECT  213.8 211.4 214.6 212.2 ;
      RECT  218.6 211.4 219.4 212.2 ;
      RECT  223.4 211.4 224.2 212.2 ;
      RECT  26.6 216.2 27.4 217.0 ;
      RECT  31.4 216.2 32.2 217.0 ;
      RECT  36.2 216.2 37.0 217.0 ;
      RECT  41.0 216.2 41.8 217.0 ;
      RECT  45.8 216.2 46.6 217.0 ;
      RECT  50.6 216.2 51.4 217.0 ;
      RECT  55.4 216.2 56.2 217.0 ;
      RECT  60.2 216.2 61.0 217.0 ;
      RECT  65.0 216.2 65.8 217.0 ;
      RECT  69.8 216.2 70.6 217.0 ;
      RECT  74.6 216.2 75.4 217.0 ;
      RECT  79.4 216.2 80.2 217.0 ;
      RECT  84.2 216.2 85.0 217.0 ;
      RECT  137.0 216.2 137.8 217.0 ;
      RECT  141.8 216.2 142.6 217.0 ;
      RECT  146.6 216.2 147.4 217.0 ;
      RECT  151.4 216.2 152.2 217.0 ;
      RECT  156.2 216.2 157.0 217.0 ;
      RECT  161.0 216.2 161.8 217.0 ;
      RECT  165.8 216.2 166.6 217.0 ;
      RECT  170.6 216.2 171.4 217.0 ;
      RECT  175.4 216.2 176.2 217.0 ;
      RECT  180.2 216.2 181.0 217.0 ;
      RECT  185.0 216.2 185.8 217.0 ;
      RECT  189.8 216.2 190.6 217.0 ;
      RECT  194.6 216.2 195.4 217.0 ;
      RECT  199.4 216.2 200.2 217.0 ;
      RECT  204.2 216.2 205.0 217.0 ;
      RECT  209.0 216.2 209.8 217.0 ;
      RECT  213.8 216.2 214.6 217.0 ;
      RECT  218.6 216.2 219.4 217.0 ;
      RECT  223.4 216.2 224.2 217.0 ;
      RECT  36.2 221.0 37.0 221.8 ;
      RECT  41.0 221.0 41.8 221.8 ;
      RECT  45.8 221.0 46.6 221.8 ;
      RECT  50.6 221.0 51.4 221.8 ;
      RECT  55.4 221.0 56.2 221.8 ;
      RECT  60.2 221.0 61.0 221.8 ;
      RECT  65.0 221.0 65.8 221.8 ;
      RECT  69.8 221.0 70.6 221.8 ;
      RECT  74.6 221.0 75.4 221.8 ;
      RECT  79.4 221.0 80.2 221.8 ;
      RECT  84.2 221.0 85.0 221.8 ;
      RECT  89.0 221.0 89.8 221.8 ;
      RECT  93.8 221.0 94.6 221.8 ;
      RECT  98.6 221.0 99.4 221.8 ;
      RECT  103.4 221.0 104.2 221.8 ;
      RECT  108.2 221.0 109.0 221.8 ;
      RECT  113.0 221.0 113.8 221.8 ;
      RECT  117.8 221.0 118.6 221.8 ;
      RECT  122.6 221.0 123.4 221.8 ;
      RECT  127.4 221.0 128.2 221.8 ;
      RECT  132.2 221.0 133.0 221.8 ;
      RECT  137.0 221.0 137.8 221.8 ;
      RECT  141.8 221.0 142.6 221.8 ;
      RECT  146.6 221.0 147.4 221.8 ;
      RECT  151.4 221.0 152.2 221.8 ;
      RECT  156.2 221.0 157.0 221.8 ;
      RECT  161.0 221.0 161.8 221.8 ;
      RECT  165.8 221.0 166.6 221.8 ;
      RECT  170.6 221.0 171.4 221.8 ;
      RECT  175.4 221.0 176.2 221.8 ;
      RECT  180.2 221.0 181.0 221.8 ;
      RECT  185.0 221.0 185.8 221.8 ;
      RECT  189.8 221.0 190.6 221.8 ;
      RECT  194.6 221.0 195.4 221.8 ;
      RECT  199.4 221.0 200.2 221.8 ;
      RECT  204.2 221.0 205.0 221.8 ;
      RECT  209.0 221.0 209.8 221.8 ;
      RECT  213.8 221.0 214.6 221.8 ;
      RECT  218.6 221.0 219.4 221.8 ;
      RECT  223.4 221.0 224.2 221.8 ;
      RECT  2.6 225.8 3.4 226.6 ;
      RECT  7.4 225.8 8.2 226.6 ;
      RECT  12.2 225.8 13.0 226.6 ;
      RECT  17.0 225.8 17.8 226.6 ;
      RECT  21.8 225.8 22.6 226.6 ;
      RECT  26.6 225.8 27.4 226.6 ;
      RECT  31.4 225.8 32.2 226.6 ;
      RECT  36.2 225.8 37.0 226.6 ;
      RECT  41.0 225.8 41.8 226.6 ;
      RECT  45.8 225.8 46.6 226.6 ;
      RECT  50.6 225.8 51.4 226.6 ;
      RECT  55.4 225.8 56.2 226.6 ;
      RECT  60.2 225.8 61.0 226.6 ;
      RECT  65.0 225.8 65.8 226.6 ;
      RECT  69.8 225.8 70.6 226.6 ;
      RECT  74.6 225.8 75.4 226.6 ;
      RECT  79.4 225.8 80.2 226.6 ;
      RECT  84.2 225.8 85.0 226.6 ;
      RECT  89.0 225.8 89.8 226.6 ;
      RECT  93.8 225.8 94.6 226.6 ;
      RECT  98.6 225.8 99.4 226.6 ;
      RECT  36.2 230.6 37.0 231.4 ;
      RECT  41.0 230.6 41.8 231.4 ;
      RECT  45.8 230.6 46.6 231.4 ;
      RECT  50.6 230.6 51.4 231.4 ;
      RECT  55.4 230.6 56.2 231.4 ;
      RECT  60.2 230.6 61.0 231.4 ;
      RECT  65.0 230.6 65.8 231.4 ;
      RECT  69.8 230.6 70.6 231.4 ;
      RECT  74.6 230.6 75.4 231.4 ;
      RECT  79.4 230.6 80.2 231.4 ;
      RECT  84.2 230.6 85.0 231.4 ;
      RECT  89.0 230.6 89.8 231.4 ;
      RECT  93.8 230.6 94.6 231.4 ;
      RECT  98.6 230.6 99.4 231.4 ;
      RECT  103.4 230.6 104.2 231.4 ;
      RECT  108.2 230.6 109.0 231.4 ;
      RECT  113.0 230.6 113.8 231.4 ;
      RECT  117.8 230.6 118.6 231.4 ;
      RECT  122.6 230.6 123.4 231.4 ;
      RECT  127.4 230.6 128.2 231.4 ;
      RECT  132.2 230.6 133.0 231.4 ;
      RECT  137.0 230.6 137.8 231.4 ;
      RECT  141.8 230.6 142.6 231.4 ;
      RECT  146.6 230.6 147.4 231.4 ;
      RECT  151.4 230.6 152.2 231.4 ;
      RECT  156.2 230.6 157.0 231.4 ;
      RECT  161.0 230.6 161.8 231.4 ;
      RECT  165.8 230.6 166.6 231.4 ;
      RECT  170.6 230.6 171.4 231.4 ;
      RECT  175.4 230.6 176.2 231.4 ;
      RECT  180.2 230.6 181.0 231.4 ;
      RECT  185.0 230.6 185.8 231.4 ;
      RECT  189.8 230.6 190.6 231.4 ;
      RECT  194.6 230.6 195.4 231.4 ;
      RECT  199.4 230.6 200.2 231.4 ;
      RECT  204.2 230.6 205.0 231.4 ;
      RECT  209.0 230.6 209.8 231.4 ;
      RECT  213.8 230.6 214.6 231.4 ;
      RECT  218.6 230.6 219.4 231.4 ;
      RECT  223.4 230.6 224.2 231.4 ;
      RECT  21.8 235.4 22.6 236.2 ;
      RECT  26.6 235.4 27.4 236.2 ;
      RECT  31.4 235.4 32.2 236.2 ;
      RECT  36.2 235.4 37.0 236.2 ;
      RECT  41.0 235.4 41.8 236.2 ;
      RECT  45.8 235.4 46.6 236.2 ;
      RECT  50.6 235.4 51.4 236.2 ;
      RECT  55.4 235.4 56.2 236.2 ;
      RECT  60.2 235.4 61.0 236.2 ;
      RECT  65.0 235.4 65.8 236.2 ;
      RECT  69.8 235.4 70.6 236.2 ;
      RECT  74.6 235.4 75.4 236.2 ;
      RECT  79.4 235.4 80.2 236.2 ;
      RECT  84.2 235.4 85.0 236.2 ;
      RECT  89.0 235.4 89.8 236.2 ;
      RECT  93.8 235.4 94.6 236.2 ;
      RECT  98.6 235.4 99.4 236.2 ;
      RECT  103.4 235.4 104.2 236.2 ;
      RECT  108.2 235.4 109.0 236.2 ;
      RECT  113.0 235.4 113.8 236.2 ;
      RECT  117.8 235.4 118.6 236.2 ;
      RECT  141.8 235.4 142.6 236.2 ;
      RECT  146.6 235.4 147.4 236.2 ;
      RECT  151.4 235.4 152.2 236.2 ;
      RECT  156.2 235.4 157.0 236.2 ;
      RECT  161.0 235.4 161.8 236.2 ;
      RECT  165.8 235.4 166.6 236.2 ;
      RECT  170.6 235.4 171.4 236.2 ;
      RECT  175.4 235.4 176.2 236.2 ;
      RECT  180.2 235.4 181.0 236.2 ;
      RECT  185.0 235.4 185.8 236.2 ;
      RECT  189.8 235.4 190.6 236.2 ;
      RECT  194.6 235.4 195.4 236.2 ;
      RECT  199.4 235.4 200.2 236.2 ;
      RECT  204.2 235.4 205.0 236.2 ;
      RECT  209.0 235.4 209.8 236.2 ;
      RECT  213.8 235.4 214.6 236.2 ;
      RECT  218.6 235.4 219.4 236.2 ;
      RECT  223.4 235.4 224.2 236.2 ;
      RECT  2.6 240.2 3.4 241.0 ;
      RECT  7.4 240.2 8.2 241.0 ;
      RECT  12.2 240.2 13.0 241.0 ;
      RECT  17.0 240.2 17.8 241.0 ;
      RECT  21.8 240.2 22.6 241.0 ;
      RECT  26.6 240.2 27.4 241.0 ;
      RECT  31.4 240.2 32.2 241.0 ;
      RECT  36.2 240.2 37.0 241.0 ;
      RECT  41.0 240.2 41.8 241.0 ;
      RECT  45.8 240.2 46.6 241.0 ;
      RECT  50.6 240.2 51.4 241.0 ;
      RECT  55.4 240.2 56.2 241.0 ;
      RECT  60.2 240.2 61.0 241.0 ;
      RECT  65.0 240.2 65.8 241.0 ;
      RECT  69.8 240.2 70.6 241.0 ;
      RECT  74.6 240.2 75.4 241.0 ;
      RECT  79.4 240.2 80.2 241.0 ;
      RECT  84.2 240.2 85.0 241.0 ;
      RECT  89.0 240.2 89.8 241.0 ;
      RECT  93.8 240.2 94.6 241.0 ;
      RECT  98.6 240.2 99.4 241.0 ;
      RECT  103.4 240.2 104.2 241.0 ;
      RECT  108.2 240.2 109.0 241.0 ;
      RECT  113.0 240.2 113.8 241.0 ;
      RECT  117.8 240.2 118.6 241.0 ;
      RECT  122.6 240.2 123.4 241.0 ;
      RECT  127.4 240.2 128.2 241.0 ;
      RECT  132.2 240.2 133.0 241.0 ;
      RECT  137.0 240.2 137.8 241.0 ;
      RECT  141.8 240.2 142.6 241.0 ;
      RECT  146.6 240.2 147.4 241.0 ;
      RECT  151.4 240.2 152.2 241.0 ;
      RECT  156.2 240.2 157.0 241.0 ;
      RECT  161.0 240.2 161.8 241.0 ;
      RECT  165.8 240.2 166.6 241.0 ;
      RECT  170.6 240.2 171.4 241.0 ;
      RECT  175.4 240.2 176.2 241.0 ;
      RECT  180.2 240.2 181.0 241.0 ;
      RECT  185.0 240.2 185.8 241.0 ;
      RECT  189.8 240.2 190.6 241.0 ;
      RECT  194.6 240.2 195.4 241.0 ;
      RECT  199.4 240.2 200.2 241.0 ;
      RECT  204.2 240.2 205.0 241.0 ;
      RECT  209.0 240.2 209.8 241.0 ;
      RECT  213.8 240.2 214.6 241.0 ;
      RECT  218.6 240.2 219.4 241.0 ;
      RECT  223.4 240.2 224.2 241.0 ;
      RECT  2.6 245.0 3.4 245.8 ;
      RECT  7.4 245.0 8.2 245.8 ;
      RECT  12.2 245.0 13.0 245.8 ;
      RECT  17.0 245.0 17.8 245.8 ;
      RECT  21.8 245.0 22.6 245.8 ;
      RECT  26.6 245.0 27.4 245.8 ;
      RECT  31.4 245.0 32.2 245.8 ;
      RECT  36.2 245.0 37.0 245.8 ;
      RECT  41.0 245.0 41.8 245.8 ;
      RECT  45.8 245.0 46.6 245.8 ;
      RECT  50.6 245.0 51.4 245.8 ;
      RECT  55.4 245.0 56.2 245.8 ;
      RECT  60.2 245.0 61.0 245.8 ;
      RECT  65.0 245.0 65.8 245.8 ;
      RECT  69.8 245.0 70.6 245.8 ;
      RECT  74.6 245.0 75.4 245.8 ;
      RECT  79.4 245.0 80.2 245.8 ;
      RECT  84.2 245.0 85.0 245.8 ;
      RECT  89.0 245.0 89.8 245.8 ;
      RECT  93.8 245.0 94.6 245.8 ;
      RECT  98.6 245.0 99.4 245.8 ;
      RECT  2.6 249.8 3.4 250.6 ;
      RECT  7.4 249.8 8.2 250.6 ;
      RECT  12.2 249.8 13.0 250.6 ;
      RECT  17.0 249.8 17.8 250.6 ;
      RECT  21.8 249.8 22.6 250.6 ;
      RECT  26.6 249.8 27.4 250.6 ;
      RECT  31.4 249.8 32.2 250.6 ;
      RECT  36.2 249.8 37.0 250.6 ;
      RECT  41.0 249.8 41.8 250.6 ;
      RECT  45.8 249.8 46.6 250.6 ;
      RECT  50.6 249.8 51.4 250.6 ;
      RECT  55.4 249.8 56.2 250.6 ;
      RECT  60.2 249.8 61.0 250.6 ;
      RECT  65.0 249.8 65.8 250.6 ;
      RECT  69.8 249.8 70.6 250.6 ;
      RECT  74.6 249.8 75.4 250.6 ;
      RECT  79.4 249.8 80.2 250.6 ;
      RECT  84.2 249.8 85.0 250.6 ;
      RECT  89.0 249.8 89.8 250.6 ;
      RECT  93.8 249.8 94.6 250.6 ;
      RECT  98.6 249.8 99.4 250.6 ;
      RECT  103.4 249.8 104.2 250.6 ;
      RECT  108.2 249.8 109.0 250.6 ;
      RECT  113.0 249.8 113.8 250.6 ;
      RECT  117.8 249.8 118.6 250.6 ;
      RECT  122.6 249.8 123.4 250.6 ;
      RECT  127.4 249.8 128.2 250.6 ;
      RECT  132.2 249.8 133.0 250.6 ;
      RECT  137.0 249.8 137.8 250.6 ;
      RECT  141.8 249.8 142.6 250.6 ;
      RECT  146.6 249.8 147.4 250.6 ;
      RECT  151.4 249.8 152.2 250.6 ;
      RECT  156.2 249.8 157.0 250.6 ;
      RECT  161.0 249.8 161.8 250.6 ;
      RECT  165.8 249.8 166.6 250.6 ;
      RECT  170.6 249.8 171.4 250.6 ;
      RECT  175.4 249.8 176.2 250.6 ;
      RECT  180.2 249.8 181.0 250.6 ;
      RECT  185.0 249.8 185.8 250.6 ;
      RECT  189.8 249.8 190.6 250.6 ;
      RECT  194.6 249.8 195.4 250.6 ;
      RECT  199.4 249.8 200.2 250.6 ;
      RECT  204.2 249.8 205.0 250.6 ;
      RECT  209.0 249.8 209.8 250.6 ;
      RECT  213.8 249.8 214.6 250.6 ;
      RECT  218.6 249.8 219.4 250.6 ;
      RECT  223.4 249.8 224.2 250.6 ;
      RECT  36.2 254.6 37.0 255.4 ;
      RECT  41.0 254.6 41.8 255.4 ;
      RECT  45.8 254.6 46.6 255.4 ;
      RECT  50.6 254.6 51.4 255.4 ;
      RECT  55.4 254.6 56.2 255.4 ;
      RECT  60.2 254.6 61.0 255.4 ;
      RECT  65.0 254.6 65.8 255.4 ;
      RECT  69.8 254.6 70.6 255.4 ;
      RECT  74.6 254.6 75.4 255.4 ;
      RECT  79.4 254.6 80.2 255.4 ;
      RECT  84.2 254.6 85.0 255.4 ;
      RECT  89.0 254.6 89.8 255.4 ;
      RECT  93.8 254.6 94.6 255.4 ;
      RECT  98.6 254.6 99.4 255.4 ;
      RECT  103.4 254.6 104.2 255.4 ;
      RECT  108.2 254.6 109.0 255.4 ;
      RECT  113.0 254.6 113.8 255.4 ;
      RECT  117.8 254.6 118.6 255.4 ;
      RECT  122.6 254.6 123.4 255.4 ;
      RECT  127.4 254.6 128.2 255.4 ;
      RECT  132.2 254.6 133.0 255.4 ;
      RECT  137.0 254.6 137.8 255.4 ;
      RECT  141.8 254.6 142.6 255.4 ;
      RECT  146.6 254.6 147.4 255.4 ;
      RECT  151.4 254.6 152.2 255.4 ;
      RECT  156.2 254.6 157.0 255.4 ;
      RECT  161.0 254.6 161.8 255.4 ;
      RECT  165.8 254.6 166.6 255.4 ;
      RECT  170.6 254.6 171.4 255.4 ;
      RECT  175.4 254.6 176.2 255.4 ;
      RECT  180.2 254.6 181.0 255.4 ;
      RECT  185.0 254.6 185.8 255.4 ;
      RECT  189.8 254.6 190.6 255.4 ;
      RECT  194.6 254.6 195.4 255.4 ;
      RECT  199.4 254.6 200.2 255.4 ;
      RECT  204.2 254.6 205.0 255.4 ;
      RECT  209.0 254.6 209.8 255.4 ;
      RECT  213.8 254.6 214.6 255.4 ;
      RECT  218.6 254.6 219.4 255.4 ;
      RECT  223.4 254.6 224.2 255.4 ;
      RECT  26.6 259.4 27.4 260.2 ;
      RECT  31.4 259.4 32.2 260.2 ;
      RECT  36.2 259.4 37.0 260.2 ;
      RECT  41.0 259.4 41.8 260.2 ;
      RECT  45.8 259.4 46.6 260.2 ;
      RECT  50.6 259.4 51.4 260.2 ;
      RECT  55.4 259.4 56.2 260.2 ;
      RECT  60.2 259.4 61.0 260.2 ;
      RECT  65.0 259.4 65.8 260.2 ;
      RECT  69.8 259.4 70.6 260.2 ;
      RECT  74.6 259.4 75.4 260.2 ;
      RECT  79.4 259.4 80.2 260.2 ;
      RECT  84.2 259.4 85.0 260.2 ;
      RECT  89.0 259.4 89.8 260.2 ;
      RECT  103.4 259.4 104.2 260.2 ;
      RECT  108.2 259.4 109.0 260.2 ;
      RECT  113.0 259.4 113.8 260.2 ;
      RECT  117.8 259.4 118.6 260.2 ;
      RECT  122.6 259.4 123.4 260.2 ;
      RECT  127.4 259.4 128.2 260.2 ;
      RECT  132.2 259.4 133.0 260.2 ;
      RECT  137.0 259.4 137.8 260.2 ;
      RECT  141.8 259.4 142.6 260.2 ;
      RECT  146.6 259.4 147.4 260.2 ;
      RECT  151.4 259.4 152.2 260.2 ;
      RECT  156.2 259.4 157.0 260.2 ;
      RECT  161.0 259.4 161.8 260.2 ;
      RECT  165.8 259.4 166.6 260.2 ;
      RECT  170.6 259.4 171.4 260.2 ;
      RECT  175.4 259.4 176.2 260.2 ;
      RECT  180.2 259.4 181.0 260.2 ;
      RECT  185.0 259.4 185.8 260.2 ;
      RECT  189.8 259.4 190.6 260.2 ;
      RECT  194.6 259.4 195.4 260.2 ;
      RECT  199.4 259.4 200.2 260.2 ;
      RECT  204.2 259.4 205.0 260.2 ;
      RECT  209.0 259.4 209.8 260.2 ;
      RECT  213.8 259.4 214.6 260.2 ;
      RECT  218.6 259.4 219.4 260.2 ;
      RECT  223.4 259.4 224.2 260.2 ;
      RECT  2.6 264.2 3.4 265.0 ;
      RECT  7.4 264.2 8.2 265.0 ;
      RECT  12.2 264.2 13.0 265.0 ;
      RECT  17.0 264.2 17.8 265.0 ;
      RECT  21.8 264.2 22.6 265.0 ;
      RECT  26.6 264.2 27.4 265.0 ;
      RECT  31.4 264.2 32.2 265.0 ;
      RECT  36.2 264.2 37.0 265.0 ;
      RECT  41.0 264.2 41.8 265.0 ;
      RECT  45.8 264.2 46.6 265.0 ;
      RECT  50.6 264.2 51.4 265.0 ;
      RECT  55.4 264.2 56.2 265.0 ;
      RECT  60.2 264.2 61.0 265.0 ;
      RECT  65.0 264.2 65.8 265.0 ;
      RECT  69.8 264.2 70.6 265.0 ;
      RECT  74.6 264.2 75.4 265.0 ;
      RECT  79.4 264.2 80.2 265.0 ;
      RECT  84.2 264.2 85.0 265.0 ;
      RECT  89.0 264.2 89.8 265.0 ;
      RECT  93.8 264.2 94.6 265.0 ;
      RECT  98.6 264.2 99.4 265.0 ;
      RECT  103.4 264.2 104.2 265.0 ;
      RECT  108.2 264.2 109.0 265.0 ;
      RECT  113.0 264.2 113.8 265.0 ;
      RECT  117.8 264.2 118.6 265.0 ;
      RECT  122.6 264.2 123.4 265.0 ;
      RECT  127.4 264.2 128.2 265.0 ;
      RECT  132.2 264.2 133.0 265.0 ;
      RECT  137.0 264.2 137.8 265.0 ;
      RECT  141.8 264.2 142.6 265.0 ;
      RECT  146.6 264.2 147.4 265.0 ;
      RECT  151.4 264.2 152.2 265.0 ;
      RECT  156.2 264.2 157.0 265.0 ;
      RECT  161.0 264.2 161.8 265.0 ;
      RECT  165.8 264.2 166.6 265.0 ;
      RECT  170.6 264.2 171.4 265.0 ;
      RECT  175.4 264.2 176.2 265.0 ;
      RECT  180.2 264.2 181.0 265.0 ;
      RECT  185.0 264.2 185.8 265.0 ;
      RECT  189.8 264.2 190.6 265.0 ;
      RECT  194.6 264.2 195.4 265.0 ;
      RECT  199.4 264.2 200.2 265.0 ;
      RECT  204.2 264.2 205.0 265.0 ;
      RECT  209.0 264.2 209.8 265.0 ;
      RECT  213.8 264.2 214.6 265.0 ;
      RECT  218.6 264.2 219.4 265.0 ;
      RECT  223.4 264.2 224.2 265.0 ;
      RECT  2.6 269.0 3.4 269.8 ;
      RECT  7.4 269.0 8.2 269.8 ;
      RECT  12.2 269.0 13.0 269.8 ;
      RECT  17.0 269.0 17.8 269.8 ;
      RECT  21.8 269.0 22.6 269.8 ;
      RECT  26.6 269.0 27.4 269.8 ;
      RECT  31.4 269.0 32.2 269.8 ;
      RECT  36.2 269.0 37.0 269.8 ;
      RECT  41.0 269.0 41.8 269.8 ;
      RECT  45.8 269.0 46.6 269.8 ;
      RECT  50.6 269.0 51.4 269.8 ;
      RECT  55.4 269.0 56.2 269.8 ;
      RECT  60.2 269.0 61.0 269.8 ;
      RECT  65.0 269.0 65.8 269.8 ;
      RECT  69.8 269.0 70.6 269.8 ;
      RECT  74.6 269.0 75.4 269.8 ;
      RECT  79.4 269.0 80.2 269.8 ;
      RECT  84.2 269.0 85.0 269.8 ;
      RECT  89.0 269.0 89.8 269.8 ;
      RECT  93.8 269.0 94.6 269.8 ;
      RECT  98.6 269.0 99.4 269.8 ;
      RECT  180.2 269.0 181.0 269.8 ;
      RECT  185.0 269.0 185.8 269.8 ;
      RECT  189.8 269.0 190.6 269.8 ;
      RECT  194.6 269.0 195.4 269.8 ;
      RECT  199.4 269.0 200.2 269.8 ;
      RECT  204.2 269.0 205.0 269.8 ;
      RECT  209.0 269.0 209.8 269.8 ;
      RECT  213.8 269.0 214.6 269.8 ;
      RECT  218.6 269.0 219.4 269.8 ;
      RECT  223.4 269.0 224.2 269.8 ;
      RECT  2.6 273.8 3.4 274.6 ;
      RECT  7.4 273.8 8.2 274.6 ;
      RECT  12.2 273.8 13.0 274.6 ;
      RECT  17.0 273.8 17.8 274.6 ;
      RECT  21.8 273.8 22.6 274.6 ;
      RECT  26.6 273.8 27.4 274.6 ;
      RECT  31.4 273.8 32.2 274.6 ;
      RECT  36.2 273.8 37.0 274.6 ;
      RECT  41.0 273.8 41.8 274.6 ;
      RECT  45.8 273.8 46.6 274.6 ;
      RECT  50.6 273.8 51.4 274.6 ;
      RECT  55.4 273.8 56.2 274.6 ;
      RECT  60.2 273.8 61.0 274.6 ;
      RECT  65.0 273.8 65.8 274.6 ;
      RECT  69.8 273.8 70.6 274.6 ;
      RECT  74.6 273.8 75.4 274.6 ;
      RECT  79.4 273.8 80.2 274.6 ;
      RECT  84.2 273.8 85.0 274.6 ;
      RECT  89.0 273.8 89.8 274.6 ;
      RECT  93.8 273.8 94.6 274.6 ;
      RECT  98.6 273.8 99.4 274.6 ;
      RECT  103.4 273.8 104.2 274.6 ;
      RECT  108.2 273.8 109.0 274.6 ;
      RECT  113.0 273.8 113.8 274.6 ;
      RECT  117.8 273.8 118.6 274.6 ;
      RECT  122.6 273.8 123.4 274.6 ;
      RECT  127.4 273.8 128.2 274.6 ;
      RECT  132.2 273.8 133.0 274.6 ;
      RECT  137.0 273.8 137.8 274.6 ;
      RECT  141.8 273.8 142.6 274.6 ;
      RECT  146.6 273.8 147.4 274.6 ;
      RECT  151.4 273.8 152.2 274.6 ;
      RECT  156.2 273.8 157.0 274.6 ;
      RECT  161.0 273.8 161.8 274.6 ;
      RECT  165.8 273.8 166.6 274.6 ;
      RECT  170.6 273.8 171.4 274.6 ;
      RECT  175.4 273.8 176.2 274.6 ;
      RECT  180.2 273.8 181.0 274.6 ;
      RECT  185.0 273.8 185.8 274.6 ;
      RECT  189.8 273.8 190.6 274.6 ;
      RECT  194.6 273.8 195.4 274.6 ;
      RECT  199.4 273.8 200.2 274.6 ;
      RECT  204.2 273.8 205.0 274.6 ;
      RECT  209.0 273.8 209.8 274.6 ;
      RECT  213.8 273.8 214.6 274.6 ;
      RECT  218.6 273.8 219.4 274.6 ;
      RECT  223.4 273.8 224.2 274.6 ;
      RECT  2.6 278.6 3.4 279.4 ;
      RECT  7.4 278.6 8.2 279.4 ;
      RECT  12.2 278.6 13.0 279.4 ;
      RECT  17.0 278.6 17.8 279.4 ;
      RECT  21.8 278.6 22.6 279.4 ;
      RECT  26.6 278.6 27.4 279.4 ;
      RECT  31.4 278.6 32.2 279.4 ;
      RECT  36.2 278.6 37.0 279.4 ;
      RECT  41.0 278.6 41.8 279.4 ;
      RECT  45.8 278.6 46.6 279.4 ;
      RECT  50.6 278.6 51.4 279.4 ;
      RECT  55.4 278.6 56.2 279.4 ;
      RECT  60.2 278.6 61.0 279.4 ;
      RECT  65.0 278.6 65.8 279.4 ;
      RECT  69.8 278.6 70.6 279.4 ;
      RECT  74.6 278.6 75.4 279.4 ;
      RECT  79.4 278.6 80.2 279.4 ;
      RECT  84.2 278.6 85.0 279.4 ;
      RECT  89.0 278.6 89.8 279.4 ;
      RECT  93.8 278.6 94.6 279.4 ;
      RECT  98.6 278.6 99.4 279.4 ;
      RECT  103.4 278.6 104.2 279.4 ;
      RECT  108.2 278.6 109.0 279.4 ;
      RECT  113.0 278.6 113.8 279.4 ;
      RECT  117.8 278.6 118.6 279.4 ;
      RECT  146.6 278.6 147.4 279.4 ;
      RECT  151.4 278.6 152.2 279.4 ;
      RECT  156.2 278.6 157.0 279.4 ;
      RECT  161.0 278.6 161.8 279.4 ;
      RECT  165.8 278.6 166.6 279.4 ;
      RECT  170.6 278.6 171.4 279.4 ;
      RECT  175.4 278.6 176.2 279.4 ;
      RECT  180.2 278.6 181.0 279.4 ;
      RECT  185.0 278.6 185.8 279.4 ;
      RECT  189.8 278.6 190.6 279.4 ;
      RECT  194.6 278.6 195.4 279.4 ;
      RECT  199.4 278.6 200.2 279.4 ;
      RECT  204.2 278.6 205.0 279.4 ;
      RECT  209.0 278.6 209.8 279.4 ;
      RECT  213.8 278.6 214.6 279.4 ;
      RECT  218.6 278.6 219.4 279.4 ;
      RECT  223.4 278.6 224.2 279.4 ;
      RECT  2.6 283.4 3.4 284.2 ;
      RECT  7.4 283.4 8.2 284.2 ;
      RECT  12.2 283.4 13.0 284.2 ;
      RECT  17.0 283.4 17.8 284.2 ;
      RECT  21.8 283.4 22.6 284.2 ;
      RECT  26.6 283.4 27.4 284.2 ;
      RECT  31.4 283.4 32.2 284.2 ;
      RECT  36.2 283.4 37.0 284.2 ;
      RECT  41.0 283.4 41.8 284.2 ;
      RECT  45.8 283.4 46.6 284.2 ;
      RECT  50.6 283.4 51.4 284.2 ;
      RECT  55.4 283.4 56.2 284.2 ;
      RECT  60.2 283.4 61.0 284.2 ;
      RECT  65.0 283.4 65.8 284.2 ;
      RECT  69.8 283.4 70.6 284.2 ;
      RECT  74.6 283.4 75.4 284.2 ;
      RECT  79.4 283.4 80.2 284.2 ;
      RECT  84.2 283.4 85.0 284.2 ;
      RECT  89.0 283.4 89.8 284.2 ;
      RECT  93.8 283.4 94.6 284.2 ;
      RECT  98.6 283.4 99.4 284.2 ;
      RECT  103.4 283.4 104.2 284.2 ;
      RECT  108.2 283.4 109.0 284.2 ;
      RECT  113.0 283.4 113.8 284.2 ;
      RECT  117.8 283.4 118.6 284.2 ;
      RECT  122.6 283.4 123.4 284.2 ;
      RECT  127.4 283.4 128.2 284.2 ;
      RECT  132.2 283.4 133.0 284.2 ;
      RECT  137.0 283.4 137.8 284.2 ;
      RECT  141.8 283.4 142.6 284.2 ;
      RECT  146.6 283.4 147.4 284.2 ;
      RECT  151.4 283.4 152.2 284.2 ;
      RECT  156.2 283.4 157.0 284.2 ;
      RECT  161.0 283.4 161.8 284.2 ;
      RECT  165.8 283.4 166.6 284.2 ;
      RECT  170.6 283.4 171.4 284.2 ;
      RECT  175.4 283.4 176.2 284.2 ;
      RECT  180.2 283.4 181.0 284.2 ;
      RECT  185.0 283.4 185.8 284.2 ;
      RECT  189.8 283.4 190.6 284.2 ;
      RECT  194.6 283.4 195.4 284.2 ;
      RECT  199.4 283.4 200.2 284.2 ;
      RECT  204.2 283.4 205.0 284.2 ;
      RECT  209.0 283.4 209.8 284.2 ;
      RECT  213.8 283.4 214.6 284.2 ;
      RECT  218.6 283.4 219.4 284.2 ;
      RECT  223.4 283.4 224.2 284.2 ;
      RECT  2.6 288.2 3.4 289.0 ;
      RECT  7.4 288.2 8.2 289.0 ;
      RECT  12.2 288.2 13.0 289.0 ;
      RECT  17.0 288.2 17.8 289.0 ;
      RECT  21.8 288.2 22.6 289.0 ;
      RECT  26.6 288.2 27.4 289.0 ;
      RECT  31.4 288.2 32.2 289.0 ;
      RECT  36.2 288.2 37.0 289.0 ;
      RECT  41.0 288.2 41.8 289.0 ;
      RECT  45.8 288.2 46.6 289.0 ;
      RECT  50.6 288.2 51.4 289.0 ;
      RECT  55.4 288.2 56.2 289.0 ;
      RECT  60.2 288.2 61.0 289.0 ;
      RECT  65.0 288.2 65.8 289.0 ;
      RECT  69.8 288.2 70.6 289.0 ;
      RECT  74.6 288.2 75.4 289.0 ;
      RECT  79.4 288.2 80.2 289.0 ;
      RECT  84.2 288.2 85.0 289.0 ;
      RECT  89.0 288.2 89.8 289.0 ;
      RECT  93.8 288.2 94.6 289.0 ;
      RECT  98.6 288.2 99.4 289.0 ;
      RECT  103.4 288.2 104.2 289.0 ;
      RECT  108.2 288.2 109.0 289.0 ;
      RECT  113.0 288.2 113.8 289.0 ;
      RECT  117.8 288.2 118.6 289.0 ;
      RECT  122.6 288.2 123.4 289.0 ;
      RECT  127.4 288.2 128.2 289.0 ;
      RECT  132.2 288.2 133.0 289.0 ;
      RECT  137.0 288.2 137.8 289.0 ;
      RECT  2.6 293.0 3.4 293.8 ;
      RECT  7.4 293.0 8.2 293.8 ;
      RECT  12.2 293.0 13.0 293.8 ;
      RECT  17.0 293.0 17.8 293.8 ;
      RECT  21.8 293.0 22.6 293.8 ;
      RECT  26.6 293.0 27.4 293.8 ;
      RECT  31.4 293.0 32.2 293.8 ;
      RECT  36.2 293.0 37.0 293.8 ;
      RECT  41.0 293.0 41.8 293.8 ;
      RECT  45.8 293.0 46.6 293.8 ;
      RECT  50.6 293.0 51.4 293.8 ;
      RECT  55.4 293.0 56.2 293.8 ;
      RECT  60.2 293.0 61.0 293.8 ;
      RECT  65.0 293.0 65.8 293.8 ;
      RECT  69.8 293.0 70.6 293.8 ;
      RECT  74.6 293.0 75.4 293.8 ;
      RECT  79.4 293.0 80.2 293.8 ;
      RECT  84.2 293.0 85.0 293.8 ;
      RECT  89.0 293.0 89.8 293.8 ;
      RECT  93.8 293.0 94.6 293.8 ;
      RECT  98.6 293.0 99.4 293.8 ;
      RECT  103.4 293.0 104.2 293.8 ;
      RECT  108.2 293.0 109.0 293.8 ;
      RECT  113.0 293.0 113.8 293.8 ;
      RECT  117.8 293.0 118.6 293.8 ;
      RECT  122.6 293.0 123.4 293.8 ;
      RECT  127.4 293.0 128.2 293.8 ;
      RECT  132.2 293.0 133.0 293.8 ;
      RECT  137.0 293.0 137.8 293.8 ;
      RECT  141.8 293.0 142.6 293.8 ;
      RECT  146.6 293.0 147.4 293.8 ;
      RECT  151.4 293.0 152.2 293.8 ;
      RECT  156.2 293.0 157.0 293.8 ;
      RECT  161.0 293.0 161.8 293.8 ;
      RECT  165.8 293.0 166.6 293.8 ;
      RECT  170.6 293.0 171.4 293.8 ;
      RECT  175.4 293.0 176.2 293.8 ;
      RECT  180.2 293.0 181.0 293.8 ;
      RECT  185.0 293.0 185.8 293.8 ;
      RECT  189.8 293.0 190.6 293.8 ;
      RECT  194.6 293.0 195.4 293.8 ;
      RECT  199.4 293.0 200.2 293.8 ;
      RECT  204.2 293.0 205.0 293.8 ;
      RECT  209.0 293.0 209.8 293.8 ;
      RECT  213.8 293.0 214.6 293.8 ;
      RECT  218.6 293.0 219.4 293.8 ;
      RECT  223.4 293.0 224.2 293.8 ;
      RECT  2.6 297.8 3.4 298.6 ;
      RECT  7.4 297.8 8.2 298.6 ;
      RECT  12.2 297.8 13.0 298.6 ;
      RECT  17.0 297.8 17.8 298.6 ;
      RECT  21.8 297.8 22.6 298.6 ;
      RECT  26.6 297.8 27.4 298.6 ;
      RECT  31.4 297.8 32.2 298.6 ;
      RECT  36.2 297.8 37.0 298.6 ;
      RECT  41.0 297.8 41.8 298.6 ;
      RECT  45.8 297.8 46.6 298.6 ;
      RECT  50.6 297.8 51.4 298.6 ;
      RECT  55.4 297.8 56.2 298.6 ;
      RECT  60.2 297.8 61.0 298.6 ;
      RECT  93.8 297.8 94.6 298.6 ;
      RECT  98.6 297.8 99.4 298.6 ;
      RECT  103.4 297.8 104.2 298.6 ;
      RECT  108.2 297.8 109.0 298.6 ;
      RECT  113.0 297.8 113.8 298.6 ;
      RECT  117.8 297.8 118.6 298.6 ;
      RECT  122.6 297.8 123.4 298.6 ;
      RECT  127.4 297.8 128.2 298.6 ;
      RECT  132.2 297.8 133.0 298.6 ;
      RECT  137.0 297.8 137.8 298.6 ;
      RECT  141.8 297.8 142.6 298.6 ;
      RECT  146.6 297.8 147.4 298.6 ;
      RECT  151.4 297.8 152.2 298.6 ;
      RECT  156.2 297.8 157.0 298.6 ;
      RECT  161.0 297.8 161.8 298.6 ;
      RECT  165.8 297.8 166.6 298.6 ;
      RECT  170.6 297.8 171.4 298.6 ;
      RECT  175.4 297.8 176.2 298.6 ;
      RECT  180.2 297.8 181.0 298.6 ;
      RECT  185.0 297.8 185.8 298.6 ;
      RECT  189.8 297.8 190.6 298.6 ;
      RECT  194.6 297.8 195.4 298.6 ;
      RECT  199.4 297.8 200.2 298.6 ;
      RECT  204.2 297.8 205.0 298.6 ;
      RECT  209.0 297.8 209.8 298.6 ;
      RECT  213.8 297.8 214.6 298.6 ;
      RECT  218.6 297.8 219.4 298.6 ;
      RECT  223.4 297.8 224.2 298.6 ;
      RECT  2.6 302.6 3.4 303.4 ;
      RECT  7.4 302.6 8.2 303.4 ;
      RECT  12.2 302.6 13.0 303.4 ;
      RECT  17.0 302.6 17.8 303.4 ;
      RECT  21.8 302.6 22.6 303.4 ;
      RECT  26.6 302.6 27.4 303.4 ;
      RECT  31.4 302.6 32.2 303.4 ;
      RECT  36.2 302.6 37.0 303.4 ;
      RECT  41.0 302.6 41.8 303.4 ;
      RECT  45.8 302.6 46.6 303.4 ;
      RECT  50.6 302.6 51.4 303.4 ;
      RECT  55.4 302.6 56.2 303.4 ;
      RECT  60.2 302.6 61.0 303.4 ;
      RECT  65.0 302.6 65.8 303.4 ;
      RECT  69.8 302.6 70.6 303.4 ;
      RECT  74.6 302.6 75.4 303.4 ;
      RECT  93.8 302.6 94.6 303.4 ;
      RECT  98.6 302.6 99.4 303.4 ;
      RECT  103.4 302.6 104.2 303.4 ;
      RECT  108.2 302.6 109.0 303.4 ;
      RECT  113.0 302.6 113.8 303.4 ;
      RECT  117.8 302.6 118.6 303.4 ;
      RECT  122.6 302.6 123.4 303.4 ;
      RECT  127.4 302.6 128.2 303.4 ;
      RECT  132.2 302.6 133.0 303.4 ;
      RECT  137.0 302.6 137.8 303.4 ;
      RECT  141.8 302.6 142.6 303.4 ;
      RECT  146.6 302.6 147.4 303.4 ;
      RECT  151.4 302.6 152.2 303.4 ;
      RECT  156.2 302.6 157.0 303.4 ;
      RECT  161.0 302.6 161.8 303.4 ;
      RECT  165.8 302.6 166.6 303.4 ;
      RECT  170.6 302.6 171.4 303.4 ;
      RECT  175.4 302.6 176.2 303.4 ;
      RECT  180.2 302.6 181.0 303.4 ;
      RECT  185.0 302.6 185.8 303.4 ;
      RECT  189.8 302.6 190.6 303.4 ;
      RECT  194.6 302.6 195.4 303.4 ;
      RECT  199.4 302.6 200.2 303.4 ;
      RECT  204.2 302.6 205.0 303.4 ;
      RECT  209.0 302.6 209.8 303.4 ;
      RECT  213.8 302.6 214.6 303.4 ;
      RECT  218.6 302.6 219.4 303.4 ;
      RECT  223.4 302.6 224.2 303.4 ;
      RECT  2.6 307.4 3.4 308.2 ;
      RECT  7.4 307.4 8.2 308.2 ;
      RECT  12.2 307.4 13.0 308.2 ;
      RECT  17.0 307.4 17.8 308.2 ;
      RECT  21.8 307.4 22.6 308.2 ;
      RECT  26.6 307.4 27.4 308.2 ;
      RECT  31.4 307.4 32.2 308.2 ;
      RECT  36.2 307.4 37.0 308.2 ;
      RECT  41.0 307.4 41.8 308.2 ;
      RECT  45.8 307.4 46.6 308.2 ;
      RECT  50.6 307.4 51.4 308.2 ;
      RECT  55.4 307.4 56.2 308.2 ;
      RECT  60.2 307.4 61.0 308.2 ;
      RECT  65.0 307.4 65.8 308.2 ;
      RECT  69.8 307.4 70.6 308.2 ;
      RECT  74.6 307.4 75.4 308.2 ;
      RECT  79.4 307.4 80.2 308.2 ;
      RECT  84.2 307.4 85.0 308.2 ;
      RECT  89.0 307.4 89.8 308.2 ;
      RECT  93.8 307.4 94.6 308.2 ;
      RECT  98.6 307.4 99.4 308.2 ;
      RECT  103.4 307.4 104.2 308.2 ;
      RECT  108.2 307.4 109.0 308.2 ;
      RECT  113.0 307.4 113.8 308.2 ;
      RECT  117.8 307.4 118.6 308.2 ;
      RECT  122.6 307.4 123.4 308.2 ;
      RECT  127.4 307.4 128.2 308.2 ;
      RECT  132.2 307.4 133.0 308.2 ;
      RECT  137.0 307.4 137.8 308.2 ;
      RECT  2.6 312.2 3.4 313.0 ;
      RECT  7.4 312.2 8.2 313.0 ;
      RECT  12.2 312.2 13.0 313.0 ;
      RECT  17.0 312.2 17.8 313.0 ;
      RECT  21.8 312.2 22.6 313.0 ;
      RECT  26.6 312.2 27.4 313.0 ;
      RECT  31.4 312.2 32.2 313.0 ;
      RECT  36.2 312.2 37.0 313.0 ;
      RECT  41.0 312.2 41.8 313.0 ;
      RECT  45.8 312.2 46.6 313.0 ;
      RECT  50.6 312.2 51.4 313.0 ;
      RECT  55.4 312.2 56.2 313.0 ;
      RECT  60.2 312.2 61.0 313.0 ;
      RECT  65.0 312.2 65.8 313.0 ;
      RECT  69.8 312.2 70.6 313.0 ;
      RECT  79.4 312.2 80.2 313.0 ;
      RECT  84.2 312.2 85.0 313.0 ;
      RECT  89.0 312.2 89.8 313.0 ;
      RECT  93.8 312.2 94.6 313.0 ;
      RECT  98.6 312.2 99.4 313.0 ;
      RECT  103.4 312.2 104.2 313.0 ;
      RECT  108.2 312.2 109.0 313.0 ;
      RECT  113.0 312.2 113.8 313.0 ;
      RECT  117.8 312.2 118.6 313.0 ;
      RECT  122.6 312.2 123.4 313.0 ;
      RECT  127.4 312.2 128.2 313.0 ;
      RECT  132.2 312.2 133.0 313.0 ;
      RECT  137.0 312.2 137.8 313.0 ;
      RECT  141.8 312.2 142.6 313.0 ;
      RECT  146.6 312.2 147.4 313.0 ;
      RECT  151.4 312.2 152.2 313.0 ;
      RECT  156.2 312.2 157.0 313.0 ;
      RECT  161.0 312.2 161.8 313.0 ;
      RECT  165.8 312.2 166.6 313.0 ;
      RECT  170.6 312.2 171.4 313.0 ;
      RECT  175.4 312.2 176.2 313.0 ;
      RECT  180.2 312.2 181.0 313.0 ;
      RECT  185.0 312.2 185.8 313.0 ;
      RECT  189.8 312.2 190.6 313.0 ;
      RECT  194.6 312.2 195.4 313.0 ;
      RECT  199.4 312.2 200.2 313.0 ;
      RECT  204.2 312.2 205.0 313.0 ;
      RECT  209.0 312.2 209.8 313.0 ;
      RECT  213.8 312.2 214.6 313.0 ;
      RECT  218.6 312.2 219.4 313.0 ;
      RECT  223.4 312.2 224.2 313.0 ;
      RECT  2.6 317.0 3.4 317.8 ;
      RECT  7.4 317.0 8.2 317.8 ;
      RECT  12.2 317.0 13.0 317.8 ;
      RECT  17.0 317.0 17.8 317.8 ;
      RECT  21.8 317.0 22.6 317.8 ;
      RECT  26.6 317.0 27.4 317.8 ;
      RECT  31.4 317.0 32.2 317.8 ;
      RECT  36.2 317.0 37.0 317.8 ;
      RECT  41.0 317.0 41.8 317.8 ;
      RECT  45.8 317.0 46.6 317.8 ;
      RECT  50.6 317.0 51.4 317.8 ;
      RECT  55.4 317.0 56.2 317.8 ;
      RECT  60.2 317.0 61.0 317.8 ;
      RECT  65.0 317.0 65.8 317.8 ;
      RECT  69.8 317.0 70.6 317.8 ;
      RECT  74.6 317.0 75.4 317.8 ;
      RECT  79.4 317.0 80.2 317.8 ;
      RECT  84.2 317.0 85.0 317.8 ;
      RECT  89.0 317.0 89.8 317.8 ;
      RECT  93.8 317.0 94.6 317.8 ;
      RECT  98.6 317.0 99.4 317.8 ;
      RECT  103.4 317.0 104.2 317.8 ;
      RECT  108.2 317.0 109.0 317.8 ;
      RECT  113.0 317.0 113.8 317.8 ;
      RECT  117.8 317.0 118.6 317.8 ;
      RECT  122.6 317.0 123.4 317.8 ;
      RECT  127.4 317.0 128.2 317.8 ;
      RECT  132.2 317.0 133.0 317.8 ;
      RECT  137.0 317.0 137.8 317.8 ;
      RECT  141.8 317.0 142.6 317.8 ;
      RECT  146.6 317.0 147.4 317.8 ;
      RECT  151.4 317.0 152.2 317.8 ;
      RECT  156.2 317.0 157.0 317.8 ;
      RECT  161.0 317.0 161.8 317.8 ;
      RECT  165.8 317.0 166.6 317.8 ;
      RECT  170.6 317.0 171.4 317.8 ;
      RECT  175.4 317.0 176.2 317.8 ;
      RECT  180.2 317.0 181.0 317.8 ;
      RECT  185.0 317.0 185.8 317.8 ;
      RECT  189.8 317.0 190.6 317.8 ;
      RECT  194.6 317.0 195.4 317.8 ;
      RECT  199.4 317.0 200.2 317.8 ;
      RECT  204.2 317.0 205.0 317.8 ;
      RECT  209.0 317.0 209.8 317.8 ;
      RECT  213.8 317.0 214.6 317.8 ;
      RECT  218.6 317.0 219.4 317.8 ;
      RECT  223.4 317.0 224.2 317.8 ;
      RECT  2.6 321.8 3.4 322.6 ;
      RECT  7.4 321.8 8.2 322.6 ;
      RECT  12.2 321.8 13.0 322.6 ;
      RECT  17.0 321.8 17.8 322.6 ;
      RECT  21.8 321.8 22.6 322.6 ;
      RECT  26.6 321.8 27.4 322.6 ;
      RECT  31.4 321.8 32.2 322.6 ;
      RECT  36.2 321.8 37.0 322.6 ;
      RECT  41.0 321.8 41.8 322.6 ;
      RECT  45.8 321.8 46.6 322.6 ;
      RECT  50.6 321.8 51.4 322.6 ;
      RECT  55.4 321.8 56.2 322.6 ;
      RECT  60.2 321.8 61.0 322.6 ;
      RECT  65.0 321.8 65.8 322.6 ;
      RECT  69.8 321.8 70.6 322.6 ;
      RECT  74.6 321.8 75.4 322.6 ;
      RECT  98.6 321.8 99.4 322.6 ;
      RECT  103.4 321.8 104.2 322.6 ;
      RECT  108.2 321.8 109.0 322.6 ;
      RECT  113.0 321.8 113.8 322.6 ;
      RECT  117.8 321.8 118.6 322.6 ;
      RECT  122.6 321.8 123.4 322.6 ;
      RECT  127.4 321.8 128.2 322.6 ;
      RECT  132.2 321.8 133.0 322.6 ;
      RECT  137.0 321.8 137.8 322.6 ;
      RECT  141.8 321.8 142.6 322.6 ;
      RECT  146.6 321.8 147.4 322.6 ;
      RECT  151.4 321.8 152.2 322.6 ;
      RECT  156.2 321.8 157.0 322.6 ;
      RECT  161.0 321.8 161.8 322.6 ;
      RECT  165.8 321.8 166.6 322.6 ;
      RECT  170.6 321.8 171.4 322.6 ;
      RECT  175.4 321.8 176.2 322.6 ;
      RECT  180.2 321.8 181.0 322.6 ;
      RECT  185.0 321.8 185.8 322.6 ;
      RECT  189.8 321.8 190.6 322.6 ;
      RECT  194.6 321.8 195.4 322.6 ;
      RECT  199.4 321.8 200.2 322.6 ;
      RECT  204.2 321.8 205.0 322.6 ;
      RECT  209.0 321.8 209.8 322.6 ;
      RECT  213.8 321.8 214.6 322.6 ;
      RECT  218.6 321.8 219.4 322.6 ;
      RECT  223.4 321.8 224.2 322.6 ;
      RECT  2.6 326.6 3.4 327.4 ;
      RECT  7.4 326.6 8.2 327.4 ;
      RECT  12.2 326.6 13.0 327.4 ;
      RECT  17.0 326.6 17.8 327.4 ;
      RECT  21.8 326.6 22.6 327.4 ;
      RECT  26.6 326.6 27.4 327.4 ;
      RECT  31.4 326.6 32.2 327.4 ;
      RECT  36.2 326.6 37.0 327.4 ;
      RECT  41.0 326.6 41.8 327.4 ;
      RECT  45.8 326.6 46.6 327.4 ;
      RECT  50.6 326.6 51.4 327.4 ;
      RECT  55.4 326.6 56.2 327.4 ;
      RECT  60.2 326.6 61.0 327.4 ;
      RECT  65.0 326.6 65.8 327.4 ;
      RECT  69.8 326.6 70.6 327.4 ;
      RECT  74.6 326.6 75.4 327.4 ;
      RECT  79.4 326.6 80.2 327.4 ;
      RECT  84.2 326.6 85.0 327.4 ;
      RECT  89.0 326.6 89.8 327.4 ;
      RECT  93.8 326.6 94.6 327.4 ;
      RECT  98.6 326.6 99.4 327.4 ;
      RECT  103.4 326.6 104.2 327.4 ;
      RECT  108.2 326.6 109.0 327.4 ;
      RECT  113.0 326.6 113.8 327.4 ;
      RECT  117.8 326.6 118.6 327.4 ;
      RECT  122.6 326.6 123.4 327.4 ;
      RECT  127.4 326.6 128.2 327.4 ;
      RECT  132.2 326.6 133.0 327.4 ;
      RECT  137.0 326.6 137.8 327.4 ;
      RECT  141.8 326.6 142.6 327.4 ;
      RECT  146.6 326.6 147.4 327.4 ;
      RECT  151.4 326.6 152.2 327.4 ;
      RECT  156.2 326.6 157.0 327.4 ;
      RECT  161.0 326.6 161.8 327.4 ;
      RECT  165.8 326.6 166.6 327.4 ;
      RECT  170.6 326.6 171.4 327.4 ;
      RECT  175.4 326.6 176.2 327.4 ;
      RECT  180.2 326.6 181.0 327.4 ;
      RECT  185.0 326.6 185.8 327.4 ;
      RECT  189.8 326.6 190.6 327.4 ;
      RECT  194.6 326.6 195.4 327.4 ;
      RECT  199.4 326.6 200.2 327.4 ;
      RECT  204.2 326.6 205.0 327.4 ;
      RECT  209.0 326.6 209.8 327.4 ;
      RECT  213.8 326.6 214.6 327.4 ;
      RECT  218.6 326.6 219.4 327.4 ;
      RECT  223.4 326.6 224.2 327.4 ;
      RECT  2.6 331.4 3.4 332.2 ;
      RECT  7.4 331.4 8.2 332.2 ;
      RECT  12.2 331.4 13.0 332.2 ;
      RECT  17.0 331.4 17.8 332.2 ;
      RECT  21.8 331.4 22.6 332.2 ;
      RECT  26.6 331.4 27.4 332.2 ;
      RECT  31.4 331.4 32.2 332.2 ;
      RECT  36.2 331.4 37.0 332.2 ;
      RECT  41.0 331.4 41.8 332.2 ;
      RECT  45.8 331.4 46.6 332.2 ;
      RECT  50.6 331.4 51.4 332.2 ;
      RECT  55.4 331.4 56.2 332.2 ;
      RECT  60.2 331.4 61.0 332.2 ;
      RECT  65.0 331.4 65.8 332.2 ;
      RECT  69.8 331.4 70.6 332.2 ;
      RECT  74.6 331.4 75.4 332.2 ;
      RECT  79.4 331.4 80.2 332.2 ;
      RECT  84.2 331.4 85.0 332.2 ;
      RECT  89.0 331.4 89.8 332.2 ;
      RECT  93.8 331.4 94.6 332.2 ;
      RECT  98.6 331.4 99.4 332.2 ;
      RECT  103.4 331.4 104.2 332.2 ;
      RECT  108.2 331.4 109.0 332.2 ;
      RECT  113.0 331.4 113.8 332.2 ;
      RECT  117.8 331.4 118.6 332.2 ;
      RECT  122.6 331.4 123.4 332.2 ;
      RECT  127.4 331.4 128.2 332.2 ;
      RECT  132.2 331.4 133.0 332.2 ;
      RECT  137.0 331.4 137.8 332.2 ;
      RECT  180.2 331.4 181.0 332.2 ;
      RECT  185.0 331.4 185.8 332.2 ;
      RECT  189.8 331.4 190.6 332.2 ;
      RECT  194.6 331.4 195.4 332.2 ;
      RECT  199.4 331.4 200.2 332.2 ;
      RECT  204.2 331.4 205.0 332.2 ;
      RECT  209.0 331.4 209.8 332.2 ;
      RECT  213.8 331.4 214.6 332.2 ;
      RECT  218.6 331.4 219.4 332.2 ;
      RECT  223.4 331.4 224.2 332.2 ;
      RECT  2.6 336.2 3.4 337.0 ;
      RECT  7.4 336.2 8.2 337.0 ;
      RECT  12.2 336.2 13.0 337.0 ;
      RECT  17.0 336.2 17.8 337.0 ;
      RECT  21.8 336.2 22.6 337.0 ;
      RECT  26.6 336.2 27.4 337.0 ;
      RECT  31.4 336.2 32.2 337.0 ;
      RECT  36.2 336.2 37.0 337.0 ;
      RECT  41.0 336.2 41.8 337.0 ;
      RECT  45.8 336.2 46.6 337.0 ;
      RECT  50.6 336.2 51.4 337.0 ;
      RECT  55.4 336.2 56.2 337.0 ;
      RECT  60.2 336.2 61.0 337.0 ;
      RECT  65.0 336.2 65.8 337.0 ;
      RECT  69.8 336.2 70.6 337.0 ;
      RECT  74.6 336.2 75.4 337.0 ;
      RECT  79.4 336.2 80.2 337.0 ;
      RECT  84.2 336.2 85.0 337.0 ;
      RECT  89.0 336.2 89.8 337.0 ;
      RECT  93.8 336.2 94.6 337.0 ;
      RECT  98.6 336.2 99.4 337.0 ;
      RECT  103.4 336.2 104.2 337.0 ;
      RECT  108.2 336.2 109.0 337.0 ;
      RECT  113.0 336.2 113.8 337.0 ;
      RECT  117.8 336.2 118.6 337.0 ;
      RECT  122.6 336.2 123.4 337.0 ;
      RECT  127.4 336.2 128.2 337.0 ;
      RECT  132.2 336.2 133.0 337.0 ;
      RECT  137.0 336.2 137.8 337.0 ;
      RECT  141.8 336.2 142.6 337.0 ;
      RECT  146.6 336.2 147.4 337.0 ;
      RECT  151.4 336.2 152.2 337.0 ;
      RECT  156.2 336.2 157.0 337.0 ;
      RECT  161.0 336.2 161.8 337.0 ;
      RECT  165.8 336.2 166.6 337.0 ;
      RECT  170.6 336.2 171.4 337.0 ;
      RECT  175.4 336.2 176.2 337.0 ;
      RECT  180.2 336.2 181.0 337.0 ;
      RECT  185.0 336.2 185.8 337.0 ;
      RECT  189.8 336.2 190.6 337.0 ;
      RECT  194.6 336.2 195.4 337.0 ;
      RECT  199.4 336.2 200.2 337.0 ;
      RECT  204.2 336.2 205.0 337.0 ;
      RECT  209.0 336.2 209.8 337.0 ;
      RECT  213.8 336.2 214.6 337.0 ;
      RECT  218.6 336.2 219.4 337.0 ;
      RECT  223.4 336.2 224.2 337.0 ;
      RECT  2.6 341.0 3.4 341.8 ;
      RECT  7.4 341.0 8.2 341.8 ;
      RECT  12.2 341.0 13.0 341.8 ;
      RECT  17.0 341.0 17.8 341.8 ;
      RECT  21.8 341.0 22.6 341.8 ;
      RECT  26.6 341.0 27.4 341.8 ;
      RECT  31.4 341.0 32.2 341.8 ;
      RECT  36.2 341.0 37.0 341.8 ;
      RECT  41.0 341.0 41.8 341.8 ;
      RECT  45.8 341.0 46.6 341.8 ;
      RECT  50.6 341.0 51.4 341.8 ;
      RECT  55.4 341.0 56.2 341.8 ;
      RECT  60.2 341.0 61.0 341.8 ;
      RECT  65.0 341.0 65.8 341.8 ;
      RECT  69.8 341.0 70.6 341.8 ;
      RECT  74.6 341.0 75.4 341.8 ;
      RECT  98.6 341.0 99.4 341.8 ;
      RECT  103.4 341.0 104.2 341.8 ;
      RECT  108.2 341.0 109.0 341.8 ;
      RECT  113.0 341.0 113.8 341.8 ;
      RECT  117.8 341.0 118.6 341.8 ;
      RECT  122.6 341.0 123.4 341.8 ;
      RECT  127.4 341.0 128.2 341.8 ;
      RECT  132.2 341.0 133.0 341.8 ;
      RECT  137.0 341.0 137.8 341.8 ;
      RECT  141.8 341.0 142.6 341.8 ;
      RECT  146.6 341.0 147.4 341.8 ;
      RECT  151.4 341.0 152.2 341.8 ;
      RECT  156.2 341.0 157.0 341.8 ;
      RECT  161.0 341.0 161.8 341.8 ;
      RECT  165.8 341.0 166.6 341.8 ;
      RECT  170.6 341.0 171.4 341.8 ;
      RECT  175.4 341.0 176.2 341.8 ;
      RECT  180.2 341.0 181.0 341.8 ;
      RECT  185.0 341.0 185.8 341.8 ;
      RECT  189.8 341.0 190.6 341.8 ;
      RECT  194.6 341.0 195.4 341.8 ;
      RECT  199.4 341.0 200.2 341.8 ;
      RECT  204.2 341.0 205.0 341.8 ;
      RECT  209.0 341.0 209.8 341.8 ;
      RECT  213.8 341.0 214.6 341.8 ;
      RECT  218.6 341.0 219.4 341.8 ;
      RECT  223.4 341.0 224.2 341.8 ;
      RECT  2.6 345.8 3.4 346.6 ;
      RECT  7.4 345.8 8.2 346.6 ;
      RECT  12.2 345.8 13.0 346.6 ;
      RECT  17.0 345.8 17.8 346.6 ;
      RECT  21.8 345.8 22.6 346.6 ;
      RECT  26.6 345.8 27.4 346.6 ;
      RECT  31.4 345.8 32.2 346.6 ;
      RECT  36.2 345.8 37.0 346.6 ;
      RECT  41.0 345.8 41.8 346.6 ;
      RECT  45.8 345.8 46.6 346.6 ;
      RECT  50.6 345.8 51.4 346.6 ;
      RECT  55.4 345.8 56.2 346.6 ;
      RECT  60.2 345.8 61.0 346.6 ;
      RECT  65.0 345.8 65.8 346.6 ;
      RECT  69.8 345.8 70.6 346.6 ;
      RECT  74.6 345.8 75.4 346.6 ;
      RECT  79.4 345.8 80.2 346.6 ;
      RECT  84.2 345.8 85.0 346.6 ;
      RECT  89.0 345.8 89.8 346.6 ;
      RECT  93.8 345.8 94.6 346.6 ;
      RECT  98.6 345.8 99.4 346.6 ;
      RECT  103.4 345.8 104.2 346.6 ;
      RECT  108.2 345.8 109.0 346.6 ;
      RECT  113.0 345.8 113.8 346.6 ;
      RECT  117.8 345.8 118.6 346.6 ;
      RECT  122.6 345.8 123.4 346.6 ;
      RECT  127.4 345.8 128.2 346.6 ;
      RECT  132.2 345.8 133.0 346.6 ;
      RECT  137.0 345.8 137.8 346.6 ;
      RECT  141.8 345.8 142.6 346.6 ;
      RECT  146.6 345.8 147.4 346.6 ;
      RECT  151.4 345.8 152.2 346.6 ;
      RECT  156.2 345.8 157.0 346.6 ;
      RECT  161.0 345.8 161.8 346.6 ;
      RECT  165.8 345.8 166.6 346.6 ;
      RECT  170.6 345.8 171.4 346.6 ;
      RECT  175.4 345.8 176.2 346.6 ;
      RECT  180.2 345.8 181.0 346.6 ;
      RECT  185.0 345.8 185.8 346.6 ;
      RECT  189.8 345.8 190.6 346.6 ;
      RECT  194.6 345.8 195.4 346.6 ;
      RECT  199.4 345.8 200.2 346.6 ;
      RECT  204.2 345.8 205.0 346.6 ;
      RECT  209.0 345.8 209.8 346.6 ;
      RECT  213.8 345.8 214.6 346.6 ;
      RECT  218.6 345.8 219.4 346.6 ;
      RECT  223.4 345.8 224.2 346.6 ;
      RECT  2.6 350.6 3.4 351.4 ;
      RECT  7.4 350.6 8.2 351.4 ;
      RECT  12.2 350.6 13.0 351.4 ;
      RECT  17.0 350.6 17.8 351.4 ;
      RECT  21.8 350.6 22.6 351.4 ;
      RECT  26.6 350.6 27.4 351.4 ;
      RECT  31.4 350.6 32.2 351.4 ;
      RECT  36.2 350.6 37.0 351.4 ;
      RECT  41.0 350.6 41.8 351.4 ;
      RECT  45.8 350.6 46.6 351.4 ;
      RECT  50.6 350.6 51.4 351.4 ;
      RECT  55.4 350.6 56.2 351.4 ;
      RECT  60.2 350.6 61.0 351.4 ;
      RECT  65.0 350.6 65.8 351.4 ;
      RECT  69.8 350.6 70.6 351.4 ;
      RECT  79.4 350.6 80.2 351.4 ;
      RECT  84.2 350.6 85.0 351.4 ;
      RECT  89.0 350.6 89.8 351.4 ;
      RECT  93.8 350.6 94.6 351.4 ;
      RECT  98.6 350.6 99.4 351.4 ;
      RECT  103.4 350.6 104.2 351.4 ;
      RECT  108.2 350.6 109.0 351.4 ;
      RECT  113.0 350.6 113.8 351.4 ;
      RECT  117.8 350.6 118.6 351.4 ;
      RECT  122.6 350.6 123.4 351.4 ;
      RECT  127.4 350.6 128.2 351.4 ;
      RECT  132.2 350.6 133.0 351.4 ;
      RECT  137.0 350.6 137.8 351.4 ;
      RECT  2.6 355.4 3.4 356.2 ;
      RECT  7.4 355.4 8.2 356.2 ;
      RECT  12.2 355.4 13.0 356.2 ;
      RECT  17.0 355.4 17.8 356.2 ;
      RECT  21.8 355.4 22.6 356.2 ;
      RECT  26.6 355.4 27.4 356.2 ;
      RECT  31.4 355.4 32.2 356.2 ;
      RECT  36.2 355.4 37.0 356.2 ;
      RECT  41.0 355.4 41.8 356.2 ;
      RECT  45.8 355.4 46.6 356.2 ;
      RECT  50.6 355.4 51.4 356.2 ;
      RECT  55.4 355.4 56.2 356.2 ;
      RECT  60.2 355.4 61.0 356.2 ;
      RECT  65.0 355.4 65.8 356.2 ;
      RECT  69.8 355.4 70.6 356.2 ;
      RECT  74.6 355.4 75.4 356.2 ;
      RECT  79.4 355.4 80.2 356.2 ;
      RECT  84.2 355.4 85.0 356.2 ;
      RECT  89.0 355.4 89.8 356.2 ;
      RECT  93.8 355.4 94.6 356.2 ;
      RECT  98.6 355.4 99.4 356.2 ;
      RECT  103.4 355.4 104.2 356.2 ;
      RECT  108.2 355.4 109.0 356.2 ;
      RECT  113.0 355.4 113.8 356.2 ;
      RECT  117.8 355.4 118.6 356.2 ;
      RECT  122.6 355.4 123.4 356.2 ;
      RECT  127.4 355.4 128.2 356.2 ;
      RECT  132.2 355.4 133.0 356.2 ;
      RECT  137.0 355.4 137.8 356.2 ;
      RECT  141.8 355.4 142.6 356.2 ;
      RECT  146.6 355.4 147.4 356.2 ;
      RECT  151.4 355.4 152.2 356.2 ;
      RECT  156.2 355.4 157.0 356.2 ;
      RECT  161.0 355.4 161.8 356.2 ;
      RECT  165.8 355.4 166.6 356.2 ;
      RECT  170.6 355.4 171.4 356.2 ;
      RECT  175.4 355.4 176.2 356.2 ;
      RECT  180.2 355.4 181.0 356.2 ;
      RECT  185.0 355.4 185.8 356.2 ;
      RECT  189.8 355.4 190.6 356.2 ;
      RECT  194.6 355.4 195.4 356.2 ;
      RECT  199.4 355.4 200.2 356.2 ;
      RECT  204.2 355.4 205.0 356.2 ;
      RECT  209.0 355.4 209.8 356.2 ;
      RECT  213.8 355.4 214.6 356.2 ;
      RECT  218.6 355.4 219.4 356.2 ;
      RECT  223.4 355.4 224.2 356.2 ;
      RECT  2.6 360.2 3.4 361.0 ;
      RECT  7.4 360.2 8.2 361.0 ;
      RECT  12.2 360.2 13.0 361.0 ;
      RECT  17.0 360.2 17.8 361.0 ;
      RECT  21.8 360.2 22.6 361.0 ;
      RECT  26.6 360.2 27.4 361.0 ;
      RECT  31.4 360.2 32.2 361.0 ;
      RECT  36.2 360.2 37.0 361.0 ;
      RECT  41.0 360.2 41.8 361.0 ;
      RECT  45.8 360.2 46.6 361.0 ;
      RECT  50.6 360.2 51.4 361.0 ;
      RECT  55.4 360.2 56.2 361.0 ;
      RECT  60.2 360.2 61.0 361.0 ;
      RECT  65.0 360.2 65.8 361.0 ;
      RECT  69.8 360.2 70.6 361.0 ;
      RECT  74.6 360.2 75.4 361.0 ;
      RECT  79.4 360.2 80.2 361.0 ;
      RECT  84.2 360.2 85.0 361.0 ;
      RECT  89.0 360.2 89.8 361.0 ;
      RECT  93.8 360.2 94.6 361.0 ;
      RECT  98.6 360.2 99.4 361.0 ;
      RECT  103.4 360.2 104.2 361.0 ;
      RECT  108.2 360.2 109.0 361.0 ;
      RECT  113.0 360.2 113.8 361.0 ;
      RECT  117.8 360.2 118.6 361.0 ;
      RECT  122.6 360.2 123.4 361.0 ;
      RECT  127.4 360.2 128.2 361.0 ;
      RECT  132.2 360.2 133.0 361.0 ;
      RECT  137.0 360.2 137.8 361.0 ;
      RECT  141.8 360.2 142.6 361.0 ;
      RECT  146.6 360.2 147.4 361.0 ;
      RECT  151.4 360.2 152.2 361.0 ;
      RECT  156.2 360.2 157.0 361.0 ;
      RECT  161.0 360.2 161.8 361.0 ;
      RECT  165.8 360.2 166.6 361.0 ;
      RECT  170.6 360.2 171.4 361.0 ;
      RECT  175.4 360.2 176.2 361.0 ;
      RECT  180.2 360.2 181.0 361.0 ;
      RECT  185.0 360.2 185.8 361.0 ;
      RECT  189.8 360.2 190.6 361.0 ;
      RECT  194.6 360.2 195.4 361.0 ;
      RECT  199.4 360.2 200.2 361.0 ;
      RECT  204.2 360.2 205.0 361.0 ;
      RECT  209.0 360.2 209.8 361.0 ;
      RECT  213.8 360.2 214.6 361.0 ;
      RECT  218.6 360.2 219.4 361.0 ;
      RECT  223.4 360.2 224.2 361.0 ;
      RECT  2.6 365.0 3.4 365.8 ;
      RECT  7.4 365.0 8.2 365.8 ;
      RECT  12.2 365.0 13.0 365.8 ;
      RECT  17.0 365.0 17.8 365.8 ;
      RECT  21.8 365.0 22.6 365.8 ;
      RECT  26.6 365.0 27.4 365.8 ;
      RECT  31.4 365.0 32.2 365.8 ;
      RECT  36.2 365.0 37.0 365.8 ;
      RECT  41.0 365.0 41.8 365.8 ;
      RECT  45.8 365.0 46.6 365.8 ;
      RECT  50.6 365.0 51.4 365.8 ;
      RECT  55.4 365.0 56.2 365.8 ;
      RECT  60.2 365.0 61.0 365.8 ;
      RECT  65.0 365.0 65.8 365.8 ;
      RECT  69.8 365.0 70.6 365.8 ;
      RECT  74.6 365.0 75.4 365.8 ;
      RECT  79.4 365.0 80.2 365.8 ;
      RECT  84.2 365.0 85.0 365.8 ;
      RECT  89.0 365.0 89.8 365.8 ;
      RECT  93.8 365.0 94.6 365.8 ;
      RECT  98.6 365.0 99.4 365.8 ;
      RECT  103.4 365.0 104.2 365.8 ;
      RECT  108.2 365.0 109.0 365.8 ;
      RECT  113.0 365.0 113.8 365.8 ;
      RECT  117.8 365.0 118.6 365.8 ;
      RECT  122.6 365.0 123.4 365.8 ;
      RECT  127.4 365.0 128.2 365.8 ;
      RECT  132.2 365.0 133.0 365.8 ;
      RECT  137.0 365.0 137.8 365.8 ;
      RECT  141.8 365.0 142.6 365.8 ;
      RECT  146.6 365.0 147.4 365.8 ;
      RECT  151.4 365.0 152.2 365.8 ;
      RECT  156.2 365.0 157.0 365.8 ;
      RECT  161.0 365.0 161.8 365.8 ;
      RECT  165.8 365.0 166.6 365.8 ;
      RECT  170.6 365.0 171.4 365.8 ;
      RECT  175.4 365.0 176.2 365.8 ;
      RECT  180.2 365.0 181.0 365.8 ;
      RECT  185.0 365.0 185.8 365.8 ;
      RECT  189.8 365.0 190.6 365.8 ;
      RECT  194.6 365.0 195.4 365.8 ;
      RECT  199.4 365.0 200.2 365.8 ;
      RECT  204.2 365.0 205.0 365.8 ;
      RECT  209.0 365.0 209.8 365.8 ;
      RECT  213.8 365.0 214.6 365.8 ;
      RECT  218.6 365.0 219.4 365.8 ;
      RECT  223.4 365.0 224.2 365.8 ;
      RECT  2.6 369.8 3.4 370.6 ;
      RECT  7.4 369.8 8.2 370.6 ;
      RECT  12.2 369.8 13.0 370.6 ;
      RECT  17.0 369.8 17.8 370.6 ;
      RECT  21.8 369.8 22.6 370.6 ;
      RECT  26.6 369.8 27.4 370.6 ;
      RECT  31.4 369.8 32.2 370.6 ;
      RECT  36.2 369.8 37.0 370.6 ;
      RECT  41.0 369.8 41.8 370.6 ;
      RECT  45.8 369.8 46.6 370.6 ;
      RECT  50.6 369.8 51.4 370.6 ;
      RECT  55.4 369.8 56.2 370.6 ;
      RECT  60.2 369.8 61.0 370.6 ;
      RECT  65.0 369.8 65.8 370.6 ;
      RECT  69.8 369.8 70.6 370.6 ;
      RECT  74.6 369.8 75.4 370.6 ;
      RECT  79.4 369.8 80.2 370.6 ;
      RECT  84.2 369.8 85.0 370.6 ;
      RECT  89.0 369.8 89.8 370.6 ;
      RECT  93.8 369.8 94.6 370.6 ;
      RECT  98.6 369.8 99.4 370.6 ;
      RECT  103.4 369.8 104.2 370.6 ;
      RECT  108.2 369.8 109.0 370.6 ;
      RECT  113.0 369.8 113.8 370.6 ;
      RECT  117.8 369.8 118.6 370.6 ;
      RECT  122.6 369.8 123.4 370.6 ;
      RECT  127.4 369.8 128.2 370.6 ;
      RECT  132.2 369.8 133.0 370.6 ;
      RECT  137.0 369.8 137.8 370.6 ;
      RECT  141.8 369.8 142.6 370.6 ;
      RECT  146.6 369.8 147.4 370.6 ;
      RECT  151.4 369.8 152.2 370.6 ;
      RECT  156.2 369.8 157.0 370.6 ;
      RECT  161.0 369.8 161.8 370.6 ;
      RECT  165.8 369.8 166.6 370.6 ;
      RECT  170.6 369.8 171.4 370.6 ;
      RECT  175.4 369.8 176.2 370.6 ;
      RECT  180.2 369.8 181.0 370.6 ;
      RECT  5.0 2.6 5.8 3.4 ;
      RECT  9.8 2.6 10.6 3.4 ;
      RECT  14.6 2.6 15.4 3.4 ;
      RECT  19.4 2.6 20.2 3.4 ;
      RECT  24.2 2.6 25.0 3.4 ;
      RECT  29.0 2.6 29.8 3.4 ;
      RECT  33.8 2.6 34.6 3.4 ;
      RECT  38.6 2.6 39.4 3.4 ;
      RECT  43.4 2.6 44.2 3.4 ;
      RECT  48.2 2.6 49.0 3.4 ;
      RECT  53.0 2.6 53.8 3.4 ;
      RECT  57.8 2.6 58.6 3.4 ;
      RECT  62.6 2.6 63.4 3.4 ;
      RECT  67.4 2.6 68.2 3.4 ;
      RECT  72.2 2.6 73.0 3.4 ;
      RECT  77.0 2.6 77.8 3.4 ;
      RECT  91.4 2.6 92.2 3.4 ;
      RECT  96.2 2.6 97.0 3.4 ;
      RECT  101.0 2.6 101.8 3.4 ;
      RECT  105.8 2.6 106.6 3.4 ;
      RECT  110.6 2.6 111.4 3.4 ;
      RECT  115.4 2.6 116.2 3.4 ;
      RECT  120.2 2.6 121.0 3.4 ;
      RECT  125.0 2.6 125.8 3.4 ;
      RECT  129.8 2.6 130.6 3.4 ;
      RECT  134.6 2.6 135.4 3.4 ;
      RECT  139.4 2.6 140.2 3.4 ;
      RECT  144.2 2.6 145.0 3.4 ;
      RECT  149.0 2.6 149.8 3.4 ;
      RECT  153.8 2.6 154.6 3.4 ;
      RECT  158.6 2.6 159.4 3.4 ;
      RECT  163.4 2.6 164.2 3.4 ;
      RECT  168.2 2.6 169.0 3.4 ;
      RECT  173.0 2.6 173.8 3.4 ;
      RECT  177.8 2.6 178.6 3.4 ;
      RECT  182.6 2.6 183.4 3.4 ;
      RECT  187.4 2.6 188.2 3.4 ;
      RECT  192.2 2.6 193.0 3.4 ;
      RECT  197.0 2.6 197.8 3.4 ;
      RECT  201.8 2.6 202.6 3.4 ;
      RECT  206.6 2.6 207.4 3.4 ;
      RECT  211.4 2.6 212.2 3.4 ;
      RECT  216.2 2.6 217.0 3.4 ;
      RECT  221.0 2.6 221.8 3.4 ;
      RECT  225.8 2.6 226.6 3.4 ;
      RECT  5.0 7.4 5.8 8.2 ;
      RECT  9.8 7.4 10.6 8.2 ;
      RECT  14.6 7.4 15.4 8.2 ;
      RECT  19.4 7.4 20.2 8.2 ;
      RECT  24.2 7.4 25.0 8.2 ;
      RECT  29.0 7.4 29.8 8.2 ;
      RECT  33.8 7.4 34.6 8.2 ;
      RECT  38.6 7.4 39.4 8.2 ;
      RECT  43.4 7.4 44.2 8.2 ;
      RECT  48.2 7.4 49.0 8.2 ;
      RECT  53.0 7.4 53.8 8.2 ;
      RECT  57.8 7.4 58.6 8.2 ;
      RECT  62.6 7.4 63.4 8.2 ;
      RECT  67.4 7.4 68.2 8.2 ;
      RECT  72.2 7.4 73.0 8.2 ;
      RECT  77.0 7.4 77.8 8.2 ;
      RECT  81.8 7.4 82.6 8.2 ;
      RECT  86.6 7.4 87.4 8.2 ;
      RECT  91.4 7.4 92.2 8.2 ;
      RECT  96.2 7.4 97.0 8.2 ;
      RECT  101.0 7.4 101.8 8.2 ;
      RECT  105.8 7.4 106.6 8.2 ;
      RECT  110.6 7.4 111.4 8.2 ;
      RECT  115.4 7.4 116.2 8.2 ;
      RECT  120.2 7.4 121.0 8.2 ;
      RECT  125.0 7.4 125.8 8.2 ;
      RECT  129.8 7.4 130.6 8.2 ;
      RECT  134.6 7.4 135.4 8.2 ;
      RECT  139.4 7.4 140.2 8.2 ;
      RECT  144.2 7.4 145.0 8.2 ;
      RECT  149.0 7.4 149.8 8.2 ;
      RECT  153.8 7.4 154.6 8.2 ;
      RECT  158.6 7.4 159.4 8.2 ;
      RECT  163.4 7.4 164.2 8.2 ;
      RECT  168.2 7.4 169.0 8.2 ;
      RECT  173.0 7.4 173.8 8.2 ;
      RECT  177.8 7.4 178.6 8.2 ;
      RECT  182.6 7.4 183.4 8.2 ;
      RECT  187.4 7.4 188.2 8.2 ;
      RECT  192.2 7.4 193.0 8.2 ;
      RECT  197.0 7.4 197.8 8.2 ;
      RECT  201.8 7.4 202.6 8.2 ;
      RECT  206.6 7.4 207.4 8.2 ;
      RECT  211.4 7.4 212.2 8.2 ;
      RECT  216.2 7.4 217.0 8.2 ;
      RECT  221.0 7.4 221.8 8.2 ;
      RECT  225.8 7.4 226.6 8.2 ;
      RECT  53.0 12.2 53.8 13.0 ;
      RECT  57.8 12.2 58.6 13.0 ;
      RECT  62.6 12.2 63.4 13.0 ;
      RECT  67.4 12.2 68.2 13.0 ;
      RECT  72.2 12.2 73.0 13.0 ;
      RECT  77.0 12.2 77.8 13.0 ;
      RECT  81.8 12.2 82.6 13.0 ;
      RECT  86.6 12.2 87.4 13.0 ;
      RECT  91.4 12.2 92.2 13.0 ;
      RECT  96.2 12.2 97.0 13.0 ;
      RECT  101.0 12.2 101.8 13.0 ;
      RECT  105.8 12.2 106.6 13.0 ;
      RECT  110.6 12.2 111.4 13.0 ;
      RECT  115.4 12.2 116.2 13.0 ;
      RECT  120.2 12.2 121.0 13.0 ;
      RECT  125.0 12.2 125.8 13.0 ;
      RECT  129.8 12.2 130.6 13.0 ;
      RECT  134.6 12.2 135.4 13.0 ;
      RECT  139.4 12.2 140.2 13.0 ;
      RECT  144.2 12.2 145.0 13.0 ;
      RECT  149.0 12.2 149.8 13.0 ;
      RECT  153.8 12.2 154.6 13.0 ;
      RECT  158.6 12.2 159.4 13.0 ;
      RECT  163.4 12.2 164.2 13.0 ;
      RECT  168.2 12.2 169.0 13.0 ;
      RECT  173.0 12.2 173.8 13.0 ;
      RECT  177.8 12.2 178.6 13.0 ;
      RECT  182.6 12.2 183.4 13.0 ;
      RECT  187.4 12.2 188.2 13.0 ;
      RECT  192.2 12.2 193.0 13.0 ;
      RECT  197.0 12.2 197.8 13.0 ;
      RECT  201.8 12.2 202.6 13.0 ;
      RECT  206.6 12.2 207.4 13.0 ;
      RECT  211.4 12.2 212.2 13.0 ;
      RECT  216.2 12.2 217.0 13.0 ;
      RECT  221.0 12.2 221.8 13.0 ;
      RECT  225.8 12.2 226.6 13.0 ;
      RECT  5.0 17.0 5.8 17.8 ;
      RECT  9.8 17.0 10.6 17.8 ;
      RECT  14.6 17.0 15.4 17.8 ;
      RECT  19.4 17.0 20.2 17.8 ;
      RECT  24.2 17.0 25.0 17.8 ;
      RECT  29.0 17.0 29.8 17.8 ;
      RECT  33.8 17.0 34.6 17.8 ;
      RECT  38.6 17.0 39.4 17.8 ;
      RECT  43.4 17.0 44.2 17.8 ;
      RECT  48.2 17.0 49.0 17.8 ;
      RECT  53.0 17.0 53.8 17.8 ;
      RECT  57.8 17.0 58.6 17.8 ;
      RECT  62.6 17.0 63.4 17.8 ;
      RECT  67.4 17.0 68.2 17.8 ;
      RECT  72.2 17.0 73.0 17.8 ;
      RECT  77.0 17.0 77.8 17.8 ;
      RECT  81.8 17.0 82.6 17.8 ;
      RECT  86.6 17.0 87.4 17.8 ;
      RECT  91.4 17.0 92.2 17.8 ;
      RECT  96.2 17.0 97.0 17.8 ;
      RECT  101.0 17.0 101.8 17.8 ;
      RECT  105.8 17.0 106.6 17.8 ;
      RECT  110.6 17.0 111.4 17.8 ;
      RECT  115.4 17.0 116.2 17.8 ;
      RECT  120.2 17.0 121.0 17.8 ;
      RECT  125.0 17.0 125.8 17.8 ;
      RECT  129.8 17.0 130.6 17.8 ;
      RECT  134.6 17.0 135.4 17.8 ;
      RECT  139.4 17.0 140.2 17.8 ;
      RECT  144.2 17.0 145.0 17.8 ;
      RECT  149.0 17.0 149.8 17.8 ;
      RECT  153.8 17.0 154.6 17.8 ;
      RECT  158.6 17.0 159.4 17.8 ;
      RECT  163.4 17.0 164.2 17.8 ;
      RECT  168.2 17.0 169.0 17.8 ;
      RECT  173.0 17.0 173.8 17.8 ;
      RECT  177.8 17.0 178.6 17.8 ;
      RECT  182.6 17.0 183.4 17.8 ;
      RECT  187.4 17.0 188.2 17.8 ;
      RECT  192.2 17.0 193.0 17.8 ;
      RECT  197.0 17.0 197.8 17.8 ;
      RECT  201.8 17.0 202.6 17.8 ;
      RECT  206.6 17.0 207.4 17.8 ;
      RECT  211.4 17.0 212.2 17.8 ;
      RECT  216.2 17.0 217.0 17.8 ;
      RECT  221.0 17.0 221.8 17.8 ;
      RECT  225.8 17.0 226.6 17.8 ;
      RECT  5.0 21.8 5.8 22.6 ;
      RECT  9.8 21.8 10.6 22.6 ;
      RECT  14.6 21.8 15.4 22.6 ;
      RECT  19.4 21.8 20.2 22.6 ;
      RECT  24.2 21.8 25.0 22.6 ;
      RECT  29.0 21.8 29.8 22.6 ;
      RECT  33.8 21.8 34.6 22.6 ;
      RECT  38.6 21.8 39.4 22.6 ;
      RECT  43.4 21.8 44.2 22.6 ;
      RECT  48.2 21.8 49.0 22.6 ;
      RECT  53.0 21.8 53.8 22.6 ;
      RECT  57.8 21.8 58.6 22.6 ;
      RECT  62.6 21.8 63.4 22.6 ;
      RECT  67.4 21.8 68.2 22.6 ;
      RECT  72.2 21.8 73.0 22.6 ;
      RECT  77.0 21.8 77.8 22.6 ;
      RECT  81.8 21.8 82.6 22.6 ;
      RECT  86.6 21.8 87.4 22.6 ;
      RECT  91.4 21.8 92.2 22.6 ;
      RECT  96.2 21.8 97.0 22.6 ;
      RECT  101.0 21.8 101.8 22.6 ;
      RECT  105.8 21.8 106.6 22.6 ;
      RECT  110.6 21.8 111.4 22.6 ;
      RECT  115.4 21.8 116.2 22.6 ;
      RECT  120.2 21.8 121.0 22.6 ;
      RECT  125.0 21.8 125.8 22.6 ;
      RECT  129.8 21.8 130.6 22.6 ;
      RECT  134.6 21.8 135.4 22.6 ;
      RECT  139.4 21.8 140.2 22.6 ;
      RECT  144.2 21.8 145.0 22.6 ;
      RECT  149.0 21.8 149.8 22.6 ;
      RECT  153.8 21.8 154.6 22.6 ;
      RECT  158.6 21.8 159.4 22.6 ;
      RECT  163.4 21.8 164.2 22.6 ;
      RECT  168.2 21.8 169.0 22.6 ;
      RECT  173.0 21.8 173.8 22.6 ;
      RECT  177.8 21.8 178.6 22.6 ;
      RECT  182.6 21.8 183.4 22.6 ;
      RECT  187.4 21.8 188.2 22.6 ;
      RECT  192.2 21.8 193.0 22.6 ;
      RECT  197.0 21.8 197.8 22.6 ;
      RECT  201.8 21.8 202.6 22.6 ;
      RECT  206.6 21.8 207.4 22.6 ;
      RECT  211.4 21.8 212.2 22.6 ;
      RECT  216.2 21.8 217.0 22.6 ;
      RECT  221.0 21.8 221.8 22.6 ;
      RECT  225.8 21.8 226.6 22.6 ;
      RECT  5.0 26.6 5.8 27.4 ;
      RECT  9.8 26.6 10.6 27.4 ;
      RECT  14.6 26.6 15.4 27.4 ;
      RECT  19.4 26.6 20.2 27.4 ;
      RECT  24.2 26.6 25.0 27.4 ;
      RECT  29.0 26.6 29.8 27.4 ;
      RECT  33.8 26.6 34.6 27.4 ;
      RECT  38.6 26.6 39.4 27.4 ;
      RECT  43.4 26.6 44.2 27.4 ;
      RECT  48.2 26.6 49.0 27.4 ;
      RECT  53.0 26.6 53.8 27.4 ;
      RECT  57.8 26.6 58.6 27.4 ;
      RECT  62.6 26.6 63.4 27.4 ;
      RECT  67.4 26.6 68.2 27.4 ;
      RECT  72.2 26.6 73.0 27.4 ;
      RECT  77.0 26.6 77.8 27.4 ;
      RECT  81.8 26.6 82.6 27.4 ;
      RECT  86.6 26.6 87.4 27.4 ;
      RECT  91.4 26.6 92.2 27.4 ;
      RECT  96.2 26.6 97.0 27.4 ;
      RECT  101.0 26.6 101.8 27.4 ;
      RECT  105.8 26.6 106.6 27.4 ;
      RECT  110.6 26.6 111.4 27.4 ;
      RECT  115.4 26.6 116.2 27.4 ;
      RECT  120.2 26.6 121.0 27.4 ;
      RECT  125.0 26.6 125.8 27.4 ;
      RECT  129.8 26.6 130.6 27.4 ;
      RECT  134.6 26.6 135.4 27.4 ;
      RECT  139.4 26.6 140.2 27.4 ;
      RECT  144.2 26.6 145.0 27.4 ;
      RECT  149.0 26.6 149.8 27.4 ;
      RECT  153.8 26.6 154.6 27.4 ;
      RECT  158.6 26.6 159.4 27.4 ;
      RECT  163.4 26.6 164.2 27.4 ;
      RECT  168.2 26.6 169.0 27.4 ;
      RECT  173.0 26.6 173.8 27.4 ;
      RECT  177.8 26.6 178.6 27.4 ;
      RECT  182.6 26.6 183.4 27.4 ;
      RECT  187.4 26.6 188.2 27.4 ;
      RECT  192.2 26.6 193.0 27.4 ;
      RECT  197.0 26.6 197.8 27.4 ;
      RECT  201.8 26.6 202.6 27.4 ;
      RECT  206.6 26.6 207.4 27.4 ;
      RECT  211.4 26.6 212.2 27.4 ;
      RECT  216.2 26.6 217.0 27.4 ;
      RECT  221.0 26.6 221.8 27.4 ;
      RECT  225.8 26.6 226.6 27.4 ;
      RECT  86.6 31.4 87.4 32.2 ;
      RECT  91.4 31.4 92.2 32.2 ;
      RECT  96.2 31.4 97.0 32.2 ;
      RECT  101.0 31.4 101.8 32.2 ;
      RECT  105.8 31.4 106.6 32.2 ;
      RECT  110.6 31.4 111.4 32.2 ;
      RECT  115.4 31.4 116.2 32.2 ;
      RECT  120.2 31.4 121.0 32.2 ;
      RECT  125.0 31.4 125.8 32.2 ;
      RECT  129.8 31.4 130.6 32.2 ;
      RECT  134.6 31.4 135.4 32.2 ;
      RECT  139.4 31.4 140.2 32.2 ;
      RECT  144.2 31.4 145.0 32.2 ;
      RECT  149.0 31.4 149.8 32.2 ;
      RECT  153.8 31.4 154.6 32.2 ;
      RECT  158.6 31.4 159.4 32.2 ;
      RECT  163.4 31.4 164.2 32.2 ;
      RECT  168.2 31.4 169.0 32.2 ;
      RECT  173.0 31.4 173.8 32.2 ;
      RECT  177.8 31.4 178.6 32.2 ;
      RECT  182.6 31.4 183.4 32.2 ;
      RECT  187.4 31.4 188.2 32.2 ;
      RECT  192.2 31.4 193.0 32.2 ;
      RECT  197.0 31.4 197.8 32.2 ;
      RECT  201.8 31.4 202.6 32.2 ;
      RECT  206.6 31.4 207.4 32.2 ;
      RECT  211.4 31.4 212.2 32.2 ;
      RECT  216.2 31.4 217.0 32.2 ;
      RECT  221.0 31.4 221.8 32.2 ;
      RECT  225.8 31.4 226.6 32.2 ;
      RECT  5.0 36.2 5.8 37.0 ;
      RECT  9.8 36.2 10.6 37.0 ;
      RECT  14.6 36.2 15.4 37.0 ;
      RECT  19.4 36.2 20.2 37.0 ;
      RECT  24.2 36.2 25.0 37.0 ;
      RECT  29.0 36.2 29.8 37.0 ;
      RECT  33.8 36.2 34.6 37.0 ;
      RECT  38.6 36.2 39.4 37.0 ;
      RECT  62.6 36.2 63.4 37.0 ;
      RECT  67.4 36.2 68.2 37.0 ;
      RECT  72.2 36.2 73.0 37.0 ;
      RECT  77.0 36.2 77.8 37.0 ;
      RECT  81.8 36.2 82.6 37.0 ;
      RECT  86.6 36.2 87.4 37.0 ;
      RECT  91.4 36.2 92.2 37.0 ;
      RECT  96.2 36.2 97.0 37.0 ;
      RECT  101.0 36.2 101.8 37.0 ;
      RECT  105.8 36.2 106.6 37.0 ;
      RECT  110.6 36.2 111.4 37.0 ;
      RECT  115.4 36.2 116.2 37.0 ;
      RECT  120.2 36.2 121.0 37.0 ;
      RECT  125.0 36.2 125.8 37.0 ;
      RECT  129.8 36.2 130.6 37.0 ;
      RECT  134.6 36.2 135.4 37.0 ;
      RECT  139.4 36.2 140.2 37.0 ;
      RECT  144.2 36.2 145.0 37.0 ;
      RECT  149.0 36.2 149.8 37.0 ;
      RECT  153.8 36.2 154.6 37.0 ;
      RECT  158.6 36.2 159.4 37.0 ;
      RECT  163.4 36.2 164.2 37.0 ;
      RECT  168.2 36.2 169.0 37.0 ;
      RECT  173.0 36.2 173.8 37.0 ;
      RECT  177.8 36.2 178.6 37.0 ;
      RECT  182.6 36.2 183.4 37.0 ;
      RECT  187.4 36.2 188.2 37.0 ;
      RECT  192.2 36.2 193.0 37.0 ;
      RECT  197.0 36.2 197.8 37.0 ;
      RECT  201.8 36.2 202.6 37.0 ;
      RECT  206.6 36.2 207.4 37.0 ;
      RECT  211.4 36.2 212.2 37.0 ;
      RECT  216.2 36.2 217.0 37.0 ;
      RECT  221.0 36.2 221.8 37.0 ;
      RECT  225.8 36.2 226.6 37.0 ;
      RECT  5.0 41.0 5.8 41.8 ;
      RECT  9.8 41.0 10.6 41.8 ;
      RECT  14.6 41.0 15.4 41.8 ;
      RECT  19.4 41.0 20.2 41.8 ;
      RECT  24.2 41.0 25.0 41.8 ;
      RECT  29.0 41.0 29.8 41.8 ;
      RECT  33.8 41.0 34.6 41.8 ;
      RECT  38.6 41.0 39.4 41.8 ;
      RECT  43.4 41.0 44.2 41.8 ;
      RECT  48.2 41.0 49.0 41.8 ;
      RECT  53.0 41.0 53.8 41.8 ;
      RECT  57.8 41.0 58.6 41.8 ;
      RECT  62.6 41.0 63.4 41.8 ;
      RECT  67.4 41.0 68.2 41.8 ;
      RECT  72.2 41.0 73.0 41.8 ;
      RECT  77.0 41.0 77.8 41.8 ;
      RECT  91.4 41.0 92.2 41.8 ;
      RECT  96.2 41.0 97.0 41.8 ;
      RECT  101.0 41.0 101.8 41.8 ;
      RECT  105.8 41.0 106.6 41.8 ;
      RECT  110.6 41.0 111.4 41.8 ;
      RECT  115.4 41.0 116.2 41.8 ;
      RECT  120.2 41.0 121.0 41.8 ;
      RECT  125.0 41.0 125.8 41.8 ;
      RECT  129.8 41.0 130.6 41.8 ;
      RECT  134.6 41.0 135.4 41.8 ;
      RECT  139.4 41.0 140.2 41.8 ;
      RECT  144.2 41.0 145.0 41.8 ;
      RECT  149.0 41.0 149.8 41.8 ;
      RECT  153.8 41.0 154.6 41.8 ;
      RECT  158.6 41.0 159.4 41.8 ;
      RECT  163.4 41.0 164.2 41.8 ;
      RECT  168.2 41.0 169.0 41.8 ;
      RECT  173.0 41.0 173.8 41.8 ;
      RECT  177.8 41.0 178.6 41.8 ;
      RECT  182.6 41.0 183.4 41.8 ;
      RECT  187.4 41.0 188.2 41.8 ;
      RECT  192.2 41.0 193.0 41.8 ;
      RECT  197.0 41.0 197.8 41.8 ;
      RECT  201.8 41.0 202.6 41.8 ;
      RECT  206.6 41.0 207.4 41.8 ;
      RECT  211.4 41.0 212.2 41.8 ;
      RECT  216.2 41.0 217.0 41.8 ;
      RECT  221.0 41.0 221.8 41.8 ;
      RECT  225.8 41.0 226.6 41.8 ;
      RECT  5.0 45.8 5.8 46.6 ;
      RECT  9.8 45.8 10.6 46.6 ;
      RECT  14.6 45.8 15.4 46.6 ;
      RECT  19.4 45.8 20.2 46.6 ;
      RECT  24.2 45.8 25.0 46.6 ;
      RECT  29.0 45.8 29.8 46.6 ;
      RECT  33.8 45.8 34.6 46.6 ;
      RECT  38.6 45.8 39.4 46.6 ;
      RECT  43.4 45.8 44.2 46.6 ;
      RECT  48.2 45.8 49.0 46.6 ;
      RECT  53.0 45.8 53.8 46.6 ;
      RECT  57.8 45.8 58.6 46.6 ;
      RECT  62.6 45.8 63.4 46.6 ;
      RECT  67.4 45.8 68.2 46.6 ;
      RECT  72.2 45.8 73.0 46.6 ;
      RECT  77.0 45.8 77.8 46.6 ;
      RECT  81.8 45.8 82.6 46.6 ;
      RECT  86.6 45.8 87.4 46.6 ;
      RECT  91.4 45.8 92.2 46.6 ;
      RECT  96.2 45.8 97.0 46.6 ;
      RECT  101.0 45.8 101.8 46.6 ;
      RECT  105.8 45.8 106.6 46.6 ;
      RECT  110.6 45.8 111.4 46.6 ;
      RECT  115.4 45.8 116.2 46.6 ;
      RECT  120.2 45.8 121.0 46.6 ;
      RECT  125.0 45.8 125.8 46.6 ;
      RECT  129.8 45.8 130.6 46.6 ;
      RECT  134.6 45.8 135.4 46.6 ;
      RECT  139.4 45.8 140.2 46.6 ;
      RECT  144.2 45.8 145.0 46.6 ;
      RECT  149.0 45.8 149.8 46.6 ;
      RECT  153.8 45.8 154.6 46.6 ;
      RECT  158.6 45.8 159.4 46.6 ;
      RECT  163.4 45.8 164.2 46.6 ;
      RECT  168.2 45.8 169.0 46.6 ;
      RECT  173.0 45.8 173.8 46.6 ;
      RECT  177.8 45.8 178.6 46.6 ;
      RECT  182.6 45.8 183.4 46.6 ;
      RECT  187.4 45.8 188.2 46.6 ;
      RECT  5.0 50.6 5.8 51.4 ;
      RECT  9.8 50.6 10.6 51.4 ;
      RECT  14.6 50.6 15.4 51.4 ;
      RECT  19.4 50.6 20.2 51.4 ;
      RECT  24.2 50.6 25.0 51.4 ;
      RECT  29.0 50.6 29.8 51.4 ;
      RECT  33.8 50.6 34.6 51.4 ;
      RECT  81.8 50.6 82.6 51.4 ;
      RECT  86.6 50.6 87.4 51.4 ;
      RECT  91.4 50.6 92.2 51.4 ;
      RECT  96.2 50.6 97.0 51.4 ;
      RECT  101.0 50.6 101.8 51.4 ;
      RECT  105.8 50.6 106.6 51.4 ;
      RECT  110.6 50.6 111.4 51.4 ;
      RECT  115.4 50.6 116.2 51.4 ;
      RECT  120.2 50.6 121.0 51.4 ;
      RECT  125.0 50.6 125.8 51.4 ;
      RECT  129.8 50.6 130.6 51.4 ;
      RECT  134.6 50.6 135.4 51.4 ;
      RECT  139.4 50.6 140.2 51.4 ;
      RECT  144.2 50.6 145.0 51.4 ;
      RECT  149.0 50.6 149.8 51.4 ;
      RECT  153.8 50.6 154.6 51.4 ;
      RECT  158.6 50.6 159.4 51.4 ;
      RECT  163.4 50.6 164.2 51.4 ;
      RECT  168.2 50.6 169.0 51.4 ;
      RECT  173.0 50.6 173.8 51.4 ;
      RECT  177.8 50.6 178.6 51.4 ;
      RECT  182.6 50.6 183.4 51.4 ;
      RECT  187.4 50.6 188.2 51.4 ;
      RECT  192.2 50.6 193.0 51.4 ;
      RECT  197.0 50.6 197.8 51.4 ;
      RECT  201.8 50.6 202.6 51.4 ;
      RECT  206.6 50.6 207.4 51.4 ;
      RECT  211.4 50.6 212.2 51.4 ;
      RECT  216.2 50.6 217.0 51.4 ;
      RECT  221.0 50.6 221.8 51.4 ;
      RECT  225.8 50.6 226.6 51.4 ;
      RECT  5.0 55.4 5.8 56.2 ;
      RECT  9.8 55.4 10.6 56.2 ;
      RECT  14.6 55.4 15.4 56.2 ;
      RECT  19.4 55.4 20.2 56.2 ;
      RECT  24.2 55.4 25.0 56.2 ;
      RECT  29.0 55.4 29.8 56.2 ;
      RECT  33.8 55.4 34.6 56.2 ;
      RECT  38.6 55.4 39.4 56.2 ;
      RECT  43.4 55.4 44.2 56.2 ;
      RECT  48.2 55.4 49.0 56.2 ;
      RECT  53.0 55.4 53.8 56.2 ;
      RECT  57.8 55.4 58.6 56.2 ;
      RECT  62.6 55.4 63.4 56.2 ;
      RECT  67.4 55.4 68.2 56.2 ;
      RECT  72.2 55.4 73.0 56.2 ;
      RECT  77.0 55.4 77.8 56.2 ;
      RECT  81.8 55.4 82.6 56.2 ;
      RECT  86.6 55.4 87.4 56.2 ;
      RECT  91.4 55.4 92.2 56.2 ;
      RECT  96.2 55.4 97.0 56.2 ;
      RECT  101.0 55.4 101.8 56.2 ;
      RECT  105.8 55.4 106.6 56.2 ;
      RECT  110.6 55.4 111.4 56.2 ;
      RECT  115.4 55.4 116.2 56.2 ;
      RECT  120.2 55.4 121.0 56.2 ;
      RECT  125.0 55.4 125.8 56.2 ;
      RECT  129.8 55.4 130.6 56.2 ;
      RECT  134.6 55.4 135.4 56.2 ;
      RECT  139.4 55.4 140.2 56.2 ;
      RECT  144.2 55.4 145.0 56.2 ;
      RECT  149.0 55.4 149.8 56.2 ;
      RECT  153.8 55.4 154.6 56.2 ;
      RECT  158.6 55.4 159.4 56.2 ;
      RECT  163.4 55.4 164.2 56.2 ;
      RECT  168.2 55.4 169.0 56.2 ;
      RECT  173.0 55.4 173.8 56.2 ;
      RECT  177.8 55.4 178.6 56.2 ;
      RECT  182.6 55.4 183.4 56.2 ;
      RECT  187.4 55.4 188.2 56.2 ;
      RECT  192.2 55.4 193.0 56.2 ;
      RECT  197.0 55.4 197.8 56.2 ;
      RECT  201.8 55.4 202.6 56.2 ;
      RECT  206.6 55.4 207.4 56.2 ;
      RECT  211.4 55.4 212.2 56.2 ;
      RECT  216.2 55.4 217.0 56.2 ;
      RECT  221.0 55.4 221.8 56.2 ;
      RECT  225.8 55.4 226.6 56.2 ;
      RECT  5.0 60.2 5.8 61.0 ;
      RECT  9.8 60.2 10.6 61.0 ;
      RECT  14.6 60.2 15.4 61.0 ;
      RECT  19.4 60.2 20.2 61.0 ;
      RECT  24.2 60.2 25.0 61.0 ;
      RECT  29.0 60.2 29.8 61.0 ;
      RECT  33.8 60.2 34.6 61.0 ;
      RECT  38.6 60.2 39.4 61.0 ;
      RECT  43.4 60.2 44.2 61.0 ;
      RECT  48.2 60.2 49.0 61.0 ;
      RECT  53.0 60.2 53.8 61.0 ;
      RECT  57.8 60.2 58.6 61.0 ;
      RECT  62.6 60.2 63.4 61.0 ;
      RECT  67.4 60.2 68.2 61.0 ;
      RECT  72.2 60.2 73.0 61.0 ;
      RECT  77.0 60.2 77.8 61.0 ;
      RECT  81.8 60.2 82.6 61.0 ;
      RECT  86.6 60.2 87.4 61.0 ;
      RECT  91.4 60.2 92.2 61.0 ;
      RECT  96.2 60.2 97.0 61.0 ;
      RECT  101.0 60.2 101.8 61.0 ;
      RECT  105.8 60.2 106.6 61.0 ;
      RECT  110.6 60.2 111.4 61.0 ;
      RECT  115.4 60.2 116.2 61.0 ;
      RECT  120.2 60.2 121.0 61.0 ;
      RECT  125.0 60.2 125.8 61.0 ;
      RECT  129.8 60.2 130.6 61.0 ;
      RECT  134.6 60.2 135.4 61.0 ;
      RECT  139.4 60.2 140.2 61.0 ;
      RECT  144.2 60.2 145.0 61.0 ;
      RECT  149.0 60.2 149.8 61.0 ;
      RECT  153.8 60.2 154.6 61.0 ;
      RECT  158.6 60.2 159.4 61.0 ;
      RECT  163.4 60.2 164.2 61.0 ;
      RECT  168.2 60.2 169.0 61.0 ;
      RECT  173.0 60.2 173.8 61.0 ;
      RECT  177.8 60.2 178.6 61.0 ;
      RECT  182.6 60.2 183.4 61.0 ;
      RECT  187.4 60.2 188.2 61.0 ;
      RECT  192.2 60.2 193.0 61.0 ;
      RECT  197.0 60.2 197.8 61.0 ;
      RECT  201.8 60.2 202.6 61.0 ;
      RECT  206.6 60.2 207.4 61.0 ;
      RECT  211.4 60.2 212.2 61.0 ;
      RECT  216.2 60.2 217.0 61.0 ;
      RECT  221.0 60.2 221.8 61.0 ;
      RECT  225.8 60.2 226.6 61.0 ;
      RECT  5.0 65.0 5.8 65.8 ;
      RECT  9.8 65.0 10.6 65.8 ;
      RECT  14.6 65.0 15.4 65.8 ;
      RECT  19.4 65.0 20.2 65.8 ;
      RECT  24.2 65.0 25.0 65.8 ;
      RECT  29.0 65.0 29.8 65.8 ;
      RECT  33.8 65.0 34.6 65.8 ;
      RECT  38.6 65.0 39.4 65.8 ;
      RECT  43.4 65.0 44.2 65.8 ;
      RECT  48.2 65.0 49.0 65.8 ;
      RECT  53.0 65.0 53.8 65.8 ;
      RECT  57.8 65.0 58.6 65.8 ;
      RECT  62.6 65.0 63.4 65.8 ;
      RECT  67.4 65.0 68.2 65.8 ;
      RECT  72.2 65.0 73.0 65.8 ;
      RECT  77.0 65.0 77.8 65.8 ;
      RECT  81.8 65.0 82.6 65.8 ;
      RECT  86.6 65.0 87.4 65.8 ;
      RECT  91.4 65.0 92.2 65.8 ;
      RECT  96.2 65.0 97.0 65.8 ;
      RECT  101.0 65.0 101.8 65.8 ;
      RECT  105.8 65.0 106.6 65.8 ;
      RECT  110.6 65.0 111.4 65.8 ;
      RECT  115.4 65.0 116.2 65.8 ;
      RECT  120.2 65.0 121.0 65.8 ;
      RECT  125.0 65.0 125.8 65.8 ;
      RECT  129.8 65.0 130.6 65.8 ;
      RECT  134.6 65.0 135.4 65.8 ;
      RECT  139.4 65.0 140.2 65.8 ;
      RECT  144.2 65.0 145.0 65.8 ;
      RECT  149.0 65.0 149.8 65.8 ;
      RECT  153.8 65.0 154.6 65.8 ;
      RECT  158.6 65.0 159.4 65.8 ;
      RECT  163.4 65.0 164.2 65.8 ;
      RECT  168.2 65.0 169.0 65.8 ;
      RECT  173.0 65.0 173.8 65.8 ;
      RECT  177.8 65.0 178.6 65.8 ;
      RECT  182.6 65.0 183.4 65.8 ;
      RECT  187.4 65.0 188.2 65.8 ;
      RECT  192.2 65.0 193.0 65.8 ;
      RECT  197.0 65.0 197.8 65.8 ;
      RECT  201.8 65.0 202.6 65.8 ;
      RECT  206.6 65.0 207.4 65.8 ;
      RECT  211.4 65.0 212.2 65.8 ;
      RECT  216.2 65.0 217.0 65.8 ;
      RECT  221.0 65.0 221.8 65.8 ;
      RECT  225.8 65.0 226.6 65.8 ;
      RECT  5.0 69.8 5.8 70.6 ;
      RECT  9.8 69.8 10.6 70.6 ;
      RECT  14.6 69.8 15.4 70.6 ;
      RECT  19.4 69.8 20.2 70.6 ;
      RECT  24.2 69.8 25.0 70.6 ;
      RECT  29.0 69.8 29.8 70.6 ;
      RECT  33.8 69.8 34.6 70.6 ;
      RECT  38.6 69.8 39.4 70.6 ;
      RECT  43.4 69.8 44.2 70.6 ;
      RECT  48.2 69.8 49.0 70.6 ;
      RECT  53.0 69.8 53.8 70.6 ;
      RECT  57.8 69.8 58.6 70.6 ;
      RECT  62.6 69.8 63.4 70.6 ;
      RECT  67.4 69.8 68.2 70.6 ;
      RECT  72.2 69.8 73.0 70.6 ;
      RECT  77.0 69.8 77.8 70.6 ;
      RECT  81.8 69.8 82.6 70.6 ;
      RECT  86.6 69.8 87.4 70.6 ;
      RECT  91.4 69.8 92.2 70.6 ;
      RECT  96.2 69.8 97.0 70.6 ;
      RECT  101.0 69.8 101.8 70.6 ;
      RECT  105.8 69.8 106.6 70.6 ;
      RECT  110.6 69.8 111.4 70.6 ;
      RECT  115.4 69.8 116.2 70.6 ;
      RECT  120.2 69.8 121.0 70.6 ;
      RECT  125.0 69.8 125.8 70.6 ;
      RECT  129.8 69.8 130.6 70.6 ;
      RECT  134.6 69.8 135.4 70.6 ;
      RECT  139.4 69.8 140.2 70.6 ;
      RECT  144.2 69.8 145.0 70.6 ;
      RECT  149.0 69.8 149.8 70.6 ;
      RECT  153.8 69.8 154.6 70.6 ;
      RECT  158.6 69.8 159.4 70.6 ;
      RECT  163.4 69.8 164.2 70.6 ;
      RECT  168.2 69.8 169.0 70.6 ;
      RECT  173.0 69.8 173.8 70.6 ;
      RECT  177.8 69.8 178.6 70.6 ;
      RECT  182.6 69.8 183.4 70.6 ;
      RECT  187.4 69.8 188.2 70.6 ;
      RECT  192.2 69.8 193.0 70.6 ;
      RECT  197.0 69.8 197.8 70.6 ;
      RECT  201.8 69.8 202.6 70.6 ;
      RECT  206.6 69.8 207.4 70.6 ;
      RECT  211.4 69.8 212.2 70.6 ;
      RECT  216.2 69.8 217.0 70.6 ;
      RECT  221.0 69.8 221.8 70.6 ;
      RECT  225.8 69.8 226.6 70.6 ;
      RECT  5.0 74.6 5.8 75.4 ;
      RECT  9.8 74.6 10.6 75.4 ;
      RECT  14.6 74.6 15.4 75.4 ;
      RECT  19.4 74.6 20.2 75.4 ;
      RECT  24.2 74.6 25.0 75.4 ;
      RECT  29.0 74.6 29.8 75.4 ;
      RECT  33.8 74.6 34.6 75.4 ;
      RECT  38.6 74.6 39.4 75.4 ;
      RECT  43.4 74.6 44.2 75.4 ;
      RECT  48.2 74.6 49.0 75.4 ;
      RECT  53.0 74.6 53.8 75.4 ;
      RECT  57.8 74.6 58.6 75.4 ;
      RECT  62.6 74.6 63.4 75.4 ;
      RECT  67.4 74.6 68.2 75.4 ;
      RECT  72.2 74.6 73.0 75.4 ;
      RECT  77.0 74.6 77.8 75.4 ;
      RECT  81.8 74.6 82.6 75.4 ;
      RECT  187.4 74.6 188.2 75.4 ;
      RECT  192.2 74.6 193.0 75.4 ;
      RECT  197.0 74.6 197.8 75.4 ;
      RECT  201.8 74.6 202.6 75.4 ;
      RECT  206.6 74.6 207.4 75.4 ;
      RECT  211.4 74.6 212.2 75.4 ;
      RECT  216.2 74.6 217.0 75.4 ;
      RECT  221.0 74.6 221.8 75.4 ;
      RECT  225.8 74.6 226.6 75.4 ;
      RECT  5.0 79.4 5.8 80.2 ;
      RECT  9.8 79.4 10.6 80.2 ;
      RECT  14.6 79.4 15.4 80.2 ;
      RECT  19.4 79.4 20.2 80.2 ;
      RECT  24.2 79.4 25.0 80.2 ;
      RECT  29.0 79.4 29.8 80.2 ;
      RECT  33.8 79.4 34.6 80.2 ;
      RECT  38.6 79.4 39.4 80.2 ;
      RECT  43.4 79.4 44.2 80.2 ;
      RECT  48.2 79.4 49.0 80.2 ;
      RECT  53.0 79.4 53.8 80.2 ;
      RECT  57.8 79.4 58.6 80.2 ;
      RECT  62.6 79.4 63.4 80.2 ;
      RECT  67.4 79.4 68.2 80.2 ;
      RECT  72.2 79.4 73.0 80.2 ;
      RECT  77.0 79.4 77.8 80.2 ;
      RECT  81.8 79.4 82.6 80.2 ;
      RECT  86.6 79.4 87.4 80.2 ;
      RECT  91.4 79.4 92.2 80.2 ;
      RECT  96.2 79.4 97.0 80.2 ;
      RECT  101.0 79.4 101.8 80.2 ;
      RECT  105.8 79.4 106.6 80.2 ;
      RECT  110.6 79.4 111.4 80.2 ;
      RECT  115.4 79.4 116.2 80.2 ;
      RECT  120.2 79.4 121.0 80.2 ;
      RECT  125.0 79.4 125.8 80.2 ;
      RECT  129.8 79.4 130.6 80.2 ;
      RECT  134.6 79.4 135.4 80.2 ;
      RECT  139.4 79.4 140.2 80.2 ;
      RECT  144.2 79.4 145.0 80.2 ;
      RECT  149.0 79.4 149.8 80.2 ;
      RECT  153.8 79.4 154.6 80.2 ;
      RECT  158.6 79.4 159.4 80.2 ;
      RECT  163.4 79.4 164.2 80.2 ;
      RECT  168.2 79.4 169.0 80.2 ;
      RECT  173.0 79.4 173.8 80.2 ;
      RECT  177.8 79.4 178.6 80.2 ;
      RECT  182.6 79.4 183.4 80.2 ;
      RECT  187.4 79.4 188.2 80.2 ;
      RECT  192.2 79.4 193.0 80.2 ;
      RECT  197.0 79.4 197.8 80.2 ;
      RECT  201.8 79.4 202.6 80.2 ;
      RECT  206.6 79.4 207.4 80.2 ;
      RECT  211.4 79.4 212.2 80.2 ;
      RECT  216.2 79.4 217.0 80.2 ;
      RECT  221.0 79.4 221.8 80.2 ;
      RECT  225.8 79.4 226.6 80.2 ;
      RECT  5.0 84.2 5.8 85.0 ;
      RECT  9.8 84.2 10.6 85.0 ;
      RECT  14.6 84.2 15.4 85.0 ;
      RECT  19.4 84.2 20.2 85.0 ;
      RECT  24.2 84.2 25.0 85.0 ;
      RECT  29.0 84.2 29.8 85.0 ;
      RECT  33.8 84.2 34.6 85.0 ;
      RECT  38.6 84.2 39.4 85.0 ;
      RECT  43.4 84.2 44.2 85.0 ;
      RECT  48.2 84.2 49.0 85.0 ;
      RECT  53.0 84.2 53.8 85.0 ;
      RECT  57.8 84.2 58.6 85.0 ;
      RECT  62.6 84.2 63.4 85.0 ;
      RECT  67.4 84.2 68.2 85.0 ;
      RECT  72.2 84.2 73.0 85.0 ;
      RECT  77.0 84.2 77.8 85.0 ;
      RECT  81.8 84.2 82.6 85.0 ;
      RECT  86.6 84.2 87.4 85.0 ;
      RECT  91.4 84.2 92.2 85.0 ;
      RECT  96.2 84.2 97.0 85.0 ;
      RECT  101.0 84.2 101.8 85.0 ;
      RECT  105.8 84.2 106.6 85.0 ;
      RECT  110.6 84.2 111.4 85.0 ;
      RECT  115.4 84.2 116.2 85.0 ;
      RECT  120.2 84.2 121.0 85.0 ;
      RECT  125.0 84.2 125.8 85.0 ;
      RECT  129.8 84.2 130.6 85.0 ;
      RECT  134.6 84.2 135.4 85.0 ;
      RECT  139.4 84.2 140.2 85.0 ;
      RECT  144.2 84.2 145.0 85.0 ;
      RECT  149.0 84.2 149.8 85.0 ;
      RECT  153.8 84.2 154.6 85.0 ;
      RECT  158.6 84.2 159.4 85.0 ;
      RECT  163.4 84.2 164.2 85.0 ;
      RECT  168.2 84.2 169.0 85.0 ;
      RECT  173.0 84.2 173.8 85.0 ;
      RECT  177.8 84.2 178.6 85.0 ;
      RECT  182.6 84.2 183.4 85.0 ;
      RECT  187.4 84.2 188.2 85.0 ;
      RECT  192.2 84.2 193.0 85.0 ;
      RECT  197.0 84.2 197.8 85.0 ;
      RECT  201.8 84.2 202.6 85.0 ;
      RECT  206.6 84.2 207.4 85.0 ;
      RECT  211.4 84.2 212.2 85.0 ;
      RECT  216.2 84.2 217.0 85.0 ;
      RECT  221.0 84.2 221.8 85.0 ;
      RECT  225.8 84.2 226.6 85.0 ;
      RECT  5.0 89.0 5.8 89.8 ;
      RECT  9.8 89.0 10.6 89.8 ;
      RECT  14.6 89.0 15.4 89.8 ;
      RECT  19.4 89.0 20.2 89.8 ;
      RECT  24.2 89.0 25.0 89.8 ;
      RECT  29.0 89.0 29.8 89.8 ;
      RECT  33.8 89.0 34.6 89.8 ;
      RECT  38.6 89.0 39.4 89.8 ;
      RECT  43.4 89.0 44.2 89.8 ;
      RECT  48.2 89.0 49.0 89.8 ;
      RECT  53.0 89.0 53.8 89.8 ;
      RECT  57.8 89.0 58.6 89.8 ;
      RECT  62.6 89.0 63.4 89.8 ;
      RECT  67.4 89.0 68.2 89.8 ;
      RECT  72.2 89.0 73.0 89.8 ;
      RECT  77.0 89.0 77.8 89.8 ;
      RECT  81.8 89.0 82.6 89.8 ;
      RECT  5.0 93.8 5.8 94.6 ;
      RECT  9.8 93.8 10.6 94.6 ;
      RECT  14.6 93.8 15.4 94.6 ;
      RECT  19.4 93.8 20.2 94.6 ;
      RECT  24.2 93.8 25.0 94.6 ;
      RECT  29.0 93.8 29.8 94.6 ;
      RECT  33.8 93.8 34.6 94.6 ;
      RECT  38.6 93.8 39.4 94.6 ;
      RECT  43.4 93.8 44.2 94.6 ;
      RECT  48.2 93.8 49.0 94.6 ;
      RECT  53.0 93.8 53.8 94.6 ;
      RECT  57.8 93.8 58.6 94.6 ;
      RECT  62.6 93.8 63.4 94.6 ;
      RECT  67.4 93.8 68.2 94.6 ;
      RECT  72.2 93.8 73.0 94.6 ;
      RECT  77.0 93.8 77.8 94.6 ;
      RECT  81.8 93.8 82.6 94.6 ;
      RECT  86.6 93.8 87.4 94.6 ;
      RECT  91.4 93.8 92.2 94.6 ;
      RECT  96.2 93.8 97.0 94.6 ;
      RECT  101.0 93.8 101.8 94.6 ;
      RECT  105.8 93.8 106.6 94.6 ;
      RECT  110.6 93.8 111.4 94.6 ;
      RECT  115.4 93.8 116.2 94.6 ;
      RECT  120.2 93.8 121.0 94.6 ;
      RECT  125.0 93.8 125.8 94.6 ;
      RECT  129.8 93.8 130.6 94.6 ;
      RECT  134.6 93.8 135.4 94.6 ;
      RECT  139.4 93.8 140.2 94.6 ;
      RECT  144.2 93.8 145.0 94.6 ;
      RECT  149.0 93.8 149.8 94.6 ;
      RECT  153.8 93.8 154.6 94.6 ;
      RECT  158.6 93.8 159.4 94.6 ;
      RECT  163.4 93.8 164.2 94.6 ;
      RECT  168.2 93.8 169.0 94.6 ;
      RECT  173.0 93.8 173.8 94.6 ;
      RECT  177.8 93.8 178.6 94.6 ;
      RECT  182.6 93.8 183.4 94.6 ;
      RECT  187.4 93.8 188.2 94.6 ;
      RECT  192.2 93.8 193.0 94.6 ;
      RECT  197.0 93.8 197.8 94.6 ;
      RECT  5.0 98.6 5.8 99.4 ;
      RECT  9.8 98.6 10.6 99.4 ;
      RECT  14.6 98.6 15.4 99.4 ;
      RECT  19.4 98.6 20.2 99.4 ;
      RECT  24.2 98.6 25.0 99.4 ;
      RECT  29.0 98.6 29.8 99.4 ;
      RECT  33.8 98.6 34.6 99.4 ;
      RECT  38.6 98.6 39.4 99.4 ;
      RECT  43.4 98.6 44.2 99.4 ;
      RECT  48.2 98.6 49.0 99.4 ;
      RECT  53.0 98.6 53.8 99.4 ;
      RECT  57.8 98.6 58.6 99.4 ;
      RECT  62.6 98.6 63.4 99.4 ;
      RECT  67.4 98.6 68.2 99.4 ;
      RECT  72.2 98.6 73.0 99.4 ;
      RECT  77.0 98.6 77.8 99.4 ;
      RECT  81.8 98.6 82.6 99.4 ;
      RECT  86.6 98.6 87.4 99.4 ;
      RECT  91.4 98.6 92.2 99.4 ;
      RECT  96.2 98.6 97.0 99.4 ;
      RECT  101.0 98.6 101.8 99.4 ;
      RECT  105.8 98.6 106.6 99.4 ;
      RECT  110.6 98.6 111.4 99.4 ;
      RECT  115.4 98.6 116.2 99.4 ;
      RECT  120.2 98.6 121.0 99.4 ;
      RECT  125.0 98.6 125.8 99.4 ;
      RECT  129.8 98.6 130.6 99.4 ;
      RECT  134.6 98.6 135.4 99.4 ;
      RECT  139.4 98.6 140.2 99.4 ;
      RECT  144.2 98.6 145.0 99.4 ;
      RECT  149.0 98.6 149.8 99.4 ;
      RECT  153.8 98.6 154.6 99.4 ;
      RECT  158.6 98.6 159.4 99.4 ;
      RECT  163.4 98.6 164.2 99.4 ;
      RECT  168.2 98.6 169.0 99.4 ;
      RECT  173.0 98.6 173.8 99.4 ;
      RECT  177.8 98.6 178.6 99.4 ;
      RECT  182.6 98.6 183.4 99.4 ;
      RECT  187.4 98.6 188.2 99.4 ;
      RECT  192.2 98.6 193.0 99.4 ;
      RECT  197.0 98.6 197.8 99.4 ;
      RECT  201.8 98.6 202.6 99.4 ;
      RECT  206.6 98.6 207.4 99.4 ;
      RECT  211.4 98.6 212.2 99.4 ;
      RECT  216.2 98.6 217.0 99.4 ;
      RECT  221.0 98.6 221.8 99.4 ;
      RECT  225.8 98.6 226.6 99.4 ;
      RECT  5.0 103.4 5.8 104.2 ;
      RECT  9.8 103.4 10.6 104.2 ;
      RECT  14.6 103.4 15.4 104.2 ;
      RECT  19.4 103.4 20.2 104.2 ;
      RECT  24.2 103.4 25.0 104.2 ;
      RECT  29.0 103.4 29.8 104.2 ;
      RECT  33.8 103.4 34.6 104.2 ;
      RECT  38.6 103.4 39.4 104.2 ;
      RECT  43.4 103.4 44.2 104.2 ;
      RECT  48.2 103.4 49.0 104.2 ;
      RECT  53.0 103.4 53.8 104.2 ;
      RECT  57.8 103.4 58.6 104.2 ;
      RECT  62.6 103.4 63.4 104.2 ;
      RECT  67.4 103.4 68.2 104.2 ;
      RECT  72.2 103.4 73.0 104.2 ;
      RECT  77.0 103.4 77.8 104.2 ;
      RECT  81.8 103.4 82.6 104.2 ;
      RECT  86.6 103.4 87.4 104.2 ;
      RECT  91.4 103.4 92.2 104.2 ;
      RECT  96.2 103.4 97.0 104.2 ;
      RECT  101.0 103.4 101.8 104.2 ;
      RECT  105.8 103.4 106.6 104.2 ;
      RECT  110.6 103.4 111.4 104.2 ;
      RECT  115.4 103.4 116.2 104.2 ;
      RECT  120.2 103.4 121.0 104.2 ;
      RECT  125.0 103.4 125.8 104.2 ;
      RECT  129.8 103.4 130.6 104.2 ;
      RECT  134.6 103.4 135.4 104.2 ;
      RECT  139.4 103.4 140.2 104.2 ;
      RECT  144.2 103.4 145.0 104.2 ;
      RECT  149.0 103.4 149.8 104.2 ;
      RECT  153.8 103.4 154.6 104.2 ;
      RECT  158.6 103.4 159.4 104.2 ;
      RECT  163.4 103.4 164.2 104.2 ;
      RECT  168.2 103.4 169.0 104.2 ;
      RECT  173.0 103.4 173.8 104.2 ;
      RECT  177.8 103.4 178.6 104.2 ;
      RECT  182.6 103.4 183.4 104.2 ;
      RECT  187.4 103.4 188.2 104.2 ;
      RECT  192.2 103.4 193.0 104.2 ;
      RECT  197.0 103.4 197.8 104.2 ;
      RECT  201.8 103.4 202.6 104.2 ;
      RECT  206.6 103.4 207.4 104.2 ;
      RECT  211.4 103.4 212.2 104.2 ;
      RECT  216.2 103.4 217.0 104.2 ;
      RECT  221.0 103.4 221.8 104.2 ;
      RECT  225.8 103.4 226.6 104.2 ;
      RECT  5.0 108.2 5.8 109.0 ;
      RECT  9.8 108.2 10.6 109.0 ;
      RECT  14.6 108.2 15.4 109.0 ;
      RECT  19.4 108.2 20.2 109.0 ;
      RECT  24.2 108.2 25.0 109.0 ;
      RECT  29.0 108.2 29.8 109.0 ;
      RECT  33.8 108.2 34.6 109.0 ;
      RECT  38.6 108.2 39.4 109.0 ;
      RECT  43.4 108.2 44.2 109.0 ;
      RECT  48.2 108.2 49.0 109.0 ;
      RECT  53.0 108.2 53.8 109.0 ;
      RECT  57.8 108.2 58.6 109.0 ;
      RECT  62.6 108.2 63.4 109.0 ;
      RECT  67.4 108.2 68.2 109.0 ;
      RECT  72.2 108.2 73.0 109.0 ;
      RECT  77.0 108.2 77.8 109.0 ;
      RECT  81.8 108.2 82.6 109.0 ;
      RECT  86.6 108.2 87.4 109.0 ;
      RECT  91.4 108.2 92.2 109.0 ;
      RECT  96.2 108.2 97.0 109.0 ;
      RECT  101.0 108.2 101.8 109.0 ;
      RECT  105.8 108.2 106.6 109.0 ;
      RECT  110.6 108.2 111.4 109.0 ;
      RECT  115.4 108.2 116.2 109.0 ;
      RECT  120.2 108.2 121.0 109.0 ;
      RECT  125.0 108.2 125.8 109.0 ;
      RECT  129.8 108.2 130.6 109.0 ;
      RECT  134.6 108.2 135.4 109.0 ;
      RECT  139.4 108.2 140.2 109.0 ;
      RECT  144.2 108.2 145.0 109.0 ;
      RECT  149.0 108.2 149.8 109.0 ;
      RECT  153.8 108.2 154.6 109.0 ;
      RECT  158.6 108.2 159.4 109.0 ;
      RECT  163.4 108.2 164.2 109.0 ;
      RECT  168.2 108.2 169.0 109.0 ;
      RECT  173.0 108.2 173.8 109.0 ;
      RECT  177.8 108.2 178.6 109.0 ;
      RECT  182.6 108.2 183.4 109.0 ;
      RECT  187.4 108.2 188.2 109.0 ;
      RECT  192.2 108.2 193.0 109.0 ;
      RECT  197.0 108.2 197.8 109.0 ;
      RECT  5.0 113.0 5.8 113.8 ;
      RECT  9.8 113.0 10.6 113.8 ;
      RECT  14.6 113.0 15.4 113.8 ;
      RECT  19.4 113.0 20.2 113.8 ;
      RECT  24.2 113.0 25.0 113.8 ;
      RECT  29.0 113.0 29.8 113.8 ;
      RECT  33.8 113.0 34.6 113.8 ;
      RECT  38.6 113.0 39.4 113.8 ;
      RECT  43.4 113.0 44.2 113.8 ;
      RECT  48.2 113.0 49.0 113.8 ;
      RECT  53.0 113.0 53.8 113.8 ;
      RECT  57.8 113.0 58.6 113.8 ;
      RECT  62.6 113.0 63.4 113.8 ;
      RECT  67.4 113.0 68.2 113.8 ;
      RECT  72.2 113.0 73.0 113.8 ;
      RECT  77.0 113.0 77.8 113.8 ;
      RECT  81.8 113.0 82.6 113.8 ;
      RECT  187.4 113.0 188.2 113.8 ;
      RECT  192.2 113.0 193.0 113.8 ;
      RECT  197.0 113.0 197.8 113.8 ;
      RECT  201.8 113.0 202.6 113.8 ;
      RECT  206.6 113.0 207.4 113.8 ;
      RECT  211.4 113.0 212.2 113.8 ;
      RECT  216.2 113.0 217.0 113.8 ;
      RECT  221.0 113.0 221.8 113.8 ;
      RECT  225.8 113.0 226.6 113.8 ;
      RECT  5.0 117.8 5.8 118.6 ;
      RECT  9.8 117.8 10.6 118.6 ;
      RECT  14.6 117.8 15.4 118.6 ;
      RECT  19.4 117.8 20.2 118.6 ;
      RECT  24.2 117.8 25.0 118.6 ;
      RECT  29.0 117.8 29.8 118.6 ;
      RECT  33.8 117.8 34.6 118.6 ;
      RECT  38.6 117.8 39.4 118.6 ;
      RECT  43.4 117.8 44.2 118.6 ;
      RECT  48.2 117.8 49.0 118.6 ;
      RECT  53.0 117.8 53.8 118.6 ;
      RECT  57.8 117.8 58.6 118.6 ;
      RECT  62.6 117.8 63.4 118.6 ;
      RECT  67.4 117.8 68.2 118.6 ;
      RECT  72.2 117.8 73.0 118.6 ;
      RECT  77.0 117.8 77.8 118.6 ;
      RECT  81.8 117.8 82.6 118.6 ;
      RECT  86.6 117.8 87.4 118.6 ;
      RECT  91.4 117.8 92.2 118.6 ;
      RECT  96.2 117.8 97.0 118.6 ;
      RECT  101.0 117.8 101.8 118.6 ;
      RECT  105.8 117.8 106.6 118.6 ;
      RECT  110.6 117.8 111.4 118.6 ;
      RECT  115.4 117.8 116.2 118.6 ;
      RECT  120.2 117.8 121.0 118.6 ;
      RECT  125.0 117.8 125.8 118.6 ;
      RECT  129.8 117.8 130.6 118.6 ;
      RECT  134.6 117.8 135.4 118.6 ;
      RECT  139.4 117.8 140.2 118.6 ;
      RECT  144.2 117.8 145.0 118.6 ;
      RECT  149.0 117.8 149.8 118.6 ;
      RECT  153.8 117.8 154.6 118.6 ;
      RECT  158.6 117.8 159.4 118.6 ;
      RECT  163.4 117.8 164.2 118.6 ;
      RECT  168.2 117.8 169.0 118.6 ;
      RECT  173.0 117.8 173.8 118.6 ;
      RECT  177.8 117.8 178.6 118.6 ;
      RECT  182.6 117.8 183.4 118.6 ;
      RECT  187.4 117.8 188.2 118.6 ;
      RECT  192.2 117.8 193.0 118.6 ;
      RECT  197.0 117.8 197.8 118.6 ;
      RECT  201.8 117.8 202.6 118.6 ;
      RECT  206.6 117.8 207.4 118.6 ;
      RECT  211.4 117.8 212.2 118.6 ;
      RECT  216.2 117.8 217.0 118.6 ;
      RECT  221.0 117.8 221.8 118.6 ;
      RECT  225.8 117.8 226.6 118.6 ;
      RECT  5.0 122.6 5.8 123.4 ;
      RECT  9.8 122.6 10.6 123.4 ;
      RECT  14.6 122.6 15.4 123.4 ;
      RECT  19.4 122.6 20.2 123.4 ;
      RECT  24.2 122.6 25.0 123.4 ;
      RECT  29.0 122.6 29.8 123.4 ;
      RECT  33.8 122.6 34.6 123.4 ;
      RECT  38.6 122.6 39.4 123.4 ;
      RECT  43.4 122.6 44.2 123.4 ;
      RECT  48.2 122.6 49.0 123.4 ;
      RECT  53.0 122.6 53.8 123.4 ;
      RECT  57.8 122.6 58.6 123.4 ;
      RECT  62.6 122.6 63.4 123.4 ;
      RECT  67.4 122.6 68.2 123.4 ;
      RECT  72.2 122.6 73.0 123.4 ;
      RECT  77.0 122.6 77.8 123.4 ;
      RECT  91.4 122.6 92.2 123.4 ;
      RECT  96.2 122.6 97.0 123.4 ;
      RECT  101.0 122.6 101.8 123.4 ;
      RECT  105.8 122.6 106.6 123.4 ;
      RECT  110.6 122.6 111.4 123.4 ;
      RECT  115.4 122.6 116.2 123.4 ;
      RECT  120.2 122.6 121.0 123.4 ;
      RECT  125.0 122.6 125.8 123.4 ;
      RECT  129.8 122.6 130.6 123.4 ;
      RECT  134.6 122.6 135.4 123.4 ;
      RECT  139.4 122.6 140.2 123.4 ;
      RECT  144.2 122.6 145.0 123.4 ;
      RECT  149.0 122.6 149.8 123.4 ;
      RECT  153.8 122.6 154.6 123.4 ;
      RECT  158.6 122.6 159.4 123.4 ;
      RECT  163.4 122.6 164.2 123.4 ;
      RECT  168.2 122.6 169.0 123.4 ;
      RECT  173.0 122.6 173.8 123.4 ;
      RECT  177.8 122.6 178.6 123.4 ;
      RECT  182.6 122.6 183.4 123.4 ;
      RECT  187.4 122.6 188.2 123.4 ;
      RECT  192.2 122.6 193.0 123.4 ;
      RECT  197.0 122.6 197.8 123.4 ;
      RECT  201.8 122.6 202.6 123.4 ;
      RECT  206.6 122.6 207.4 123.4 ;
      RECT  211.4 122.6 212.2 123.4 ;
      RECT  216.2 122.6 217.0 123.4 ;
      RECT  221.0 122.6 221.8 123.4 ;
      RECT  225.8 122.6 226.6 123.4 ;
      RECT  5.0 127.4 5.8 128.2 ;
      RECT  9.8 127.4 10.6 128.2 ;
      RECT  14.6 127.4 15.4 128.2 ;
      RECT  19.4 127.4 20.2 128.2 ;
      RECT  24.2 127.4 25.0 128.2 ;
      RECT  29.0 127.4 29.8 128.2 ;
      RECT  33.8 127.4 34.6 128.2 ;
      RECT  38.6 127.4 39.4 128.2 ;
      RECT  43.4 127.4 44.2 128.2 ;
      RECT  48.2 127.4 49.0 128.2 ;
      RECT  53.0 127.4 53.8 128.2 ;
      RECT  57.8 127.4 58.6 128.2 ;
      RECT  62.6 127.4 63.4 128.2 ;
      RECT  67.4 127.4 68.2 128.2 ;
      RECT  72.2 127.4 73.0 128.2 ;
      RECT  77.0 127.4 77.8 128.2 ;
      RECT  81.8 127.4 82.6 128.2 ;
      RECT  86.6 127.4 87.4 128.2 ;
      RECT  91.4 127.4 92.2 128.2 ;
      RECT  96.2 127.4 97.0 128.2 ;
      RECT  101.0 127.4 101.8 128.2 ;
      RECT  105.8 127.4 106.6 128.2 ;
      RECT  110.6 127.4 111.4 128.2 ;
      RECT  115.4 127.4 116.2 128.2 ;
      RECT  120.2 127.4 121.0 128.2 ;
      RECT  125.0 127.4 125.8 128.2 ;
      RECT  129.8 127.4 130.6 128.2 ;
      RECT  134.6 127.4 135.4 128.2 ;
      RECT  139.4 127.4 140.2 128.2 ;
      RECT  144.2 127.4 145.0 128.2 ;
      RECT  149.0 127.4 149.8 128.2 ;
      RECT  153.8 127.4 154.6 128.2 ;
      RECT  158.6 127.4 159.4 128.2 ;
      RECT  163.4 127.4 164.2 128.2 ;
      RECT  168.2 127.4 169.0 128.2 ;
      RECT  173.0 127.4 173.8 128.2 ;
      RECT  177.8 127.4 178.6 128.2 ;
      RECT  182.6 127.4 183.4 128.2 ;
      RECT  187.4 127.4 188.2 128.2 ;
      RECT  192.2 127.4 193.0 128.2 ;
      RECT  197.0 127.4 197.8 128.2 ;
      RECT  201.8 127.4 202.6 128.2 ;
      RECT  206.6 127.4 207.4 128.2 ;
      RECT  211.4 127.4 212.2 128.2 ;
      RECT  216.2 127.4 217.0 128.2 ;
      RECT  221.0 127.4 221.8 128.2 ;
      RECT  225.8 127.4 226.6 128.2 ;
      RECT  5.0 132.2 5.8 133.0 ;
      RECT  9.8 132.2 10.6 133.0 ;
      RECT  14.6 132.2 15.4 133.0 ;
      RECT  19.4 132.2 20.2 133.0 ;
      RECT  24.2 132.2 25.0 133.0 ;
      RECT  29.0 132.2 29.8 133.0 ;
      RECT  57.8 132.2 58.6 133.0 ;
      RECT  62.6 132.2 63.4 133.0 ;
      RECT  67.4 132.2 68.2 133.0 ;
      RECT  72.2 132.2 73.0 133.0 ;
      RECT  77.0 132.2 77.8 133.0 ;
      RECT  81.8 132.2 82.6 133.0 ;
      RECT  86.6 132.2 87.4 133.0 ;
      RECT  91.4 132.2 92.2 133.0 ;
      RECT  96.2 132.2 97.0 133.0 ;
      RECT  101.0 132.2 101.8 133.0 ;
      RECT  105.8 132.2 106.6 133.0 ;
      RECT  110.6 132.2 111.4 133.0 ;
      RECT  115.4 132.2 116.2 133.0 ;
      RECT  120.2 132.2 121.0 133.0 ;
      RECT  125.0 132.2 125.8 133.0 ;
      RECT  129.8 132.2 130.6 133.0 ;
      RECT  134.6 132.2 135.4 133.0 ;
      RECT  139.4 132.2 140.2 133.0 ;
      RECT  144.2 132.2 145.0 133.0 ;
      RECT  149.0 132.2 149.8 133.0 ;
      RECT  153.8 132.2 154.6 133.0 ;
      RECT  158.6 132.2 159.4 133.0 ;
      RECT  163.4 132.2 164.2 133.0 ;
      RECT  168.2 132.2 169.0 133.0 ;
      RECT  173.0 132.2 173.8 133.0 ;
      RECT  177.8 132.2 178.6 133.0 ;
      RECT  182.6 132.2 183.4 133.0 ;
      RECT  187.4 132.2 188.2 133.0 ;
      RECT  192.2 132.2 193.0 133.0 ;
      RECT  197.0 132.2 197.8 133.0 ;
      RECT  201.8 132.2 202.6 133.0 ;
      RECT  206.6 132.2 207.4 133.0 ;
      RECT  211.4 132.2 212.2 133.0 ;
      RECT  216.2 132.2 217.0 133.0 ;
      RECT  221.0 132.2 221.8 133.0 ;
      RECT  225.8 132.2 226.6 133.0 ;
      RECT  5.0 137.0 5.8 137.8 ;
      RECT  9.8 137.0 10.6 137.8 ;
      RECT  14.6 137.0 15.4 137.8 ;
      RECT  19.4 137.0 20.2 137.8 ;
      RECT  24.2 137.0 25.0 137.8 ;
      RECT  29.0 137.0 29.8 137.8 ;
      RECT  33.8 137.0 34.6 137.8 ;
      RECT  38.6 137.0 39.4 137.8 ;
      RECT  43.4 137.0 44.2 137.8 ;
      RECT  48.2 137.0 49.0 137.8 ;
      RECT  53.0 137.0 53.8 137.8 ;
      RECT  57.8 137.0 58.6 137.8 ;
      RECT  62.6 137.0 63.4 137.8 ;
      RECT  67.4 137.0 68.2 137.8 ;
      RECT  72.2 137.0 73.0 137.8 ;
      RECT  77.0 137.0 77.8 137.8 ;
      RECT  81.8 137.0 82.6 137.8 ;
      RECT  86.6 137.0 87.4 137.8 ;
      RECT  91.4 137.0 92.2 137.8 ;
      RECT  96.2 137.0 97.0 137.8 ;
      RECT  101.0 137.0 101.8 137.8 ;
      RECT  105.8 137.0 106.6 137.8 ;
      RECT  110.6 137.0 111.4 137.8 ;
      RECT  115.4 137.0 116.2 137.8 ;
      RECT  120.2 137.0 121.0 137.8 ;
      RECT  125.0 137.0 125.8 137.8 ;
      RECT  129.8 137.0 130.6 137.8 ;
      RECT  134.6 137.0 135.4 137.8 ;
      RECT  139.4 137.0 140.2 137.8 ;
      RECT  144.2 137.0 145.0 137.8 ;
      RECT  149.0 137.0 149.8 137.8 ;
      RECT  153.8 137.0 154.6 137.8 ;
      RECT  158.6 137.0 159.4 137.8 ;
      RECT  163.4 137.0 164.2 137.8 ;
      RECT  168.2 137.0 169.0 137.8 ;
      RECT  173.0 137.0 173.8 137.8 ;
      RECT  177.8 137.0 178.6 137.8 ;
      RECT  182.6 137.0 183.4 137.8 ;
      RECT  187.4 137.0 188.2 137.8 ;
      RECT  192.2 137.0 193.0 137.8 ;
      RECT  197.0 137.0 197.8 137.8 ;
      RECT  201.8 137.0 202.6 137.8 ;
      RECT  206.6 137.0 207.4 137.8 ;
      RECT  211.4 137.0 212.2 137.8 ;
      RECT  216.2 137.0 217.0 137.8 ;
      RECT  221.0 137.0 221.8 137.8 ;
      RECT  225.8 137.0 226.6 137.8 ;
      RECT  5.0 141.8 5.8 142.6 ;
      RECT  9.8 141.8 10.6 142.6 ;
      RECT  14.6 141.8 15.4 142.6 ;
      RECT  19.4 141.8 20.2 142.6 ;
      RECT  24.2 141.8 25.0 142.6 ;
      RECT  29.0 141.8 29.8 142.6 ;
      RECT  33.8 141.8 34.6 142.6 ;
      RECT  38.6 141.8 39.4 142.6 ;
      RECT  43.4 141.8 44.2 142.6 ;
      RECT  48.2 141.8 49.0 142.6 ;
      RECT  53.0 141.8 53.8 142.6 ;
      RECT  57.8 141.8 58.6 142.6 ;
      RECT  62.6 141.8 63.4 142.6 ;
      RECT  67.4 141.8 68.2 142.6 ;
      RECT  72.2 141.8 73.0 142.6 ;
      RECT  77.0 141.8 77.8 142.6 ;
      RECT  81.8 141.8 82.6 142.6 ;
      RECT  86.6 141.8 87.4 142.6 ;
      RECT  91.4 141.8 92.2 142.6 ;
      RECT  96.2 141.8 97.0 142.6 ;
      RECT  101.0 141.8 101.8 142.6 ;
      RECT  105.8 141.8 106.6 142.6 ;
      RECT  110.6 141.8 111.4 142.6 ;
      RECT  115.4 141.8 116.2 142.6 ;
      RECT  120.2 141.8 121.0 142.6 ;
      RECT  125.0 141.8 125.8 142.6 ;
      RECT  129.8 141.8 130.6 142.6 ;
      RECT  134.6 141.8 135.4 142.6 ;
      RECT  139.4 141.8 140.2 142.6 ;
      RECT  144.2 141.8 145.0 142.6 ;
      RECT  149.0 141.8 149.8 142.6 ;
      RECT  153.8 141.8 154.6 142.6 ;
      RECT  158.6 141.8 159.4 142.6 ;
      RECT  163.4 141.8 164.2 142.6 ;
      RECT  168.2 141.8 169.0 142.6 ;
      RECT  173.0 141.8 173.8 142.6 ;
      RECT  177.8 141.8 178.6 142.6 ;
      RECT  182.6 141.8 183.4 142.6 ;
      RECT  187.4 141.8 188.2 142.6 ;
      RECT  192.2 141.8 193.0 142.6 ;
      RECT  197.0 141.8 197.8 142.6 ;
      RECT  201.8 141.8 202.6 142.6 ;
      RECT  206.6 141.8 207.4 142.6 ;
      RECT  211.4 141.8 212.2 142.6 ;
      RECT  216.2 141.8 217.0 142.6 ;
      RECT  221.0 141.8 221.8 142.6 ;
      RECT  225.8 141.8 226.6 142.6 ;
      RECT  5.0 146.6 5.8 147.4 ;
      RECT  9.8 146.6 10.6 147.4 ;
      RECT  14.6 146.6 15.4 147.4 ;
      RECT  19.4 146.6 20.2 147.4 ;
      RECT  24.2 146.6 25.0 147.4 ;
      RECT  29.0 146.6 29.8 147.4 ;
      RECT  33.8 146.6 34.6 147.4 ;
      RECT  38.6 146.6 39.4 147.4 ;
      RECT  43.4 146.6 44.2 147.4 ;
      RECT  48.2 146.6 49.0 147.4 ;
      RECT  53.0 146.6 53.8 147.4 ;
      RECT  57.8 146.6 58.6 147.4 ;
      RECT  62.6 146.6 63.4 147.4 ;
      RECT  67.4 146.6 68.2 147.4 ;
      RECT  72.2 146.6 73.0 147.4 ;
      RECT  77.0 146.6 77.8 147.4 ;
      RECT  81.8 146.6 82.6 147.4 ;
      RECT  86.6 146.6 87.4 147.4 ;
      RECT  91.4 146.6 92.2 147.4 ;
      RECT  96.2 146.6 97.0 147.4 ;
      RECT  101.0 146.6 101.8 147.4 ;
      RECT  105.8 146.6 106.6 147.4 ;
      RECT  110.6 146.6 111.4 147.4 ;
      RECT  115.4 146.6 116.2 147.4 ;
      RECT  120.2 146.6 121.0 147.4 ;
      RECT  125.0 146.6 125.8 147.4 ;
      RECT  129.8 146.6 130.6 147.4 ;
      RECT  134.6 146.6 135.4 147.4 ;
      RECT  139.4 146.6 140.2 147.4 ;
      RECT  144.2 146.6 145.0 147.4 ;
      RECT  149.0 146.6 149.8 147.4 ;
      RECT  153.8 146.6 154.6 147.4 ;
      RECT  158.6 146.6 159.4 147.4 ;
      RECT  163.4 146.6 164.2 147.4 ;
      RECT  168.2 146.6 169.0 147.4 ;
      RECT  173.0 146.6 173.8 147.4 ;
      RECT  177.8 146.6 178.6 147.4 ;
      RECT  182.6 146.6 183.4 147.4 ;
      RECT  187.4 146.6 188.2 147.4 ;
      RECT  192.2 146.6 193.0 147.4 ;
      RECT  197.0 146.6 197.8 147.4 ;
      RECT  5.0 151.4 5.8 152.2 ;
      RECT  9.8 151.4 10.6 152.2 ;
      RECT  14.6 151.4 15.4 152.2 ;
      RECT  19.4 151.4 20.2 152.2 ;
      RECT  24.2 151.4 25.0 152.2 ;
      RECT  29.0 151.4 29.8 152.2 ;
      RECT  33.8 151.4 34.6 152.2 ;
      RECT  38.6 151.4 39.4 152.2 ;
      RECT  43.4 151.4 44.2 152.2 ;
      RECT  48.2 151.4 49.0 152.2 ;
      RECT  53.0 151.4 53.8 152.2 ;
      RECT  57.8 151.4 58.6 152.2 ;
      RECT  62.6 151.4 63.4 152.2 ;
      RECT  67.4 151.4 68.2 152.2 ;
      RECT  72.2 151.4 73.0 152.2 ;
      RECT  77.0 151.4 77.8 152.2 ;
      RECT  81.8 151.4 82.6 152.2 ;
      RECT  187.4 151.4 188.2 152.2 ;
      RECT  192.2 151.4 193.0 152.2 ;
      RECT  197.0 151.4 197.8 152.2 ;
      RECT  201.8 151.4 202.6 152.2 ;
      RECT  206.6 151.4 207.4 152.2 ;
      RECT  211.4 151.4 212.2 152.2 ;
      RECT  216.2 151.4 217.0 152.2 ;
      RECT  221.0 151.4 221.8 152.2 ;
      RECT  225.8 151.4 226.6 152.2 ;
      RECT  5.0 156.2 5.8 157.0 ;
      RECT  9.8 156.2 10.6 157.0 ;
      RECT  14.6 156.2 15.4 157.0 ;
      RECT  19.4 156.2 20.2 157.0 ;
      RECT  24.2 156.2 25.0 157.0 ;
      RECT  29.0 156.2 29.8 157.0 ;
      RECT  33.8 156.2 34.6 157.0 ;
      RECT  38.6 156.2 39.4 157.0 ;
      RECT  43.4 156.2 44.2 157.0 ;
      RECT  48.2 156.2 49.0 157.0 ;
      RECT  53.0 156.2 53.8 157.0 ;
      RECT  57.8 156.2 58.6 157.0 ;
      RECT  62.6 156.2 63.4 157.0 ;
      RECT  67.4 156.2 68.2 157.0 ;
      RECT  72.2 156.2 73.0 157.0 ;
      RECT  77.0 156.2 77.8 157.0 ;
      RECT  81.8 156.2 82.6 157.0 ;
      RECT  86.6 156.2 87.4 157.0 ;
      RECT  91.4 156.2 92.2 157.0 ;
      RECT  96.2 156.2 97.0 157.0 ;
      RECT  101.0 156.2 101.8 157.0 ;
      RECT  105.8 156.2 106.6 157.0 ;
      RECT  110.6 156.2 111.4 157.0 ;
      RECT  115.4 156.2 116.2 157.0 ;
      RECT  120.2 156.2 121.0 157.0 ;
      RECT  125.0 156.2 125.8 157.0 ;
      RECT  129.8 156.2 130.6 157.0 ;
      RECT  134.6 156.2 135.4 157.0 ;
      RECT  139.4 156.2 140.2 157.0 ;
      RECT  144.2 156.2 145.0 157.0 ;
      RECT  149.0 156.2 149.8 157.0 ;
      RECT  153.8 156.2 154.6 157.0 ;
      RECT  158.6 156.2 159.4 157.0 ;
      RECT  163.4 156.2 164.2 157.0 ;
      RECT  168.2 156.2 169.0 157.0 ;
      RECT  173.0 156.2 173.8 157.0 ;
      RECT  177.8 156.2 178.6 157.0 ;
      RECT  182.6 156.2 183.4 157.0 ;
      RECT  187.4 156.2 188.2 157.0 ;
      RECT  192.2 156.2 193.0 157.0 ;
      RECT  197.0 156.2 197.8 157.0 ;
      RECT  201.8 156.2 202.6 157.0 ;
      RECT  206.6 156.2 207.4 157.0 ;
      RECT  211.4 156.2 212.2 157.0 ;
      RECT  216.2 156.2 217.0 157.0 ;
      RECT  221.0 156.2 221.8 157.0 ;
      RECT  225.8 156.2 226.6 157.0 ;
      RECT  5.0 161.0 5.8 161.8 ;
      RECT  9.8 161.0 10.6 161.8 ;
      RECT  14.6 161.0 15.4 161.8 ;
      RECT  19.4 161.0 20.2 161.8 ;
      RECT  24.2 161.0 25.0 161.8 ;
      RECT  29.0 161.0 29.8 161.8 ;
      RECT  33.8 161.0 34.6 161.8 ;
      RECT  38.6 161.0 39.4 161.8 ;
      RECT  43.4 161.0 44.2 161.8 ;
      RECT  48.2 161.0 49.0 161.8 ;
      RECT  53.0 161.0 53.8 161.8 ;
      RECT  57.8 161.0 58.6 161.8 ;
      RECT  62.6 161.0 63.4 161.8 ;
      RECT  67.4 161.0 68.2 161.8 ;
      RECT  72.2 161.0 73.0 161.8 ;
      RECT  77.0 161.0 77.8 161.8 ;
      RECT  91.4 161.0 92.2 161.8 ;
      RECT  96.2 161.0 97.0 161.8 ;
      RECT  101.0 161.0 101.8 161.8 ;
      RECT  105.8 161.0 106.6 161.8 ;
      RECT  110.6 161.0 111.4 161.8 ;
      RECT  115.4 161.0 116.2 161.8 ;
      RECT  120.2 161.0 121.0 161.8 ;
      RECT  125.0 161.0 125.8 161.8 ;
      RECT  129.8 161.0 130.6 161.8 ;
      RECT  134.6 161.0 135.4 161.8 ;
      RECT  139.4 161.0 140.2 161.8 ;
      RECT  144.2 161.0 145.0 161.8 ;
      RECT  149.0 161.0 149.8 161.8 ;
      RECT  153.8 161.0 154.6 161.8 ;
      RECT  158.6 161.0 159.4 161.8 ;
      RECT  163.4 161.0 164.2 161.8 ;
      RECT  168.2 161.0 169.0 161.8 ;
      RECT  173.0 161.0 173.8 161.8 ;
      RECT  177.8 161.0 178.6 161.8 ;
      RECT  182.6 161.0 183.4 161.8 ;
      RECT  187.4 161.0 188.2 161.8 ;
      RECT  192.2 161.0 193.0 161.8 ;
      RECT  197.0 161.0 197.8 161.8 ;
      RECT  201.8 161.0 202.6 161.8 ;
      RECT  206.6 161.0 207.4 161.8 ;
      RECT  211.4 161.0 212.2 161.8 ;
      RECT  216.2 161.0 217.0 161.8 ;
      RECT  221.0 161.0 221.8 161.8 ;
      RECT  225.8 161.0 226.6 161.8 ;
      RECT  201.8 165.8 202.6 166.6 ;
      RECT  206.6 165.8 207.4 166.6 ;
      RECT  211.4 165.8 212.2 166.6 ;
      RECT  216.2 165.8 217.0 166.6 ;
      RECT  221.0 165.8 221.8 166.6 ;
      RECT  225.8 165.8 226.6 166.6 ;
      RECT  33.8 170.6 34.6 171.4 ;
      RECT  38.6 170.6 39.4 171.4 ;
      RECT  43.4 170.6 44.2 171.4 ;
      RECT  48.2 170.6 49.0 171.4 ;
      RECT  53.0 170.6 53.8 171.4 ;
      RECT  57.8 170.6 58.6 171.4 ;
      RECT  62.6 170.6 63.4 171.4 ;
      RECT  67.4 170.6 68.2 171.4 ;
      RECT  72.2 170.6 73.0 171.4 ;
      RECT  77.0 170.6 77.8 171.4 ;
      RECT  81.8 170.6 82.6 171.4 ;
      RECT  86.6 170.6 87.4 171.4 ;
      RECT  91.4 170.6 92.2 171.4 ;
      RECT  96.2 170.6 97.0 171.4 ;
      RECT  101.0 170.6 101.8 171.4 ;
      RECT  105.8 170.6 106.6 171.4 ;
      RECT  110.6 170.6 111.4 171.4 ;
      RECT  115.4 170.6 116.2 171.4 ;
      RECT  120.2 170.6 121.0 171.4 ;
      RECT  125.0 170.6 125.8 171.4 ;
      RECT  129.8 170.6 130.6 171.4 ;
      RECT  134.6 170.6 135.4 171.4 ;
      RECT  139.4 170.6 140.2 171.4 ;
      RECT  144.2 170.6 145.0 171.4 ;
      RECT  149.0 170.6 149.8 171.4 ;
      RECT  153.8 170.6 154.6 171.4 ;
      RECT  158.6 170.6 159.4 171.4 ;
      RECT  163.4 170.6 164.2 171.4 ;
      RECT  168.2 170.6 169.0 171.4 ;
      RECT  173.0 170.6 173.8 171.4 ;
      RECT  177.8 170.6 178.6 171.4 ;
      RECT  182.6 170.6 183.4 171.4 ;
      RECT  187.4 170.6 188.2 171.4 ;
      RECT  192.2 170.6 193.0 171.4 ;
      RECT  197.0 170.6 197.8 171.4 ;
      RECT  201.8 170.6 202.6 171.4 ;
      RECT  206.6 170.6 207.4 171.4 ;
      RECT  211.4 170.6 212.2 171.4 ;
      RECT  216.2 170.6 217.0 171.4 ;
      RECT  221.0 170.6 221.8 171.4 ;
      RECT  225.8 170.6 226.6 171.4 ;
      RECT  5.0 175.4 5.8 176.2 ;
      RECT  9.8 175.4 10.6 176.2 ;
      RECT  14.6 175.4 15.4 176.2 ;
      RECT  19.4 175.4 20.2 176.2 ;
      RECT  24.2 175.4 25.0 176.2 ;
      RECT  29.0 175.4 29.8 176.2 ;
      RECT  33.8 175.4 34.6 176.2 ;
      RECT  38.6 175.4 39.4 176.2 ;
      RECT  43.4 175.4 44.2 176.2 ;
      RECT  48.2 175.4 49.0 176.2 ;
      RECT  53.0 175.4 53.8 176.2 ;
      RECT  57.8 175.4 58.6 176.2 ;
      RECT  62.6 175.4 63.4 176.2 ;
      RECT  67.4 175.4 68.2 176.2 ;
      RECT  72.2 175.4 73.0 176.2 ;
      RECT  77.0 175.4 77.8 176.2 ;
      RECT  81.8 175.4 82.6 176.2 ;
      RECT  86.6 175.4 87.4 176.2 ;
      RECT  91.4 175.4 92.2 176.2 ;
      RECT  96.2 175.4 97.0 176.2 ;
      RECT  101.0 175.4 101.8 176.2 ;
      RECT  105.8 175.4 106.6 176.2 ;
      RECT  110.6 175.4 111.4 176.2 ;
      RECT  115.4 175.4 116.2 176.2 ;
      RECT  120.2 175.4 121.0 176.2 ;
      RECT  125.0 175.4 125.8 176.2 ;
      RECT  129.8 175.4 130.6 176.2 ;
      RECT  134.6 175.4 135.4 176.2 ;
      RECT  139.4 175.4 140.2 176.2 ;
      RECT  144.2 175.4 145.0 176.2 ;
      RECT  149.0 175.4 149.8 176.2 ;
      RECT  153.8 175.4 154.6 176.2 ;
      RECT  158.6 175.4 159.4 176.2 ;
      RECT  163.4 175.4 164.2 176.2 ;
      RECT  168.2 175.4 169.0 176.2 ;
      RECT  173.0 175.4 173.8 176.2 ;
      RECT  177.8 175.4 178.6 176.2 ;
      RECT  182.6 175.4 183.4 176.2 ;
      RECT  187.4 175.4 188.2 176.2 ;
      RECT  192.2 175.4 193.0 176.2 ;
      RECT  197.0 175.4 197.8 176.2 ;
      RECT  201.8 175.4 202.6 176.2 ;
      RECT  206.6 175.4 207.4 176.2 ;
      RECT  211.4 175.4 212.2 176.2 ;
      RECT  216.2 175.4 217.0 176.2 ;
      RECT  221.0 175.4 221.8 176.2 ;
      RECT  225.8 175.4 226.6 176.2 ;
      RECT  33.8 180.2 34.6 181.0 ;
      RECT  38.6 180.2 39.4 181.0 ;
      RECT  43.4 180.2 44.2 181.0 ;
      RECT  48.2 180.2 49.0 181.0 ;
      RECT  53.0 180.2 53.8 181.0 ;
      RECT  57.8 180.2 58.6 181.0 ;
      RECT  62.6 180.2 63.4 181.0 ;
      RECT  67.4 180.2 68.2 181.0 ;
      RECT  72.2 180.2 73.0 181.0 ;
      RECT  77.0 180.2 77.8 181.0 ;
      RECT  81.8 180.2 82.6 181.0 ;
      RECT  86.6 180.2 87.4 181.0 ;
      RECT  91.4 180.2 92.2 181.0 ;
      RECT  96.2 180.2 97.0 181.0 ;
      RECT  101.0 180.2 101.8 181.0 ;
      RECT  105.8 180.2 106.6 181.0 ;
      RECT  110.6 180.2 111.4 181.0 ;
      RECT  115.4 180.2 116.2 181.0 ;
      RECT  120.2 180.2 121.0 181.0 ;
      RECT  125.0 180.2 125.8 181.0 ;
      RECT  129.8 180.2 130.6 181.0 ;
      RECT  134.6 180.2 135.4 181.0 ;
      RECT  139.4 180.2 140.2 181.0 ;
      RECT  144.2 180.2 145.0 181.0 ;
      RECT  149.0 180.2 149.8 181.0 ;
      RECT  153.8 180.2 154.6 181.0 ;
      RECT  158.6 180.2 159.4 181.0 ;
      RECT  163.4 180.2 164.2 181.0 ;
      RECT  168.2 180.2 169.0 181.0 ;
      RECT  173.0 180.2 173.8 181.0 ;
      RECT  177.8 180.2 178.6 181.0 ;
      RECT  24.2 185.0 25.0 185.8 ;
      RECT  29.0 185.0 29.8 185.8 ;
      RECT  33.8 185.0 34.6 185.8 ;
      RECT  38.6 185.0 39.4 185.8 ;
      RECT  43.4 185.0 44.2 185.8 ;
      RECT  48.2 185.0 49.0 185.8 ;
      RECT  53.0 185.0 53.8 185.8 ;
      RECT  57.8 185.0 58.6 185.8 ;
      RECT  62.6 185.0 63.4 185.8 ;
      RECT  67.4 185.0 68.2 185.8 ;
      RECT  72.2 185.0 73.0 185.8 ;
      RECT  77.0 185.0 77.8 185.8 ;
      RECT  81.8 185.0 82.6 185.8 ;
      RECT  86.6 185.0 87.4 185.8 ;
      RECT  91.4 185.0 92.2 185.8 ;
      RECT  96.2 185.0 97.0 185.8 ;
      RECT  101.0 185.0 101.8 185.8 ;
      RECT  105.8 185.0 106.6 185.8 ;
      RECT  110.6 185.0 111.4 185.8 ;
      RECT  115.4 185.0 116.2 185.8 ;
      RECT  120.2 185.0 121.0 185.8 ;
      RECT  125.0 185.0 125.8 185.8 ;
      RECT  129.8 185.0 130.6 185.8 ;
      RECT  134.6 185.0 135.4 185.8 ;
      RECT  139.4 185.0 140.2 185.8 ;
      RECT  144.2 185.0 145.0 185.8 ;
      RECT  149.0 185.0 149.8 185.8 ;
      RECT  153.8 185.0 154.6 185.8 ;
      RECT  158.6 185.0 159.4 185.8 ;
      RECT  163.4 185.0 164.2 185.8 ;
      RECT  168.2 185.0 169.0 185.8 ;
      RECT  173.0 185.0 173.8 185.8 ;
      RECT  177.8 185.0 178.6 185.8 ;
      RECT  182.6 185.0 183.4 185.8 ;
      RECT  187.4 185.0 188.2 185.8 ;
      RECT  192.2 185.0 193.0 185.8 ;
      RECT  197.0 185.0 197.8 185.8 ;
      RECT  201.8 185.0 202.6 185.8 ;
      RECT  206.6 185.0 207.4 185.8 ;
      RECT  211.4 185.0 212.2 185.8 ;
      RECT  216.2 185.0 217.0 185.8 ;
      RECT  221.0 185.0 221.8 185.8 ;
      RECT  225.8 185.0 226.6 185.8 ;
      RECT  33.8 189.8 34.6 190.6 ;
      RECT  38.6 189.8 39.4 190.6 ;
      RECT  43.4 189.8 44.2 190.6 ;
      RECT  48.2 189.8 49.0 190.6 ;
      RECT  53.0 189.8 53.8 190.6 ;
      RECT  57.8 189.8 58.6 190.6 ;
      RECT  62.6 189.8 63.4 190.6 ;
      RECT  67.4 189.8 68.2 190.6 ;
      RECT  72.2 189.8 73.0 190.6 ;
      RECT  77.0 189.8 77.8 190.6 ;
      RECT  81.8 189.8 82.6 190.6 ;
      RECT  86.6 189.8 87.4 190.6 ;
      RECT  91.4 189.8 92.2 190.6 ;
      RECT  96.2 189.8 97.0 190.6 ;
      RECT  101.0 189.8 101.8 190.6 ;
      RECT  105.8 189.8 106.6 190.6 ;
      RECT  110.6 189.8 111.4 190.6 ;
      RECT  115.4 189.8 116.2 190.6 ;
      RECT  120.2 189.8 121.0 190.6 ;
      RECT  125.0 189.8 125.8 190.6 ;
      RECT  129.8 189.8 130.6 190.6 ;
      RECT  134.6 189.8 135.4 190.6 ;
      RECT  139.4 189.8 140.2 190.6 ;
      RECT  144.2 189.8 145.0 190.6 ;
      RECT  149.0 189.8 149.8 190.6 ;
      RECT  153.8 189.8 154.6 190.6 ;
      RECT  158.6 189.8 159.4 190.6 ;
      RECT  163.4 189.8 164.2 190.6 ;
      RECT  168.2 189.8 169.0 190.6 ;
      RECT  173.0 189.8 173.8 190.6 ;
      RECT  177.8 189.8 178.6 190.6 ;
      RECT  5.0 194.6 5.8 195.4 ;
      RECT  9.8 194.6 10.6 195.4 ;
      RECT  14.6 194.6 15.4 195.4 ;
      RECT  19.4 194.6 20.2 195.4 ;
      RECT  24.2 194.6 25.0 195.4 ;
      RECT  29.0 194.6 29.8 195.4 ;
      RECT  33.8 194.6 34.6 195.4 ;
      RECT  38.6 194.6 39.4 195.4 ;
      RECT  43.4 194.6 44.2 195.4 ;
      RECT  48.2 194.6 49.0 195.4 ;
      RECT  53.0 194.6 53.8 195.4 ;
      RECT  57.8 194.6 58.6 195.4 ;
      RECT  62.6 194.6 63.4 195.4 ;
      RECT  67.4 194.6 68.2 195.4 ;
      RECT  72.2 194.6 73.0 195.4 ;
      RECT  77.0 194.6 77.8 195.4 ;
      RECT  81.8 194.6 82.6 195.4 ;
      RECT  86.6 194.6 87.4 195.4 ;
      RECT  91.4 194.6 92.2 195.4 ;
      RECT  96.2 194.6 97.0 195.4 ;
      RECT  177.8 194.6 178.6 195.4 ;
      RECT  182.6 194.6 183.4 195.4 ;
      RECT  187.4 194.6 188.2 195.4 ;
      RECT  192.2 194.6 193.0 195.4 ;
      RECT  197.0 194.6 197.8 195.4 ;
      RECT  201.8 194.6 202.6 195.4 ;
      RECT  206.6 194.6 207.4 195.4 ;
      RECT  211.4 194.6 212.2 195.4 ;
      RECT  216.2 194.6 217.0 195.4 ;
      RECT  221.0 194.6 221.8 195.4 ;
      RECT  225.8 194.6 226.6 195.4 ;
      RECT  33.8 199.4 34.6 200.2 ;
      RECT  38.6 199.4 39.4 200.2 ;
      RECT  43.4 199.4 44.2 200.2 ;
      RECT  48.2 199.4 49.0 200.2 ;
      RECT  53.0 199.4 53.8 200.2 ;
      RECT  57.8 199.4 58.6 200.2 ;
      RECT  62.6 199.4 63.4 200.2 ;
      RECT  67.4 199.4 68.2 200.2 ;
      RECT  72.2 199.4 73.0 200.2 ;
      RECT  77.0 199.4 77.8 200.2 ;
      RECT  81.8 199.4 82.6 200.2 ;
      RECT  86.6 199.4 87.4 200.2 ;
      RECT  91.4 199.4 92.2 200.2 ;
      RECT  96.2 199.4 97.0 200.2 ;
      RECT  101.0 199.4 101.8 200.2 ;
      RECT  105.8 199.4 106.6 200.2 ;
      RECT  110.6 199.4 111.4 200.2 ;
      RECT  115.4 199.4 116.2 200.2 ;
      RECT  120.2 199.4 121.0 200.2 ;
      RECT  125.0 199.4 125.8 200.2 ;
      RECT  129.8 199.4 130.6 200.2 ;
      RECT  134.6 199.4 135.4 200.2 ;
      RECT  139.4 199.4 140.2 200.2 ;
      RECT  144.2 199.4 145.0 200.2 ;
      RECT  149.0 199.4 149.8 200.2 ;
      RECT  153.8 199.4 154.6 200.2 ;
      RECT  158.6 199.4 159.4 200.2 ;
      RECT  163.4 199.4 164.2 200.2 ;
      RECT  168.2 199.4 169.0 200.2 ;
      RECT  173.0 199.4 173.8 200.2 ;
      RECT  177.8 199.4 178.6 200.2 ;
      RECT  24.2 204.2 25.0 205.0 ;
      RECT  29.0 204.2 29.8 205.0 ;
      RECT  33.8 204.2 34.6 205.0 ;
      RECT  38.6 204.2 39.4 205.0 ;
      RECT  43.4 204.2 44.2 205.0 ;
      RECT  48.2 204.2 49.0 205.0 ;
      RECT  53.0 204.2 53.8 205.0 ;
      RECT  57.8 204.2 58.6 205.0 ;
      RECT  62.6 204.2 63.4 205.0 ;
      RECT  67.4 204.2 68.2 205.0 ;
      RECT  72.2 204.2 73.0 205.0 ;
      RECT  77.0 204.2 77.8 205.0 ;
      RECT  81.8 204.2 82.6 205.0 ;
      RECT  139.4 204.2 140.2 205.0 ;
      RECT  144.2 204.2 145.0 205.0 ;
      RECT  149.0 204.2 149.8 205.0 ;
      RECT  153.8 204.2 154.6 205.0 ;
      RECT  158.6 204.2 159.4 205.0 ;
      RECT  163.4 204.2 164.2 205.0 ;
      RECT  168.2 204.2 169.0 205.0 ;
      RECT  173.0 204.2 173.8 205.0 ;
      RECT  177.8 204.2 178.6 205.0 ;
      RECT  182.6 204.2 183.4 205.0 ;
      RECT  187.4 204.2 188.2 205.0 ;
      RECT  192.2 204.2 193.0 205.0 ;
      RECT  197.0 204.2 197.8 205.0 ;
      RECT  201.8 204.2 202.6 205.0 ;
      RECT  206.6 204.2 207.4 205.0 ;
      RECT  211.4 204.2 212.2 205.0 ;
      RECT  216.2 204.2 217.0 205.0 ;
      RECT  221.0 204.2 221.8 205.0 ;
      RECT  225.8 204.2 226.6 205.0 ;
      RECT  5.0 209.0 5.8 209.8 ;
      RECT  9.8 209.0 10.6 209.8 ;
      RECT  14.6 209.0 15.4 209.8 ;
      RECT  19.4 209.0 20.2 209.8 ;
      RECT  24.2 209.0 25.0 209.8 ;
      RECT  29.0 209.0 29.8 209.8 ;
      RECT  33.8 209.0 34.6 209.8 ;
      RECT  38.6 209.0 39.4 209.8 ;
      RECT  43.4 209.0 44.2 209.8 ;
      RECT  48.2 209.0 49.0 209.8 ;
      RECT  53.0 209.0 53.8 209.8 ;
      RECT  57.8 209.0 58.6 209.8 ;
      RECT  62.6 209.0 63.4 209.8 ;
      RECT  67.4 209.0 68.2 209.8 ;
      RECT  72.2 209.0 73.0 209.8 ;
      RECT  77.0 209.0 77.8 209.8 ;
      RECT  81.8 209.0 82.6 209.8 ;
      RECT  86.6 209.0 87.4 209.8 ;
      RECT  91.4 209.0 92.2 209.8 ;
      RECT  96.2 209.0 97.0 209.8 ;
      RECT  101.0 209.0 101.8 209.8 ;
      RECT  105.8 209.0 106.6 209.8 ;
      RECT  110.6 209.0 111.4 209.8 ;
      RECT  115.4 209.0 116.2 209.8 ;
      RECT  120.2 209.0 121.0 209.8 ;
      RECT  125.0 209.0 125.8 209.8 ;
      RECT  129.8 209.0 130.6 209.8 ;
      RECT  134.6 209.0 135.4 209.8 ;
      RECT  139.4 209.0 140.2 209.8 ;
      RECT  144.2 209.0 145.0 209.8 ;
      RECT  149.0 209.0 149.8 209.8 ;
      RECT  153.8 209.0 154.6 209.8 ;
      RECT  158.6 209.0 159.4 209.8 ;
      RECT  163.4 209.0 164.2 209.8 ;
      RECT  168.2 209.0 169.0 209.8 ;
      RECT  173.0 209.0 173.8 209.8 ;
      RECT  177.8 209.0 178.6 209.8 ;
      RECT  5.0 213.8 5.8 214.6 ;
      RECT  9.8 213.8 10.6 214.6 ;
      RECT  14.6 213.8 15.4 214.6 ;
      RECT  19.4 213.8 20.2 214.6 ;
      RECT  24.2 213.8 25.0 214.6 ;
      RECT  29.0 213.8 29.8 214.6 ;
      RECT  33.8 213.8 34.6 214.6 ;
      RECT  38.6 213.8 39.4 214.6 ;
      RECT  43.4 213.8 44.2 214.6 ;
      RECT  48.2 213.8 49.0 214.6 ;
      RECT  53.0 213.8 53.8 214.6 ;
      RECT  57.8 213.8 58.6 214.6 ;
      RECT  62.6 213.8 63.4 214.6 ;
      RECT  67.4 213.8 68.2 214.6 ;
      RECT  72.2 213.8 73.0 214.6 ;
      RECT  77.0 213.8 77.8 214.6 ;
      RECT  81.8 213.8 82.6 214.6 ;
      RECT  86.6 213.8 87.4 214.6 ;
      RECT  91.4 213.8 92.2 214.6 ;
      RECT  96.2 213.8 97.0 214.6 ;
      RECT  177.8 213.8 178.6 214.6 ;
      RECT  182.6 213.8 183.4 214.6 ;
      RECT  187.4 213.8 188.2 214.6 ;
      RECT  192.2 213.8 193.0 214.6 ;
      RECT  197.0 213.8 197.8 214.6 ;
      RECT  201.8 213.8 202.6 214.6 ;
      RECT  206.6 213.8 207.4 214.6 ;
      RECT  211.4 213.8 212.2 214.6 ;
      RECT  216.2 213.8 217.0 214.6 ;
      RECT  221.0 213.8 221.8 214.6 ;
      RECT  225.8 213.8 226.6 214.6 ;
      RECT  5.0 218.6 5.8 219.4 ;
      RECT  9.8 218.6 10.6 219.4 ;
      RECT  14.6 218.6 15.4 219.4 ;
      RECT  19.4 218.6 20.2 219.4 ;
      RECT  24.2 218.6 25.0 219.4 ;
      RECT  29.0 218.6 29.8 219.4 ;
      RECT  33.8 218.6 34.6 219.4 ;
      RECT  38.6 218.6 39.4 219.4 ;
      RECT  43.4 218.6 44.2 219.4 ;
      RECT  48.2 218.6 49.0 219.4 ;
      RECT  53.0 218.6 53.8 219.4 ;
      RECT  57.8 218.6 58.6 219.4 ;
      RECT  62.6 218.6 63.4 219.4 ;
      RECT  67.4 218.6 68.2 219.4 ;
      RECT  72.2 218.6 73.0 219.4 ;
      RECT  77.0 218.6 77.8 219.4 ;
      RECT  81.8 218.6 82.6 219.4 ;
      RECT  86.6 218.6 87.4 219.4 ;
      RECT  91.4 218.6 92.2 219.4 ;
      RECT  96.2 218.6 97.0 219.4 ;
      RECT  101.0 218.6 101.8 219.4 ;
      RECT  105.8 218.6 106.6 219.4 ;
      RECT  110.6 218.6 111.4 219.4 ;
      RECT  115.4 218.6 116.2 219.4 ;
      RECT  120.2 218.6 121.0 219.4 ;
      RECT  125.0 218.6 125.8 219.4 ;
      RECT  129.8 218.6 130.6 219.4 ;
      RECT  134.6 218.6 135.4 219.4 ;
      RECT  139.4 218.6 140.2 219.4 ;
      RECT  144.2 218.6 145.0 219.4 ;
      RECT  149.0 218.6 149.8 219.4 ;
      RECT  153.8 218.6 154.6 219.4 ;
      RECT  158.6 218.6 159.4 219.4 ;
      RECT  163.4 218.6 164.2 219.4 ;
      RECT  168.2 218.6 169.0 219.4 ;
      RECT  173.0 218.6 173.8 219.4 ;
      RECT  177.8 218.6 178.6 219.4 ;
      RECT  33.8 223.4 34.6 224.2 ;
      RECT  38.6 223.4 39.4 224.2 ;
      RECT  43.4 223.4 44.2 224.2 ;
      RECT  48.2 223.4 49.0 224.2 ;
      RECT  53.0 223.4 53.8 224.2 ;
      RECT  57.8 223.4 58.6 224.2 ;
      RECT  62.6 223.4 63.4 224.2 ;
      RECT  67.4 223.4 68.2 224.2 ;
      RECT  72.2 223.4 73.0 224.2 ;
      RECT  77.0 223.4 77.8 224.2 ;
      RECT  81.8 223.4 82.6 224.2 ;
      RECT  86.6 223.4 87.4 224.2 ;
      RECT  91.4 223.4 92.2 224.2 ;
      RECT  96.2 223.4 97.0 224.2 ;
      RECT  101.0 223.4 101.8 224.2 ;
      RECT  105.8 223.4 106.6 224.2 ;
      RECT  110.6 223.4 111.4 224.2 ;
      RECT  115.4 223.4 116.2 224.2 ;
      RECT  120.2 223.4 121.0 224.2 ;
      RECT  139.4 223.4 140.2 224.2 ;
      RECT  144.2 223.4 145.0 224.2 ;
      RECT  149.0 223.4 149.8 224.2 ;
      RECT  153.8 223.4 154.6 224.2 ;
      RECT  158.6 223.4 159.4 224.2 ;
      RECT  163.4 223.4 164.2 224.2 ;
      RECT  168.2 223.4 169.0 224.2 ;
      RECT  173.0 223.4 173.8 224.2 ;
      RECT  177.8 223.4 178.6 224.2 ;
      RECT  182.6 223.4 183.4 224.2 ;
      RECT  187.4 223.4 188.2 224.2 ;
      RECT  192.2 223.4 193.0 224.2 ;
      RECT  197.0 223.4 197.8 224.2 ;
      RECT  201.8 223.4 202.6 224.2 ;
      RECT  206.6 223.4 207.4 224.2 ;
      RECT  211.4 223.4 212.2 224.2 ;
      RECT  216.2 223.4 217.0 224.2 ;
      RECT  221.0 223.4 221.8 224.2 ;
      RECT  225.8 223.4 226.6 224.2 ;
      RECT  24.2 228.2 25.0 229.0 ;
      RECT  29.0 228.2 29.8 229.0 ;
      RECT  33.8 228.2 34.6 229.0 ;
      RECT  38.6 228.2 39.4 229.0 ;
      RECT  43.4 228.2 44.2 229.0 ;
      RECT  48.2 228.2 49.0 229.0 ;
      RECT  53.0 228.2 53.8 229.0 ;
      RECT  57.8 228.2 58.6 229.0 ;
      RECT  62.6 228.2 63.4 229.0 ;
      RECT  67.4 228.2 68.2 229.0 ;
      RECT  72.2 228.2 73.0 229.0 ;
      RECT  77.0 228.2 77.8 229.0 ;
      RECT  81.8 228.2 82.6 229.0 ;
      RECT  86.6 228.2 87.4 229.0 ;
      RECT  91.4 228.2 92.2 229.0 ;
      RECT  96.2 228.2 97.0 229.0 ;
      RECT  101.0 228.2 101.8 229.0 ;
      RECT  105.8 228.2 106.6 229.0 ;
      RECT  110.6 228.2 111.4 229.0 ;
      RECT  115.4 228.2 116.2 229.0 ;
      RECT  120.2 228.2 121.0 229.0 ;
      RECT  125.0 228.2 125.8 229.0 ;
      RECT  129.8 228.2 130.6 229.0 ;
      RECT  134.6 228.2 135.4 229.0 ;
      RECT  139.4 228.2 140.2 229.0 ;
      RECT  144.2 228.2 145.0 229.0 ;
      RECT  149.0 228.2 149.8 229.0 ;
      RECT  153.8 228.2 154.6 229.0 ;
      RECT  158.6 228.2 159.4 229.0 ;
      RECT  163.4 228.2 164.2 229.0 ;
      RECT  168.2 228.2 169.0 229.0 ;
      RECT  173.0 228.2 173.8 229.0 ;
      RECT  177.8 228.2 178.6 229.0 ;
      RECT  33.8 233.0 34.6 233.8 ;
      RECT  38.6 233.0 39.4 233.8 ;
      RECT  43.4 233.0 44.2 233.8 ;
      RECT  48.2 233.0 49.0 233.8 ;
      RECT  53.0 233.0 53.8 233.8 ;
      RECT  57.8 233.0 58.6 233.8 ;
      RECT  62.6 233.0 63.4 233.8 ;
      RECT  67.4 233.0 68.2 233.8 ;
      RECT  72.2 233.0 73.0 233.8 ;
      RECT  77.0 233.0 77.8 233.8 ;
      RECT  81.8 233.0 82.6 233.8 ;
      RECT  86.6 233.0 87.4 233.8 ;
      RECT  91.4 233.0 92.2 233.8 ;
      RECT  96.2 233.0 97.0 233.8 ;
      RECT  101.0 233.0 101.8 233.8 ;
      RECT  105.8 233.0 106.6 233.8 ;
      RECT  110.6 233.0 111.4 233.8 ;
      RECT  115.4 233.0 116.2 233.8 ;
      RECT  120.2 233.0 121.0 233.8 ;
      RECT  125.0 233.0 125.8 233.8 ;
      RECT  129.8 233.0 130.6 233.8 ;
      RECT  134.6 233.0 135.4 233.8 ;
      RECT  139.4 233.0 140.2 233.8 ;
      RECT  144.2 233.0 145.0 233.8 ;
      RECT  149.0 233.0 149.8 233.8 ;
      RECT  153.8 233.0 154.6 233.8 ;
      RECT  158.6 233.0 159.4 233.8 ;
      RECT  163.4 233.0 164.2 233.8 ;
      RECT  168.2 233.0 169.0 233.8 ;
      RECT  173.0 233.0 173.8 233.8 ;
      RECT  177.8 233.0 178.6 233.8 ;
      RECT  182.6 233.0 183.4 233.8 ;
      RECT  187.4 233.0 188.2 233.8 ;
      RECT  192.2 233.0 193.0 233.8 ;
      RECT  197.0 233.0 197.8 233.8 ;
      RECT  201.8 233.0 202.6 233.8 ;
      RECT  206.6 233.0 207.4 233.8 ;
      RECT  211.4 233.0 212.2 233.8 ;
      RECT  216.2 233.0 217.0 233.8 ;
      RECT  221.0 233.0 221.8 233.8 ;
      RECT  225.8 233.0 226.6 233.8 ;
      RECT  5.0 237.8 5.8 238.6 ;
      RECT  9.8 237.8 10.6 238.6 ;
      RECT  14.6 237.8 15.4 238.6 ;
      RECT  19.4 237.8 20.2 238.6 ;
      RECT  24.2 237.8 25.0 238.6 ;
      RECT  29.0 237.8 29.8 238.6 ;
      RECT  33.8 237.8 34.6 238.6 ;
      RECT  38.6 237.8 39.4 238.6 ;
      RECT  43.4 237.8 44.2 238.6 ;
      RECT  48.2 237.8 49.0 238.6 ;
      RECT  53.0 237.8 53.8 238.6 ;
      RECT  57.8 237.8 58.6 238.6 ;
      RECT  62.6 237.8 63.4 238.6 ;
      RECT  67.4 237.8 68.2 238.6 ;
      RECT  72.2 237.8 73.0 238.6 ;
      RECT  77.0 237.8 77.8 238.6 ;
      RECT  81.8 237.8 82.6 238.6 ;
      RECT  86.6 237.8 87.4 238.6 ;
      RECT  91.4 237.8 92.2 238.6 ;
      RECT  96.2 237.8 97.0 238.6 ;
      RECT  177.8 237.8 178.6 238.6 ;
      RECT  182.6 237.8 183.4 238.6 ;
      RECT  187.4 237.8 188.2 238.6 ;
      RECT  192.2 237.8 193.0 238.6 ;
      RECT  197.0 237.8 197.8 238.6 ;
      RECT  201.8 237.8 202.6 238.6 ;
      RECT  206.6 237.8 207.4 238.6 ;
      RECT  211.4 237.8 212.2 238.6 ;
      RECT  216.2 237.8 217.0 238.6 ;
      RECT  221.0 237.8 221.8 238.6 ;
      RECT  225.8 237.8 226.6 238.6 ;
      RECT  33.8 242.6 34.6 243.4 ;
      RECT  38.6 242.6 39.4 243.4 ;
      RECT  43.4 242.6 44.2 243.4 ;
      RECT  48.2 242.6 49.0 243.4 ;
      RECT  53.0 242.6 53.8 243.4 ;
      RECT  57.8 242.6 58.6 243.4 ;
      RECT  62.6 242.6 63.4 243.4 ;
      RECT  67.4 242.6 68.2 243.4 ;
      RECT  72.2 242.6 73.0 243.4 ;
      RECT  77.0 242.6 77.8 243.4 ;
      RECT  81.8 242.6 82.6 243.4 ;
      RECT  86.6 242.6 87.4 243.4 ;
      RECT  91.4 242.6 92.2 243.4 ;
      RECT  96.2 242.6 97.0 243.4 ;
      RECT  101.0 242.6 101.8 243.4 ;
      RECT  105.8 242.6 106.6 243.4 ;
      RECT  110.6 242.6 111.4 243.4 ;
      RECT  115.4 242.6 116.2 243.4 ;
      RECT  120.2 242.6 121.0 243.4 ;
      RECT  125.0 242.6 125.8 243.4 ;
      RECT  129.8 242.6 130.6 243.4 ;
      RECT  134.6 242.6 135.4 243.4 ;
      RECT  139.4 242.6 140.2 243.4 ;
      RECT  144.2 242.6 145.0 243.4 ;
      RECT  149.0 242.6 149.8 243.4 ;
      RECT  153.8 242.6 154.6 243.4 ;
      RECT  158.6 242.6 159.4 243.4 ;
      RECT  163.4 242.6 164.2 243.4 ;
      RECT  168.2 242.6 169.0 243.4 ;
      RECT  173.0 242.6 173.8 243.4 ;
      RECT  177.8 242.6 178.6 243.4 ;
      RECT  24.2 247.4 25.0 248.2 ;
      RECT  29.0 247.4 29.8 248.2 ;
      RECT  33.8 247.4 34.6 248.2 ;
      RECT  38.6 247.4 39.4 248.2 ;
      RECT  43.4 247.4 44.2 248.2 ;
      RECT  48.2 247.4 49.0 248.2 ;
      RECT  53.0 247.4 53.8 248.2 ;
      RECT  57.8 247.4 58.6 248.2 ;
      RECT  62.6 247.4 63.4 248.2 ;
      RECT  67.4 247.4 68.2 248.2 ;
      RECT  72.2 247.4 73.0 248.2 ;
      RECT  77.0 247.4 77.8 248.2 ;
      RECT  81.8 247.4 82.6 248.2 ;
      RECT  86.6 247.4 87.4 248.2 ;
      RECT  144.2 247.4 145.0 248.2 ;
      RECT  149.0 247.4 149.8 248.2 ;
      RECT  153.8 247.4 154.6 248.2 ;
      RECT  158.6 247.4 159.4 248.2 ;
      RECT  163.4 247.4 164.2 248.2 ;
      RECT  168.2 247.4 169.0 248.2 ;
      RECT  173.0 247.4 173.8 248.2 ;
      RECT  177.8 247.4 178.6 248.2 ;
      RECT  182.6 247.4 183.4 248.2 ;
      RECT  187.4 247.4 188.2 248.2 ;
      RECT  192.2 247.4 193.0 248.2 ;
      RECT  197.0 247.4 197.8 248.2 ;
      RECT  201.8 247.4 202.6 248.2 ;
      RECT  206.6 247.4 207.4 248.2 ;
      RECT  211.4 247.4 212.2 248.2 ;
      RECT  216.2 247.4 217.0 248.2 ;
      RECT  221.0 247.4 221.8 248.2 ;
      RECT  225.8 247.4 226.6 248.2 ;
      RECT  33.8 252.2 34.6 253.0 ;
      RECT  38.6 252.2 39.4 253.0 ;
      RECT  43.4 252.2 44.2 253.0 ;
      RECT  48.2 252.2 49.0 253.0 ;
      RECT  53.0 252.2 53.8 253.0 ;
      RECT  57.8 252.2 58.6 253.0 ;
      RECT  62.6 252.2 63.4 253.0 ;
      RECT  67.4 252.2 68.2 253.0 ;
      RECT  72.2 252.2 73.0 253.0 ;
      RECT  77.0 252.2 77.8 253.0 ;
      RECT  81.8 252.2 82.6 253.0 ;
      RECT  86.6 252.2 87.4 253.0 ;
      RECT  91.4 252.2 92.2 253.0 ;
      RECT  96.2 252.2 97.0 253.0 ;
      RECT  101.0 252.2 101.8 253.0 ;
      RECT  105.8 252.2 106.6 253.0 ;
      RECT  110.6 252.2 111.4 253.0 ;
      RECT  115.4 252.2 116.2 253.0 ;
      RECT  120.2 252.2 121.0 253.0 ;
      RECT  125.0 252.2 125.8 253.0 ;
      RECT  129.8 252.2 130.6 253.0 ;
      RECT  134.6 252.2 135.4 253.0 ;
      RECT  139.4 252.2 140.2 253.0 ;
      RECT  144.2 252.2 145.0 253.0 ;
      RECT  149.0 252.2 149.8 253.0 ;
      RECT  153.8 252.2 154.6 253.0 ;
      RECT  158.6 252.2 159.4 253.0 ;
      RECT  163.4 252.2 164.2 253.0 ;
      RECT  168.2 252.2 169.0 253.0 ;
      RECT  173.0 252.2 173.8 253.0 ;
      RECT  177.8 252.2 178.6 253.0 ;
      RECT  5.0 257.0 5.8 257.8 ;
      RECT  9.8 257.0 10.6 257.8 ;
      RECT  14.6 257.0 15.4 257.8 ;
      RECT  19.4 257.0 20.2 257.8 ;
      RECT  24.2 257.0 25.0 257.8 ;
      RECT  29.0 257.0 29.8 257.8 ;
      RECT  33.8 257.0 34.6 257.8 ;
      RECT  38.6 257.0 39.4 257.8 ;
      RECT  43.4 257.0 44.2 257.8 ;
      RECT  48.2 257.0 49.0 257.8 ;
      RECT  53.0 257.0 53.8 257.8 ;
      RECT  57.8 257.0 58.6 257.8 ;
      RECT  62.6 257.0 63.4 257.8 ;
      RECT  67.4 257.0 68.2 257.8 ;
      RECT  72.2 257.0 73.0 257.8 ;
      RECT  77.0 257.0 77.8 257.8 ;
      RECT  81.8 257.0 82.6 257.8 ;
      RECT  86.6 257.0 87.4 257.8 ;
      RECT  177.8 257.0 178.6 257.8 ;
      RECT  182.6 257.0 183.4 257.8 ;
      RECT  187.4 257.0 188.2 257.8 ;
      RECT  192.2 257.0 193.0 257.8 ;
      RECT  197.0 257.0 197.8 257.8 ;
      RECT  201.8 257.0 202.6 257.8 ;
      RECT  206.6 257.0 207.4 257.8 ;
      RECT  211.4 257.0 212.2 257.8 ;
      RECT  216.2 257.0 217.0 257.8 ;
      RECT  221.0 257.0 221.8 257.8 ;
      RECT  225.8 257.0 226.6 257.8 ;
      RECT  5.0 261.8 5.8 262.6 ;
      RECT  9.8 261.8 10.6 262.6 ;
      RECT  14.6 261.8 15.4 262.6 ;
      RECT  19.4 261.8 20.2 262.6 ;
      RECT  24.2 261.8 25.0 262.6 ;
      RECT  29.0 261.8 29.8 262.6 ;
      RECT  33.8 261.8 34.6 262.6 ;
      RECT  38.6 261.8 39.4 262.6 ;
      RECT  43.4 261.8 44.2 262.6 ;
      RECT  48.2 261.8 49.0 262.6 ;
      RECT  53.0 261.8 53.8 262.6 ;
      RECT  57.8 261.8 58.6 262.6 ;
      RECT  62.6 261.8 63.4 262.6 ;
      RECT  67.4 261.8 68.2 262.6 ;
      RECT  72.2 261.8 73.0 262.6 ;
      RECT  77.0 261.8 77.8 262.6 ;
      RECT  81.8 261.8 82.6 262.6 ;
      RECT  86.6 261.8 87.4 262.6 ;
      RECT  91.4 261.8 92.2 262.6 ;
      RECT  96.2 261.8 97.0 262.6 ;
      RECT  101.0 261.8 101.8 262.6 ;
      RECT  105.8 261.8 106.6 262.6 ;
      RECT  110.6 261.8 111.4 262.6 ;
      RECT  115.4 261.8 116.2 262.6 ;
      RECT  120.2 261.8 121.0 262.6 ;
      RECT  125.0 261.8 125.8 262.6 ;
      RECT  129.8 261.8 130.6 262.6 ;
      RECT  134.6 261.8 135.4 262.6 ;
      RECT  139.4 261.8 140.2 262.6 ;
      RECT  144.2 261.8 145.0 262.6 ;
      RECT  149.0 261.8 149.8 262.6 ;
      RECT  153.8 261.8 154.6 262.6 ;
      RECT  158.6 261.8 159.4 262.6 ;
      RECT  163.4 261.8 164.2 262.6 ;
      RECT  168.2 261.8 169.0 262.6 ;
      RECT  173.0 261.8 173.8 262.6 ;
      RECT  177.8 261.8 178.6 262.6 ;
      RECT  5.0 266.6 5.8 267.4 ;
      RECT  9.8 266.6 10.6 267.4 ;
      RECT  14.6 266.6 15.4 267.4 ;
      RECT  19.4 266.6 20.2 267.4 ;
      RECT  24.2 266.6 25.0 267.4 ;
      RECT  29.0 266.6 29.8 267.4 ;
      RECT  33.8 266.6 34.6 267.4 ;
      RECT  38.6 266.6 39.4 267.4 ;
      RECT  43.4 266.6 44.2 267.4 ;
      RECT  48.2 266.6 49.0 267.4 ;
      RECT  53.0 266.6 53.8 267.4 ;
      RECT  57.8 266.6 58.6 267.4 ;
      RECT  62.6 266.6 63.4 267.4 ;
      RECT  67.4 266.6 68.2 267.4 ;
      RECT  72.2 266.6 73.0 267.4 ;
      RECT  77.0 266.6 77.8 267.4 ;
      RECT  81.8 266.6 82.6 267.4 ;
      RECT  86.6 266.6 87.4 267.4 ;
      RECT  91.4 266.6 92.2 267.4 ;
      RECT  96.2 266.6 97.0 267.4 ;
      RECT  101.0 266.6 101.8 267.4 ;
      RECT  105.8 266.6 106.6 267.4 ;
      RECT  110.6 266.6 111.4 267.4 ;
      RECT  115.4 266.6 116.2 267.4 ;
      RECT  120.2 266.6 121.0 267.4 ;
      RECT  144.2 266.6 145.0 267.4 ;
      RECT  149.0 266.6 149.8 267.4 ;
      RECT  153.8 266.6 154.6 267.4 ;
      RECT  158.6 266.6 159.4 267.4 ;
      RECT  163.4 266.6 164.2 267.4 ;
      RECT  168.2 266.6 169.0 267.4 ;
      RECT  173.0 266.6 173.8 267.4 ;
      RECT  177.8 266.6 178.6 267.4 ;
      RECT  182.6 266.6 183.4 267.4 ;
      RECT  187.4 266.6 188.2 267.4 ;
      RECT  192.2 266.6 193.0 267.4 ;
      RECT  197.0 266.6 197.8 267.4 ;
      RECT  201.8 266.6 202.6 267.4 ;
      RECT  206.6 266.6 207.4 267.4 ;
      RECT  211.4 266.6 212.2 267.4 ;
      RECT  216.2 266.6 217.0 267.4 ;
      RECT  221.0 266.6 221.8 267.4 ;
      RECT  225.8 266.6 226.6 267.4 ;
      RECT  5.0 271.4 5.8 272.2 ;
      RECT  9.8 271.4 10.6 272.2 ;
      RECT  14.6 271.4 15.4 272.2 ;
      RECT  19.4 271.4 20.2 272.2 ;
      RECT  24.2 271.4 25.0 272.2 ;
      RECT  29.0 271.4 29.8 272.2 ;
      RECT  33.8 271.4 34.6 272.2 ;
      RECT  38.6 271.4 39.4 272.2 ;
      RECT  43.4 271.4 44.2 272.2 ;
      RECT  48.2 271.4 49.0 272.2 ;
      RECT  53.0 271.4 53.8 272.2 ;
      RECT  57.8 271.4 58.6 272.2 ;
      RECT  62.6 271.4 63.4 272.2 ;
      RECT  67.4 271.4 68.2 272.2 ;
      RECT  72.2 271.4 73.0 272.2 ;
      RECT  77.0 271.4 77.8 272.2 ;
      RECT  81.8 271.4 82.6 272.2 ;
      RECT  86.6 271.4 87.4 272.2 ;
      RECT  91.4 271.4 92.2 272.2 ;
      RECT  96.2 271.4 97.0 272.2 ;
      RECT  101.0 271.4 101.8 272.2 ;
      RECT  105.8 271.4 106.6 272.2 ;
      RECT  110.6 271.4 111.4 272.2 ;
      RECT  115.4 271.4 116.2 272.2 ;
      RECT  120.2 271.4 121.0 272.2 ;
      RECT  125.0 271.4 125.8 272.2 ;
      RECT  129.8 271.4 130.6 272.2 ;
      RECT  134.6 271.4 135.4 272.2 ;
      RECT  139.4 271.4 140.2 272.2 ;
      RECT  144.2 271.4 145.0 272.2 ;
      RECT  149.0 271.4 149.8 272.2 ;
      RECT  153.8 271.4 154.6 272.2 ;
      RECT  158.6 271.4 159.4 272.2 ;
      RECT  163.4 271.4 164.2 272.2 ;
      RECT  168.2 271.4 169.0 272.2 ;
      RECT  173.0 271.4 173.8 272.2 ;
      RECT  177.8 271.4 178.6 272.2 ;
      RECT  5.0 276.2 5.8 277.0 ;
      RECT  9.8 276.2 10.6 277.0 ;
      RECT  14.6 276.2 15.4 277.0 ;
      RECT  19.4 276.2 20.2 277.0 ;
      RECT  24.2 276.2 25.0 277.0 ;
      RECT  29.0 276.2 29.8 277.0 ;
      RECT  33.8 276.2 34.6 277.0 ;
      RECT  38.6 276.2 39.4 277.0 ;
      RECT  43.4 276.2 44.2 277.0 ;
      RECT  48.2 276.2 49.0 277.0 ;
      RECT  53.0 276.2 53.8 277.0 ;
      RECT  57.8 276.2 58.6 277.0 ;
      RECT  62.6 276.2 63.4 277.0 ;
      RECT  67.4 276.2 68.2 277.0 ;
      RECT  72.2 276.2 73.0 277.0 ;
      RECT  77.0 276.2 77.8 277.0 ;
      RECT  81.8 276.2 82.6 277.0 ;
      RECT  86.6 276.2 87.4 277.0 ;
      RECT  91.4 276.2 92.2 277.0 ;
      RECT  96.2 276.2 97.0 277.0 ;
      RECT  177.8 276.2 178.6 277.0 ;
      RECT  182.6 276.2 183.4 277.0 ;
      RECT  187.4 276.2 188.2 277.0 ;
      RECT  192.2 276.2 193.0 277.0 ;
      RECT  197.0 276.2 197.8 277.0 ;
      RECT  201.8 276.2 202.6 277.0 ;
      RECT  206.6 276.2 207.4 277.0 ;
      RECT  211.4 276.2 212.2 277.0 ;
      RECT  216.2 276.2 217.0 277.0 ;
      RECT  221.0 276.2 221.8 277.0 ;
      RECT  225.8 276.2 226.6 277.0 ;
      RECT  5.0 281.0 5.8 281.8 ;
      RECT  9.8 281.0 10.6 281.8 ;
      RECT  14.6 281.0 15.4 281.8 ;
      RECT  19.4 281.0 20.2 281.8 ;
      RECT  24.2 281.0 25.0 281.8 ;
      RECT  29.0 281.0 29.8 281.8 ;
      RECT  33.8 281.0 34.6 281.8 ;
      RECT  38.6 281.0 39.4 281.8 ;
      RECT  43.4 281.0 44.2 281.8 ;
      RECT  48.2 281.0 49.0 281.8 ;
      RECT  53.0 281.0 53.8 281.8 ;
      RECT  57.8 281.0 58.6 281.8 ;
      RECT  62.6 281.0 63.4 281.8 ;
      RECT  67.4 281.0 68.2 281.8 ;
      RECT  72.2 281.0 73.0 281.8 ;
      RECT  77.0 281.0 77.8 281.8 ;
      RECT  81.8 281.0 82.6 281.8 ;
      RECT  86.6 281.0 87.4 281.8 ;
      RECT  91.4 281.0 92.2 281.8 ;
      RECT  96.2 281.0 97.0 281.8 ;
      RECT  101.0 281.0 101.8 281.8 ;
      RECT  105.8 281.0 106.6 281.8 ;
      RECT  110.6 281.0 111.4 281.8 ;
      RECT  115.4 281.0 116.2 281.8 ;
      RECT  120.2 281.0 121.0 281.8 ;
      RECT  125.0 281.0 125.8 281.8 ;
      RECT  129.8 281.0 130.6 281.8 ;
      RECT  134.6 281.0 135.4 281.8 ;
      RECT  139.4 281.0 140.2 281.8 ;
      RECT  144.2 281.0 145.0 281.8 ;
      RECT  149.0 281.0 149.8 281.8 ;
      RECT  153.8 281.0 154.6 281.8 ;
      RECT  158.6 281.0 159.4 281.8 ;
      RECT  163.4 281.0 164.2 281.8 ;
      RECT  168.2 281.0 169.0 281.8 ;
      RECT  173.0 281.0 173.8 281.8 ;
      RECT  177.8 281.0 178.6 281.8 ;
      RECT  5.0 285.8 5.8 286.6 ;
      RECT  9.8 285.8 10.6 286.6 ;
      RECT  14.6 285.8 15.4 286.6 ;
      RECT  19.4 285.8 20.2 286.6 ;
      RECT  24.2 285.8 25.0 286.6 ;
      RECT  29.0 285.8 29.8 286.6 ;
      RECT  33.8 285.8 34.6 286.6 ;
      RECT  38.6 285.8 39.4 286.6 ;
      RECT  43.4 285.8 44.2 286.6 ;
      RECT  48.2 285.8 49.0 286.6 ;
      RECT  53.0 285.8 53.8 286.6 ;
      RECT  57.8 285.8 58.6 286.6 ;
      RECT  62.6 285.8 63.4 286.6 ;
      RECT  67.4 285.8 68.2 286.6 ;
      RECT  72.2 285.8 73.0 286.6 ;
      RECT  77.0 285.8 77.8 286.6 ;
      RECT  81.8 285.8 82.6 286.6 ;
      RECT  86.6 285.8 87.4 286.6 ;
      RECT  91.4 285.8 92.2 286.6 ;
      RECT  96.2 285.8 97.0 286.6 ;
      RECT  101.0 285.8 101.8 286.6 ;
      RECT  105.8 285.8 106.6 286.6 ;
      RECT  110.6 285.8 111.4 286.6 ;
      RECT  115.4 285.8 116.2 286.6 ;
      RECT  120.2 285.8 121.0 286.6 ;
      RECT  125.0 285.8 125.8 286.6 ;
      RECT  129.8 285.8 130.6 286.6 ;
      RECT  134.6 285.8 135.4 286.6 ;
      RECT  139.4 285.8 140.2 286.6 ;
      RECT  144.2 285.8 145.0 286.6 ;
      RECT  149.0 285.8 149.8 286.6 ;
      RECT  153.8 285.8 154.6 286.6 ;
      RECT  158.6 285.8 159.4 286.6 ;
      RECT  163.4 285.8 164.2 286.6 ;
      RECT  168.2 285.8 169.0 286.6 ;
      RECT  173.0 285.8 173.8 286.6 ;
      RECT  177.8 285.8 178.6 286.6 ;
      RECT  182.6 285.8 183.4 286.6 ;
      RECT  187.4 285.8 188.2 286.6 ;
      RECT  192.2 285.8 193.0 286.6 ;
      RECT  197.0 285.8 197.8 286.6 ;
      RECT  201.8 285.8 202.6 286.6 ;
      RECT  206.6 285.8 207.4 286.6 ;
      RECT  211.4 285.8 212.2 286.6 ;
      RECT  216.2 285.8 217.0 286.6 ;
      RECT  221.0 285.8 221.8 286.6 ;
      RECT  225.8 285.8 226.6 286.6 ;
      RECT  5.0 290.6 5.8 291.4 ;
      RECT  9.8 290.6 10.6 291.4 ;
      RECT  14.6 290.6 15.4 291.4 ;
      RECT  19.4 290.6 20.2 291.4 ;
      RECT  24.2 290.6 25.0 291.4 ;
      RECT  29.0 290.6 29.8 291.4 ;
      RECT  33.8 290.6 34.6 291.4 ;
      RECT  38.6 290.6 39.4 291.4 ;
      RECT  43.4 290.6 44.2 291.4 ;
      RECT  48.2 290.6 49.0 291.4 ;
      RECT  53.0 290.6 53.8 291.4 ;
      RECT  57.8 290.6 58.6 291.4 ;
      RECT  62.6 290.6 63.4 291.4 ;
      RECT  67.4 290.6 68.2 291.4 ;
      RECT  81.8 290.6 82.6 291.4 ;
      RECT  86.6 290.6 87.4 291.4 ;
      RECT  91.4 290.6 92.2 291.4 ;
      RECT  96.2 290.6 97.0 291.4 ;
      RECT  101.0 290.6 101.8 291.4 ;
      RECT  105.8 290.6 106.6 291.4 ;
      RECT  110.6 290.6 111.4 291.4 ;
      RECT  115.4 290.6 116.2 291.4 ;
      RECT  120.2 290.6 121.0 291.4 ;
      RECT  125.0 290.6 125.8 291.4 ;
      RECT  129.8 290.6 130.6 291.4 ;
      RECT  134.6 290.6 135.4 291.4 ;
      RECT  139.4 290.6 140.2 291.4 ;
      RECT  144.2 290.6 145.0 291.4 ;
      RECT  149.0 290.6 149.8 291.4 ;
      RECT  153.8 290.6 154.6 291.4 ;
      RECT  158.6 290.6 159.4 291.4 ;
      RECT  163.4 290.6 164.2 291.4 ;
      RECT  168.2 290.6 169.0 291.4 ;
      RECT  173.0 290.6 173.8 291.4 ;
      RECT  177.8 290.6 178.6 291.4 ;
      RECT  5.0 295.4 5.8 296.2 ;
      RECT  9.8 295.4 10.6 296.2 ;
      RECT  14.6 295.4 15.4 296.2 ;
      RECT  19.4 295.4 20.2 296.2 ;
      RECT  24.2 295.4 25.0 296.2 ;
      RECT  29.0 295.4 29.8 296.2 ;
      RECT  33.8 295.4 34.6 296.2 ;
      RECT  38.6 295.4 39.4 296.2 ;
      RECT  43.4 295.4 44.2 296.2 ;
      RECT  48.2 295.4 49.0 296.2 ;
      RECT  53.0 295.4 53.8 296.2 ;
      RECT  57.8 295.4 58.6 296.2 ;
      RECT  62.6 295.4 63.4 296.2 ;
      RECT  67.4 295.4 68.2 296.2 ;
      RECT  72.2 295.4 73.0 296.2 ;
      RECT  77.0 295.4 77.8 296.2 ;
      RECT  81.8 295.4 82.6 296.2 ;
      RECT  86.6 295.4 87.4 296.2 ;
      RECT  91.4 295.4 92.2 296.2 ;
      RECT  96.2 295.4 97.0 296.2 ;
      RECT  101.0 295.4 101.8 296.2 ;
      RECT  105.8 295.4 106.6 296.2 ;
      RECT  110.6 295.4 111.4 296.2 ;
      RECT  115.4 295.4 116.2 296.2 ;
      RECT  120.2 295.4 121.0 296.2 ;
      RECT  125.0 295.4 125.8 296.2 ;
      RECT  129.8 295.4 130.6 296.2 ;
      RECT  134.6 295.4 135.4 296.2 ;
      RECT  139.4 295.4 140.2 296.2 ;
      RECT  144.2 295.4 145.0 296.2 ;
      RECT  149.0 295.4 149.8 296.2 ;
      RECT  153.8 295.4 154.6 296.2 ;
      RECT  158.6 295.4 159.4 296.2 ;
      RECT  163.4 295.4 164.2 296.2 ;
      RECT  168.2 295.4 169.0 296.2 ;
      RECT  173.0 295.4 173.8 296.2 ;
      RECT  177.8 295.4 178.6 296.2 ;
      RECT  182.6 295.4 183.4 296.2 ;
      RECT  187.4 295.4 188.2 296.2 ;
      RECT  192.2 295.4 193.0 296.2 ;
      RECT  197.0 295.4 197.8 296.2 ;
      RECT  201.8 295.4 202.6 296.2 ;
      RECT  206.6 295.4 207.4 296.2 ;
      RECT  211.4 295.4 212.2 296.2 ;
      RECT  216.2 295.4 217.0 296.2 ;
      RECT  221.0 295.4 221.8 296.2 ;
      RECT  225.8 295.4 226.6 296.2 ;
      RECT  5.0 300.2 5.8 301.0 ;
      RECT  9.8 300.2 10.6 301.0 ;
      RECT  14.6 300.2 15.4 301.0 ;
      RECT  19.4 300.2 20.2 301.0 ;
      RECT  24.2 300.2 25.0 301.0 ;
      RECT  29.0 300.2 29.8 301.0 ;
      RECT  33.8 300.2 34.6 301.0 ;
      RECT  38.6 300.2 39.4 301.0 ;
      RECT  43.4 300.2 44.2 301.0 ;
      RECT  48.2 300.2 49.0 301.0 ;
      RECT  53.0 300.2 53.8 301.0 ;
      RECT  57.8 300.2 58.6 301.0 ;
      RECT  62.6 300.2 63.4 301.0 ;
      RECT  67.4 300.2 68.2 301.0 ;
      RECT  72.2 300.2 73.0 301.0 ;
      RECT  77.0 300.2 77.8 301.0 ;
      RECT  81.8 300.2 82.6 301.0 ;
      RECT  86.6 300.2 87.4 301.0 ;
      RECT  91.4 300.2 92.2 301.0 ;
      RECT  96.2 300.2 97.0 301.0 ;
      RECT  101.0 300.2 101.8 301.0 ;
      RECT  105.8 300.2 106.6 301.0 ;
      RECT  110.6 300.2 111.4 301.0 ;
      RECT  115.4 300.2 116.2 301.0 ;
      RECT  120.2 300.2 121.0 301.0 ;
      RECT  125.0 300.2 125.8 301.0 ;
      RECT  129.8 300.2 130.6 301.0 ;
      RECT  134.6 300.2 135.4 301.0 ;
      RECT  139.4 300.2 140.2 301.0 ;
      RECT  177.8 300.2 178.6 301.0 ;
      RECT  182.6 300.2 183.4 301.0 ;
      RECT  187.4 300.2 188.2 301.0 ;
      RECT  192.2 300.2 193.0 301.0 ;
      RECT  197.0 300.2 197.8 301.0 ;
      RECT  201.8 300.2 202.6 301.0 ;
      RECT  206.6 300.2 207.4 301.0 ;
      RECT  211.4 300.2 212.2 301.0 ;
      RECT  216.2 300.2 217.0 301.0 ;
      RECT  221.0 300.2 221.8 301.0 ;
      RECT  225.8 300.2 226.6 301.0 ;
      RECT  5.0 305.0 5.8 305.8 ;
      RECT  9.8 305.0 10.6 305.8 ;
      RECT  14.6 305.0 15.4 305.8 ;
      RECT  19.4 305.0 20.2 305.8 ;
      RECT  24.2 305.0 25.0 305.8 ;
      RECT  29.0 305.0 29.8 305.8 ;
      RECT  33.8 305.0 34.6 305.8 ;
      RECT  38.6 305.0 39.4 305.8 ;
      RECT  43.4 305.0 44.2 305.8 ;
      RECT  48.2 305.0 49.0 305.8 ;
      RECT  53.0 305.0 53.8 305.8 ;
      RECT  57.8 305.0 58.6 305.8 ;
      RECT  62.6 305.0 63.4 305.8 ;
      RECT  67.4 305.0 68.2 305.8 ;
      RECT  72.2 305.0 73.0 305.8 ;
      RECT  77.0 305.0 77.8 305.8 ;
      RECT  81.8 305.0 82.6 305.8 ;
      RECT  86.6 305.0 87.4 305.8 ;
      RECT  91.4 305.0 92.2 305.8 ;
      RECT  96.2 305.0 97.0 305.8 ;
      RECT  101.0 305.0 101.8 305.8 ;
      RECT  105.8 305.0 106.6 305.8 ;
      RECT  110.6 305.0 111.4 305.8 ;
      RECT  115.4 305.0 116.2 305.8 ;
      RECT  120.2 305.0 121.0 305.8 ;
      RECT  125.0 305.0 125.8 305.8 ;
      RECT  129.8 305.0 130.6 305.8 ;
      RECT  134.6 305.0 135.4 305.8 ;
      RECT  139.4 305.0 140.2 305.8 ;
      RECT  144.2 305.0 145.0 305.8 ;
      RECT  149.0 305.0 149.8 305.8 ;
      RECT  153.8 305.0 154.6 305.8 ;
      RECT  158.6 305.0 159.4 305.8 ;
      RECT  163.4 305.0 164.2 305.8 ;
      RECT  168.2 305.0 169.0 305.8 ;
      RECT  173.0 305.0 173.8 305.8 ;
      RECT  177.8 305.0 178.6 305.8 ;
      RECT  5.0 309.8 5.8 310.6 ;
      RECT  9.8 309.8 10.6 310.6 ;
      RECT  14.6 309.8 15.4 310.6 ;
      RECT  19.4 309.8 20.2 310.6 ;
      RECT  24.2 309.8 25.0 310.6 ;
      RECT  29.0 309.8 29.8 310.6 ;
      RECT  33.8 309.8 34.6 310.6 ;
      RECT  38.6 309.8 39.4 310.6 ;
      RECT  43.4 309.8 44.2 310.6 ;
      RECT  48.2 309.8 49.0 310.6 ;
      RECT  53.0 309.8 53.8 310.6 ;
      RECT  57.8 309.8 58.6 310.6 ;
      RECT  62.6 309.8 63.4 310.6 ;
      RECT  67.4 309.8 68.2 310.6 ;
      RECT  72.2 309.8 73.0 310.6 ;
      RECT  77.0 309.8 77.8 310.6 ;
      RECT  81.8 309.8 82.6 310.6 ;
      RECT  86.6 309.8 87.4 310.6 ;
      RECT  91.4 309.8 92.2 310.6 ;
      RECT  96.2 309.8 97.0 310.6 ;
      RECT  101.0 309.8 101.8 310.6 ;
      RECT  105.8 309.8 106.6 310.6 ;
      RECT  110.6 309.8 111.4 310.6 ;
      RECT  115.4 309.8 116.2 310.6 ;
      RECT  120.2 309.8 121.0 310.6 ;
      RECT  125.0 309.8 125.8 310.6 ;
      RECT  129.8 309.8 130.6 310.6 ;
      RECT  134.6 309.8 135.4 310.6 ;
      RECT  139.4 309.8 140.2 310.6 ;
      RECT  144.2 309.8 145.0 310.6 ;
      RECT  149.0 309.8 149.8 310.6 ;
      RECT  153.8 309.8 154.6 310.6 ;
      RECT  158.6 309.8 159.4 310.6 ;
      RECT  163.4 309.8 164.2 310.6 ;
      RECT  168.2 309.8 169.0 310.6 ;
      RECT  173.0 309.8 173.8 310.6 ;
      RECT  177.8 309.8 178.6 310.6 ;
      RECT  182.6 309.8 183.4 310.6 ;
      RECT  187.4 309.8 188.2 310.6 ;
      RECT  192.2 309.8 193.0 310.6 ;
      RECT  197.0 309.8 197.8 310.6 ;
      RECT  201.8 309.8 202.6 310.6 ;
      RECT  206.6 309.8 207.4 310.6 ;
      RECT  211.4 309.8 212.2 310.6 ;
      RECT  216.2 309.8 217.0 310.6 ;
      RECT  221.0 309.8 221.8 310.6 ;
      RECT  225.8 309.8 226.6 310.6 ;
      RECT  5.0 314.6 5.8 315.4 ;
      RECT  9.8 314.6 10.6 315.4 ;
      RECT  14.6 314.6 15.4 315.4 ;
      RECT  19.4 314.6 20.2 315.4 ;
      RECT  24.2 314.6 25.0 315.4 ;
      RECT  29.0 314.6 29.8 315.4 ;
      RECT  33.8 314.6 34.6 315.4 ;
      RECT  38.6 314.6 39.4 315.4 ;
      RECT  43.4 314.6 44.2 315.4 ;
      RECT  48.2 314.6 49.0 315.4 ;
      RECT  53.0 314.6 53.8 315.4 ;
      RECT  57.8 314.6 58.6 315.4 ;
      RECT  62.6 314.6 63.4 315.4 ;
      RECT  67.4 314.6 68.2 315.4 ;
      RECT  72.2 314.6 73.0 315.4 ;
      RECT  77.0 314.6 77.8 315.4 ;
      RECT  81.8 314.6 82.6 315.4 ;
      RECT  86.6 314.6 87.4 315.4 ;
      RECT  91.4 314.6 92.2 315.4 ;
      RECT  96.2 314.6 97.0 315.4 ;
      RECT  101.0 314.6 101.8 315.4 ;
      RECT  105.8 314.6 106.6 315.4 ;
      RECT  110.6 314.6 111.4 315.4 ;
      RECT  115.4 314.6 116.2 315.4 ;
      RECT  120.2 314.6 121.0 315.4 ;
      RECT  125.0 314.6 125.8 315.4 ;
      RECT  129.8 314.6 130.6 315.4 ;
      RECT  134.6 314.6 135.4 315.4 ;
      RECT  139.4 314.6 140.2 315.4 ;
      RECT  144.2 314.6 145.0 315.4 ;
      RECT  149.0 314.6 149.8 315.4 ;
      RECT  153.8 314.6 154.6 315.4 ;
      RECT  158.6 314.6 159.4 315.4 ;
      RECT  163.4 314.6 164.2 315.4 ;
      RECT  168.2 314.6 169.0 315.4 ;
      RECT  173.0 314.6 173.8 315.4 ;
      RECT  177.8 314.6 178.6 315.4 ;
      RECT  5.0 319.4 5.8 320.2 ;
      RECT  9.8 319.4 10.6 320.2 ;
      RECT  14.6 319.4 15.4 320.2 ;
      RECT  19.4 319.4 20.2 320.2 ;
      RECT  24.2 319.4 25.0 320.2 ;
      RECT  29.0 319.4 29.8 320.2 ;
      RECT  33.8 319.4 34.6 320.2 ;
      RECT  38.6 319.4 39.4 320.2 ;
      RECT  43.4 319.4 44.2 320.2 ;
      RECT  48.2 319.4 49.0 320.2 ;
      RECT  53.0 319.4 53.8 320.2 ;
      RECT  57.8 319.4 58.6 320.2 ;
      RECT  62.6 319.4 63.4 320.2 ;
      RECT  67.4 319.4 68.2 320.2 ;
      RECT  72.2 319.4 73.0 320.2 ;
      RECT  77.0 319.4 77.8 320.2 ;
      RECT  81.8 319.4 82.6 320.2 ;
      RECT  86.6 319.4 87.4 320.2 ;
      RECT  91.4 319.4 92.2 320.2 ;
      RECT  96.2 319.4 97.0 320.2 ;
      RECT  101.0 319.4 101.8 320.2 ;
      RECT  105.8 319.4 106.6 320.2 ;
      RECT  110.6 319.4 111.4 320.2 ;
      RECT  115.4 319.4 116.2 320.2 ;
      RECT  120.2 319.4 121.0 320.2 ;
      RECT  125.0 319.4 125.8 320.2 ;
      RECT  129.8 319.4 130.6 320.2 ;
      RECT  134.6 319.4 135.4 320.2 ;
      RECT  139.4 319.4 140.2 320.2 ;
      RECT  177.8 319.4 178.6 320.2 ;
      RECT  182.6 319.4 183.4 320.2 ;
      RECT  187.4 319.4 188.2 320.2 ;
      RECT  192.2 319.4 193.0 320.2 ;
      RECT  197.0 319.4 197.8 320.2 ;
      RECT  201.8 319.4 202.6 320.2 ;
      RECT  206.6 319.4 207.4 320.2 ;
      RECT  211.4 319.4 212.2 320.2 ;
      RECT  216.2 319.4 217.0 320.2 ;
      RECT  221.0 319.4 221.8 320.2 ;
      RECT  225.8 319.4 226.6 320.2 ;
      RECT  5.0 324.2 5.8 325.0 ;
      RECT  9.8 324.2 10.6 325.0 ;
      RECT  14.6 324.2 15.4 325.0 ;
      RECT  19.4 324.2 20.2 325.0 ;
      RECT  24.2 324.2 25.0 325.0 ;
      RECT  29.0 324.2 29.8 325.0 ;
      RECT  33.8 324.2 34.6 325.0 ;
      RECT  38.6 324.2 39.4 325.0 ;
      RECT  43.4 324.2 44.2 325.0 ;
      RECT  48.2 324.2 49.0 325.0 ;
      RECT  53.0 324.2 53.8 325.0 ;
      RECT  57.8 324.2 58.6 325.0 ;
      RECT  62.6 324.2 63.4 325.0 ;
      RECT  67.4 324.2 68.2 325.0 ;
      RECT  72.2 324.2 73.0 325.0 ;
      RECT  77.0 324.2 77.8 325.0 ;
      RECT  96.2 324.2 97.0 325.0 ;
      RECT  101.0 324.2 101.8 325.0 ;
      RECT  105.8 324.2 106.6 325.0 ;
      RECT  110.6 324.2 111.4 325.0 ;
      RECT  115.4 324.2 116.2 325.0 ;
      RECT  120.2 324.2 121.0 325.0 ;
      RECT  125.0 324.2 125.8 325.0 ;
      RECT  129.8 324.2 130.6 325.0 ;
      RECT  134.6 324.2 135.4 325.0 ;
      RECT  139.4 324.2 140.2 325.0 ;
      RECT  144.2 324.2 145.0 325.0 ;
      RECT  149.0 324.2 149.8 325.0 ;
      RECT  153.8 324.2 154.6 325.0 ;
      RECT  158.6 324.2 159.4 325.0 ;
      RECT  163.4 324.2 164.2 325.0 ;
      RECT  168.2 324.2 169.0 325.0 ;
      RECT  173.0 324.2 173.8 325.0 ;
      RECT  177.8 324.2 178.6 325.0 ;
      RECT  5.0 329.0 5.8 329.8 ;
      RECT  9.8 329.0 10.6 329.8 ;
      RECT  14.6 329.0 15.4 329.8 ;
      RECT  19.4 329.0 20.2 329.8 ;
      RECT  24.2 329.0 25.0 329.8 ;
      RECT  29.0 329.0 29.8 329.8 ;
      RECT  33.8 329.0 34.6 329.8 ;
      RECT  38.6 329.0 39.4 329.8 ;
      RECT  43.4 329.0 44.2 329.8 ;
      RECT  48.2 329.0 49.0 329.8 ;
      RECT  53.0 329.0 53.8 329.8 ;
      RECT  57.8 329.0 58.6 329.8 ;
      RECT  62.6 329.0 63.4 329.8 ;
      RECT  67.4 329.0 68.2 329.8 ;
      RECT  72.2 329.0 73.0 329.8 ;
      RECT  77.0 329.0 77.8 329.8 ;
      RECT  81.8 329.0 82.6 329.8 ;
      RECT  86.6 329.0 87.4 329.8 ;
      RECT  91.4 329.0 92.2 329.8 ;
      RECT  96.2 329.0 97.0 329.8 ;
      RECT  101.0 329.0 101.8 329.8 ;
      RECT  105.8 329.0 106.6 329.8 ;
      RECT  110.6 329.0 111.4 329.8 ;
      RECT  115.4 329.0 116.2 329.8 ;
      RECT  120.2 329.0 121.0 329.8 ;
      RECT  125.0 329.0 125.8 329.8 ;
      RECT  129.8 329.0 130.6 329.8 ;
      RECT  134.6 329.0 135.4 329.8 ;
      RECT  139.4 329.0 140.2 329.8 ;
      RECT  144.2 329.0 145.0 329.8 ;
      RECT  149.0 329.0 149.8 329.8 ;
      RECT  153.8 329.0 154.6 329.8 ;
      RECT  158.6 329.0 159.4 329.8 ;
      RECT  163.4 329.0 164.2 329.8 ;
      RECT  168.2 329.0 169.0 329.8 ;
      RECT  173.0 329.0 173.8 329.8 ;
      RECT  177.8 329.0 178.6 329.8 ;
      RECT  182.6 329.0 183.4 329.8 ;
      RECT  187.4 329.0 188.2 329.8 ;
      RECT  192.2 329.0 193.0 329.8 ;
      RECT  197.0 329.0 197.8 329.8 ;
      RECT  201.8 329.0 202.6 329.8 ;
      RECT  206.6 329.0 207.4 329.8 ;
      RECT  211.4 329.0 212.2 329.8 ;
      RECT  216.2 329.0 217.0 329.8 ;
      RECT  221.0 329.0 221.8 329.8 ;
      RECT  225.8 329.0 226.6 329.8 ;
      RECT  5.0 333.8 5.8 334.6 ;
      RECT  9.8 333.8 10.6 334.6 ;
      RECT  14.6 333.8 15.4 334.6 ;
      RECT  19.4 333.8 20.2 334.6 ;
      RECT  24.2 333.8 25.0 334.6 ;
      RECT  29.0 333.8 29.8 334.6 ;
      RECT  33.8 333.8 34.6 334.6 ;
      RECT  38.6 333.8 39.4 334.6 ;
      RECT  43.4 333.8 44.2 334.6 ;
      RECT  48.2 333.8 49.0 334.6 ;
      RECT  53.0 333.8 53.8 334.6 ;
      RECT  57.8 333.8 58.6 334.6 ;
      RECT  62.6 333.8 63.4 334.6 ;
      RECT  67.4 333.8 68.2 334.6 ;
      RECT  81.8 333.8 82.6 334.6 ;
      RECT  86.6 333.8 87.4 334.6 ;
      RECT  91.4 333.8 92.2 334.6 ;
      RECT  96.2 333.8 97.0 334.6 ;
      RECT  101.0 333.8 101.8 334.6 ;
      RECT  105.8 333.8 106.6 334.6 ;
      RECT  110.6 333.8 111.4 334.6 ;
      RECT  115.4 333.8 116.2 334.6 ;
      RECT  120.2 333.8 121.0 334.6 ;
      RECT  125.0 333.8 125.8 334.6 ;
      RECT  129.8 333.8 130.6 334.6 ;
      RECT  134.6 333.8 135.4 334.6 ;
      RECT  139.4 333.8 140.2 334.6 ;
      RECT  144.2 333.8 145.0 334.6 ;
      RECT  149.0 333.8 149.8 334.6 ;
      RECT  153.8 333.8 154.6 334.6 ;
      RECT  158.6 333.8 159.4 334.6 ;
      RECT  163.4 333.8 164.2 334.6 ;
      RECT  168.2 333.8 169.0 334.6 ;
      RECT  173.0 333.8 173.8 334.6 ;
      RECT  177.8 333.8 178.6 334.6 ;
      RECT  5.0 338.6 5.8 339.4 ;
      RECT  9.8 338.6 10.6 339.4 ;
      RECT  14.6 338.6 15.4 339.4 ;
      RECT  19.4 338.6 20.2 339.4 ;
      RECT  24.2 338.6 25.0 339.4 ;
      RECT  29.0 338.6 29.8 339.4 ;
      RECT  33.8 338.6 34.6 339.4 ;
      RECT  38.6 338.6 39.4 339.4 ;
      RECT  43.4 338.6 44.2 339.4 ;
      RECT  48.2 338.6 49.0 339.4 ;
      RECT  53.0 338.6 53.8 339.4 ;
      RECT  57.8 338.6 58.6 339.4 ;
      RECT  62.6 338.6 63.4 339.4 ;
      RECT  67.4 338.6 68.2 339.4 ;
      RECT  72.2 338.6 73.0 339.4 ;
      RECT  77.0 338.6 77.8 339.4 ;
      RECT  81.8 338.6 82.6 339.4 ;
      RECT  86.6 338.6 87.4 339.4 ;
      RECT  91.4 338.6 92.2 339.4 ;
      RECT  96.2 338.6 97.0 339.4 ;
      RECT  101.0 338.6 101.8 339.4 ;
      RECT  105.8 338.6 106.6 339.4 ;
      RECT  110.6 338.6 111.4 339.4 ;
      RECT  115.4 338.6 116.2 339.4 ;
      RECT  120.2 338.6 121.0 339.4 ;
      RECT  125.0 338.6 125.8 339.4 ;
      RECT  129.8 338.6 130.6 339.4 ;
      RECT  134.6 338.6 135.4 339.4 ;
      RECT  139.4 338.6 140.2 339.4 ;
      RECT  177.8 338.6 178.6 339.4 ;
      RECT  182.6 338.6 183.4 339.4 ;
      RECT  187.4 338.6 188.2 339.4 ;
      RECT  192.2 338.6 193.0 339.4 ;
      RECT  197.0 338.6 197.8 339.4 ;
      RECT  201.8 338.6 202.6 339.4 ;
      RECT  206.6 338.6 207.4 339.4 ;
      RECT  211.4 338.6 212.2 339.4 ;
      RECT  216.2 338.6 217.0 339.4 ;
      RECT  221.0 338.6 221.8 339.4 ;
      RECT  225.8 338.6 226.6 339.4 ;
      RECT  5.0 343.4 5.8 344.2 ;
      RECT  9.8 343.4 10.6 344.2 ;
      RECT  14.6 343.4 15.4 344.2 ;
      RECT  19.4 343.4 20.2 344.2 ;
      RECT  24.2 343.4 25.0 344.2 ;
      RECT  29.0 343.4 29.8 344.2 ;
      RECT  33.8 343.4 34.6 344.2 ;
      RECT  38.6 343.4 39.4 344.2 ;
      RECT  43.4 343.4 44.2 344.2 ;
      RECT  48.2 343.4 49.0 344.2 ;
      RECT  53.0 343.4 53.8 344.2 ;
      RECT  57.8 343.4 58.6 344.2 ;
      RECT  62.6 343.4 63.4 344.2 ;
      RECT  67.4 343.4 68.2 344.2 ;
      RECT  72.2 343.4 73.0 344.2 ;
      RECT  77.0 343.4 77.8 344.2 ;
      RECT  101.0 343.4 101.8 344.2 ;
      RECT  105.8 343.4 106.6 344.2 ;
      RECT  110.6 343.4 111.4 344.2 ;
      RECT  115.4 343.4 116.2 344.2 ;
      RECT  120.2 343.4 121.0 344.2 ;
      RECT  125.0 343.4 125.8 344.2 ;
      RECT  129.8 343.4 130.6 344.2 ;
      RECT  134.6 343.4 135.4 344.2 ;
      RECT  139.4 343.4 140.2 344.2 ;
      RECT  144.2 343.4 145.0 344.2 ;
      RECT  149.0 343.4 149.8 344.2 ;
      RECT  153.8 343.4 154.6 344.2 ;
      RECT  158.6 343.4 159.4 344.2 ;
      RECT  163.4 343.4 164.2 344.2 ;
      RECT  168.2 343.4 169.0 344.2 ;
      RECT  173.0 343.4 173.8 344.2 ;
      RECT  177.8 343.4 178.6 344.2 ;
      RECT  5.0 348.2 5.8 349.0 ;
      RECT  9.8 348.2 10.6 349.0 ;
      RECT  14.6 348.2 15.4 349.0 ;
      RECT  19.4 348.2 20.2 349.0 ;
      RECT  24.2 348.2 25.0 349.0 ;
      RECT  29.0 348.2 29.8 349.0 ;
      RECT  33.8 348.2 34.6 349.0 ;
      RECT  38.6 348.2 39.4 349.0 ;
      RECT  43.4 348.2 44.2 349.0 ;
      RECT  48.2 348.2 49.0 349.0 ;
      RECT  53.0 348.2 53.8 349.0 ;
      RECT  57.8 348.2 58.6 349.0 ;
      RECT  62.6 348.2 63.4 349.0 ;
      RECT  67.4 348.2 68.2 349.0 ;
      RECT  72.2 348.2 73.0 349.0 ;
      RECT  77.0 348.2 77.8 349.0 ;
      RECT  81.8 348.2 82.6 349.0 ;
      RECT  86.6 348.2 87.4 349.0 ;
      RECT  91.4 348.2 92.2 349.0 ;
      RECT  96.2 348.2 97.0 349.0 ;
      RECT  101.0 348.2 101.8 349.0 ;
      RECT  105.8 348.2 106.6 349.0 ;
      RECT  110.6 348.2 111.4 349.0 ;
      RECT  115.4 348.2 116.2 349.0 ;
      RECT  120.2 348.2 121.0 349.0 ;
      RECT  125.0 348.2 125.8 349.0 ;
      RECT  129.8 348.2 130.6 349.0 ;
      RECT  134.6 348.2 135.4 349.0 ;
      RECT  139.4 348.2 140.2 349.0 ;
      RECT  144.2 348.2 145.0 349.0 ;
      RECT  149.0 348.2 149.8 349.0 ;
      RECT  153.8 348.2 154.6 349.0 ;
      RECT  158.6 348.2 159.4 349.0 ;
      RECT  163.4 348.2 164.2 349.0 ;
      RECT  168.2 348.2 169.0 349.0 ;
      RECT  173.0 348.2 173.8 349.0 ;
      RECT  177.8 348.2 178.6 349.0 ;
      RECT  182.6 348.2 183.4 349.0 ;
      RECT  187.4 348.2 188.2 349.0 ;
      RECT  192.2 348.2 193.0 349.0 ;
      RECT  197.0 348.2 197.8 349.0 ;
      RECT  201.8 348.2 202.6 349.0 ;
      RECT  206.6 348.2 207.4 349.0 ;
      RECT  211.4 348.2 212.2 349.0 ;
      RECT  216.2 348.2 217.0 349.0 ;
      RECT  221.0 348.2 221.8 349.0 ;
      RECT  225.8 348.2 226.6 349.0 ;
      RECT  5.0 353.0 5.8 353.8 ;
      RECT  9.8 353.0 10.6 353.8 ;
      RECT  14.6 353.0 15.4 353.8 ;
      RECT  19.4 353.0 20.2 353.8 ;
      RECT  24.2 353.0 25.0 353.8 ;
      RECT  29.0 353.0 29.8 353.8 ;
      RECT  33.8 353.0 34.6 353.8 ;
      RECT  38.6 353.0 39.4 353.8 ;
      RECT  43.4 353.0 44.2 353.8 ;
      RECT  48.2 353.0 49.0 353.8 ;
      RECT  53.0 353.0 53.8 353.8 ;
      RECT  57.8 353.0 58.6 353.8 ;
      RECT  62.6 353.0 63.4 353.8 ;
      RECT  67.4 353.0 68.2 353.8 ;
      RECT  72.2 353.0 73.0 353.8 ;
      RECT  77.0 353.0 77.8 353.8 ;
      RECT  81.8 353.0 82.6 353.8 ;
      RECT  86.6 353.0 87.4 353.8 ;
      RECT  91.4 353.0 92.2 353.8 ;
      RECT  96.2 353.0 97.0 353.8 ;
      RECT  101.0 353.0 101.8 353.8 ;
      RECT  105.8 353.0 106.6 353.8 ;
      RECT  110.6 353.0 111.4 353.8 ;
      RECT  115.4 353.0 116.2 353.8 ;
      RECT  120.2 353.0 121.0 353.8 ;
      RECT  125.0 353.0 125.8 353.8 ;
      RECT  129.8 353.0 130.6 353.8 ;
      RECT  134.6 353.0 135.4 353.8 ;
      RECT  139.4 353.0 140.2 353.8 ;
      RECT  144.2 353.0 145.0 353.8 ;
      RECT  149.0 353.0 149.8 353.8 ;
      RECT  153.8 353.0 154.6 353.8 ;
      RECT  158.6 353.0 159.4 353.8 ;
      RECT  163.4 353.0 164.2 353.8 ;
      RECT  168.2 353.0 169.0 353.8 ;
      RECT  173.0 353.0 173.8 353.8 ;
      RECT  177.8 353.0 178.6 353.8 ;
      RECT  5.0 357.8 5.8 358.6 ;
      RECT  9.8 357.8 10.6 358.6 ;
      RECT  14.6 357.8 15.4 358.6 ;
      RECT  19.4 357.8 20.2 358.6 ;
      RECT  24.2 357.8 25.0 358.6 ;
      RECT  29.0 357.8 29.8 358.6 ;
      RECT  33.8 357.8 34.6 358.6 ;
      RECT  38.6 357.8 39.4 358.6 ;
      RECT  43.4 357.8 44.2 358.6 ;
      RECT  48.2 357.8 49.0 358.6 ;
      RECT  53.0 357.8 53.8 358.6 ;
      RECT  57.8 357.8 58.6 358.6 ;
      RECT  62.6 357.8 63.4 358.6 ;
      RECT  67.4 357.8 68.2 358.6 ;
      RECT  72.2 357.8 73.0 358.6 ;
      RECT  77.0 357.8 77.8 358.6 ;
      RECT  81.8 357.8 82.6 358.6 ;
      RECT  86.6 357.8 87.4 358.6 ;
      RECT  91.4 357.8 92.2 358.6 ;
      RECT  96.2 357.8 97.0 358.6 ;
      RECT  101.0 357.8 101.8 358.6 ;
      RECT  105.8 357.8 106.6 358.6 ;
      RECT  110.6 357.8 111.4 358.6 ;
      RECT  115.4 357.8 116.2 358.6 ;
      RECT  120.2 357.8 121.0 358.6 ;
      RECT  125.0 357.8 125.8 358.6 ;
      RECT  129.8 357.8 130.6 358.6 ;
      RECT  134.6 357.8 135.4 358.6 ;
      RECT  139.4 357.8 140.2 358.6 ;
      RECT  144.2 357.8 145.0 358.6 ;
      RECT  149.0 357.8 149.8 358.6 ;
      RECT  153.8 357.8 154.6 358.6 ;
      RECT  158.6 357.8 159.4 358.6 ;
      RECT  163.4 357.8 164.2 358.6 ;
      RECT  168.2 357.8 169.0 358.6 ;
      RECT  173.0 357.8 173.8 358.6 ;
      RECT  177.8 357.8 178.6 358.6 ;
      RECT  182.6 357.8 183.4 358.6 ;
      RECT  187.4 357.8 188.2 358.6 ;
      RECT  192.2 357.8 193.0 358.6 ;
      RECT  197.0 357.8 197.8 358.6 ;
      RECT  201.8 357.8 202.6 358.6 ;
      RECT  206.6 357.8 207.4 358.6 ;
      RECT  211.4 357.8 212.2 358.6 ;
      RECT  216.2 357.8 217.0 358.6 ;
      RECT  221.0 357.8 221.8 358.6 ;
      RECT  225.8 357.8 226.6 358.6 ;
      RECT  5.0 362.6 5.8 363.4 ;
      RECT  9.8 362.6 10.6 363.4 ;
      RECT  14.6 362.6 15.4 363.4 ;
      RECT  19.4 362.6 20.2 363.4 ;
      RECT  24.2 362.6 25.0 363.4 ;
      RECT  29.0 362.6 29.8 363.4 ;
      RECT  33.8 362.6 34.6 363.4 ;
      RECT  38.6 362.6 39.4 363.4 ;
      RECT  43.4 362.6 44.2 363.4 ;
      RECT  48.2 362.6 49.0 363.4 ;
      RECT  53.0 362.6 53.8 363.4 ;
      RECT  57.8 362.6 58.6 363.4 ;
      RECT  62.6 362.6 63.4 363.4 ;
      RECT  67.4 362.6 68.2 363.4 ;
      RECT  72.2 362.6 73.0 363.4 ;
      RECT  77.0 362.6 77.8 363.4 ;
      RECT  101.0 362.6 101.8 363.4 ;
      RECT  105.8 362.6 106.6 363.4 ;
      RECT  110.6 362.6 111.4 363.4 ;
      RECT  115.4 362.6 116.2 363.4 ;
      RECT  120.2 362.6 121.0 363.4 ;
      RECT  125.0 362.6 125.8 363.4 ;
      RECT  129.8 362.6 130.6 363.4 ;
      RECT  134.6 362.6 135.4 363.4 ;
      RECT  139.4 362.6 140.2 363.4 ;
      RECT  177.8 362.6 178.6 363.4 ;
      RECT  182.6 362.6 183.4 363.4 ;
      RECT  187.4 362.6 188.2 363.4 ;
      RECT  192.2 362.6 193.0 363.4 ;
      RECT  197.0 362.6 197.8 363.4 ;
      RECT  201.8 362.6 202.6 363.4 ;
      RECT  206.6 362.6 207.4 363.4 ;
      RECT  211.4 362.6 212.2 363.4 ;
      RECT  216.2 362.6 217.0 363.4 ;
      RECT  221.0 362.6 221.8 363.4 ;
      RECT  225.8 362.6 226.6 363.4 ;
      RECT  5.0 367.4 5.8 368.2 ;
      RECT  9.8 367.4 10.6 368.2 ;
      RECT  14.6 367.4 15.4 368.2 ;
      RECT  19.4 367.4 20.2 368.2 ;
      RECT  24.2 367.4 25.0 368.2 ;
      RECT  29.0 367.4 29.8 368.2 ;
      RECT  33.8 367.4 34.6 368.2 ;
      RECT  38.6 367.4 39.4 368.2 ;
      RECT  43.4 367.4 44.2 368.2 ;
      RECT  48.2 367.4 49.0 368.2 ;
      RECT  53.0 367.4 53.8 368.2 ;
      RECT  57.8 367.4 58.6 368.2 ;
      RECT  62.6 367.4 63.4 368.2 ;
      RECT  67.4 367.4 68.2 368.2 ;
      RECT  72.2 367.4 73.0 368.2 ;
      RECT  77.0 367.4 77.8 368.2 ;
      RECT  81.8 367.4 82.6 368.2 ;
      RECT  86.6 367.4 87.4 368.2 ;
      RECT  91.4 367.4 92.2 368.2 ;
      RECT  96.2 367.4 97.0 368.2 ;
      RECT  101.0 367.4 101.8 368.2 ;
      RECT  105.8 367.4 106.6 368.2 ;
      RECT  110.6 367.4 111.4 368.2 ;
      RECT  115.4 367.4 116.2 368.2 ;
      RECT  120.2 367.4 121.0 368.2 ;
      RECT  125.0 367.4 125.8 368.2 ;
      RECT  129.8 367.4 130.6 368.2 ;
      RECT  134.6 367.4 135.4 368.2 ;
      RECT  139.4 367.4 140.2 368.2 ;
      RECT  144.2 367.4 145.0 368.2 ;
      RECT  149.0 367.4 149.8 368.2 ;
      RECT  153.8 367.4 154.6 368.2 ;
      RECT  158.6 367.4 159.4 368.2 ;
      RECT  163.4 367.4 164.2 368.2 ;
      RECT  168.2 367.4 169.0 368.2 ;
      RECT  173.0 367.4 173.8 368.2 ;
      RECT  177.8 367.4 178.6 368.2 ;
      RECT  105.8 247.4 106.6 248.2 ;
      RECT  105.8 204.2 106.6 205.0 ;
      RECT  187.4 369.8 188.2 370.6 ;
      RECT  197.0 369.8 197.8 370.6 ;
      RECT  201.8 369.8 202.6 370.6 ;
      RECT  211.4 369.8 212.2 370.6 ;
      RECT  216.2 369.8 217.0 370.6 ;
   LAYER  metal4 ;
      RECT  105.6 247.2 106.8 248.4 ;
      RECT  105.6 204.0 106.8 205.2 ;
      RECT  187.2 369.6 188.4 370.8 ;
      RECT  196.8 369.6 198.0 370.8 ;
      RECT  201.6 369.6 202.8 370.8 ;
      RECT  211.2 369.6 212.4 370.8 ;
      RECT  216.0 369.6 217.2 370.8 ;
      RECT  2.4 0.0 3.6 1.2 ;
      RECT  7.2 0.0 8.4 1.2 ;
      RECT  12.0 0.0 13.2 1.2 ;
      RECT  16.8 0.0 18.0 1.2 ;
      RECT  21.6 0.0 22.8 1.2 ;
      RECT  26.4 0.0 27.6 1.2 ;
      RECT  31.2 0.0 32.4 1.2 ;
      RECT  36.0 0.0 37.2 1.2 ;
      RECT  40.8 0.0 42.0 1.2 ;
      RECT  45.6 0.0 46.8 1.2 ;
      RECT  50.4 0.0 51.6 1.2 ;
      RECT  55.2 0.0 56.4 1.2 ;
      RECT  60.0 0.0 61.2 1.2 ;
      RECT  64.8 0.0 66.0 1.2 ;
      RECT  69.6 0.0 70.8 1.2 ;
      RECT  74.4 0.0 75.6 1.2 ;
      RECT  79.2 0.0 80.4 1.2 ;
      RECT  84.0 0.0 85.2 1.2 ;
      RECT  88.8 0.0 90.0 1.2 ;
      RECT  93.6 0.0 94.8 1.2 ;
      RECT  98.4 0.0 99.6 1.2 ;
      RECT  103.2 0.0 104.4 1.2 ;
      RECT  108.0 0.0 109.2 1.2 ;
      RECT  112.8 0.0 114.0 1.2 ;
      RECT  117.6 0.0 118.8 1.2 ;
      RECT  122.4 0.0 123.6 1.2 ;
      RECT  127.2 0.0 128.4 1.2 ;
      RECT  132.0 0.0 133.2 1.2 ;
      RECT  136.8 0.0 138.0 1.2 ;
      RECT  141.6 0.0 142.8 1.2 ;
      RECT  146.4 0.0 147.6 1.2 ;
      RECT  151.2 0.0 152.4 1.2 ;
      RECT  156.0 0.0 157.2 1.2 ;
      RECT  160.8 0.0 162.0 1.2 ;
      RECT  165.6 0.0 166.8 1.2 ;
      RECT  170.4 0.0 171.6 1.2 ;
      RECT  175.2 0.0 176.4 1.2 ;
      RECT  180.0 0.0 181.2 1.2 ;
      RECT  184.8 0.0 186.0 1.2 ;
      RECT  189.6 0.0 190.8 1.2 ;
      RECT  194.4 0.0 195.6 1.2 ;
      RECT  199.2 0.0 200.4 1.2 ;
      RECT  204.0 0.0 205.2 1.2 ;
      RECT  208.8 0.0 210.0 1.2 ;
      RECT  213.6 0.0 214.8 1.2 ;
      RECT  218.4 0.0 219.6 1.2 ;
      RECT  223.2 0.0 224.4 1.2 ;
      RECT  2.4 4.8 3.6 6.0 ;
      RECT  7.2 4.8 8.4 6.0 ;
      RECT  12.0 4.8 13.2 6.0 ;
      RECT  16.8 4.8 18.0 6.0 ;
      RECT  21.6 4.8 22.8 6.0 ;
      RECT  26.4 4.8 27.6 6.0 ;
      RECT  31.2 4.8 32.4 6.0 ;
      RECT  36.0 4.8 37.2 6.0 ;
      RECT  79.2 4.8 80.4 6.0 ;
      RECT  84.0 4.8 85.2 6.0 ;
      RECT  88.8 4.8 90.0 6.0 ;
      RECT  93.6 4.8 94.8 6.0 ;
      RECT  98.4 4.8 99.6 6.0 ;
      RECT  103.2 4.8 104.4 6.0 ;
      RECT  108.0 4.8 109.2 6.0 ;
      RECT  112.8 4.8 114.0 6.0 ;
      RECT  117.6 4.8 118.8 6.0 ;
      RECT  122.4 4.8 123.6 6.0 ;
      RECT  127.2 4.8 128.4 6.0 ;
      RECT  132.0 4.8 133.2 6.0 ;
      RECT  136.8 4.8 138.0 6.0 ;
      RECT  141.6 4.8 142.8 6.0 ;
      RECT  146.4 4.8 147.6 6.0 ;
      RECT  151.2 4.8 152.4 6.0 ;
      RECT  156.0 4.8 157.2 6.0 ;
      RECT  160.8 4.8 162.0 6.0 ;
      RECT  165.6 4.8 166.8 6.0 ;
      RECT  170.4 4.8 171.6 6.0 ;
      RECT  175.2 4.8 176.4 6.0 ;
      RECT  180.0 4.8 181.2 6.0 ;
      RECT  184.8 4.8 186.0 6.0 ;
      RECT  189.6 4.8 190.8 6.0 ;
      RECT  194.4 4.8 195.6 6.0 ;
      RECT  199.2 4.8 200.4 6.0 ;
      RECT  204.0 4.8 205.2 6.0 ;
      RECT  208.8 4.8 210.0 6.0 ;
      RECT  213.6 4.8 214.8 6.0 ;
      RECT  218.4 4.8 219.6 6.0 ;
      RECT  223.2 4.8 224.4 6.0 ;
      RECT  31.2 9.6 32.4 10.8 ;
      RECT  36.0 9.6 37.2 10.8 ;
      RECT  40.8 9.6 42.0 10.8 ;
      RECT  45.6 9.6 46.8 10.8 ;
      RECT  50.4 9.6 51.6 10.8 ;
      RECT  55.2 9.6 56.4 10.8 ;
      RECT  60.0 9.6 61.2 10.8 ;
      RECT  64.8 9.6 66.0 10.8 ;
      RECT  69.6 9.6 70.8 10.8 ;
      RECT  74.4 9.6 75.6 10.8 ;
      RECT  79.2 9.6 80.4 10.8 ;
      RECT  84.0 9.6 85.2 10.8 ;
      RECT  88.8 9.6 90.0 10.8 ;
      RECT  93.6 9.6 94.8 10.8 ;
      RECT  98.4 9.6 99.6 10.8 ;
      RECT  103.2 9.6 104.4 10.8 ;
      RECT  108.0 9.6 109.2 10.8 ;
      RECT  112.8 9.6 114.0 10.8 ;
      RECT  117.6 9.6 118.8 10.8 ;
      RECT  122.4 9.6 123.6 10.8 ;
      RECT  127.2 9.6 128.4 10.8 ;
      RECT  132.0 9.6 133.2 10.8 ;
      RECT  136.8 9.6 138.0 10.8 ;
      RECT  141.6 9.6 142.8 10.8 ;
      RECT  146.4 9.6 147.6 10.8 ;
      RECT  151.2 9.6 152.4 10.8 ;
      RECT  156.0 9.6 157.2 10.8 ;
      RECT  160.8 9.6 162.0 10.8 ;
      RECT  165.6 9.6 166.8 10.8 ;
      RECT  170.4 9.6 171.6 10.8 ;
      RECT  175.2 9.6 176.4 10.8 ;
      RECT  180.0 9.6 181.2 10.8 ;
      RECT  184.8 9.6 186.0 10.8 ;
      RECT  189.6 9.6 190.8 10.8 ;
      RECT  194.4 9.6 195.6 10.8 ;
      RECT  199.2 9.6 200.4 10.8 ;
      RECT  204.0 9.6 205.2 10.8 ;
      RECT  208.8 9.6 210.0 10.8 ;
      RECT  213.6 9.6 214.8 10.8 ;
      RECT  218.4 9.6 219.6 10.8 ;
      RECT  223.2 9.6 224.4 10.8 ;
      RECT  50.4 14.4 51.6 15.6 ;
      RECT  55.2 14.4 56.4 15.6 ;
      RECT  60.0 14.4 61.2 15.6 ;
      RECT  64.8 14.4 66.0 15.6 ;
      RECT  69.6 14.4 70.8 15.6 ;
      RECT  74.4 14.4 75.6 15.6 ;
      RECT  79.2 14.4 80.4 15.6 ;
      RECT  84.0 14.4 85.2 15.6 ;
      RECT  88.8 14.4 90.0 15.6 ;
      RECT  93.6 14.4 94.8 15.6 ;
      RECT  98.4 14.4 99.6 15.6 ;
      RECT  103.2 14.4 104.4 15.6 ;
      RECT  108.0 14.4 109.2 15.6 ;
      RECT  112.8 14.4 114.0 15.6 ;
      RECT  117.6 14.4 118.8 15.6 ;
      RECT  122.4 14.4 123.6 15.6 ;
      RECT  127.2 14.4 128.4 15.6 ;
      RECT  132.0 14.4 133.2 15.6 ;
      RECT  136.8 14.4 138.0 15.6 ;
      RECT  141.6 14.4 142.8 15.6 ;
      RECT  146.4 14.4 147.6 15.6 ;
      RECT  151.2 14.4 152.4 15.6 ;
      RECT  156.0 14.4 157.2 15.6 ;
      RECT  160.8 14.4 162.0 15.6 ;
      RECT  165.6 14.4 166.8 15.6 ;
      RECT  170.4 14.4 171.6 15.6 ;
      RECT  175.2 14.4 176.4 15.6 ;
      RECT  180.0 14.4 181.2 15.6 ;
      RECT  184.8 14.4 186.0 15.6 ;
      RECT  189.6 14.4 190.8 15.6 ;
      RECT  194.4 14.4 195.6 15.6 ;
      RECT  199.2 14.4 200.4 15.6 ;
      RECT  204.0 14.4 205.2 15.6 ;
      RECT  208.8 14.4 210.0 15.6 ;
      RECT  213.6 14.4 214.8 15.6 ;
      RECT  218.4 14.4 219.6 15.6 ;
      RECT  223.2 14.4 224.4 15.6 ;
      RECT  2.4 19.2 3.6 20.4 ;
      RECT  7.2 19.2 8.4 20.4 ;
      RECT  12.0 19.2 13.2 20.4 ;
      RECT  16.8 19.2 18.0 20.4 ;
      RECT  21.6 19.2 22.8 20.4 ;
      RECT  26.4 19.2 27.6 20.4 ;
      RECT  31.2 19.2 32.4 20.4 ;
      RECT  36.0 19.2 37.2 20.4 ;
      RECT  40.8 19.2 42.0 20.4 ;
      RECT  45.6 19.2 46.8 20.4 ;
      RECT  50.4 19.2 51.6 20.4 ;
      RECT  55.2 19.2 56.4 20.4 ;
      RECT  60.0 19.2 61.2 20.4 ;
      RECT  64.8 19.2 66.0 20.4 ;
      RECT  69.6 19.2 70.8 20.4 ;
      RECT  74.4 19.2 75.6 20.4 ;
      RECT  79.2 19.2 80.4 20.4 ;
      RECT  84.0 19.2 85.2 20.4 ;
      RECT  88.8 19.2 90.0 20.4 ;
      RECT  93.6 19.2 94.8 20.4 ;
      RECT  98.4 19.2 99.6 20.4 ;
      RECT  103.2 19.2 104.4 20.4 ;
      RECT  108.0 19.2 109.2 20.4 ;
      RECT  112.8 19.2 114.0 20.4 ;
      RECT  117.6 19.2 118.8 20.4 ;
      RECT  122.4 19.2 123.6 20.4 ;
      RECT  127.2 19.2 128.4 20.4 ;
      RECT  132.0 19.2 133.2 20.4 ;
      RECT  136.8 19.2 138.0 20.4 ;
      RECT  141.6 19.2 142.8 20.4 ;
      RECT  146.4 19.2 147.6 20.4 ;
      RECT  151.2 19.2 152.4 20.4 ;
      RECT  156.0 19.2 157.2 20.4 ;
      RECT  160.8 19.2 162.0 20.4 ;
      RECT  165.6 19.2 166.8 20.4 ;
      RECT  170.4 19.2 171.6 20.4 ;
      RECT  175.2 19.2 176.4 20.4 ;
      RECT  180.0 19.2 181.2 20.4 ;
      RECT  184.8 19.2 186.0 20.4 ;
      RECT  189.6 19.2 190.8 20.4 ;
      RECT  194.4 19.2 195.6 20.4 ;
      RECT  199.2 19.2 200.4 20.4 ;
      RECT  204.0 19.2 205.2 20.4 ;
      RECT  208.8 19.2 210.0 20.4 ;
      RECT  213.6 19.2 214.8 20.4 ;
      RECT  218.4 19.2 219.6 20.4 ;
      RECT  223.2 19.2 224.4 20.4 ;
      RECT  2.4 24.0 3.6 25.2 ;
      RECT  7.2 24.0 8.4 25.2 ;
      RECT  12.0 24.0 13.2 25.2 ;
      RECT  16.8 24.0 18.0 25.2 ;
      RECT  21.6 24.0 22.8 25.2 ;
      RECT  26.4 24.0 27.6 25.2 ;
      RECT  31.2 24.0 32.4 25.2 ;
      RECT  36.0 24.0 37.2 25.2 ;
      RECT  40.8 24.0 42.0 25.2 ;
      RECT  45.6 24.0 46.8 25.2 ;
      RECT  50.4 24.0 51.6 25.2 ;
      RECT  55.2 24.0 56.4 25.2 ;
      RECT  60.0 24.0 61.2 25.2 ;
      RECT  64.8 24.0 66.0 25.2 ;
      RECT  69.6 24.0 70.8 25.2 ;
      RECT  74.4 24.0 75.6 25.2 ;
      RECT  79.2 24.0 80.4 25.2 ;
      RECT  84.0 24.0 85.2 25.2 ;
      RECT  88.8 24.0 90.0 25.2 ;
      RECT  93.6 24.0 94.8 25.2 ;
      RECT  98.4 24.0 99.6 25.2 ;
      RECT  103.2 24.0 104.4 25.2 ;
      RECT  108.0 24.0 109.2 25.2 ;
      RECT  112.8 24.0 114.0 25.2 ;
      RECT  117.6 24.0 118.8 25.2 ;
      RECT  122.4 24.0 123.6 25.2 ;
      RECT  127.2 24.0 128.4 25.2 ;
      RECT  132.0 24.0 133.2 25.2 ;
      RECT  136.8 24.0 138.0 25.2 ;
      RECT  141.6 24.0 142.8 25.2 ;
      RECT  146.4 24.0 147.6 25.2 ;
      RECT  151.2 24.0 152.4 25.2 ;
      RECT  156.0 24.0 157.2 25.2 ;
      RECT  160.8 24.0 162.0 25.2 ;
      RECT  165.6 24.0 166.8 25.2 ;
      RECT  170.4 24.0 171.6 25.2 ;
      RECT  175.2 24.0 176.4 25.2 ;
      RECT  180.0 24.0 181.2 25.2 ;
      RECT  184.8 24.0 186.0 25.2 ;
      RECT  189.6 24.0 190.8 25.2 ;
      RECT  194.4 24.0 195.6 25.2 ;
      RECT  199.2 24.0 200.4 25.2 ;
      RECT  204.0 24.0 205.2 25.2 ;
      RECT  208.8 24.0 210.0 25.2 ;
      RECT  213.6 24.0 214.8 25.2 ;
      RECT  218.4 24.0 219.6 25.2 ;
      RECT  223.2 24.0 224.4 25.2 ;
      RECT  45.6 28.8 46.8 30.0 ;
      RECT  50.4 28.8 51.6 30.0 ;
      RECT  55.2 28.8 56.4 30.0 ;
      RECT  60.0 28.8 61.2 30.0 ;
      RECT  64.8 28.8 66.0 30.0 ;
      RECT  69.6 28.8 70.8 30.0 ;
      RECT  74.4 28.8 75.6 30.0 ;
      RECT  79.2 28.8 80.4 30.0 ;
      RECT  84.0 28.8 85.2 30.0 ;
      RECT  88.8 28.8 90.0 30.0 ;
      RECT  93.6 28.8 94.8 30.0 ;
      RECT  98.4 28.8 99.6 30.0 ;
      RECT  103.2 28.8 104.4 30.0 ;
      RECT  108.0 28.8 109.2 30.0 ;
      RECT  112.8 28.8 114.0 30.0 ;
      RECT  117.6 28.8 118.8 30.0 ;
      RECT  122.4 28.8 123.6 30.0 ;
      RECT  127.2 28.8 128.4 30.0 ;
      RECT  132.0 28.8 133.2 30.0 ;
      RECT  136.8 28.8 138.0 30.0 ;
      RECT  141.6 28.8 142.8 30.0 ;
      RECT  146.4 28.8 147.6 30.0 ;
      RECT  151.2 28.8 152.4 30.0 ;
      RECT  156.0 28.8 157.2 30.0 ;
      RECT  160.8 28.8 162.0 30.0 ;
      RECT  165.6 28.8 166.8 30.0 ;
      RECT  170.4 28.8 171.6 30.0 ;
      RECT  175.2 28.8 176.4 30.0 ;
      RECT  180.0 28.8 181.2 30.0 ;
      RECT  184.8 28.8 186.0 30.0 ;
      RECT  189.6 28.8 190.8 30.0 ;
      RECT  194.4 28.8 195.6 30.0 ;
      RECT  199.2 28.8 200.4 30.0 ;
      RECT  204.0 28.8 205.2 30.0 ;
      RECT  208.8 28.8 210.0 30.0 ;
      RECT  213.6 28.8 214.8 30.0 ;
      RECT  218.4 28.8 219.6 30.0 ;
      RECT  223.2 28.8 224.4 30.0 ;
      RECT  84.0 33.6 85.2 34.8 ;
      RECT  88.8 33.6 90.0 34.8 ;
      RECT  93.6 33.6 94.8 34.8 ;
      RECT  98.4 33.6 99.6 34.8 ;
      RECT  103.2 33.6 104.4 34.8 ;
      RECT  108.0 33.6 109.2 34.8 ;
      RECT  112.8 33.6 114.0 34.8 ;
      RECT  117.6 33.6 118.8 34.8 ;
      RECT  122.4 33.6 123.6 34.8 ;
      RECT  127.2 33.6 128.4 34.8 ;
      RECT  132.0 33.6 133.2 34.8 ;
      RECT  136.8 33.6 138.0 34.8 ;
      RECT  141.6 33.6 142.8 34.8 ;
      RECT  146.4 33.6 147.6 34.8 ;
      RECT  151.2 33.6 152.4 34.8 ;
      RECT  156.0 33.6 157.2 34.8 ;
      RECT  160.8 33.6 162.0 34.8 ;
      RECT  165.6 33.6 166.8 34.8 ;
      RECT  170.4 33.6 171.6 34.8 ;
      RECT  175.2 33.6 176.4 34.8 ;
      RECT  180.0 33.6 181.2 34.8 ;
      RECT  184.8 33.6 186.0 34.8 ;
      RECT  189.6 33.6 190.8 34.8 ;
      RECT  194.4 33.6 195.6 34.8 ;
      RECT  199.2 33.6 200.4 34.8 ;
      RECT  204.0 33.6 205.2 34.8 ;
      RECT  208.8 33.6 210.0 34.8 ;
      RECT  213.6 33.6 214.8 34.8 ;
      RECT  218.4 33.6 219.6 34.8 ;
      RECT  223.2 33.6 224.4 34.8 ;
      RECT  2.4 38.4 3.6 39.6 ;
      RECT  7.2 38.4 8.4 39.6 ;
      RECT  12.0 38.4 13.2 39.6 ;
      RECT  16.8 38.4 18.0 39.6 ;
      RECT  21.6 38.4 22.8 39.6 ;
      RECT  26.4 38.4 27.6 39.6 ;
      RECT  31.2 38.4 32.4 39.6 ;
      RECT  36.0 38.4 37.2 39.6 ;
      RECT  40.8 38.4 42.0 39.6 ;
      RECT  60.0 38.4 61.2 39.6 ;
      RECT  64.8 38.4 66.0 39.6 ;
      RECT  69.6 38.4 70.8 39.6 ;
      RECT  74.4 38.4 75.6 39.6 ;
      RECT  79.2 38.4 80.4 39.6 ;
      RECT  84.0 38.4 85.2 39.6 ;
      RECT  88.8 38.4 90.0 39.6 ;
      RECT  93.6 38.4 94.8 39.6 ;
      RECT  98.4 38.4 99.6 39.6 ;
      RECT  103.2 38.4 104.4 39.6 ;
      RECT  108.0 38.4 109.2 39.6 ;
      RECT  112.8 38.4 114.0 39.6 ;
      RECT  117.6 38.4 118.8 39.6 ;
      RECT  122.4 38.4 123.6 39.6 ;
      RECT  127.2 38.4 128.4 39.6 ;
      RECT  132.0 38.4 133.2 39.6 ;
      RECT  136.8 38.4 138.0 39.6 ;
      RECT  141.6 38.4 142.8 39.6 ;
      RECT  146.4 38.4 147.6 39.6 ;
      RECT  151.2 38.4 152.4 39.6 ;
      RECT  156.0 38.4 157.2 39.6 ;
      RECT  160.8 38.4 162.0 39.6 ;
      RECT  165.6 38.4 166.8 39.6 ;
      RECT  170.4 38.4 171.6 39.6 ;
      RECT  175.2 38.4 176.4 39.6 ;
      RECT  180.0 38.4 181.2 39.6 ;
      RECT  184.8 38.4 186.0 39.6 ;
      RECT  189.6 38.4 190.8 39.6 ;
      RECT  194.4 38.4 195.6 39.6 ;
      RECT  199.2 38.4 200.4 39.6 ;
      RECT  204.0 38.4 205.2 39.6 ;
      RECT  208.8 38.4 210.0 39.6 ;
      RECT  213.6 38.4 214.8 39.6 ;
      RECT  218.4 38.4 219.6 39.6 ;
      RECT  223.2 38.4 224.4 39.6 ;
      RECT  2.4 43.2 3.6 44.4 ;
      RECT  7.2 43.2 8.4 44.4 ;
      RECT  12.0 43.2 13.2 44.4 ;
      RECT  16.8 43.2 18.0 44.4 ;
      RECT  21.6 43.2 22.8 44.4 ;
      RECT  26.4 43.2 27.6 44.4 ;
      RECT  31.2 43.2 32.4 44.4 ;
      RECT  36.0 43.2 37.2 44.4 ;
      RECT  40.8 43.2 42.0 44.4 ;
      RECT  45.6 43.2 46.8 44.4 ;
      RECT  50.4 43.2 51.6 44.4 ;
      RECT  55.2 43.2 56.4 44.4 ;
      RECT  60.0 43.2 61.2 44.4 ;
      RECT  64.8 43.2 66.0 44.4 ;
      RECT  69.6 43.2 70.8 44.4 ;
      RECT  74.4 43.2 75.6 44.4 ;
      RECT  79.2 43.2 80.4 44.4 ;
      RECT  84.0 43.2 85.2 44.4 ;
      RECT  88.8 43.2 90.0 44.4 ;
      RECT  93.6 43.2 94.8 44.4 ;
      RECT  98.4 43.2 99.6 44.4 ;
      RECT  103.2 43.2 104.4 44.4 ;
      RECT  108.0 43.2 109.2 44.4 ;
      RECT  112.8 43.2 114.0 44.4 ;
      RECT  117.6 43.2 118.8 44.4 ;
      RECT  122.4 43.2 123.6 44.4 ;
      RECT  127.2 43.2 128.4 44.4 ;
      RECT  132.0 43.2 133.2 44.4 ;
      RECT  136.8 43.2 138.0 44.4 ;
      RECT  141.6 43.2 142.8 44.4 ;
      RECT  146.4 43.2 147.6 44.4 ;
      RECT  151.2 43.2 152.4 44.4 ;
      RECT  156.0 43.2 157.2 44.4 ;
      RECT  160.8 43.2 162.0 44.4 ;
      RECT  165.6 43.2 166.8 44.4 ;
      RECT  170.4 43.2 171.6 44.4 ;
      RECT  175.2 43.2 176.4 44.4 ;
      RECT  180.0 43.2 181.2 44.4 ;
      RECT  184.8 43.2 186.0 44.4 ;
      RECT  189.6 43.2 190.8 44.4 ;
      RECT  194.4 43.2 195.6 44.4 ;
      RECT  199.2 43.2 200.4 44.4 ;
      RECT  204.0 43.2 205.2 44.4 ;
      RECT  208.8 43.2 210.0 44.4 ;
      RECT  213.6 43.2 214.8 44.4 ;
      RECT  218.4 43.2 219.6 44.4 ;
      RECT  223.2 43.2 224.4 44.4 ;
      RECT  2.4 48.0 3.6 49.2 ;
      RECT  7.2 48.0 8.4 49.2 ;
      RECT  12.0 48.0 13.2 49.2 ;
      RECT  16.8 48.0 18.0 49.2 ;
      RECT  21.6 48.0 22.8 49.2 ;
      RECT  26.4 48.0 27.6 49.2 ;
      RECT  31.2 48.0 32.4 49.2 ;
      RECT  36.0 48.0 37.2 49.2 ;
      RECT  40.8 48.0 42.0 49.2 ;
      RECT  45.6 48.0 46.8 49.2 ;
      RECT  50.4 48.0 51.6 49.2 ;
      RECT  55.2 48.0 56.4 49.2 ;
      RECT  60.0 48.0 61.2 49.2 ;
      RECT  64.8 48.0 66.0 49.2 ;
      RECT  69.6 48.0 70.8 49.2 ;
      RECT  74.4 48.0 75.6 49.2 ;
      RECT  79.2 48.0 80.4 49.2 ;
      RECT  84.0 48.0 85.2 49.2 ;
      RECT  88.8 48.0 90.0 49.2 ;
      RECT  93.6 48.0 94.8 49.2 ;
      RECT  98.4 48.0 99.6 49.2 ;
      RECT  103.2 48.0 104.4 49.2 ;
      RECT  108.0 48.0 109.2 49.2 ;
      RECT  112.8 48.0 114.0 49.2 ;
      RECT  117.6 48.0 118.8 49.2 ;
      RECT  122.4 48.0 123.6 49.2 ;
      RECT  127.2 48.0 128.4 49.2 ;
      RECT  132.0 48.0 133.2 49.2 ;
      RECT  136.8 48.0 138.0 49.2 ;
      RECT  141.6 48.0 142.8 49.2 ;
      RECT  146.4 48.0 147.6 49.2 ;
      RECT  151.2 48.0 152.4 49.2 ;
      RECT  156.0 48.0 157.2 49.2 ;
      RECT  160.8 48.0 162.0 49.2 ;
      RECT  165.6 48.0 166.8 49.2 ;
      RECT  170.4 48.0 171.6 49.2 ;
      RECT  175.2 48.0 176.4 49.2 ;
      RECT  180.0 48.0 181.2 49.2 ;
      RECT  184.8 48.0 186.0 49.2 ;
      RECT  189.6 48.0 190.8 49.2 ;
      RECT  194.4 48.0 195.6 49.2 ;
      RECT  199.2 48.0 200.4 49.2 ;
      RECT  204.0 48.0 205.2 49.2 ;
      RECT  208.8 48.0 210.0 49.2 ;
      RECT  213.6 48.0 214.8 49.2 ;
      RECT  218.4 48.0 219.6 49.2 ;
      RECT  223.2 48.0 224.4 49.2 ;
      RECT  2.4 52.8 3.6 54.0 ;
      RECT  7.2 52.8 8.4 54.0 ;
      RECT  12.0 52.8 13.2 54.0 ;
      RECT  16.8 52.8 18.0 54.0 ;
      RECT  21.6 52.8 22.8 54.0 ;
      RECT  26.4 52.8 27.6 54.0 ;
      RECT  31.2 52.8 32.4 54.0 ;
      RECT  36.0 52.8 37.2 54.0 ;
      RECT  40.8 52.8 42.0 54.0 ;
      RECT  45.6 52.8 46.8 54.0 ;
      RECT  50.4 52.8 51.6 54.0 ;
      RECT  55.2 52.8 56.4 54.0 ;
      RECT  60.0 52.8 61.2 54.0 ;
      RECT  64.8 52.8 66.0 54.0 ;
      RECT  69.6 52.8 70.8 54.0 ;
      RECT  74.4 52.8 75.6 54.0 ;
      RECT  79.2 52.8 80.4 54.0 ;
      RECT  2.4 57.6 3.6 58.8 ;
      RECT  7.2 57.6 8.4 58.8 ;
      RECT  12.0 57.6 13.2 58.8 ;
      RECT  16.8 57.6 18.0 58.8 ;
      RECT  21.6 57.6 22.8 58.8 ;
      RECT  26.4 57.6 27.6 58.8 ;
      RECT  31.2 57.6 32.4 58.8 ;
      RECT  36.0 57.6 37.2 58.8 ;
      RECT  40.8 57.6 42.0 58.8 ;
      RECT  45.6 57.6 46.8 58.8 ;
      RECT  50.4 57.6 51.6 58.8 ;
      RECT  55.2 57.6 56.4 58.8 ;
      RECT  60.0 57.6 61.2 58.8 ;
      RECT  64.8 57.6 66.0 58.8 ;
      RECT  69.6 57.6 70.8 58.8 ;
      RECT  74.4 57.6 75.6 58.8 ;
      RECT  79.2 57.6 80.4 58.8 ;
      RECT  84.0 57.6 85.2 58.8 ;
      RECT  88.8 57.6 90.0 58.8 ;
      RECT  93.6 57.6 94.8 58.8 ;
      RECT  98.4 57.6 99.6 58.8 ;
      RECT  103.2 57.6 104.4 58.8 ;
      RECT  108.0 57.6 109.2 58.8 ;
      RECT  112.8 57.6 114.0 58.8 ;
      RECT  117.6 57.6 118.8 58.8 ;
      RECT  122.4 57.6 123.6 58.8 ;
      RECT  127.2 57.6 128.4 58.8 ;
      RECT  132.0 57.6 133.2 58.8 ;
      RECT  136.8 57.6 138.0 58.8 ;
      RECT  141.6 57.6 142.8 58.8 ;
      RECT  146.4 57.6 147.6 58.8 ;
      RECT  151.2 57.6 152.4 58.8 ;
      RECT  156.0 57.6 157.2 58.8 ;
      RECT  160.8 57.6 162.0 58.8 ;
      RECT  165.6 57.6 166.8 58.8 ;
      RECT  170.4 57.6 171.6 58.8 ;
      RECT  175.2 57.6 176.4 58.8 ;
      RECT  180.0 57.6 181.2 58.8 ;
      RECT  184.8 57.6 186.0 58.8 ;
      RECT  189.6 57.6 190.8 58.8 ;
      RECT  194.4 57.6 195.6 58.8 ;
      RECT  199.2 57.6 200.4 58.8 ;
      RECT  204.0 57.6 205.2 58.8 ;
      RECT  208.8 57.6 210.0 58.8 ;
      RECT  213.6 57.6 214.8 58.8 ;
      RECT  218.4 57.6 219.6 58.8 ;
      RECT  223.2 57.6 224.4 58.8 ;
      RECT  2.4 62.4 3.6 63.6 ;
      RECT  7.2 62.4 8.4 63.6 ;
      RECT  12.0 62.4 13.2 63.6 ;
      RECT  16.8 62.4 18.0 63.6 ;
      RECT  21.6 62.4 22.8 63.6 ;
      RECT  26.4 62.4 27.6 63.6 ;
      RECT  31.2 62.4 32.4 63.6 ;
      RECT  36.0 62.4 37.2 63.6 ;
      RECT  40.8 62.4 42.0 63.6 ;
      RECT  45.6 62.4 46.8 63.6 ;
      RECT  50.4 62.4 51.6 63.6 ;
      RECT  55.2 62.4 56.4 63.6 ;
      RECT  60.0 62.4 61.2 63.6 ;
      RECT  64.8 62.4 66.0 63.6 ;
      RECT  69.6 62.4 70.8 63.6 ;
      RECT  74.4 62.4 75.6 63.6 ;
      RECT  79.2 62.4 80.4 63.6 ;
      RECT  88.8 62.4 90.0 63.6 ;
      RECT  93.6 62.4 94.8 63.6 ;
      RECT  98.4 62.4 99.6 63.6 ;
      RECT  103.2 62.4 104.4 63.6 ;
      RECT  108.0 62.4 109.2 63.6 ;
      RECT  112.8 62.4 114.0 63.6 ;
      RECT  117.6 62.4 118.8 63.6 ;
      RECT  122.4 62.4 123.6 63.6 ;
      RECT  127.2 62.4 128.4 63.6 ;
      RECT  132.0 62.4 133.2 63.6 ;
      RECT  136.8 62.4 138.0 63.6 ;
      RECT  141.6 62.4 142.8 63.6 ;
      RECT  146.4 62.4 147.6 63.6 ;
      RECT  151.2 62.4 152.4 63.6 ;
      RECT  156.0 62.4 157.2 63.6 ;
      RECT  160.8 62.4 162.0 63.6 ;
      RECT  165.6 62.4 166.8 63.6 ;
      RECT  170.4 62.4 171.6 63.6 ;
      RECT  175.2 62.4 176.4 63.6 ;
      RECT  180.0 62.4 181.2 63.6 ;
      RECT  184.8 62.4 186.0 63.6 ;
      RECT  189.6 62.4 190.8 63.6 ;
      RECT  194.4 62.4 195.6 63.6 ;
      RECT  199.2 62.4 200.4 63.6 ;
      RECT  204.0 62.4 205.2 63.6 ;
      RECT  208.8 62.4 210.0 63.6 ;
      RECT  213.6 62.4 214.8 63.6 ;
      RECT  218.4 62.4 219.6 63.6 ;
      RECT  223.2 62.4 224.4 63.6 ;
      RECT  2.4 67.2 3.6 68.4 ;
      RECT  7.2 67.2 8.4 68.4 ;
      RECT  12.0 67.2 13.2 68.4 ;
      RECT  16.8 67.2 18.0 68.4 ;
      RECT  21.6 67.2 22.8 68.4 ;
      RECT  26.4 67.2 27.6 68.4 ;
      RECT  31.2 67.2 32.4 68.4 ;
      RECT  36.0 67.2 37.2 68.4 ;
      RECT  40.8 67.2 42.0 68.4 ;
      RECT  45.6 67.2 46.8 68.4 ;
      RECT  50.4 67.2 51.6 68.4 ;
      RECT  55.2 67.2 56.4 68.4 ;
      RECT  60.0 67.2 61.2 68.4 ;
      RECT  64.8 67.2 66.0 68.4 ;
      RECT  69.6 67.2 70.8 68.4 ;
      RECT  74.4 67.2 75.6 68.4 ;
      RECT  79.2 67.2 80.4 68.4 ;
      RECT  84.0 67.2 85.2 68.4 ;
      RECT  88.8 67.2 90.0 68.4 ;
      RECT  93.6 67.2 94.8 68.4 ;
      RECT  98.4 67.2 99.6 68.4 ;
      RECT  103.2 67.2 104.4 68.4 ;
      RECT  108.0 67.2 109.2 68.4 ;
      RECT  112.8 67.2 114.0 68.4 ;
      RECT  117.6 67.2 118.8 68.4 ;
      RECT  122.4 67.2 123.6 68.4 ;
      RECT  127.2 67.2 128.4 68.4 ;
      RECT  132.0 67.2 133.2 68.4 ;
      RECT  136.8 67.2 138.0 68.4 ;
      RECT  141.6 67.2 142.8 68.4 ;
      RECT  146.4 67.2 147.6 68.4 ;
      RECT  151.2 67.2 152.4 68.4 ;
      RECT  156.0 67.2 157.2 68.4 ;
      RECT  160.8 67.2 162.0 68.4 ;
      RECT  165.6 67.2 166.8 68.4 ;
      RECT  170.4 67.2 171.6 68.4 ;
      RECT  175.2 67.2 176.4 68.4 ;
      RECT  180.0 67.2 181.2 68.4 ;
      RECT  184.8 67.2 186.0 68.4 ;
      RECT  189.6 67.2 190.8 68.4 ;
      RECT  2.4 72.0 3.6 73.2 ;
      RECT  7.2 72.0 8.4 73.2 ;
      RECT  12.0 72.0 13.2 73.2 ;
      RECT  16.8 72.0 18.0 73.2 ;
      RECT  21.6 72.0 22.8 73.2 ;
      RECT  26.4 72.0 27.6 73.2 ;
      RECT  31.2 72.0 32.4 73.2 ;
      RECT  36.0 72.0 37.2 73.2 ;
      RECT  40.8 72.0 42.0 73.2 ;
      RECT  45.6 72.0 46.8 73.2 ;
      RECT  50.4 72.0 51.6 73.2 ;
      RECT  55.2 72.0 56.4 73.2 ;
      RECT  60.0 72.0 61.2 73.2 ;
      RECT  64.8 72.0 66.0 73.2 ;
      RECT  69.6 72.0 70.8 73.2 ;
      RECT  74.4 72.0 75.6 73.2 ;
      RECT  79.2 72.0 80.4 73.2 ;
      RECT  189.6 72.0 190.8 73.2 ;
      RECT  194.4 72.0 195.6 73.2 ;
      RECT  199.2 72.0 200.4 73.2 ;
      RECT  204.0 72.0 205.2 73.2 ;
      RECT  208.8 72.0 210.0 73.2 ;
      RECT  213.6 72.0 214.8 73.2 ;
      RECT  218.4 72.0 219.6 73.2 ;
      RECT  223.2 72.0 224.4 73.2 ;
      RECT  2.4 76.8 3.6 78.0 ;
      RECT  7.2 76.8 8.4 78.0 ;
      RECT  12.0 76.8 13.2 78.0 ;
      RECT  16.8 76.8 18.0 78.0 ;
      RECT  21.6 76.8 22.8 78.0 ;
      RECT  26.4 76.8 27.6 78.0 ;
      RECT  31.2 76.8 32.4 78.0 ;
      RECT  36.0 76.8 37.2 78.0 ;
      RECT  40.8 76.8 42.0 78.0 ;
      RECT  45.6 76.8 46.8 78.0 ;
      RECT  50.4 76.8 51.6 78.0 ;
      RECT  55.2 76.8 56.4 78.0 ;
      RECT  60.0 76.8 61.2 78.0 ;
      RECT  64.8 76.8 66.0 78.0 ;
      RECT  69.6 76.8 70.8 78.0 ;
      RECT  74.4 76.8 75.6 78.0 ;
      RECT  79.2 76.8 80.4 78.0 ;
      RECT  84.0 76.8 85.2 78.0 ;
      RECT  88.8 76.8 90.0 78.0 ;
      RECT  93.6 76.8 94.8 78.0 ;
      RECT  98.4 76.8 99.6 78.0 ;
      RECT  103.2 76.8 104.4 78.0 ;
      RECT  108.0 76.8 109.2 78.0 ;
      RECT  112.8 76.8 114.0 78.0 ;
      RECT  117.6 76.8 118.8 78.0 ;
      RECT  122.4 76.8 123.6 78.0 ;
      RECT  127.2 76.8 128.4 78.0 ;
      RECT  132.0 76.8 133.2 78.0 ;
      RECT  136.8 76.8 138.0 78.0 ;
      RECT  141.6 76.8 142.8 78.0 ;
      RECT  146.4 76.8 147.6 78.0 ;
      RECT  151.2 76.8 152.4 78.0 ;
      RECT  156.0 76.8 157.2 78.0 ;
      RECT  160.8 76.8 162.0 78.0 ;
      RECT  165.6 76.8 166.8 78.0 ;
      RECT  170.4 76.8 171.6 78.0 ;
      RECT  175.2 76.8 176.4 78.0 ;
      RECT  180.0 76.8 181.2 78.0 ;
      RECT  184.8 76.8 186.0 78.0 ;
      RECT  189.6 76.8 190.8 78.0 ;
      RECT  194.4 76.8 195.6 78.0 ;
      RECT  199.2 76.8 200.4 78.0 ;
      RECT  204.0 76.8 205.2 78.0 ;
      RECT  208.8 76.8 210.0 78.0 ;
      RECT  213.6 76.8 214.8 78.0 ;
      RECT  218.4 76.8 219.6 78.0 ;
      RECT  223.2 76.8 224.4 78.0 ;
      RECT  2.4 81.6 3.6 82.8 ;
      RECT  7.2 81.6 8.4 82.8 ;
      RECT  12.0 81.6 13.2 82.8 ;
      RECT  16.8 81.6 18.0 82.8 ;
      RECT  21.6 81.6 22.8 82.8 ;
      RECT  26.4 81.6 27.6 82.8 ;
      RECT  31.2 81.6 32.4 82.8 ;
      RECT  36.0 81.6 37.2 82.8 ;
      RECT  40.8 81.6 42.0 82.8 ;
      RECT  45.6 81.6 46.8 82.8 ;
      RECT  50.4 81.6 51.6 82.8 ;
      RECT  55.2 81.6 56.4 82.8 ;
      RECT  60.0 81.6 61.2 82.8 ;
      RECT  64.8 81.6 66.0 82.8 ;
      RECT  69.6 81.6 70.8 82.8 ;
      RECT  74.4 81.6 75.6 82.8 ;
      RECT  79.2 81.6 80.4 82.8 ;
      RECT  84.0 81.6 85.2 82.8 ;
      RECT  88.8 81.6 90.0 82.8 ;
      RECT  93.6 81.6 94.8 82.8 ;
      RECT  98.4 81.6 99.6 82.8 ;
      RECT  103.2 81.6 104.4 82.8 ;
      RECT  108.0 81.6 109.2 82.8 ;
      RECT  112.8 81.6 114.0 82.8 ;
      RECT  117.6 81.6 118.8 82.8 ;
      RECT  122.4 81.6 123.6 82.8 ;
      RECT  127.2 81.6 128.4 82.8 ;
      RECT  132.0 81.6 133.2 82.8 ;
      RECT  136.8 81.6 138.0 82.8 ;
      RECT  141.6 81.6 142.8 82.8 ;
      RECT  146.4 81.6 147.6 82.8 ;
      RECT  151.2 81.6 152.4 82.8 ;
      RECT  156.0 81.6 157.2 82.8 ;
      RECT  160.8 81.6 162.0 82.8 ;
      RECT  165.6 81.6 166.8 82.8 ;
      RECT  170.4 81.6 171.6 82.8 ;
      RECT  175.2 81.6 176.4 82.8 ;
      RECT  180.0 81.6 181.2 82.8 ;
      RECT  184.8 81.6 186.0 82.8 ;
      RECT  189.6 81.6 190.8 82.8 ;
      RECT  194.4 81.6 195.6 82.8 ;
      RECT  2.4 86.4 3.6 87.6 ;
      RECT  7.2 86.4 8.4 87.6 ;
      RECT  12.0 86.4 13.2 87.6 ;
      RECT  16.8 86.4 18.0 87.6 ;
      RECT  21.6 86.4 22.8 87.6 ;
      RECT  26.4 86.4 27.6 87.6 ;
      RECT  31.2 86.4 32.4 87.6 ;
      RECT  36.0 86.4 37.2 87.6 ;
      RECT  40.8 86.4 42.0 87.6 ;
      RECT  45.6 86.4 46.8 87.6 ;
      RECT  50.4 86.4 51.6 87.6 ;
      RECT  55.2 86.4 56.4 87.6 ;
      RECT  60.0 86.4 61.2 87.6 ;
      RECT  64.8 86.4 66.0 87.6 ;
      RECT  69.6 86.4 70.8 87.6 ;
      RECT  74.4 86.4 75.6 87.6 ;
      RECT  79.2 86.4 80.4 87.6 ;
      RECT  84.0 86.4 85.2 87.6 ;
      RECT  88.8 86.4 90.0 87.6 ;
      RECT  93.6 86.4 94.8 87.6 ;
      RECT  98.4 86.4 99.6 87.6 ;
      RECT  103.2 86.4 104.4 87.6 ;
      RECT  108.0 86.4 109.2 87.6 ;
      RECT  112.8 86.4 114.0 87.6 ;
      RECT  117.6 86.4 118.8 87.6 ;
      RECT  122.4 86.4 123.6 87.6 ;
      RECT  127.2 86.4 128.4 87.6 ;
      RECT  132.0 86.4 133.2 87.6 ;
      RECT  136.8 86.4 138.0 87.6 ;
      RECT  141.6 86.4 142.8 87.6 ;
      RECT  146.4 86.4 147.6 87.6 ;
      RECT  151.2 86.4 152.4 87.6 ;
      RECT  156.0 86.4 157.2 87.6 ;
      RECT  160.8 86.4 162.0 87.6 ;
      RECT  165.6 86.4 166.8 87.6 ;
      RECT  170.4 86.4 171.6 87.6 ;
      RECT  175.2 86.4 176.4 87.6 ;
      RECT  180.0 86.4 181.2 87.6 ;
      RECT  184.8 86.4 186.0 87.6 ;
      RECT  189.6 86.4 190.8 87.6 ;
      RECT  194.4 86.4 195.6 87.6 ;
      RECT  199.2 86.4 200.4 87.6 ;
      RECT  204.0 86.4 205.2 87.6 ;
      RECT  208.8 86.4 210.0 87.6 ;
      RECT  213.6 86.4 214.8 87.6 ;
      RECT  218.4 86.4 219.6 87.6 ;
      RECT  223.2 86.4 224.4 87.6 ;
      RECT  2.4 91.2 3.6 92.4 ;
      RECT  7.2 91.2 8.4 92.4 ;
      RECT  12.0 91.2 13.2 92.4 ;
      RECT  16.8 91.2 18.0 92.4 ;
      RECT  21.6 91.2 22.8 92.4 ;
      RECT  26.4 91.2 27.6 92.4 ;
      RECT  31.2 91.2 32.4 92.4 ;
      RECT  36.0 91.2 37.2 92.4 ;
      RECT  40.8 91.2 42.0 92.4 ;
      RECT  45.6 91.2 46.8 92.4 ;
      RECT  50.4 91.2 51.6 92.4 ;
      RECT  55.2 91.2 56.4 92.4 ;
      RECT  60.0 91.2 61.2 92.4 ;
      RECT  64.8 91.2 66.0 92.4 ;
      RECT  69.6 91.2 70.8 92.4 ;
      RECT  74.4 91.2 75.6 92.4 ;
      RECT  79.2 91.2 80.4 92.4 ;
      RECT  184.8 91.2 186.0 92.4 ;
      RECT  189.6 91.2 190.8 92.4 ;
      RECT  194.4 91.2 195.6 92.4 ;
      RECT  199.2 91.2 200.4 92.4 ;
      RECT  204.0 91.2 205.2 92.4 ;
      RECT  208.8 91.2 210.0 92.4 ;
      RECT  213.6 91.2 214.8 92.4 ;
      RECT  218.4 91.2 219.6 92.4 ;
      RECT  223.2 91.2 224.4 92.4 ;
      RECT  2.4 96.0 3.6 97.2 ;
      RECT  7.2 96.0 8.4 97.2 ;
      RECT  12.0 96.0 13.2 97.2 ;
      RECT  16.8 96.0 18.0 97.2 ;
      RECT  21.6 96.0 22.8 97.2 ;
      RECT  26.4 96.0 27.6 97.2 ;
      RECT  31.2 96.0 32.4 97.2 ;
      RECT  36.0 96.0 37.2 97.2 ;
      RECT  40.8 96.0 42.0 97.2 ;
      RECT  45.6 96.0 46.8 97.2 ;
      RECT  50.4 96.0 51.6 97.2 ;
      RECT  55.2 96.0 56.4 97.2 ;
      RECT  60.0 96.0 61.2 97.2 ;
      RECT  64.8 96.0 66.0 97.2 ;
      RECT  69.6 96.0 70.8 97.2 ;
      RECT  74.4 96.0 75.6 97.2 ;
      RECT  79.2 96.0 80.4 97.2 ;
      RECT  84.0 96.0 85.2 97.2 ;
      RECT  88.8 96.0 90.0 97.2 ;
      RECT  93.6 96.0 94.8 97.2 ;
      RECT  98.4 96.0 99.6 97.2 ;
      RECT  103.2 96.0 104.4 97.2 ;
      RECT  108.0 96.0 109.2 97.2 ;
      RECT  112.8 96.0 114.0 97.2 ;
      RECT  117.6 96.0 118.8 97.2 ;
      RECT  122.4 96.0 123.6 97.2 ;
      RECT  127.2 96.0 128.4 97.2 ;
      RECT  132.0 96.0 133.2 97.2 ;
      RECT  136.8 96.0 138.0 97.2 ;
      RECT  141.6 96.0 142.8 97.2 ;
      RECT  146.4 96.0 147.6 97.2 ;
      RECT  151.2 96.0 152.4 97.2 ;
      RECT  156.0 96.0 157.2 97.2 ;
      RECT  160.8 96.0 162.0 97.2 ;
      RECT  165.6 96.0 166.8 97.2 ;
      RECT  170.4 96.0 171.6 97.2 ;
      RECT  175.2 96.0 176.4 97.2 ;
      RECT  180.0 96.0 181.2 97.2 ;
      RECT  184.8 96.0 186.0 97.2 ;
      RECT  189.6 96.0 190.8 97.2 ;
      RECT  194.4 96.0 195.6 97.2 ;
      RECT  199.2 96.0 200.4 97.2 ;
      RECT  204.0 96.0 205.2 97.2 ;
      RECT  208.8 96.0 210.0 97.2 ;
      RECT  213.6 96.0 214.8 97.2 ;
      RECT  218.4 96.0 219.6 97.2 ;
      RECT  223.2 96.0 224.4 97.2 ;
      RECT  2.4 100.8 3.6 102.0 ;
      RECT  7.2 100.8 8.4 102.0 ;
      RECT  12.0 100.8 13.2 102.0 ;
      RECT  16.8 100.8 18.0 102.0 ;
      RECT  21.6 100.8 22.8 102.0 ;
      RECT  26.4 100.8 27.6 102.0 ;
      RECT  31.2 100.8 32.4 102.0 ;
      RECT  36.0 100.8 37.2 102.0 ;
      RECT  40.8 100.8 42.0 102.0 ;
      RECT  45.6 100.8 46.8 102.0 ;
      RECT  50.4 100.8 51.6 102.0 ;
      RECT  55.2 100.8 56.4 102.0 ;
      RECT  60.0 100.8 61.2 102.0 ;
      RECT  64.8 100.8 66.0 102.0 ;
      RECT  69.6 100.8 70.8 102.0 ;
      RECT  74.4 100.8 75.6 102.0 ;
      RECT  79.2 100.8 80.4 102.0 ;
      RECT  88.8 100.8 90.0 102.0 ;
      RECT  93.6 100.8 94.8 102.0 ;
      RECT  98.4 100.8 99.6 102.0 ;
      RECT  103.2 100.8 104.4 102.0 ;
      RECT  108.0 100.8 109.2 102.0 ;
      RECT  112.8 100.8 114.0 102.0 ;
      RECT  117.6 100.8 118.8 102.0 ;
      RECT  122.4 100.8 123.6 102.0 ;
      RECT  127.2 100.8 128.4 102.0 ;
      RECT  132.0 100.8 133.2 102.0 ;
      RECT  136.8 100.8 138.0 102.0 ;
      RECT  141.6 100.8 142.8 102.0 ;
      RECT  146.4 100.8 147.6 102.0 ;
      RECT  151.2 100.8 152.4 102.0 ;
      RECT  156.0 100.8 157.2 102.0 ;
      RECT  160.8 100.8 162.0 102.0 ;
      RECT  165.6 100.8 166.8 102.0 ;
      RECT  170.4 100.8 171.6 102.0 ;
      RECT  175.2 100.8 176.4 102.0 ;
      RECT  180.0 100.8 181.2 102.0 ;
      RECT  184.8 100.8 186.0 102.0 ;
      RECT  189.6 100.8 190.8 102.0 ;
      RECT  194.4 100.8 195.6 102.0 ;
      RECT  199.2 100.8 200.4 102.0 ;
      RECT  204.0 100.8 205.2 102.0 ;
      RECT  208.8 100.8 210.0 102.0 ;
      RECT  213.6 100.8 214.8 102.0 ;
      RECT  218.4 100.8 219.6 102.0 ;
      RECT  223.2 100.8 224.4 102.0 ;
      RECT  2.4 105.6 3.6 106.8 ;
      RECT  7.2 105.6 8.4 106.8 ;
      RECT  12.0 105.6 13.2 106.8 ;
      RECT  16.8 105.6 18.0 106.8 ;
      RECT  21.6 105.6 22.8 106.8 ;
      RECT  26.4 105.6 27.6 106.8 ;
      RECT  31.2 105.6 32.4 106.8 ;
      RECT  36.0 105.6 37.2 106.8 ;
      RECT  40.8 105.6 42.0 106.8 ;
      RECT  45.6 105.6 46.8 106.8 ;
      RECT  50.4 105.6 51.6 106.8 ;
      RECT  55.2 105.6 56.4 106.8 ;
      RECT  60.0 105.6 61.2 106.8 ;
      RECT  64.8 105.6 66.0 106.8 ;
      RECT  69.6 105.6 70.8 106.8 ;
      RECT  74.4 105.6 75.6 106.8 ;
      RECT  79.2 105.6 80.4 106.8 ;
      RECT  84.0 105.6 85.2 106.8 ;
      RECT  88.8 105.6 90.0 106.8 ;
      RECT  93.6 105.6 94.8 106.8 ;
      RECT  98.4 105.6 99.6 106.8 ;
      RECT  103.2 105.6 104.4 106.8 ;
      RECT  108.0 105.6 109.2 106.8 ;
      RECT  112.8 105.6 114.0 106.8 ;
      RECT  117.6 105.6 118.8 106.8 ;
      RECT  122.4 105.6 123.6 106.8 ;
      RECT  127.2 105.6 128.4 106.8 ;
      RECT  132.0 105.6 133.2 106.8 ;
      RECT  136.8 105.6 138.0 106.8 ;
      RECT  141.6 105.6 142.8 106.8 ;
      RECT  146.4 105.6 147.6 106.8 ;
      RECT  151.2 105.6 152.4 106.8 ;
      RECT  156.0 105.6 157.2 106.8 ;
      RECT  160.8 105.6 162.0 106.8 ;
      RECT  165.6 105.6 166.8 106.8 ;
      RECT  170.4 105.6 171.6 106.8 ;
      RECT  175.2 105.6 176.4 106.8 ;
      RECT  180.0 105.6 181.2 106.8 ;
      RECT  184.8 105.6 186.0 106.8 ;
      RECT  189.6 105.6 190.8 106.8 ;
      RECT  194.4 105.6 195.6 106.8 ;
      RECT  199.2 105.6 200.4 106.8 ;
      RECT  204.0 105.6 205.2 106.8 ;
      RECT  208.8 105.6 210.0 106.8 ;
      RECT  213.6 105.6 214.8 106.8 ;
      RECT  218.4 105.6 219.6 106.8 ;
      RECT  223.2 105.6 224.4 106.8 ;
      RECT  2.4 110.4 3.6 111.6 ;
      RECT  7.2 110.4 8.4 111.6 ;
      RECT  12.0 110.4 13.2 111.6 ;
      RECT  16.8 110.4 18.0 111.6 ;
      RECT  21.6 110.4 22.8 111.6 ;
      RECT  26.4 110.4 27.6 111.6 ;
      RECT  31.2 110.4 32.4 111.6 ;
      RECT  36.0 110.4 37.2 111.6 ;
      RECT  40.8 110.4 42.0 111.6 ;
      RECT  45.6 110.4 46.8 111.6 ;
      RECT  50.4 110.4 51.6 111.6 ;
      RECT  55.2 110.4 56.4 111.6 ;
      RECT  60.0 110.4 61.2 111.6 ;
      RECT  64.8 110.4 66.0 111.6 ;
      RECT  69.6 110.4 70.8 111.6 ;
      RECT  74.4 110.4 75.6 111.6 ;
      RECT  79.2 110.4 80.4 111.6 ;
      RECT  189.6 110.4 190.8 111.6 ;
      RECT  194.4 110.4 195.6 111.6 ;
      RECT  199.2 110.4 200.4 111.6 ;
      RECT  204.0 110.4 205.2 111.6 ;
      RECT  208.8 110.4 210.0 111.6 ;
      RECT  213.6 110.4 214.8 111.6 ;
      RECT  218.4 110.4 219.6 111.6 ;
      RECT  223.2 110.4 224.4 111.6 ;
      RECT  2.4 115.2 3.6 116.4 ;
      RECT  7.2 115.2 8.4 116.4 ;
      RECT  12.0 115.2 13.2 116.4 ;
      RECT  16.8 115.2 18.0 116.4 ;
      RECT  21.6 115.2 22.8 116.4 ;
      RECT  26.4 115.2 27.6 116.4 ;
      RECT  31.2 115.2 32.4 116.4 ;
      RECT  36.0 115.2 37.2 116.4 ;
      RECT  40.8 115.2 42.0 116.4 ;
      RECT  45.6 115.2 46.8 116.4 ;
      RECT  50.4 115.2 51.6 116.4 ;
      RECT  55.2 115.2 56.4 116.4 ;
      RECT  60.0 115.2 61.2 116.4 ;
      RECT  64.8 115.2 66.0 116.4 ;
      RECT  69.6 115.2 70.8 116.4 ;
      RECT  74.4 115.2 75.6 116.4 ;
      RECT  79.2 115.2 80.4 116.4 ;
      RECT  84.0 115.2 85.2 116.4 ;
      RECT  88.8 115.2 90.0 116.4 ;
      RECT  93.6 115.2 94.8 116.4 ;
      RECT  98.4 115.2 99.6 116.4 ;
      RECT  103.2 115.2 104.4 116.4 ;
      RECT  108.0 115.2 109.2 116.4 ;
      RECT  112.8 115.2 114.0 116.4 ;
      RECT  117.6 115.2 118.8 116.4 ;
      RECT  122.4 115.2 123.6 116.4 ;
      RECT  127.2 115.2 128.4 116.4 ;
      RECT  132.0 115.2 133.2 116.4 ;
      RECT  136.8 115.2 138.0 116.4 ;
      RECT  141.6 115.2 142.8 116.4 ;
      RECT  146.4 115.2 147.6 116.4 ;
      RECT  151.2 115.2 152.4 116.4 ;
      RECT  156.0 115.2 157.2 116.4 ;
      RECT  160.8 115.2 162.0 116.4 ;
      RECT  165.6 115.2 166.8 116.4 ;
      RECT  170.4 115.2 171.6 116.4 ;
      RECT  175.2 115.2 176.4 116.4 ;
      RECT  180.0 115.2 181.2 116.4 ;
      RECT  184.8 115.2 186.0 116.4 ;
      RECT  189.6 115.2 190.8 116.4 ;
      RECT  194.4 115.2 195.6 116.4 ;
      RECT  199.2 115.2 200.4 116.4 ;
      RECT  204.0 115.2 205.2 116.4 ;
      RECT  208.8 115.2 210.0 116.4 ;
      RECT  213.6 115.2 214.8 116.4 ;
      RECT  218.4 115.2 219.6 116.4 ;
      RECT  223.2 115.2 224.4 116.4 ;
      RECT  2.4 120.0 3.6 121.2 ;
      RECT  7.2 120.0 8.4 121.2 ;
      RECT  12.0 120.0 13.2 121.2 ;
      RECT  16.8 120.0 18.0 121.2 ;
      RECT  21.6 120.0 22.8 121.2 ;
      RECT  26.4 120.0 27.6 121.2 ;
      RECT  31.2 120.0 32.4 121.2 ;
      RECT  36.0 120.0 37.2 121.2 ;
      RECT  40.8 120.0 42.0 121.2 ;
      RECT  45.6 120.0 46.8 121.2 ;
      RECT  50.4 120.0 51.6 121.2 ;
      RECT  55.2 120.0 56.4 121.2 ;
      RECT  60.0 120.0 61.2 121.2 ;
      RECT  64.8 120.0 66.0 121.2 ;
      RECT  69.6 120.0 70.8 121.2 ;
      RECT  74.4 120.0 75.6 121.2 ;
      RECT  79.2 120.0 80.4 121.2 ;
      RECT  84.0 120.0 85.2 121.2 ;
      RECT  88.8 120.0 90.0 121.2 ;
      RECT  93.6 120.0 94.8 121.2 ;
      RECT  98.4 120.0 99.6 121.2 ;
      RECT  103.2 120.0 104.4 121.2 ;
      RECT  108.0 120.0 109.2 121.2 ;
      RECT  112.8 120.0 114.0 121.2 ;
      RECT  117.6 120.0 118.8 121.2 ;
      RECT  122.4 120.0 123.6 121.2 ;
      RECT  127.2 120.0 128.4 121.2 ;
      RECT  132.0 120.0 133.2 121.2 ;
      RECT  136.8 120.0 138.0 121.2 ;
      RECT  141.6 120.0 142.8 121.2 ;
      RECT  146.4 120.0 147.6 121.2 ;
      RECT  151.2 120.0 152.4 121.2 ;
      RECT  156.0 120.0 157.2 121.2 ;
      RECT  160.8 120.0 162.0 121.2 ;
      RECT  165.6 120.0 166.8 121.2 ;
      RECT  170.4 120.0 171.6 121.2 ;
      RECT  175.2 120.0 176.4 121.2 ;
      RECT  180.0 120.0 181.2 121.2 ;
      RECT  184.8 120.0 186.0 121.2 ;
      RECT  189.6 120.0 190.8 121.2 ;
      RECT  194.4 120.0 195.6 121.2 ;
      RECT  199.2 120.0 200.4 121.2 ;
      RECT  204.0 120.0 205.2 121.2 ;
      RECT  208.8 120.0 210.0 121.2 ;
      RECT  213.6 120.0 214.8 121.2 ;
      RECT  218.4 120.0 219.6 121.2 ;
      RECT  223.2 120.0 224.4 121.2 ;
      RECT  2.4 124.8 3.6 126.0 ;
      RECT  7.2 124.8 8.4 126.0 ;
      RECT  12.0 124.8 13.2 126.0 ;
      RECT  16.8 124.8 18.0 126.0 ;
      RECT  21.6 124.8 22.8 126.0 ;
      RECT  26.4 124.8 27.6 126.0 ;
      RECT  31.2 124.8 32.4 126.0 ;
      RECT  36.0 124.8 37.2 126.0 ;
      RECT  40.8 124.8 42.0 126.0 ;
      RECT  45.6 124.8 46.8 126.0 ;
      RECT  50.4 124.8 51.6 126.0 ;
      RECT  55.2 124.8 56.4 126.0 ;
      RECT  60.0 124.8 61.2 126.0 ;
      RECT  64.8 124.8 66.0 126.0 ;
      RECT  69.6 124.8 70.8 126.0 ;
      RECT  74.4 124.8 75.6 126.0 ;
      RECT  79.2 124.8 80.4 126.0 ;
      RECT  84.0 124.8 85.2 126.0 ;
      RECT  88.8 124.8 90.0 126.0 ;
      RECT  93.6 124.8 94.8 126.0 ;
      RECT  98.4 124.8 99.6 126.0 ;
      RECT  103.2 124.8 104.4 126.0 ;
      RECT  108.0 124.8 109.2 126.0 ;
      RECT  112.8 124.8 114.0 126.0 ;
      RECT  117.6 124.8 118.8 126.0 ;
      RECT  122.4 124.8 123.6 126.0 ;
      RECT  127.2 124.8 128.4 126.0 ;
      RECT  132.0 124.8 133.2 126.0 ;
      RECT  136.8 124.8 138.0 126.0 ;
      RECT  141.6 124.8 142.8 126.0 ;
      RECT  146.4 124.8 147.6 126.0 ;
      RECT  151.2 124.8 152.4 126.0 ;
      RECT  156.0 124.8 157.2 126.0 ;
      RECT  160.8 124.8 162.0 126.0 ;
      RECT  165.6 124.8 166.8 126.0 ;
      RECT  170.4 124.8 171.6 126.0 ;
      RECT  175.2 124.8 176.4 126.0 ;
      RECT  180.0 124.8 181.2 126.0 ;
      RECT  184.8 124.8 186.0 126.0 ;
      RECT  189.6 124.8 190.8 126.0 ;
      RECT  194.4 124.8 195.6 126.0 ;
      RECT  199.2 124.8 200.4 126.0 ;
      RECT  204.0 124.8 205.2 126.0 ;
      RECT  208.8 124.8 210.0 126.0 ;
      RECT  213.6 124.8 214.8 126.0 ;
      RECT  218.4 124.8 219.6 126.0 ;
      RECT  223.2 124.8 224.4 126.0 ;
      RECT  2.4 129.6 3.6 130.8 ;
      RECT  7.2 129.6 8.4 130.8 ;
      RECT  12.0 129.6 13.2 130.8 ;
      RECT  16.8 129.6 18.0 130.8 ;
      RECT  21.6 129.6 22.8 130.8 ;
      RECT  26.4 129.6 27.6 130.8 ;
      RECT  31.2 129.6 32.4 130.8 ;
      RECT  55.2 129.6 56.4 130.8 ;
      RECT  60.0 129.6 61.2 130.8 ;
      RECT  64.8 129.6 66.0 130.8 ;
      RECT  69.6 129.6 70.8 130.8 ;
      RECT  74.4 129.6 75.6 130.8 ;
      RECT  79.2 129.6 80.4 130.8 ;
      RECT  84.0 129.6 85.2 130.8 ;
      RECT  88.8 129.6 90.0 130.8 ;
      RECT  93.6 129.6 94.8 130.8 ;
      RECT  98.4 129.6 99.6 130.8 ;
      RECT  103.2 129.6 104.4 130.8 ;
      RECT  108.0 129.6 109.2 130.8 ;
      RECT  112.8 129.6 114.0 130.8 ;
      RECT  117.6 129.6 118.8 130.8 ;
      RECT  122.4 129.6 123.6 130.8 ;
      RECT  127.2 129.6 128.4 130.8 ;
      RECT  132.0 129.6 133.2 130.8 ;
      RECT  136.8 129.6 138.0 130.8 ;
      RECT  141.6 129.6 142.8 130.8 ;
      RECT  146.4 129.6 147.6 130.8 ;
      RECT  151.2 129.6 152.4 130.8 ;
      RECT  156.0 129.6 157.2 130.8 ;
      RECT  160.8 129.6 162.0 130.8 ;
      RECT  165.6 129.6 166.8 130.8 ;
      RECT  170.4 129.6 171.6 130.8 ;
      RECT  175.2 129.6 176.4 130.8 ;
      RECT  180.0 129.6 181.2 130.8 ;
      RECT  184.8 129.6 186.0 130.8 ;
      RECT  189.6 129.6 190.8 130.8 ;
      RECT  194.4 129.6 195.6 130.8 ;
      RECT  199.2 129.6 200.4 130.8 ;
      RECT  204.0 129.6 205.2 130.8 ;
      RECT  208.8 129.6 210.0 130.8 ;
      RECT  213.6 129.6 214.8 130.8 ;
      RECT  218.4 129.6 219.6 130.8 ;
      RECT  223.2 129.6 224.4 130.8 ;
      RECT  2.4 134.4 3.6 135.6 ;
      RECT  7.2 134.4 8.4 135.6 ;
      RECT  12.0 134.4 13.2 135.6 ;
      RECT  16.8 134.4 18.0 135.6 ;
      RECT  21.6 134.4 22.8 135.6 ;
      RECT  26.4 134.4 27.6 135.6 ;
      RECT  31.2 134.4 32.4 135.6 ;
      RECT  36.0 134.4 37.2 135.6 ;
      RECT  40.8 134.4 42.0 135.6 ;
      RECT  45.6 134.4 46.8 135.6 ;
      RECT  50.4 134.4 51.6 135.6 ;
      RECT  55.2 134.4 56.4 135.6 ;
      RECT  60.0 134.4 61.2 135.6 ;
      RECT  64.8 134.4 66.0 135.6 ;
      RECT  69.6 134.4 70.8 135.6 ;
      RECT  74.4 134.4 75.6 135.6 ;
      RECT  79.2 134.4 80.4 135.6 ;
      RECT  84.0 134.4 85.2 135.6 ;
      RECT  88.8 134.4 90.0 135.6 ;
      RECT  93.6 134.4 94.8 135.6 ;
      RECT  98.4 134.4 99.6 135.6 ;
      RECT  103.2 134.4 104.4 135.6 ;
      RECT  108.0 134.4 109.2 135.6 ;
      RECT  112.8 134.4 114.0 135.6 ;
      RECT  117.6 134.4 118.8 135.6 ;
      RECT  122.4 134.4 123.6 135.6 ;
      RECT  127.2 134.4 128.4 135.6 ;
      RECT  132.0 134.4 133.2 135.6 ;
      RECT  136.8 134.4 138.0 135.6 ;
      RECT  141.6 134.4 142.8 135.6 ;
      RECT  146.4 134.4 147.6 135.6 ;
      RECT  151.2 134.4 152.4 135.6 ;
      RECT  156.0 134.4 157.2 135.6 ;
      RECT  160.8 134.4 162.0 135.6 ;
      RECT  165.6 134.4 166.8 135.6 ;
      RECT  170.4 134.4 171.6 135.6 ;
      RECT  175.2 134.4 176.4 135.6 ;
      RECT  180.0 134.4 181.2 135.6 ;
      RECT  184.8 134.4 186.0 135.6 ;
      RECT  189.6 134.4 190.8 135.6 ;
      RECT  194.4 134.4 195.6 135.6 ;
      RECT  199.2 134.4 200.4 135.6 ;
      RECT  2.4 139.2 3.6 140.4 ;
      RECT  7.2 139.2 8.4 140.4 ;
      RECT  12.0 139.2 13.2 140.4 ;
      RECT  16.8 139.2 18.0 140.4 ;
      RECT  21.6 139.2 22.8 140.4 ;
      RECT  26.4 139.2 27.6 140.4 ;
      RECT  31.2 139.2 32.4 140.4 ;
      RECT  36.0 139.2 37.2 140.4 ;
      RECT  40.8 139.2 42.0 140.4 ;
      RECT  45.6 139.2 46.8 140.4 ;
      RECT  50.4 139.2 51.6 140.4 ;
      RECT  55.2 139.2 56.4 140.4 ;
      RECT  60.0 139.2 61.2 140.4 ;
      RECT  64.8 139.2 66.0 140.4 ;
      RECT  69.6 139.2 70.8 140.4 ;
      RECT  74.4 139.2 75.6 140.4 ;
      RECT  79.2 139.2 80.4 140.4 ;
      RECT  84.0 139.2 85.2 140.4 ;
      RECT  88.8 139.2 90.0 140.4 ;
      RECT  93.6 139.2 94.8 140.4 ;
      RECT  98.4 139.2 99.6 140.4 ;
      RECT  103.2 139.2 104.4 140.4 ;
      RECT  108.0 139.2 109.2 140.4 ;
      RECT  112.8 139.2 114.0 140.4 ;
      RECT  117.6 139.2 118.8 140.4 ;
      RECT  122.4 139.2 123.6 140.4 ;
      RECT  127.2 139.2 128.4 140.4 ;
      RECT  132.0 139.2 133.2 140.4 ;
      RECT  136.8 139.2 138.0 140.4 ;
      RECT  141.6 139.2 142.8 140.4 ;
      RECT  146.4 139.2 147.6 140.4 ;
      RECT  151.2 139.2 152.4 140.4 ;
      RECT  156.0 139.2 157.2 140.4 ;
      RECT  160.8 139.2 162.0 140.4 ;
      RECT  165.6 139.2 166.8 140.4 ;
      RECT  170.4 139.2 171.6 140.4 ;
      RECT  175.2 139.2 176.4 140.4 ;
      RECT  180.0 139.2 181.2 140.4 ;
      RECT  184.8 139.2 186.0 140.4 ;
      RECT  189.6 139.2 190.8 140.4 ;
      RECT  194.4 139.2 195.6 140.4 ;
      RECT  199.2 139.2 200.4 140.4 ;
      RECT  204.0 139.2 205.2 140.4 ;
      RECT  208.8 139.2 210.0 140.4 ;
      RECT  213.6 139.2 214.8 140.4 ;
      RECT  218.4 139.2 219.6 140.4 ;
      RECT  223.2 139.2 224.4 140.4 ;
      RECT  2.4 144.0 3.6 145.2 ;
      RECT  7.2 144.0 8.4 145.2 ;
      RECT  12.0 144.0 13.2 145.2 ;
      RECT  16.8 144.0 18.0 145.2 ;
      RECT  21.6 144.0 22.8 145.2 ;
      RECT  26.4 144.0 27.6 145.2 ;
      RECT  31.2 144.0 32.4 145.2 ;
      RECT  36.0 144.0 37.2 145.2 ;
      RECT  40.8 144.0 42.0 145.2 ;
      RECT  45.6 144.0 46.8 145.2 ;
      RECT  50.4 144.0 51.6 145.2 ;
      RECT  55.2 144.0 56.4 145.2 ;
      RECT  60.0 144.0 61.2 145.2 ;
      RECT  64.8 144.0 66.0 145.2 ;
      RECT  69.6 144.0 70.8 145.2 ;
      RECT  74.4 144.0 75.6 145.2 ;
      RECT  79.2 144.0 80.4 145.2 ;
      RECT  84.0 144.0 85.2 145.2 ;
      RECT  88.8 144.0 90.0 145.2 ;
      RECT  93.6 144.0 94.8 145.2 ;
      RECT  98.4 144.0 99.6 145.2 ;
      RECT  103.2 144.0 104.4 145.2 ;
      RECT  108.0 144.0 109.2 145.2 ;
      RECT  112.8 144.0 114.0 145.2 ;
      RECT  117.6 144.0 118.8 145.2 ;
      RECT  122.4 144.0 123.6 145.2 ;
      RECT  127.2 144.0 128.4 145.2 ;
      RECT  132.0 144.0 133.2 145.2 ;
      RECT  136.8 144.0 138.0 145.2 ;
      RECT  141.6 144.0 142.8 145.2 ;
      RECT  146.4 144.0 147.6 145.2 ;
      RECT  151.2 144.0 152.4 145.2 ;
      RECT  156.0 144.0 157.2 145.2 ;
      RECT  160.8 144.0 162.0 145.2 ;
      RECT  165.6 144.0 166.8 145.2 ;
      RECT  170.4 144.0 171.6 145.2 ;
      RECT  175.2 144.0 176.4 145.2 ;
      RECT  180.0 144.0 181.2 145.2 ;
      RECT  184.8 144.0 186.0 145.2 ;
      RECT  189.6 144.0 190.8 145.2 ;
      RECT  194.4 144.0 195.6 145.2 ;
      RECT  199.2 144.0 200.4 145.2 ;
      RECT  204.0 144.0 205.2 145.2 ;
      RECT  208.8 144.0 210.0 145.2 ;
      RECT  213.6 144.0 214.8 145.2 ;
      RECT  218.4 144.0 219.6 145.2 ;
      RECT  223.2 144.0 224.4 145.2 ;
      RECT  2.4 148.8 3.6 150.0 ;
      RECT  7.2 148.8 8.4 150.0 ;
      RECT  12.0 148.8 13.2 150.0 ;
      RECT  16.8 148.8 18.0 150.0 ;
      RECT  21.6 148.8 22.8 150.0 ;
      RECT  26.4 148.8 27.6 150.0 ;
      RECT  31.2 148.8 32.4 150.0 ;
      RECT  36.0 148.8 37.2 150.0 ;
      RECT  40.8 148.8 42.0 150.0 ;
      RECT  45.6 148.8 46.8 150.0 ;
      RECT  50.4 148.8 51.6 150.0 ;
      RECT  55.2 148.8 56.4 150.0 ;
      RECT  60.0 148.8 61.2 150.0 ;
      RECT  64.8 148.8 66.0 150.0 ;
      RECT  69.6 148.8 70.8 150.0 ;
      RECT  74.4 148.8 75.6 150.0 ;
      RECT  79.2 148.8 80.4 150.0 ;
      RECT  84.0 148.8 85.2 150.0 ;
      RECT  88.8 148.8 90.0 150.0 ;
      RECT  93.6 148.8 94.8 150.0 ;
      RECT  98.4 148.8 99.6 150.0 ;
      RECT  103.2 148.8 104.4 150.0 ;
      RECT  108.0 148.8 109.2 150.0 ;
      RECT  112.8 148.8 114.0 150.0 ;
      RECT  117.6 148.8 118.8 150.0 ;
      RECT  122.4 148.8 123.6 150.0 ;
      RECT  127.2 148.8 128.4 150.0 ;
      RECT  132.0 148.8 133.2 150.0 ;
      RECT  136.8 148.8 138.0 150.0 ;
      RECT  141.6 148.8 142.8 150.0 ;
      RECT  146.4 148.8 147.6 150.0 ;
      RECT  151.2 148.8 152.4 150.0 ;
      RECT  156.0 148.8 157.2 150.0 ;
      RECT  160.8 148.8 162.0 150.0 ;
      RECT  165.6 148.8 166.8 150.0 ;
      RECT  170.4 148.8 171.6 150.0 ;
      RECT  175.2 148.8 176.4 150.0 ;
      RECT  180.0 148.8 181.2 150.0 ;
      RECT  184.8 148.8 186.0 150.0 ;
      RECT  189.6 148.8 190.8 150.0 ;
      RECT  194.4 148.8 195.6 150.0 ;
      RECT  199.2 148.8 200.4 150.0 ;
      RECT  204.0 148.8 205.2 150.0 ;
      RECT  208.8 148.8 210.0 150.0 ;
      RECT  213.6 148.8 214.8 150.0 ;
      RECT  218.4 148.8 219.6 150.0 ;
      RECT  223.2 148.8 224.4 150.0 ;
      RECT  2.4 153.6 3.6 154.8 ;
      RECT  7.2 153.6 8.4 154.8 ;
      RECT  12.0 153.6 13.2 154.8 ;
      RECT  16.8 153.6 18.0 154.8 ;
      RECT  21.6 153.6 22.8 154.8 ;
      RECT  26.4 153.6 27.6 154.8 ;
      RECT  31.2 153.6 32.4 154.8 ;
      RECT  36.0 153.6 37.2 154.8 ;
      RECT  40.8 153.6 42.0 154.8 ;
      RECT  45.6 153.6 46.8 154.8 ;
      RECT  50.4 153.6 51.6 154.8 ;
      RECT  55.2 153.6 56.4 154.8 ;
      RECT  60.0 153.6 61.2 154.8 ;
      RECT  64.8 153.6 66.0 154.8 ;
      RECT  69.6 153.6 70.8 154.8 ;
      RECT  74.4 153.6 75.6 154.8 ;
      RECT  79.2 153.6 80.4 154.8 ;
      RECT  184.8 153.6 186.0 154.8 ;
      RECT  189.6 153.6 190.8 154.8 ;
      RECT  194.4 153.6 195.6 154.8 ;
      RECT  199.2 153.6 200.4 154.8 ;
      RECT  204.0 153.6 205.2 154.8 ;
      RECT  208.8 153.6 210.0 154.8 ;
      RECT  213.6 153.6 214.8 154.8 ;
      RECT  218.4 153.6 219.6 154.8 ;
      RECT  223.2 153.6 224.4 154.8 ;
      RECT  2.4 158.4 3.6 159.6 ;
      RECT  7.2 158.4 8.4 159.6 ;
      RECT  12.0 158.4 13.2 159.6 ;
      RECT  16.8 158.4 18.0 159.6 ;
      RECT  21.6 158.4 22.8 159.6 ;
      RECT  26.4 158.4 27.6 159.6 ;
      RECT  31.2 158.4 32.4 159.6 ;
      RECT  36.0 158.4 37.2 159.6 ;
      RECT  40.8 158.4 42.0 159.6 ;
      RECT  45.6 158.4 46.8 159.6 ;
      RECT  50.4 158.4 51.6 159.6 ;
      RECT  55.2 158.4 56.4 159.6 ;
      RECT  60.0 158.4 61.2 159.6 ;
      RECT  64.8 158.4 66.0 159.6 ;
      RECT  69.6 158.4 70.8 159.6 ;
      RECT  74.4 158.4 75.6 159.6 ;
      RECT  79.2 158.4 80.4 159.6 ;
      RECT  84.0 158.4 85.2 159.6 ;
      RECT  88.8 158.4 90.0 159.6 ;
      RECT  93.6 158.4 94.8 159.6 ;
      RECT  98.4 158.4 99.6 159.6 ;
      RECT  103.2 158.4 104.4 159.6 ;
      RECT  108.0 158.4 109.2 159.6 ;
      RECT  112.8 158.4 114.0 159.6 ;
      RECT  117.6 158.4 118.8 159.6 ;
      RECT  122.4 158.4 123.6 159.6 ;
      RECT  127.2 158.4 128.4 159.6 ;
      RECT  132.0 158.4 133.2 159.6 ;
      RECT  136.8 158.4 138.0 159.6 ;
      RECT  141.6 158.4 142.8 159.6 ;
      RECT  146.4 158.4 147.6 159.6 ;
      RECT  151.2 158.4 152.4 159.6 ;
      RECT  156.0 158.4 157.2 159.6 ;
      RECT  160.8 158.4 162.0 159.6 ;
      RECT  165.6 158.4 166.8 159.6 ;
      RECT  170.4 158.4 171.6 159.6 ;
      RECT  175.2 158.4 176.4 159.6 ;
      RECT  180.0 158.4 181.2 159.6 ;
      RECT  184.8 158.4 186.0 159.6 ;
      RECT  189.6 158.4 190.8 159.6 ;
      RECT  194.4 158.4 195.6 159.6 ;
      RECT  199.2 158.4 200.4 159.6 ;
      RECT  204.0 158.4 205.2 159.6 ;
      RECT  208.8 158.4 210.0 159.6 ;
      RECT  213.6 158.4 214.8 159.6 ;
      RECT  218.4 158.4 219.6 159.6 ;
      RECT  223.2 158.4 224.4 159.6 ;
      RECT  2.4 163.2 3.6 164.4 ;
      RECT  7.2 163.2 8.4 164.4 ;
      RECT  12.0 163.2 13.2 164.4 ;
      RECT  16.8 163.2 18.0 164.4 ;
      RECT  21.6 163.2 22.8 164.4 ;
      RECT  26.4 163.2 27.6 164.4 ;
      RECT  31.2 163.2 32.4 164.4 ;
      RECT  36.0 163.2 37.2 164.4 ;
      RECT  40.8 163.2 42.0 164.4 ;
      RECT  45.6 163.2 46.8 164.4 ;
      RECT  50.4 163.2 51.6 164.4 ;
      RECT  55.2 163.2 56.4 164.4 ;
      RECT  60.0 163.2 61.2 164.4 ;
      RECT  64.8 163.2 66.0 164.4 ;
      RECT  69.6 163.2 70.8 164.4 ;
      RECT  74.4 163.2 75.6 164.4 ;
      RECT  79.2 163.2 80.4 164.4 ;
      RECT  84.0 163.2 85.2 164.4 ;
      RECT  88.8 163.2 90.0 164.4 ;
      RECT  93.6 163.2 94.8 164.4 ;
      RECT  98.4 163.2 99.6 164.4 ;
      RECT  103.2 163.2 104.4 164.4 ;
      RECT  108.0 163.2 109.2 164.4 ;
      RECT  112.8 163.2 114.0 164.4 ;
      RECT  117.6 163.2 118.8 164.4 ;
      RECT  122.4 163.2 123.6 164.4 ;
      RECT  127.2 163.2 128.4 164.4 ;
      RECT  132.0 163.2 133.2 164.4 ;
      RECT  136.8 163.2 138.0 164.4 ;
      RECT  141.6 163.2 142.8 164.4 ;
      RECT  146.4 163.2 147.6 164.4 ;
      RECT  151.2 163.2 152.4 164.4 ;
      RECT  156.0 163.2 157.2 164.4 ;
      RECT  160.8 163.2 162.0 164.4 ;
      RECT  165.6 163.2 166.8 164.4 ;
      RECT  170.4 163.2 171.6 164.4 ;
      RECT  175.2 163.2 176.4 164.4 ;
      RECT  180.0 163.2 181.2 164.4 ;
      RECT  184.8 163.2 186.0 164.4 ;
      RECT  189.6 163.2 190.8 164.4 ;
      RECT  199.2 168.0 200.4 169.2 ;
      RECT  204.0 168.0 205.2 169.2 ;
      RECT  208.8 168.0 210.0 169.2 ;
      RECT  213.6 168.0 214.8 169.2 ;
      RECT  218.4 168.0 219.6 169.2 ;
      RECT  223.2 168.0 224.4 169.2 ;
      RECT  21.6 172.8 22.8 174.0 ;
      RECT  26.4 172.8 27.6 174.0 ;
      RECT  31.2 172.8 32.4 174.0 ;
      RECT  36.0 172.8 37.2 174.0 ;
      RECT  40.8 172.8 42.0 174.0 ;
      RECT  45.6 172.8 46.8 174.0 ;
      RECT  50.4 172.8 51.6 174.0 ;
      RECT  55.2 172.8 56.4 174.0 ;
      RECT  60.0 172.8 61.2 174.0 ;
      RECT  64.8 172.8 66.0 174.0 ;
      RECT  69.6 172.8 70.8 174.0 ;
      RECT  74.4 172.8 75.6 174.0 ;
      RECT  79.2 172.8 80.4 174.0 ;
      RECT  84.0 172.8 85.2 174.0 ;
      RECT  88.8 172.8 90.0 174.0 ;
      RECT  93.6 172.8 94.8 174.0 ;
      RECT  98.4 172.8 99.6 174.0 ;
      RECT  103.2 172.8 104.4 174.0 ;
      RECT  108.0 172.8 109.2 174.0 ;
      RECT  112.8 172.8 114.0 174.0 ;
      RECT  117.6 172.8 118.8 174.0 ;
      RECT  122.4 172.8 123.6 174.0 ;
      RECT  127.2 172.8 128.4 174.0 ;
      RECT  132.0 172.8 133.2 174.0 ;
      RECT  136.8 172.8 138.0 174.0 ;
      RECT  141.6 172.8 142.8 174.0 ;
      RECT  146.4 172.8 147.6 174.0 ;
      RECT  151.2 172.8 152.4 174.0 ;
      RECT  156.0 172.8 157.2 174.0 ;
      RECT  160.8 172.8 162.0 174.0 ;
      RECT  165.6 172.8 166.8 174.0 ;
      RECT  170.4 172.8 171.6 174.0 ;
      RECT  175.2 172.8 176.4 174.0 ;
      RECT  180.0 172.8 181.2 174.0 ;
      RECT  184.8 172.8 186.0 174.0 ;
      RECT  189.6 172.8 190.8 174.0 ;
      RECT  194.4 172.8 195.6 174.0 ;
      RECT  199.2 172.8 200.4 174.0 ;
      RECT  204.0 172.8 205.2 174.0 ;
      RECT  208.8 172.8 210.0 174.0 ;
      RECT  213.6 172.8 214.8 174.0 ;
      RECT  218.4 172.8 219.6 174.0 ;
      RECT  223.2 172.8 224.4 174.0 ;
      RECT  2.4 177.6 3.6 178.8 ;
      RECT  7.2 177.6 8.4 178.8 ;
      RECT  12.0 177.6 13.2 178.8 ;
      RECT  16.8 177.6 18.0 178.8 ;
      RECT  21.6 177.6 22.8 178.8 ;
      RECT  26.4 177.6 27.6 178.8 ;
      RECT  31.2 177.6 32.4 178.8 ;
      RECT  36.0 177.6 37.2 178.8 ;
      RECT  40.8 177.6 42.0 178.8 ;
      RECT  45.6 177.6 46.8 178.8 ;
      RECT  50.4 177.6 51.6 178.8 ;
      RECT  55.2 177.6 56.4 178.8 ;
      RECT  60.0 177.6 61.2 178.8 ;
      RECT  64.8 177.6 66.0 178.8 ;
      RECT  69.6 177.6 70.8 178.8 ;
      RECT  74.4 177.6 75.6 178.8 ;
      RECT  79.2 177.6 80.4 178.8 ;
      RECT  84.0 177.6 85.2 178.8 ;
      RECT  88.8 177.6 90.0 178.8 ;
      RECT  93.6 177.6 94.8 178.8 ;
      RECT  98.4 177.6 99.6 178.8 ;
      RECT  103.2 177.6 104.4 178.8 ;
      RECT  108.0 177.6 109.2 178.8 ;
      RECT  112.8 177.6 114.0 178.8 ;
      RECT  117.6 177.6 118.8 178.8 ;
      RECT  122.4 177.6 123.6 178.8 ;
      RECT  127.2 177.6 128.4 178.8 ;
      RECT  132.0 177.6 133.2 178.8 ;
      RECT  136.8 177.6 138.0 178.8 ;
      RECT  141.6 177.6 142.8 178.8 ;
      RECT  146.4 177.6 147.6 178.8 ;
      RECT  151.2 177.6 152.4 178.8 ;
      RECT  156.0 177.6 157.2 178.8 ;
      RECT  160.8 177.6 162.0 178.8 ;
      RECT  165.6 177.6 166.8 178.8 ;
      RECT  170.4 177.6 171.6 178.8 ;
      RECT  175.2 177.6 176.4 178.8 ;
      RECT  180.0 177.6 181.2 178.8 ;
      RECT  184.8 177.6 186.0 178.8 ;
      RECT  189.6 177.6 190.8 178.8 ;
      RECT  194.4 177.6 195.6 178.8 ;
      RECT  199.2 177.6 200.4 178.8 ;
      RECT  204.0 177.6 205.2 178.8 ;
      RECT  208.8 177.6 210.0 178.8 ;
      RECT  213.6 177.6 214.8 178.8 ;
      RECT  218.4 177.6 219.6 178.8 ;
      RECT  223.2 177.6 224.4 178.8 ;
      RECT  2.4 182.4 3.6 183.6 ;
      RECT  7.2 182.4 8.4 183.6 ;
      RECT  12.0 182.4 13.2 183.6 ;
      RECT  16.8 182.4 18.0 183.6 ;
      RECT  21.6 182.4 22.8 183.6 ;
      RECT  26.4 182.4 27.6 183.6 ;
      RECT  31.2 182.4 32.4 183.6 ;
      RECT  36.0 182.4 37.2 183.6 ;
      RECT  40.8 182.4 42.0 183.6 ;
      RECT  45.6 182.4 46.8 183.6 ;
      RECT  50.4 182.4 51.6 183.6 ;
      RECT  55.2 182.4 56.4 183.6 ;
      RECT  60.0 182.4 61.2 183.6 ;
      RECT  64.8 182.4 66.0 183.6 ;
      RECT  69.6 182.4 70.8 183.6 ;
      RECT  74.4 182.4 75.6 183.6 ;
      RECT  79.2 182.4 80.4 183.6 ;
      RECT  84.0 182.4 85.2 183.6 ;
      RECT  88.8 182.4 90.0 183.6 ;
      RECT  93.6 182.4 94.8 183.6 ;
      RECT  98.4 182.4 99.6 183.6 ;
      RECT  103.2 182.4 104.4 183.6 ;
      RECT  108.0 182.4 109.2 183.6 ;
      RECT  112.8 182.4 114.0 183.6 ;
      RECT  117.6 182.4 118.8 183.6 ;
      RECT  122.4 182.4 123.6 183.6 ;
      RECT  127.2 182.4 128.4 183.6 ;
      RECT  132.0 182.4 133.2 183.6 ;
      RECT  136.8 182.4 138.0 183.6 ;
      RECT  141.6 182.4 142.8 183.6 ;
      RECT  146.4 182.4 147.6 183.6 ;
      RECT  151.2 182.4 152.4 183.6 ;
      RECT  156.0 182.4 157.2 183.6 ;
      RECT  160.8 182.4 162.0 183.6 ;
      RECT  165.6 182.4 166.8 183.6 ;
      RECT  170.4 182.4 171.6 183.6 ;
      RECT  175.2 182.4 176.4 183.6 ;
      RECT  180.0 182.4 181.2 183.6 ;
      RECT  2.4 187.2 3.6 188.4 ;
      RECT  7.2 187.2 8.4 188.4 ;
      RECT  12.0 187.2 13.2 188.4 ;
      RECT  16.8 187.2 18.0 188.4 ;
      RECT  21.6 187.2 22.8 188.4 ;
      RECT  26.4 187.2 27.6 188.4 ;
      RECT  31.2 187.2 32.4 188.4 ;
      RECT  36.0 187.2 37.2 188.4 ;
      RECT  40.8 187.2 42.0 188.4 ;
      RECT  45.6 187.2 46.8 188.4 ;
      RECT  50.4 187.2 51.6 188.4 ;
      RECT  55.2 187.2 56.4 188.4 ;
      RECT  60.0 187.2 61.2 188.4 ;
      RECT  64.8 187.2 66.0 188.4 ;
      RECT  69.6 187.2 70.8 188.4 ;
      RECT  74.4 187.2 75.6 188.4 ;
      RECT  79.2 187.2 80.4 188.4 ;
      RECT  84.0 187.2 85.2 188.4 ;
      RECT  88.8 187.2 90.0 188.4 ;
      RECT  93.6 187.2 94.8 188.4 ;
      RECT  98.4 187.2 99.6 188.4 ;
      RECT  103.2 187.2 104.4 188.4 ;
      RECT  108.0 187.2 109.2 188.4 ;
      RECT  112.8 187.2 114.0 188.4 ;
      RECT  117.6 187.2 118.8 188.4 ;
      RECT  122.4 187.2 123.6 188.4 ;
      RECT  127.2 187.2 128.4 188.4 ;
      RECT  132.0 187.2 133.2 188.4 ;
      RECT  136.8 187.2 138.0 188.4 ;
      RECT  141.6 187.2 142.8 188.4 ;
      RECT  146.4 187.2 147.6 188.4 ;
      RECT  151.2 187.2 152.4 188.4 ;
      RECT  156.0 187.2 157.2 188.4 ;
      RECT  160.8 187.2 162.0 188.4 ;
      RECT  165.6 187.2 166.8 188.4 ;
      RECT  170.4 187.2 171.6 188.4 ;
      RECT  175.2 187.2 176.4 188.4 ;
      RECT  180.0 187.2 181.2 188.4 ;
      RECT  184.8 187.2 186.0 188.4 ;
      RECT  189.6 187.2 190.8 188.4 ;
      RECT  194.4 187.2 195.6 188.4 ;
      RECT  199.2 187.2 200.4 188.4 ;
      RECT  204.0 187.2 205.2 188.4 ;
      RECT  208.8 187.2 210.0 188.4 ;
      RECT  213.6 187.2 214.8 188.4 ;
      RECT  218.4 187.2 219.6 188.4 ;
      RECT  223.2 187.2 224.4 188.4 ;
      RECT  36.0 192.0 37.2 193.2 ;
      RECT  40.8 192.0 42.0 193.2 ;
      RECT  45.6 192.0 46.8 193.2 ;
      RECT  50.4 192.0 51.6 193.2 ;
      RECT  55.2 192.0 56.4 193.2 ;
      RECT  60.0 192.0 61.2 193.2 ;
      RECT  64.8 192.0 66.0 193.2 ;
      RECT  69.6 192.0 70.8 193.2 ;
      RECT  74.4 192.0 75.6 193.2 ;
      RECT  79.2 192.0 80.4 193.2 ;
      RECT  84.0 192.0 85.2 193.2 ;
      RECT  88.8 192.0 90.0 193.2 ;
      RECT  93.6 192.0 94.8 193.2 ;
      RECT  98.4 192.0 99.6 193.2 ;
      RECT  103.2 192.0 104.4 193.2 ;
      RECT  108.0 192.0 109.2 193.2 ;
      RECT  112.8 192.0 114.0 193.2 ;
      RECT  117.6 192.0 118.8 193.2 ;
      RECT  122.4 192.0 123.6 193.2 ;
      RECT  127.2 192.0 128.4 193.2 ;
      RECT  132.0 192.0 133.2 193.2 ;
      RECT  136.8 192.0 138.0 193.2 ;
      RECT  141.6 192.0 142.8 193.2 ;
      RECT  146.4 192.0 147.6 193.2 ;
      RECT  151.2 192.0 152.4 193.2 ;
      RECT  156.0 192.0 157.2 193.2 ;
      RECT  160.8 192.0 162.0 193.2 ;
      RECT  165.6 192.0 166.8 193.2 ;
      RECT  170.4 192.0 171.6 193.2 ;
      RECT  175.2 192.0 176.4 193.2 ;
      RECT  180.0 192.0 181.2 193.2 ;
      RECT  184.8 192.0 186.0 193.2 ;
      RECT  189.6 192.0 190.8 193.2 ;
      RECT  194.4 192.0 195.6 193.2 ;
      RECT  199.2 192.0 200.4 193.2 ;
      RECT  204.0 192.0 205.2 193.2 ;
      RECT  208.8 192.0 210.0 193.2 ;
      RECT  213.6 192.0 214.8 193.2 ;
      RECT  218.4 192.0 219.6 193.2 ;
      RECT  223.2 192.0 224.4 193.2 ;
      RECT  26.4 196.8 27.6 198.0 ;
      RECT  31.2 196.8 32.4 198.0 ;
      RECT  36.0 196.8 37.2 198.0 ;
      RECT  40.8 196.8 42.0 198.0 ;
      RECT  45.6 196.8 46.8 198.0 ;
      RECT  50.4 196.8 51.6 198.0 ;
      RECT  55.2 196.8 56.4 198.0 ;
      RECT  60.0 196.8 61.2 198.0 ;
      RECT  64.8 196.8 66.0 198.0 ;
      RECT  69.6 196.8 70.8 198.0 ;
      RECT  74.4 196.8 75.6 198.0 ;
      RECT  79.2 196.8 80.4 198.0 ;
      RECT  84.0 196.8 85.2 198.0 ;
      RECT  88.8 196.8 90.0 198.0 ;
      RECT  93.6 196.8 94.8 198.0 ;
      RECT  98.4 196.8 99.6 198.0 ;
      RECT  103.2 196.8 104.4 198.0 ;
      RECT  108.0 196.8 109.2 198.0 ;
      RECT  112.8 196.8 114.0 198.0 ;
      RECT  117.6 196.8 118.8 198.0 ;
      RECT  122.4 196.8 123.6 198.0 ;
      RECT  127.2 196.8 128.4 198.0 ;
      RECT  132.0 196.8 133.2 198.0 ;
      RECT  136.8 196.8 138.0 198.0 ;
      RECT  141.6 196.8 142.8 198.0 ;
      RECT  146.4 196.8 147.6 198.0 ;
      RECT  151.2 196.8 152.4 198.0 ;
      RECT  156.0 196.8 157.2 198.0 ;
      RECT  160.8 196.8 162.0 198.0 ;
      RECT  165.6 196.8 166.8 198.0 ;
      RECT  170.4 196.8 171.6 198.0 ;
      RECT  175.2 196.8 176.4 198.0 ;
      RECT  180.0 196.8 181.2 198.0 ;
      RECT  184.8 196.8 186.0 198.0 ;
      RECT  189.6 196.8 190.8 198.0 ;
      RECT  194.4 196.8 195.6 198.0 ;
      RECT  199.2 196.8 200.4 198.0 ;
      RECT  204.0 196.8 205.2 198.0 ;
      RECT  208.8 196.8 210.0 198.0 ;
      RECT  213.6 196.8 214.8 198.0 ;
      RECT  218.4 196.8 219.6 198.0 ;
      RECT  223.2 196.8 224.4 198.0 ;
      RECT  36.0 201.6 37.2 202.8 ;
      RECT  40.8 201.6 42.0 202.8 ;
      RECT  45.6 201.6 46.8 202.8 ;
      RECT  50.4 201.6 51.6 202.8 ;
      RECT  55.2 201.6 56.4 202.8 ;
      RECT  60.0 201.6 61.2 202.8 ;
      RECT  64.8 201.6 66.0 202.8 ;
      RECT  69.6 201.6 70.8 202.8 ;
      RECT  74.4 201.6 75.6 202.8 ;
      RECT  79.2 201.6 80.4 202.8 ;
      RECT  84.0 201.6 85.2 202.8 ;
      RECT  88.8 201.6 90.0 202.8 ;
      RECT  93.6 201.6 94.8 202.8 ;
      RECT  98.4 201.6 99.6 202.8 ;
      RECT  103.2 201.6 104.4 202.8 ;
      RECT  108.0 201.6 109.2 202.8 ;
      RECT  112.8 201.6 114.0 202.8 ;
      RECT  117.6 201.6 118.8 202.8 ;
      RECT  122.4 201.6 123.6 202.8 ;
      RECT  127.2 201.6 128.4 202.8 ;
      RECT  132.0 201.6 133.2 202.8 ;
      RECT  136.8 201.6 138.0 202.8 ;
      RECT  141.6 201.6 142.8 202.8 ;
      RECT  146.4 201.6 147.6 202.8 ;
      RECT  151.2 201.6 152.4 202.8 ;
      RECT  156.0 201.6 157.2 202.8 ;
      RECT  160.8 201.6 162.0 202.8 ;
      RECT  165.6 201.6 166.8 202.8 ;
      RECT  170.4 201.6 171.6 202.8 ;
      RECT  175.2 201.6 176.4 202.8 ;
      RECT  180.0 201.6 181.2 202.8 ;
      RECT  184.8 201.6 186.0 202.8 ;
      RECT  189.6 201.6 190.8 202.8 ;
      RECT  194.4 201.6 195.6 202.8 ;
      RECT  199.2 201.6 200.4 202.8 ;
      RECT  204.0 201.6 205.2 202.8 ;
      RECT  208.8 201.6 210.0 202.8 ;
      RECT  213.6 201.6 214.8 202.8 ;
      RECT  218.4 201.6 219.6 202.8 ;
      RECT  223.2 201.6 224.4 202.8 ;
      RECT  2.4 206.4 3.6 207.6 ;
      RECT  7.2 206.4 8.4 207.6 ;
      RECT  12.0 206.4 13.2 207.6 ;
      RECT  16.8 206.4 18.0 207.6 ;
      RECT  21.6 206.4 22.8 207.6 ;
      RECT  26.4 206.4 27.6 207.6 ;
      RECT  31.2 206.4 32.4 207.6 ;
      RECT  36.0 206.4 37.2 207.6 ;
      RECT  40.8 206.4 42.0 207.6 ;
      RECT  45.6 206.4 46.8 207.6 ;
      RECT  50.4 206.4 51.6 207.6 ;
      RECT  55.2 206.4 56.4 207.6 ;
      RECT  60.0 206.4 61.2 207.6 ;
      RECT  64.8 206.4 66.0 207.6 ;
      RECT  69.6 206.4 70.8 207.6 ;
      RECT  74.4 206.4 75.6 207.6 ;
      RECT  79.2 206.4 80.4 207.6 ;
      RECT  84.0 206.4 85.2 207.6 ;
      RECT  180.0 206.4 181.2 207.6 ;
      RECT  184.8 206.4 186.0 207.6 ;
      RECT  189.6 206.4 190.8 207.6 ;
      RECT  194.4 206.4 195.6 207.6 ;
      RECT  199.2 206.4 200.4 207.6 ;
      RECT  204.0 206.4 205.2 207.6 ;
      RECT  208.8 206.4 210.0 207.6 ;
      RECT  213.6 206.4 214.8 207.6 ;
      RECT  218.4 206.4 219.6 207.6 ;
      RECT  223.2 206.4 224.4 207.6 ;
      RECT  36.0 211.2 37.2 212.4 ;
      RECT  40.8 211.2 42.0 212.4 ;
      RECT  45.6 211.2 46.8 212.4 ;
      RECT  50.4 211.2 51.6 212.4 ;
      RECT  55.2 211.2 56.4 212.4 ;
      RECT  60.0 211.2 61.2 212.4 ;
      RECT  64.8 211.2 66.0 212.4 ;
      RECT  69.6 211.2 70.8 212.4 ;
      RECT  74.4 211.2 75.6 212.4 ;
      RECT  79.2 211.2 80.4 212.4 ;
      RECT  84.0 211.2 85.2 212.4 ;
      RECT  88.8 211.2 90.0 212.4 ;
      RECT  93.6 211.2 94.8 212.4 ;
      RECT  98.4 211.2 99.6 212.4 ;
      RECT  103.2 211.2 104.4 212.4 ;
      RECT  108.0 211.2 109.2 212.4 ;
      RECT  112.8 211.2 114.0 212.4 ;
      RECT  117.6 211.2 118.8 212.4 ;
      RECT  122.4 211.2 123.6 212.4 ;
      RECT  127.2 211.2 128.4 212.4 ;
      RECT  132.0 211.2 133.2 212.4 ;
      RECT  136.8 211.2 138.0 212.4 ;
      RECT  141.6 211.2 142.8 212.4 ;
      RECT  146.4 211.2 147.6 212.4 ;
      RECT  151.2 211.2 152.4 212.4 ;
      RECT  156.0 211.2 157.2 212.4 ;
      RECT  160.8 211.2 162.0 212.4 ;
      RECT  165.6 211.2 166.8 212.4 ;
      RECT  170.4 211.2 171.6 212.4 ;
      RECT  175.2 211.2 176.4 212.4 ;
      RECT  180.0 211.2 181.2 212.4 ;
      RECT  184.8 211.2 186.0 212.4 ;
      RECT  189.6 211.2 190.8 212.4 ;
      RECT  194.4 211.2 195.6 212.4 ;
      RECT  199.2 211.2 200.4 212.4 ;
      RECT  204.0 211.2 205.2 212.4 ;
      RECT  208.8 211.2 210.0 212.4 ;
      RECT  213.6 211.2 214.8 212.4 ;
      RECT  218.4 211.2 219.6 212.4 ;
      RECT  223.2 211.2 224.4 212.4 ;
      RECT  26.4 216.0 27.6 217.2 ;
      RECT  31.2 216.0 32.4 217.2 ;
      RECT  36.0 216.0 37.2 217.2 ;
      RECT  40.8 216.0 42.0 217.2 ;
      RECT  45.6 216.0 46.8 217.2 ;
      RECT  50.4 216.0 51.6 217.2 ;
      RECT  55.2 216.0 56.4 217.2 ;
      RECT  60.0 216.0 61.2 217.2 ;
      RECT  64.8 216.0 66.0 217.2 ;
      RECT  69.6 216.0 70.8 217.2 ;
      RECT  74.4 216.0 75.6 217.2 ;
      RECT  79.2 216.0 80.4 217.2 ;
      RECT  84.0 216.0 85.2 217.2 ;
      RECT  136.8 216.0 138.0 217.2 ;
      RECT  141.6 216.0 142.8 217.2 ;
      RECT  146.4 216.0 147.6 217.2 ;
      RECT  151.2 216.0 152.4 217.2 ;
      RECT  156.0 216.0 157.2 217.2 ;
      RECT  160.8 216.0 162.0 217.2 ;
      RECT  165.6 216.0 166.8 217.2 ;
      RECT  170.4 216.0 171.6 217.2 ;
      RECT  175.2 216.0 176.4 217.2 ;
      RECT  180.0 216.0 181.2 217.2 ;
      RECT  184.8 216.0 186.0 217.2 ;
      RECT  189.6 216.0 190.8 217.2 ;
      RECT  194.4 216.0 195.6 217.2 ;
      RECT  199.2 216.0 200.4 217.2 ;
      RECT  204.0 216.0 205.2 217.2 ;
      RECT  208.8 216.0 210.0 217.2 ;
      RECT  213.6 216.0 214.8 217.2 ;
      RECT  218.4 216.0 219.6 217.2 ;
      RECT  223.2 216.0 224.4 217.2 ;
      RECT  36.0 220.8 37.2 222.0 ;
      RECT  40.8 220.8 42.0 222.0 ;
      RECT  45.6 220.8 46.8 222.0 ;
      RECT  50.4 220.8 51.6 222.0 ;
      RECT  55.2 220.8 56.4 222.0 ;
      RECT  60.0 220.8 61.2 222.0 ;
      RECT  64.8 220.8 66.0 222.0 ;
      RECT  69.6 220.8 70.8 222.0 ;
      RECT  74.4 220.8 75.6 222.0 ;
      RECT  79.2 220.8 80.4 222.0 ;
      RECT  84.0 220.8 85.2 222.0 ;
      RECT  88.8 220.8 90.0 222.0 ;
      RECT  93.6 220.8 94.8 222.0 ;
      RECT  98.4 220.8 99.6 222.0 ;
      RECT  103.2 220.8 104.4 222.0 ;
      RECT  108.0 220.8 109.2 222.0 ;
      RECT  112.8 220.8 114.0 222.0 ;
      RECT  117.6 220.8 118.8 222.0 ;
      RECT  122.4 220.8 123.6 222.0 ;
      RECT  127.2 220.8 128.4 222.0 ;
      RECT  132.0 220.8 133.2 222.0 ;
      RECT  136.8 220.8 138.0 222.0 ;
      RECT  141.6 220.8 142.8 222.0 ;
      RECT  146.4 220.8 147.6 222.0 ;
      RECT  151.2 220.8 152.4 222.0 ;
      RECT  156.0 220.8 157.2 222.0 ;
      RECT  160.8 220.8 162.0 222.0 ;
      RECT  165.6 220.8 166.8 222.0 ;
      RECT  170.4 220.8 171.6 222.0 ;
      RECT  175.2 220.8 176.4 222.0 ;
      RECT  180.0 220.8 181.2 222.0 ;
      RECT  184.8 220.8 186.0 222.0 ;
      RECT  189.6 220.8 190.8 222.0 ;
      RECT  194.4 220.8 195.6 222.0 ;
      RECT  199.2 220.8 200.4 222.0 ;
      RECT  204.0 220.8 205.2 222.0 ;
      RECT  208.8 220.8 210.0 222.0 ;
      RECT  213.6 220.8 214.8 222.0 ;
      RECT  218.4 220.8 219.6 222.0 ;
      RECT  223.2 220.8 224.4 222.0 ;
      RECT  2.4 225.6 3.6 226.8 ;
      RECT  7.2 225.6 8.4 226.8 ;
      RECT  12.0 225.6 13.2 226.8 ;
      RECT  16.8 225.6 18.0 226.8 ;
      RECT  21.6 225.6 22.8 226.8 ;
      RECT  26.4 225.6 27.6 226.8 ;
      RECT  31.2 225.6 32.4 226.8 ;
      RECT  36.0 225.6 37.2 226.8 ;
      RECT  40.8 225.6 42.0 226.8 ;
      RECT  45.6 225.6 46.8 226.8 ;
      RECT  50.4 225.6 51.6 226.8 ;
      RECT  55.2 225.6 56.4 226.8 ;
      RECT  60.0 225.6 61.2 226.8 ;
      RECT  64.8 225.6 66.0 226.8 ;
      RECT  69.6 225.6 70.8 226.8 ;
      RECT  74.4 225.6 75.6 226.8 ;
      RECT  79.2 225.6 80.4 226.8 ;
      RECT  84.0 225.6 85.2 226.8 ;
      RECT  88.8 225.6 90.0 226.8 ;
      RECT  93.6 225.6 94.8 226.8 ;
      RECT  98.4 225.6 99.6 226.8 ;
      RECT  36.0 230.4 37.2 231.6 ;
      RECT  40.8 230.4 42.0 231.6 ;
      RECT  45.6 230.4 46.8 231.6 ;
      RECT  50.4 230.4 51.6 231.6 ;
      RECT  55.2 230.4 56.4 231.6 ;
      RECT  60.0 230.4 61.2 231.6 ;
      RECT  64.8 230.4 66.0 231.6 ;
      RECT  69.6 230.4 70.8 231.6 ;
      RECT  74.4 230.4 75.6 231.6 ;
      RECT  79.2 230.4 80.4 231.6 ;
      RECT  84.0 230.4 85.2 231.6 ;
      RECT  88.8 230.4 90.0 231.6 ;
      RECT  93.6 230.4 94.8 231.6 ;
      RECT  98.4 230.4 99.6 231.6 ;
      RECT  103.2 230.4 104.4 231.6 ;
      RECT  108.0 230.4 109.2 231.6 ;
      RECT  112.8 230.4 114.0 231.6 ;
      RECT  117.6 230.4 118.8 231.6 ;
      RECT  122.4 230.4 123.6 231.6 ;
      RECT  127.2 230.4 128.4 231.6 ;
      RECT  132.0 230.4 133.2 231.6 ;
      RECT  136.8 230.4 138.0 231.6 ;
      RECT  141.6 230.4 142.8 231.6 ;
      RECT  146.4 230.4 147.6 231.6 ;
      RECT  151.2 230.4 152.4 231.6 ;
      RECT  156.0 230.4 157.2 231.6 ;
      RECT  160.8 230.4 162.0 231.6 ;
      RECT  165.6 230.4 166.8 231.6 ;
      RECT  170.4 230.4 171.6 231.6 ;
      RECT  175.2 230.4 176.4 231.6 ;
      RECT  180.0 230.4 181.2 231.6 ;
      RECT  184.8 230.4 186.0 231.6 ;
      RECT  189.6 230.4 190.8 231.6 ;
      RECT  194.4 230.4 195.6 231.6 ;
      RECT  199.2 230.4 200.4 231.6 ;
      RECT  204.0 230.4 205.2 231.6 ;
      RECT  208.8 230.4 210.0 231.6 ;
      RECT  213.6 230.4 214.8 231.6 ;
      RECT  218.4 230.4 219.6 231.6 ;
      RECT  223.2 230.4 224.4 231.6 ;
      RECT  21.6 235.2 22.8 236.4 ;
      RECT  26.4 235.2 27.6 236.4 ;
      RECT  31.2 235.2 32.4 236.4 ;
      RECT  36.0 235.2 37.2 236.4 ;
      RECT  40.8 235.2 42.0 236.4 ;
      RECT  45.6 235.2 46.8 236.4 ;
      RECT  50.4 235.2 51.6 236.4 ;
      RECT  55.2 235.2 56.4 236.4 ;
      RECT  60.0 235.2 61.2 236.4 ;
      RECT  64.8 235.2 66.0 236.4 ;
      RECT  69.6 235.2 70.8 236.4 ;
      RECT  74.4 235.2 75.6 236.4 ;
      RECT  79.2 235.2 80.4 236.4 ;
      RECT  84.0 235.2 85.2 236.4 ;
      RECT  88.8 235.2 90.0 236.4 ;
      RECT  93.6 235.2 94.8 236.4 ;
      RECT  98.4 235.2 99.6 236.4 ;
      RECT  103.2 235.2 104.4 236.4 ;
      RECT  108.0 235.2 109.2 236.4 ;
      RECT  112.8 235.2 114.0 236.4 ;
      RECT  117.6 235.2 118.8 236.4 ;
      RECT  141.6 235.2 142.8 236.4 ;
      RECT  146.4 235.2 147.6 236.4 ;
      RECT  151.2 235.2 152.4 236.4 ;
      RECT  156.0 235.2 157.2 236.4 ;
      RECT  160.8 235.2 162.0 236.4 ;
      RECT  165.6 235.2 166.8 236.4 ;
      RECT  170.4 235.2 171.6 236.4 ;
      RECT  175.2 235.2 176.4 236.4 ;
      RECT  180.0 235.2 181.2 236.4 ;
      RECT  184.8 235.2 186.0 236.4 ;
      RECT  189.6 235.2 190.8 236.4 ;
      RECT  194.4 235.2 195.6 236.4 ;
      RECT  199.2 235.2 200.4 236.4 ;
      RECT  204.0 235.2 205.2 236.4 ;
      RECT  208.8 235.2 210.0 236.4 ;
      RECT  213.6 235.2 214.8 236.4 ;
      RECT  218.4 235.2 219.6 236.4 ;
      RECT  223.2 235.2 224.4 236.4 ;
      RECT  2.4 240.0 3.6 241.2 ;
      RECT  7.2 240.0 8.4 241.2 ;
      RECT  12.0 240.0 13.2 241.2 ;
      RECT  16.8 240.0 18.0 241.2 ;
      RECT  21.6 240.0 22.8 241.2 ;
      RECT  26.4 240.0 27.6 241.2 ;
      RECT  31.2 240.0 32.4 241.2 ;
      RECT  36.0 240.0 37.2 241.2 ;
      RECT  40.8 240.0 42.0 241.2 ;
      RECT  45.6 240.0 46.8 241.2 ;
      RECT  50.4 240.0 51.6 241.2 ;
      RECT  55.2 240.0 56.4 241.2 ;
      RECT  60.0 240.0 61.2 241.2 ;
      RECT  64.8 240.0 66.0 241.2 ;
      RECT  69.6 240.0 70.8 241.2 ;
      RECT  74.4 240.0 75.6 241.2 ;
      RECT  79.2 240.0 80.4 241.2 ;
      RECT  84.0 240.0 85.2 241.2 ;
      RECT  88.8 240.0 90.0 241.2 ;
      RECT  93.6 240.0 94.8 241.2 ;
      RECT  98.4 240.0 99.6 241.2 ;
      RECT  103.2 240.0 104.4 241.2 ;
      RECT  108.0 240.0 109.2 241.2 ;
      RECT  112.8 240.0 114.0 241.2 ;
      RECT  117.6 240.0 118.8 241.2 ;
      RECT  122.4 240.0 123.6 241.2 ;
      RECT  127.2 240.0 128.4 241.2 ;
      RECT  132.0 240.0 133.2 241.2 ;
      RECT  136.8 240.0 138.0 241.2 ;
      RECT  141.6 240.0 142.8 241.2 ;
      RECT  146.4 240.0 147.6 241.2 ;
      RECT  151.2 240.0 152.4 241.2 ;
      RECT  156.0 240.0 157.2 241.2 ;
      RECT  160.8 240.0 162.0 241.2 ;
      RECT  165.6 240.0 166.8 241.2 ;
      RECT  170.4 240.0 171.6 241.2 ;
      RECT  175.2 240.0 176.4 241.2 ;
      RECT  180.0 240.0 181.2 241.2 ;
      RECT  184.8 240.0 186.0 241.2 ;
      RECT  189.6 240.0 190.8 241.2 ;
      RECT  194.4 240.0 195.6 241.2 ;
      RECT  199.2 240.0 200.4 241.2 ;
      RECT  204.0 240.0 205.2 241.2 ;
      RECT  208.8 240.0 210.0 241.2 ;
      RECT  213.6 240.0 214.8 241.2 ;
      RECT  218.4 240.0 219.6 241.2 ;
      RECT  223.2 240.0 224.4 241.2 ;
      RECT  2.4 244.8 3.6 246.0 ;
      RECT  7.2 244.8 8.4 246.0 ;
      RECT  12.0 244.8 13.2 246.0 ;
      RECT  16.8 244.8 18.0 246.0 ;
      RECT  21.6 244.8 22.8 246.0 ;
      RECT  26.4 244.8 27.6 246.0 ;
      RECT  31.2 244.8 32.4 246.0 ;
      RECT  36.0 244.8 37.2 246.0 ;
      RECT  40.8 244.8 42.0 246.0 ;
      RECT  45.6 244.8 46.8 246.0 ;
      RECT  50.4 244.8 51.6 246.0 ;
      RECT  55.2 244.8 56.4 246.0 ;
      RECT  60.0 244.8 61.2 246.0 ;
      RECT  64.8 244.8 66.0 246.0 ;
      RECT  69.6 244.8 70.8 246.0 ;
      RECT  74.4 244.8 75.6 246.0 ;
      RECT  79.2 244.8 80.4 246.0 ;
      RECT  84.0 244.8 85.2 246.0 ;
      RECT  88.8 244.8 90.0 246.0 ;
      RECT  93.6 244.8 94.8 246.0 ;
      RECT  98.4 244.8 99.6 246.0 ;
      RECT  2.4 249.6 3.6 250.8 ;
      RECT  7.2 249.6 8.4 250.8 ;
      RECT  12.0 249.6 13.2 250.8 ;
      RECT  16.8 249.6 18.0 250.8 ;
      RECT  21.6 249.6 22.8 250.8 ;
      RECT  26.4 249.6 27.6 250.8 ;
      RECT  31.2 249.6 32.4 250.8 ;
      RECT  36.0 249.6 37.2 250.8 ;
      RECT  40.8 249.6 42.0 250.8 ;
      RECT  45.6 249.6 46.8 250.8 ;
      RECT  50.4 249.6 51.6 250.8 ;
      RECT  55.2 249.6 56.4 250.8 ;
      RECT  60.0 249.6 61.2 250.8 ;
      RECT  64.8 249.6 66.0 250.8 ;
      RECT  69.6 249.6 70.8 250.8 ;
      RECT  74.4 249.6 75.6 250.8 ;
      RECT  79.2 249.6 80.4 250.8 ;
      RECT  84.0 249.6 85.2 250.8 ;
      RECT  88.8 249.6 90.0 250.8 ;
      RECT  93.6 249.6 94.8 250.8 ;
      RECT  98.4 249.6 99.6 250.8 ;
      RECT  103.2 249.6 104.4 250.8 ;
      RECT  108.0 249.6 109.2 250.8 ;
      RECT  112.8 249.6 114.0 250.8 ;
      RECT  117.6 249.6 118.8 250.8 ;
      RECT  122.4 249.6 123.6 250.8 ;
      RECT  127.2 249.6 128.4 250.8 ;
      RECT  132.0 249.6 133.2 250.8 ;
      RECT  136.8 249.6 138.0 250.8 ;
      RECT  141.6 249.6 142.8 250.8 ;
      RECT  146.4 249.6 147.6 250.8 ;
      RECT  151.2 249.6 152.4 250.8 ;
      RECT  156.0 249.6 157.2 250.8 ;
      RECT  160.8 249.6 162.0 250.8 ;
      RECT  165.6 249.6 166.8 250.8 ;
      RECT  170.4 249.6 171.6 250.8 ;
      RECT  175.2 249.6 176.4 250.8 ;
      RECT  180.0 249.6 181.2 250.8 ;
      RECT  184.8 249.6 186.0 250.8 ;
      RECT  189.6 249.6 190.8 250.8 ;
      RECT  194.4 249.6 195.6 250.8 ;
      RECT  199.2 249.6 200.4 250.8 ;
      RECT  204.0 249.6 205.2 250.8 ;
      RECT  208.8 249.6 210.0 250.8 ;
      RECT  213.6 249.6 214.8 250.8 ;
      RECT  218.4 249.6 219.6 250.8 ;
      RECT  223.2 249.6 224.4 250.8 ;
      RECT  36.0 254.4 37.2 255.6 ;
      RECT  40.8 254.4 42.0 255.6 ;
      RECT  45.6 254.4 46.8 255.6 ;
      RECT  50.4 254.4 51.6 255.6 ;
      RECT  55.2 254.4 56.4 255.6 ;
      RECT  60.0 254.4 61.2 255.6 ;
      RECT  64.8 254.4 66.0 255.6 ;
      RECT  69.6 254.4 70.8 255.6 ;
      RECT  74.4 254.4 75.6 255.6 ;
      RECT  79.2 254.4 80.4 255.6 ;
      RECT  84.0 254.4 85.2 255.6 ;
      RECT  88.8 254.4 90.0 255.6 ;
      RECT  93.6 254.4 94.8 255.6 ;
      RECT  98.4 254.4 99.6 255.6 ;
      RECT  103.2 254.4 104.4 255.6 ;
      RECT  108.0 254.4 109.2 255.6 ;
      RECT  112.8 254.4 114.0 255.6 ;
      RECT  117.6 254.4 118.8 255.6 ;
      RECT  122.4 254.4 123.6 255.6 ;
      RECT  127.2 254.4 128.4 255.6 ;
      RECT  132.0 254.4 133.2 255.6 ;
      RECT  136.8 254.4 138.0 255.6 ;
      RECT  141.6 254.4 142.8 255.6 ;
      RECT  146.4 254.4 147.6 255.6 ;
      RECT  151.2 254.4 152.4 255.6 ;
      RECT  156.0 254.4 157.2 255.6 ;
      RECT  160.8 254.4 162.0 255.6 ;
      RECT  165.6 254.4 166.8 255.6 ;
      RECT  170.4 254.4 171.6 255.6 ;
      RECT  175.2 254.4 176.4 255.6 ;
      RECT  180.0 254.4 181.2 255.6 ;
      RECT  184.8 254.4 186.0 255.6 ;
      RECT  189.6 254.4 190.8 255.6 ;
      RECT  194.4 254.4 195.6 255.6 ;
      RECT  199.2 254.4 200.4 255.6 ;
      RECT  204.0 254.4 205.2 255.6 ;
      RECT  208.8 254.4 210.0 255.6 ;
      RECT  213.6 254.4 214.8 255.6 ;
      RECT  218.4 254.4 219.6 255.6 ;
      RECT  223.2 254.4 224.4 255.6 ;
      RECT  26.4 259.2 27.6 260.4 ;
      RECT  31.2 259.2 32.4 260.4 ;
      RECT  36.0 259.2 37.2 260.4 ;
      RECT  40.8 259.2 42.0 260.4 ;
      RECT  45.6 259.2 46.8 260.4 ;
      RECT  50.4 259.2 51.6 260.4 ;
      RECT  55.2 259.2 56.4 260.4 ;
      RECT  60.0 259.2 61.2 260.4 ;
      RECT  64.8 259.2 66.0 260.4 ;
      RECT  69.6 259.2 70.8 260.4 ;
      RECT  74.4 259.2 75.6 260.4 ;
      RECT  79.2 259.2 80.4 260.4 ;
      RECT  84.0 259.2 85.2 260.4 ;
      RECT  88.8 259.2 90.0 260.4 ;
      RECT  103.2 259.2 104.4 260.4 ;
      RECT  108.0 259.2 109.2 260.4 ;
      RECT  112.8 259.2 114.0 260.4 ;
      RECT  117.6 259.2 118.8 260.4 ;
      RECT  122.4 259.2 123.6 260.4 ;
      RECT  127.2 259.2 128.4 260.4 ;
      RECT  132.0 259.2 133.2 260.4 ;
      RECT  136.8 259.2 138.0 260.4 ;
      RECT  141.6 259.2 142.8 260.4 ;
      RECT  146.4 259.2 147.6 260.4 ;
      RECT  151.2 259.2 152.4 260.4 ;
      RECT  156.0 259.2 157.2 260.4 ;
      RECT  160.8 259.2 162.0 260.4 ;
      RECT  165.6 259.2 166.8 260.4 ;
      RECT  170.4 259.2 171.6 260.4 ;
      RECT  175.2 259.2 176.4 260.4 ;
      RECT  180.0 259.2 181.2 260.4 ;
      RECT  184.8 259.2 186.0 260.4 ;
      RECT  189.6 259.2 190.8 260.4 ;
      RECT  194.4 259.2 195.6 260.4 ;
      RECT  199.2 259.2 200.4 260.4 ;
      RECT  204.0 259.2 205.2 260.4 ;
      RECT  208.8 259.2 210.0 260.4 ;
      RECT  213.6 259.2 214.8 260.4 ;
      RECT  218.4 259.2 219.6 260.4 ;
      RECT  223.2 259.2 224.4 260.4 ;
      RECT  2.4 264.0 3.6 265.2 ;
      RECT  7.2 264.0 8.4 265.2 ;
      RECT  12.0 264.0 13.2 265.2 ;
      RECT  16.8 264.0 18.0 265.2 ;
      RECT  21.6 264.0 22.8 265.2 ;
      RECT  26.4 264.0 27.6 265.2 ;
      RECT  31.2 264.0 32.4 265.2 ;
      RECT  36.0 264.0 37.2 265.2 ;
      RECT  40.8 264.0 42.0 265.2 ;
      RECT  45.6 264.0 46.8 265.2 ;
      RECT  50.4 264.0 51.6 265.2 ;
      RECT  55.2 264.0 56.4 265.2 ;
      RECT  60.0 264.0 61.2 265.2 ;
      RECT  64.8 264.0 66.0 265.2 ;
      RECT  69.6 264.0 70.8 265.2 ;
      RECT  74.4 264.0 75.6 265.2 ;
      RECT  79.2 264.0 80.4 265.2 ;
      RECT  84.0 264.0 85.2 265.2 ;
      RECT  88.8 264.0 90.0 265.2 ;
      RECT  93.6 264.0 94.8 265.2 ;
      RECT  98.4 264.0 99.6 265.2 ;
      RECT  103.2 264.0 104.4 265.2 ;
      RECT  108.0 264.0 109.2 265.2 ;
      RECT  112.8 264.0 114.0 265.2 ;
      RECT  117.6 264.0 118.8 265.2 ;
      RECT  122.4 264.0 123.6 265.2 ;
      RECT  127.2 264.0 128.4 265.2 ;
      RECT  132.0 264.0 133.2 265.2 ;
      RECT  136.8 264.0 138.0 265.2 ;
      RECT  141.6 264.0 142.8 265.2 ;
      RECT  146.4 264.0 147.6 265.2 ;
      RECT  151.2 264.0 152.4 265.2 ;
      RECT  156.0 264.0 157.2 265.2 ;
      RECT  160.8 264.0 162.0 265.2 ;
      RECT  165.6 264.0 166.8 265.2 ;
      RECT  170.4 264.0 171.6 265.2 ;
      RECT  175.2 264.0 176.4 265.2 ;
      RECT  180.0 264.0 181.2 265.2 ;
      RECT  184.8 264.0 186.0 265.2 ;
      RECT  189.6 264.0 190.8 265.2 ;
      RECT  194.4 264.0 195.6 265.2 ;
      RECT  199.2 264.0 200.4 265.2 ;
      RECT  204.0 264.0 205.2 265.2 ;
      RECT  208.8 264.0 210.0 265.2 ;
      RECT  213.6 264.0 214.8 265.2 ;
      RECT  218.4 264.0 219.6 265.2 ;
      RECT  223.2 264.0 224.4 265.2 ;
      RECT  2.4 268.8 3.6 270.0 ;
      RECT  7.2 268.8 8.4 270.0 ;
      RECT  12.0 268.8 13.2 270.0 ;
      RECT  16.8 268.8 18.0 270.0 ;
      RECT  21.6 268.8 22.8 270.0 ;
      RECT  26.4 268.8 27.6 270.0 ;
      RECT  31.2 268.8 32.4 270.0 ;
      RECT  36.0 268.8 37.2 270.0 ;
      RECT  40.8 268.8 42.0 270.0 ;
      RECT  45.6 268.8 46.8 270.0 ;
      RECT  50.4 268.8 51.6 270.0 ;
      RECT  55.2 268.8 56.4 270.0 ;
      RECT  60.0 268.8 61.2 270.0 ;
      RECT  64.8 268.8 66.0 270.0 ;
      RECT  69.6 268.8 70.8 270.0 ;
      RECT  74.4 268.8 75.6 270.0 ;
      RECT  79.2 268.8 80.4 270.0 ;
      RECT  84.0 268.8 85.2 270.0 ;
      RECT  88.8 268.8 90.0 270.0 ;
      RECT  93.6 268.8 94.8 270.0 ;
      RECT  98.4 268.8 99.6 270.0 ;
      RECT  180.0 268.8 181.2 270.0 ;
      RECT  184.8 268.8 186.0 270.0 ;
      RECT  189.6 268.8 190.8 270.0 ;
      RECT  194.4 268.8 195.6 270.0 ;
      RECT  199.2 268.8 200.4 270.0 ;
      RECT  204.0 268.8 205.2 270.0 ;
      RECT  208.8 268.8 210.0 270.0 ;
      RECT  213.6 268.8 214.8 270.0 ;
      RECT  218.4 268.8 219.6 270.0 ;
      RECT  223.2 268.8 224.4 270.0 ;
      RECT  2.4 273.6 3.6 274.8 ;
      RECT  7.2 273.6 8.4 274.8 ;
      RECT  12.0 273.6 13.2 274.8 ;
      RECT  16.8 273.6 18.0 274.8 ;
      RECT  21.6 273.6 22.8 274.8 ;
      RECT  26.4 273.6 27.6 274.8 ;
      RECT  31.2 273.6 32.4 274.8 ;
      RECT  36.0 273.6 37.2 274.8 ;
      RECT  40.8 273.6 42.0 274.8 ;
      RECT  45.6 273.6 46.8 274.8 ;
      RECT  50.4 273.6 51.6 274.8 ;
      RECT  55.2 273.6 56.4 274.8 ;
      RECT  60.0 273.6 61.2 274.8 ;
      RECT  64.8 273.6 66.0 274.8 ;
      RECT  69.6 273.6 70.8 274.8 ;
      RECT  74.4 273.6 75.6 274.8 ;
      RECT  79.2 273.6 80.4 274.8 ;
      RECT  84.0 273.6 85.2 274.8 ;
      RECT  88.8 273.6 90.0 274.8 ;
      RECT  93.6 273.6 94.8 274.8 ;
      RECT  98.4 273.6 99.6 274.8 ;
      RECT  103.2 273.6 104.4 274.8 ;
      RECT  108.0 273.6 109.2 274.8 ;
      RECT  112.8 273.6 114.0 274.8 ;
      RECT  117.6 273.6 118.8 274.8 ;
      RECT  122.4 273.6 123.6 274.8 ;
      RECT  127.2 273.6 128.4 274.8 ;
      RECT  132.0 273.6 133.2 274.8 ;
      RECT  136.8 273.6 138.0 274.8 ;
      RECT  141.6 273.6 142.8 274.8 ;
      RECT  146.4 273.6 147.6 274.8 ;
      RECT  151.2 273.6 152.4 274.8 ;
      RECT  156.0 273.6 157.2 274.8 ;
      RECT  160.8 273.6 162.0 274.8 ;
      RECT  165.6 273.6 166.8 274.8 ;
      RECT  170.4 273.6 171.6 274.8 ;
      RECT  175.2 273.6 176.4 274.8 ;
      RECT  180.0 273.6 181.2 274.8 ;
      RECT  184.8 273.6 186.0 274.8 ;
      RECT  189.6 273.6 190.8 274.8 ;
      RECT  194.4 273.6 195.6 274.8 ;
      RECT  199.2 273.6 200.4 274.8 ;
      RECT  204.0 273.6 205.2 274.8 ;
      RECT  208.8 273.6 210.0 274.8 ;
      RECT  213.6 273.6 214.8 274.8 ;
      RECT  218.4 273.6 219.6 274.8 ;
      RECT  223.2 273.6 224.4 274.8 ;
      RECT  2.4 278.4 3.6 279.6 ;
      RECT  7.2 278.4 8.4 279.6 ;
      RECT  12.0 278.4 13.2 279.6 ;
      RECT  16.8 278.4 18.0 279.6 ;
      RECT  21.6 278.4 22.8 279.6 ;
      RECT  26.4 278.4 27.6 279.6 ;
      RECT  31.2 278.4 32.4 279.6 ;
      RECT  36.0 278.4 37.2 279.6 ;
      RECT  40.8 278.4 42.0 279.6 ;
      RECT  45.6 278.4 46.8 279.6 ;
      RECT  50.4 278.4 51.6 279.6 ;
      RECT  55.2 278.4 56.4 279.6 ;
      RECT  60.0 278.4 61.2 279.6 ;
      RECT  64.8 278.4 66.0 279.6 ;
      RECT  69.6 278.4 70.8 279.6 ;
      RECT  74.4 278.4 75.6 279.6 ;
      RECT  79.2 278.4 80.4 279.6 ;
      RECT  84.0 278.4 85.2 279.6 ;
      RECT  88.8 278.4 90.0 279.6 ;
      RECT  93.6 278.4 94.8 279.6 ;
      RECT  98.4 278.4 99.6 279.6 ;
      RECT  103.2 278.4 104.4 279.6 ;
      RECT  108.0 278.4 109.2 279.6 ;
      RECT  112.8 278.4 114.0 279.6 ;
      RECT  117.6 278.4 118.8 279.6 ;
      RECT  146.4 278.4 147.6 279.6 ;
      RECT  151.2 278.4 152.4 279.6 ;
      RECT  156.0 278.4 157.2 279.6 ;
      RECT  160.8 278.4 162.0 279.6 ;
      RECT  165.6 278.4 166.8 279.6 ;
      RECT  170.4 278.4 171.6 279.6 ;
      RECT  175.2 278.4 176.4 279.6 ;
      RECT  180.0 278.4 181.2 279.6 ;
      RECT  184.8 278.4 186.0 279.6 ;
      RECT  189.6 278.4 190.8 279.6 ;
      RECT  194.4 278.4 195.6 279.6 ;
      RECT  199.2 278.4 200.4 279.6 ;
      RECT  204.0 278.4 205.2 279.6 ;
      RECT  208.8 278.4 210.0 279.6 ;
      RECT  213.6 278.4 214.8 279.6 ;
      RECT  218.4 278.4 219.6 279.6 ;
      RECT  223.2 278.4 224.4 279.6 ;
      RECT  2.4 283.2 3.6 284.4 ;
      RECT  7.2 283.2 8.4 284.4 ;
      RECT  12.0 283.2 13.2 284.4 ;
      RECT  16.8 283.2 18.0 284.4 ;
      RECT  21.6 283.2 22.8 284.4 ;
      RECT  26.4 283.2 27.6 284.4 ;
      RECT  31.2 283.2 32.4 284.4 ;
      RECT  36.0 283.2 37.2 284.4 ;
      RECT  40.8 283.2 42.0 284.4 ;
      RECT  45.6 283.2 46.8 284.4 ;
      RECT  50.4 283.2 51.6 284.4 ;
      RECT  55.2 283.2 56.4 284.4 ;
      RECT  60.0 283.2 61.2 284.4 ;
      RECT  64.8 283.2 66.0 284.4 ;
      RECT  69.6 283.2 70.8 284.4 ;
      RECT  74.4 283.2 75.6 284.4 ;
      RECT  79.2 283.2 80.4 284.4 ;
      RECT  84.0 283.2 85.2 284.4 ;
      RECT  88.8 283.2 90.0 284.4 ;
      RECT  93.6 283.2 94.8 284.4 ;
      RECT  98.4 283.2 99.6 284.4 ;
      RECT  103.2 283.2 104.4 284.4 ;
      RECT  108.0 283.2 109.2 284.4 ;
      RECT  112.8 283.2 114.0 284.4 ;
      RECT  117.6 283.2 118.8 284.4 ;
      RECT  122.4 283.2 123.6 284.4 ;
      RECT  127.2 283.2 128.4 284.4 ;
      RECT  132.0 283.2 133.2 284.4 ;
      RECT  136.8 283.2 138.0 284.4 ;
      RECT  141.6 283.2 142.8 284.4 ;
      RECT  146.4 283.2 147.6 284.4 ;
      RECT  151.2 283.2 152.4 284.4 ;
      RECT  156.0 283.2 157.2 284.4 ;
      RECT  160.8 283.2 162.0 284.4 ;
      RECT  165.6 283.2 166.8 284.4 ;
      RECT  170.4 283.2 171.6 284.4 ;
      RECT  175.2 283.2 176.4 284.4 ;
      RECT  180.0 283.2 181.2 284.4 ;
      RECT  184.8 283.2 186.0 284.4 ;
      RECT  189.6 283.2 190.8 284.4 ;
      RECT  194.4 283.2 195.6 284.4 ;
      RECT  199.2 283.2 200.4 284.4 ;
      RECT  204.0 283.2 205.2 284.4 ;
      RECT  208.8 283.2 210.0 284.4 ;
      RECT  213.6 283.2 214.8 284.4 ;
      RECT  218.4 283.2 219.6 284.4 ;
      RECT  223.2 283.2 224.4 284.4 ;
      RECT  2.4 288.0 3.6 289.2 ;
      RECT  7.2 288.0 8.4 289.2 ;
      RECT  12.0 288.0 13.2 289.2 ;
      RECT  16.8 288.0 18.0 289.2 ;
      RECT  21.6 288.0 22.8 289.2 ;
      RECT  26.4 288.0 27.6 289.2 ;
      RECT  31.2 288.0 32.4 289.2 ;
      RECT  36.0 288.0 37.2 289.2 ;
      RECT  40.8 288.0 42.0 289.2 ;
      RECT  45.6 288.0 46.8 289.2 ;
      RECT  50.4 288.0 51.6 289.2 ;
      RECT  55.2 288.0 56.4 289.2 ;
      RECT  60.0 288.0 61.2 289.2 ;
      RECT  64.8 288.0 66.0 289.2 ;
      RECT  69.6 288.0 70.8 289.2 ;
      RECT  74.4 288.0 75.6 289.2 ;
      RECT  79.2 288.0 80.4 289.2 ;
      RECT  84.0 288.0 85.2 289.2 ;
      RECT  88.8 288.0 90.0 289.2 ;
      RECT  93.6 288.0 94.8 289.2 ;
      RECT  98.4 288.0 99.6 289.2 ;
      RECT  103.2 288.0 104.4 289.2 ;
      RECT  108.0 288.0 109.2 289.2 ;
      RECT  112.8 288.0 114.0 289.2 ;
      RECT  117.6 288.0 118.8 289.2 ;
      RECT  122.4 288.0 123.6 289.2 ;
      RECT  127.2 288.0 128.4 289.2 ;
      RECT  132.0 288.0 133.2 289.2 ;
      RECT  136.8 288.0 138.0 289.2 ;
      RECT  2.4 292.8 3.6 294.0 ;
      RECT  7.2 292.8 8.4 294.0 ;
      RECT  12.0 292.8 13.2 294.0 ;
      RECT  16.8 292.8 18.0 294.0 ;
      RECT  21.6 292.8 22.8 294.0 ;
      RECT  26.4 292.8 27.6 294.0 ;
      RECT  31.2 292.8 32.4 294.0 ;
      RECT  36.0 292.8 37.2 294.0 ;
      RECT  40.8 292.8 42.0 294.0 ;
      RECT  45.6 292.8 46.8 294.0 ;
      RECT  50.4 292.8 51.6 294.0 ;
      RECT  55.2 292.8 56.4 294.0 ;
      RECT  60.0 292.8 61.2 294.0 ;
      RECT  64.8 292.8 66.0 294.0 ;
      RECT  69.6 292.8 70.8 294.0 ;
      RECT  74.4 292.8 75.6 294.0 ;
      RECT  79.2 292.8 80.4 294.0 ;
      RECT  84.0 292.8 85.2 294.0 ;
      RECT  88.8 292.8 90.0 294.0 ;
      RECT  93.6 292.8 94.8 294.0 ;
      RECT  98.4 292.8 99.6 294.0 ;
      RECT  103.2 292.8 104.4 294.0 ;
      RECT  108.0 292.8 109.2 294.0 ;
      RECT  112.8 292.8 114.0 294.0 ;
      RECT  117.6 292.8 118.8 294.0 ;
      RECT  122.4 292.8 123.6 294.0 ;
      RECT  127.2 292.8 128.4 294.0 ;
      RECT  132.0 292.8 133.2 294.0 ;
      RECT  136.8 292.8 138.0 294.0 ;
      RECT  141.6 292.8 142.8 294.0 ;
      RECT  146.4 292.8 147.6 294.0 ;
      RECT  151.2 292.8 152.4 294.0 ;
      RECT  156.0 292.8 157.2 294.0 ;
      RECT  160.8 292.8 162.0 294.0 ;
      RECT  165.6 292.8 166.8 294.0 ;
      RECT  170.4 292.8 171.6 294.0 ;
      RECT  175.2 292.8 176.4 294.0 ;
      RECT  180.0 292.8 181.2 294.0 ;
      RECT  184.8 292.8 186.0 294.0 ;
      RECT  189.6 292.8 190.8 294.0 ;
      RECT  194.4 292.8 195.6 294.0 ;
      RECT  199.2 292.8 200.4 294.0 ;
      RECT  204.0 292.8 205.2 294.0 ;
      RECT  208.8 292.8 210.0 294.0 ;
      RECT  213.6 292.8 214.8 294.0 ;
      RECT  218.4 292.8 219.6 294.0 ;
      RECT  223.2 292.8 224.4 294.0 ;
      RECT  2.4 297.6 3.6 298.8 ;
      RECT  7.2 297.6 8.4 298.8 ;
      RECT  12.0 297.6 13.2 298.8 ;
      RECT  16.8 297.6 18.0 298.8 ;
      RECT  21.6 297.6 22.8 298.8 ;
      RECT  26.4 297.6 27.6 298.8 ;
      RECT  31.2 297.6 32.4 298.8 ;
      RECT  36.0 297.6 37.2 298.8 ;
      RECT  40.8 297.6 42.0 298.8 ;
      RECT  45.6 297.6 46.8 298.8 ;
      RECT  50.4 297.6 51.6 298.8 ;
      RECT  55.2 297.6 56.4 298.8 ;
      RECT  60.0 297.6 61.2 298.8 ;
      RECT  93.6 297.6 94.8 298.8 ;
      RECT  98.4 297.6 99.6 298.8 ;
      RECT  103.2 297.6 104.4 298.8 ;
      RECT  108.0 297.6 109.2 298.8 ;
      RECT  112.8 297.6 114.0 298.8 ;
      RECT  117.6 297.6 118.8 298.8 ;
      RECT  122.4 297.6 123.6 298.8 ;
      RECT  127.2 297.6 128.4 298.8 ;
      RECT  132.0 297.6 133.2 298.8 ;
      RECT  136.8 297.6 138.0 298.8 ;
      RECT  141.6 297.6 142.8 298.8 ;
      RECT  146.4 297.6 147.6 298.8 ;
      RECT  151.2 297.6 152.4 298.8 ;
      RECT  156.0 297.6 157.2 298.8 ;
      RECT  160.8 297.6 162.0 298.8 ;
      RECT  165.6 297.6 166.8 298.8 ;
      RECT  170.4 297.6 171.6 298.8 ;
      RECT  175.2 297.6 176.4 298.8 ;
      RECT  180.0 297.6 181.2 298.8 ;
      RECT  184.8 297.6 186.0 298.8 ;
      RECT  189.6 297.6 190.8 298.8 ;
      RECT  194.4 297.6 195.6 298.8 ;
      RECT  199.2 297.6 200.4 298.8 ;
      RECT  204.0 297.6 205.2 298.8 ;
      RECT  208.8 297.6 210.0 298.8 ;
      RECT  213.6 297.6 214.8 298.8 ;
      RECT  218.4 297.6 219.6 298.8 ;
      RECT  223.2 297.6 224.4 298.8 ;
      RECT  2.4 302.4 3.6 303.6 ;
      RECT  7.2 302.4 8.4 303.6 ;
      RECT  12.0 302.4 13.2 303.6 ;
      RECT  16.8 302.4 18.0 303.6 ;
      RECT  21.6 302.4 22.8 303.6 ;
      RECT  26.4 302.4 27.6 303.6 ;
      RECT  31.2 302.4 32.4 303.6 ;
      RECT  36.0 302.4 37.2 303.6 ;
      RECT  40.8 302.4 42.0 303.6 ;
      RECT  45.6 302.4 46.8 303.6 ;
      RECT  50.4 302.4 51.6 303.6 ;
      RECT  55.2 302.4 56.4 303.6 ;
      RECT  60.0 302.4 61.2 303.6 ;
      RECT  64.8 302.4 66.0 303.6 ;
      RECT  69.6 302.4 70.8 303.6 ;
      RECT  74.4 302.4 75.6 303.6 ;
      RECT  93.6 302.4 94.8 303.6 ;
      RECT  98.4 302.4 99.6 303.6 ;
      RECT  103.2 302.4 104.4 303.6 ;
      RECT  108.0 302.4 109.2 303.6 ;
      RECT  112.8 302.4 114.0 303.6 ;
      RECT  117.6 302.4 118.8 303.6 ;
      RECT  122.4 302.4 123.6 303.6 ;
      RECT  127.2 302.4 128.4 303.6 ;
      RECT  132.0 302.4 133.2 303.6 ;
      RECT  136.8 302.4 138.0 303.6 ;
      RECT  141.6 302.4 142.8 303.6 ;
      RECT  146.4 302.4 147.6 303.6 ;
      RECT  151.2 302.4 152.4 303.6 ;
      RECT  156.0 302.4 157.2 303.6 ;
      RECT  160.8 302.4 162.0 303.6 ;
      RECT  165.6 302.4 166.8 303.6 ;
      RECT  170.4 302.4 171.6 303.6 ;
      RECT  175.2 302.4 176.4 303.6 ;
      RECT  180.0 302.4 181.2 303.6 ;
      RECT  184.8 302.4 186.0 303.6 ;
      RECT  189.6 302.4 190.8 303.6 ;
      RECT  194.4 302.4 195.6 303.6 ;
      RECT  199.2 302.4 200.4 303.6 ;
      RECT  204.0 302.4 205.2 303.6 ;
      RECT  208.8 302.4 210.0 303.6 ;
      RECT  213.6 302.4 214.8 303.6 ;
      RECT  218.4 302.4 219.6 303.6 ;
      RECT  223.2 302.4 224.4 303.6 ;
      RECT  2.4 307.2 3.6 308.4 ;
      RECT  7.2 307.2 8.4 308.4 ;
      RECT  12.0 307.2 13.2 308.4 ;
      RECT  16.8 307.2 18.0 308.4 ;
      RECT  21.6 307.2 22.8 308.4 ;
      RECT  26.4 307.2 27.6 308.4 ;
      RECT  31.2 307.2 32.4 308.4 ;
      RECT  36.0 307.2 37.2 308.4 ;
      RECT  40.8 307.2 42.0 308.4 ;
      RECT  45.6 307.2 46.8 308.4 ;
      RECT  50.4 307.2 51.6 308.4 ;
      RECT  55.2 307.2 56.4 308.4 ;
      RECT  60.0 307.2 61.2 308.4 ;
      RECT  64.8 307.2 66.0 308.4 ;
      RECT  69.6 307.2 70.8 308.4 ;
      RECT  74.4 307.2 75.6 308.4 ;
      RECT  79.2 307.2 80.4 308.4 ;
      RECT  84.0 307.2 85.2 308.4 ;
      RECT  88.8 307.2 90.0 308.4 ;
      RECT  93.6 307.2 94.8 308.4 ;
      RECT  98.4 307.2 99.6 308.4 ;
      RECT  103.2 307.2 104.4 308.4 ;
      RECT  108.0 307.2 109.2 308.4 ;
      RECT  112.8 307.2 114.0 308.4 ;
      RECT  117.6 307.2 118.8 308.4 ;
      RECT  122.4 307.2 123.6 308.4 ;
      RECT  127.2 307.2 128.4 308.4 ;
      RECT  132.0 307.2 133.2 308.4 ;
      RECT  136.8 307.2 138.0 308.4 ;
      RECT  2.4 312.0 3.6 313.2 ;
      RECT  7.2 312.0 8.4 313.2 ;
      RECT  12.0 312.0 13.2 313.2 ;
      RECT  16.8 312.0 18.0 313.2 ;
      RECT  21.6 312.0 22.8 313.2 ;
      RECT  26.4 312.0 27.6 313.2 ;
      RECT  31.2 312.0 32.4 313.2 ;
      RECT  36.0 312.0 37.2 313.2 ;
      RECT  40.8 312.0 42.0 313.2 ;
      RECT  45.6 312.0 46.8 313.2 ;
      RECT  50.4 312.0 51.6 313.2 ;
      RECT  55.2 312.0 56.4 313.2 ;
      RECT  60.0 312.0 61.2 313.2 ;
      RECT  64.8 312.0 66.0 313.2 ;
      RECT  69.6 312.0 70.8 313.2 ;
      RECT  79.2 312.0 80.4 313.2 ;
      RECT  84.0 312.0 85.2 313.2 ;
      RECT  88.8 312.0 90.0 313.2 ;
      RECT  93.6 312.0 94.8 313.2 ;
      RECT  98.4 312.0 99.6 313.2 ;
      RECT  103.2 312.0 104.4 313.2 ;
      RECT  108.0 312.0 109.2 313.2 ;
      RECT  112.8 312.0 114.0 313.2 ;
      RECT  117.6 312.0 118.8 313.2 ;
      RECT  122.4 312.0 123.6 313.2 ;
      RECT  127.2 312.0 128.4 313.2 ;
      RECT  132.0 312.0 133.2 313.2 ;
      RECT  136.8 312.0 138.0 313.2 ;
      RECT  141.6 312.0 142.8 313.2 ;
      RECT  146.4 312.0 147.6 313.2 ;
      RECT  151.2 312.0 152.4 313.2 ;
      RECT  156.0 312.0 157.2 313.2 ;
      RECT  160.8 312.0 162.0 313.2 ;
      RECT  165.6 312.0 166.8 313.2 ;
      RECT  170.4 312.0 171.6 313.2 ;
      RECT  175.2 312.0 176.4 313.2 ;
      RECT  180.0 312.0 181.2 313.2 ;
      RECT  184.8 312.0 186.0 313.2 ;
      RECT  189.6 312.0 190.8 313.2 ;
      RECT  194.4 312.0 195.6 313.2 ;
      RECT  199.2 312.0 200.4 313.2 ;
      RECT  204.0 312.0 205.2 313.2 ;
      RECT  208.8 312.0 210.0 313.2 ;
      RECT  213.6 312.0 214.8 313.2 ;
      RECT  218.4 312.0 219.6 313.2 ;
      RECT  223.2 312.0 224.4 313.2 ;
      RECT  2.4 316.8 3.6 318.0 ;
      RECT  7.2 316.8 8.4 318.0 ;
      RECT  12.0 316.8 13.2 318.0 ;
      RECT  16.8 316.8 18.0 318.0 ;
      RECT  21.6 316.8 22.8 318.0 ;
      RECT  26.4 316.8 27.6 318.0 ;
      RECT  31.2 316.8 32.4 318.0 ;
      RECT  36.0 316.8 37.2 318.0 ;
      RECT  40.8 316.8 42.0 318.0 ;
      RECT  45.6 316.8 46.8 318.0 ;
      RECT  50.4 316.8 51.6 318.0 ;
      RECT  55.2 316.8 56.4 318.0 ;
      RECT  60.0 316.8 61.2 318.0 ;
      RECT  64.8 316.8 66.0 318.0 ;
      RECT  69.6 316.8 70.8 318.0 ;
      RECT  74.4 316.8 75.6 318.0 ;
      RECT  79.2 316.8 80.4 318.0 ;
      RECT  84.0 316.8 85.2 318.0 ;
      RECT  88.8 316.8 90.0 318.0 ;
      RECT  93.6 316.8 94.8 318.0 ;
      RECT  98.4 316.8 99.6 318.0 ;
      RECT  103.2 316.8 104.4 318.0 ;
      RECT  108.0 316.8 109.2 318.0 ;
      RECT  112.8 316.8 114.0 318.0 ;
      RECT  117.6 316.8 118.8 318.0 ;
      RECT  122.4 316.8 123.6 318.0 ;
      RECT  127.2 316.8 128.4 318.0 ;
      RECT  132.0 316.8 133.2 318.0 ;
      RECT  136.8 316.8 138.0 318.0 ;
      RECT  141.6 316.8 142.8 318.0 ;
      RECT  146.4 316.8 147.6 318.0 ;
      RECT  151.2 316.8 152.4 318.0 ;
      RECT  156.0 316.8 157.2 318.0 ;
      RECT  160.8 316.8 162.0 318.0 ;
      RECT  165.6 316.8 166.8 318.0 ;
      RECT  170.4 316.8 171.6 318.0 ;
      RECT  175.2 316.8 176.4 318.0 ;
      RECT  180.0 316.8 181.2 318.0 ;
      RECT  184.8 316.8 186.0 318.0 ;
      RECT  189.6 316.8 190.8 318.0 ;
      RECT  194.4 316.8 195.6 318.0 ;
      RECT  199.2 316.8 200.4 318.0 ;
      RECT  204.0 316.8 205.2 318.0 ;
      RECT  208.8 316.8 210.0 318.0 ;
      RECT  213.6 316.8 214.8 318.0 ;
      RECT  218.4 316.8 219.6 318.0 ;
      RECT  223.2 316.8 224.4 318.0 ;
      RECT  2.4 321.6 3.6 322.8 ;
      RECT  7.2 321.6 8.4 322.8 ;
      RECT  12.0 321.6 13.2 322.8 ;
      RECT  16.8 321.6 18.0 322.8 ;
      RECT  21.6 321.6 22.8 322.8 ;
      RECT  26.4 321.6 27.6 322.8 ;
      RECT  31.2 321.6 32.4 322.8 ;
      RECT  36.0 321.6 37.2 322.8 ;
      RECT  40.8 321.6 42.0 322.8 ;
      RECT  45.6 321.6 46.8 322.8 ;
      RECT  50.4 321.6 51.6 322.8 ;
      RECT  55.2 321.6 56.4 322.8 ;
      RECT  60.0 321.6 61.2 322.8 ;
      RECT  64.8 321.6 66.0 322.8 ;
      RECT  69.6 321.6 70.8 322.8 ;
      RECT  74.4 321.6 75.6 322.8 ;
      RECT  98.4 321.6 99.6 322.8 ;
      RECT  103.2 321.6 104.4 322.8 ;
      RECT  108.0 321.6 109.2 322.8 ;
      RECT  112.8 321.6 114.0 322.8 ;
      RECT  117.6 321.6 118.8 322.8 ;
      RECT  122.4 321.6 123.6 322.8 ;
      RECT  127.2 321.6 128.4 322.8 ;
      RECT  132.0 321.6 133.2 322.8 ;
      RECT  136.8 321.6 138.0 322.8 ;
      RECT  141.6 321.6 142.8 322.8 ;
      RECT  146.4 321.6 147.6 322.8 ;
      RECT  151.2 321.6 152.4 322.8 ;
      RECT  156.0 321.6 157.2 322.8 ;
      RECT  160.8 321.6 162.0 322.8 ;
      RECT  165.6 321.6 166.8 322.8 ;
      RECT  170.4 321.6 171.6 322.8 ;
      RECT  175.2 321.6 176.4 322.8 ;
      RECT  180.0 321.6 181.2 322.8 ;
      RECT  184.8 321.6 186.0 322.8 ;
      RECT  189.6 321.6 190.8 322.8 ;
      RECT  194.4 321.6 195.6 322.8 ;
      RECT  199.2 321.6 200.4 322.8 ;
      RECT  204.0 321.6 205.2 322.8 ;
      RECT  208.8 321.6 210.0 322.8 ;
      RECT  213.6 321.6 214.8 322.8 ;
      RECT  218.4 321.6 219.6 322.8 ;
      RECT  223.2 321.6 224.4 322.8 ;
      RECT  2.4 326.4 3.6 327.6 ;
      RECT  7.2 326.4 8.4 327.6 ;
      RECT  12.0 326.4 13.2 327.6 ;
      RECT  16.8 326.4 18.0 327.6 ;
      RECT  21.6 326.4 22.8 327.6 ;
      RECT  26.4 326.4 27.6 327.6 ;
      RECT  31.2 326.4 32.4 327.6 ;
      RECT  36.0 326.4 37.2 327.6 ;
      RECT  40.8 326.4 42.0 327.6 ;
      RECT  45.6 326.4 46.8 327.6 ;
      RECT  50.4 326.4 51.6 327.6 ;
      RECT  55.2 326.4 56.4 327.6 ;
      RECT  60.0 326.4 61.2 327.6 ;
      RECT  64.8 326.4 66.0 327.6 ;
      RECT  69.6 326.4 70.8 327.6 ;
      RECT  74.4 326.4 75.6 327.6 ;
      RECT  79.2 326.4 80.4 327.6 ;
      RECT  84.0 326.4 85.2 327.6 ;
      RECT  88.8 326.4 90.0 327.6 ;
      RECT  93.6 326.4 94.8 327.6 ;
      RECT  98.4 326.4 99.6 327.6 ;
      RECT  103.2 326.4 104.4 327.6 ;
      RECT  108.0 326.4 109.2 327.6 ;
      RECT  112.8 326.4 114.0 327.6 ;
      RECT  117.6 326.4 118.8 327.6 ;
      RECT  122.4 326.4 123.6 327.6 ;
      RECT  127.2 326.4 128.4 327.6 ;
      RECT  132.0 326.4 133.2 327.6 ;
      RECT  136.8 326.4 138.0 327.6 ;
      RECT  141.6 326.4 142.8 327.6 ;
      RECT  146.4 326.4 147.6 327.6 ;
      RECT  151.2 326.4 152.4 327.6 ;
      RECT  156.0 326.4 157.2 327.6 ;
      RECT  160.8 326.4 162.0 327.6 ;
      RECT  165.6 326.4 166.8 327.6 ;
      RECT  170.4 326.4 171.6 327.6 ;
      RECT  175.2 326.4 176.4 327.6 ;
      RECT  180.0 326.4 181.2 327.6 ;
      RECT  184.8 326.4 186.0 327.6 ;
      RECT  189.6 326.4 190.8 327.6 ;
      RECT  194.4 326.4 195.6 327.6 ;
      RECT  199.2 326.4 200.4 327.6 ;
      RECT  204.0 326.4 205.2 327.6 ;
      RECT  208.8 326.4 210.0 327.6 ;
      RECT  213.6 326.4 214.8 327.6 ;
      RECT  218.4 326.4 219.6 327.6 ;
      RECT  223.2 326.4 224.4 327.6 ;
      RECT  2.4 331.2 3.6 332.4 ;
      RECT  7.2 331.2 8.4 332.4 ;
      RECT  12.0 331.2 13.2 332.4 ;
      RECT  16.8 331.2 18.0 332.4 ;
      RECT  21.6 331.2 22.8 332.4 ;
      RECT  26.4 331.2 27.6 332.4 ;
      RECT  31.2 331.2 32.4 332.4 ;
      RECT  36.0 331.2 37.2 332.4 ;
      RECT  40.8 331.2 42.0 332.4 ;
      RECT  45.6 331.2 46.8 332.4 ;
      RECT  50.4 331.2 51.6 332.4 ;
      RECT  55.2 331.2 56.4 332.4 ;
      RECT  60.0 331.2 61.2 332.4 ;
      RECT  64.8 331.2 66.0 332.4 ;
      RECT  69.6 331.2 70.8 332.4 ;
      RECT  74.4 331.2 75.6 332.4 ;
      RECT  79.2 331.2 80.4 332.4 ;
      RECT  84.0 331.2 85.2 332.4 ;
      RECT  88.8 331.2 90.0 332.4 ;
      RECT  93.6 331.2 94.8 332.4 ;
      RECT  98.4 331.2 99.6 332.4 ;
      RECT  103.2 331.2 104.4 332.4 ;
      RECT  108.0 331.2 109.2 332.4 ;
      RECT  112.8 331.2 114.0 332.4 ;
      RECT  117.6 331.2 118.8 332.4 ;
      RECT  122.4 331.2 123.6 332.4 ;
      RECT  127.2 331.2 128.4 332.4 ;
      RECT  132.0 331.2 133.2 332.4 ;
      RECT  136.8 331.2 138.0 332.4 ;
      RECT  180.0 331.2 181.2 332.4 ;
      RECT  184.8 331.2 186.0 332.4 ;
      RECT  189.6 331.2 190.8 332.4 ;
      RECT  194.4 331.2 195.6 332.4 ;
      RECT  199.2 331.2 200.4 332.4 ;
      RECT  204.0 331.2 205.2 332.4 ;
      RECT  208.8 331.2 210.0 332.4 ;
      RECT  213.6 331.2 214.8 332.4 ;
      RECT  218.4 331.2 219.6 332.4 ;
      RECT  223.2 331.2 224.4 332.4 ;
      RECT  2.4 336.0 3.6 337.2 ;
      RECT  7.2 336.0 8.4 337.2 ;
      RECT  12.0 336.0 13.2 337.2 ;
      RECT  16.8 336.0 18.0 337.2 ;
      RECT  21.6 336.0 22.8 337.2 ;
      RECT  26.4 336.0 27.6 337.2 ;
      RECT  31.2 336.0 32.4 337.2 ;
      RECT  36.0 336.0 37.2 337.2 ;
      RECT  40.8 336.0 42.0 337.2 ;
      RECT  45.6 336.0 46.8 337.2 ;
      RECT  50.4 336.0 51.6 337.2 ;
      RECT  55.2 336.0 56.4 337.2 ;
      RECT  60.0 336.0 61.2 337.2 ;
      RECT  64.8 336.0 66.0 337.2 ;
      RECT  69.6 336.0 70.8 337.2 ;
      RECT  74.4 336.0 75.6 337.2 ;
      RECT  79.2 336.0 80.4 337.2 ;
      RECT  84.0 336.0 85.2 337.2 ;
      RECT  88.8 336.0 90.0 337.2 ;
      RECT  93.6 336.0 94.8 337.2 ;
      RECT  98.4 336.0 99.6 337.2 ;
      RECT  103.2 336.0 104.4 337.2 ;
      RECT  108.0 336.0 109.2 337.2 ;
      RECT  112.8 336.0 114.0 337.2 ;
      RECT  117.6 336.0 118.8 337.2 ;
      RECT  122.4 336.0 123.6 337.2 ;
      RECT  127.2 336.0 128.4 337.2 ;
      RECT  132.0 336.0 133.2 337.2 ;
      RECT  136.8 336.0 138.0 337.2 ;
      RECT  141.6 336.0 142.8 337.2 ;
      RECT  146.4 336.0 147.6 337.2 ;
      RECT  151.2 336.0 152.4 337.2 ;
      RECT  156.0 336.0 157.2 337.2 ;
      RECT  160.8 336.0 162.0 337.2 ;
      RECT  165.6 336.0 166.8 337.2 ;
      RECT  170.4 336.0 171.6 337.2 ;
      RECT  175.2 336.0 176.4 337.2 ;
      RECT  180.0 336.0 181.2 337.2 ;
      RECT  184.8 336.0 186.0 337.2 ;
      RECT  189.6 336.0 190.8 337.2 ;
      RECT  194.4 336.0 195.6 337.2 ;
      RECT  199.2 336.0 200.4 337.2 ;
      RECT  204.0 336.0 205.2 337.2 ;
      RECT  208.8 336.0 210.0 337.2 ;
      RECT  213.6 336.0 214.8 337.2 ;
      RECT  218.4 336.0 219.6 337.2 ;
      RECT  223.2 336.0 224.4 337.2 ;
      RECT  2.4 340.8 3.6 342.0 ;
      RECT  7.2 340.8 8.4 342.0 ;
      RECT  12.0 340.8 13.2 342.0 ;
      RECT  16.8 340.8 18.0 342.0 ;
      RECT  21.6 340.8 22.8 342.0 ;
      RECT  26.4 340.8 27.6 342.0 ;
      RECT  31.2 340.8 32.4 342.0 ;
      RECT  36.0 340.8 37.2 342.0 ;
      RECT  40.8 340.8 42.0 342.0 ;
      RECT  45.6 340.8 46.8 342.0 ;
      RECT  50.4 340.8 51.6 342.0 ;
      RECT  55.2 340.8 56.4 342.0 ;
      RECT  60.0 340.8 61.2 342.0 ;
      RECT  64.8 340.8 66.0 342.0 ;
      RECT  69.6 340.8 70.8 342.0 ;
      RECT  74.4 340.8 75.6 342.0 ;
      RECT  98.4 340.8 99.6 342.0 ;
      RECT  103.2 340.8 104.4 342.0 ;
      RECT  108.0 340.8 109.2 342.0 ;
      RECT  112.8 340.8 114.0 342.0 ;
      RECT  117.6 340.8 118.8 342.0 ;
      RECT  122.4 340.8 123.6 342.0 ;
      RECT  127.2 340.8 128.4 342.0 ;
      RECT  132.0 340.8 133.2 342.0 ;
      RECT  136.8 340.8 138.0 342.0 ;
      RECT  141.6 340.8 142.8 342.0 ;
      RECT  146.4 340.8 147.6 342.0 ;
      RECT  151.2 340.8 152.4 342.0 ;
      RECT  156.0 340.8 157.2 342.0 ;
      RECT  160.8 340.8 162.0 342.0 ;
      RECT  165.6 340.8 166.8 342.0 ;
      RECT  170.4 340.8 171.6 342.0 ;
      RECT  175.2 340.8 176.4 342.0 ;
      RECT  180.0 340.8 181.2 342.0 ;
      RECT  184.8 340.8 186.0 342.0 ;
      RECT  189.6 340.8 190.8 342.0 ;
      RECT  194.4 340.8 195.6 342.0 ;
      RECT  199.2 340.8 200.4 342.0 ;
      RECT  204.0 340.8 205.2 342.0 ;
      RECT  208.8 340.8 210.0 342.0 ;
      RECT  213.6 340.8 214.8 342.0 ;
      RECT  218.4 340.8 219.6 342.0 ;
      RECT  223.2 340.8 224.4 342.0 ;
      RECT  2.4 345.6 3.6 346.8 ;
      RECT  7.2 345.6 8.4 346.8 ;
      RECT  12.0 345.6 13.2 346.8 ;
      RECT  16.8 345.6 18.0 346.8 ;
      RECT  21.6 345.6 22.8 346.8 ;
      RECT  26.4 345.6 27.6 346.8 ;
      RECT  31.2 345.6 32.4 346.8 ;
      RECT  36.0 345.6 37.2 346.8 ;
      RECT  40.8 345.6 42.0 346.8 ;
      RECT  45.6 345.6 46.8 346.8 ;
      RECT  50.4 345.6 51.6 346.8 ;
      RECT  55.2 345.6 56.4 346.8 ;
      RECT  60.0 345.6 61.2 346.8 ;
      RECT  64.8 345.6 66.0 346.8 ;
      RECT  69.6 345.6 70.8 346.8 ;
      RECT  74.4 345.6 75.6 346.8 ;
      RECT  79.2 345.6 80.4 346.8 ;
      RECT  84.0 345.6 85.2 346.8 ;
      RECT  88.8 345.6 90.0 346.8 ;
      RECT  93.6 345.6 94.8 346.8 ;
      RECT  98.4 345.6 99.6 346.8 ;
      RECT  103.2 345.6 104.4 346.8 ;
      RECT  108.0 345.6 109.2 346.8 ;
      RECT  112.8 345.6 114.0 346.8 ;
      RECT  117.6 345.6 118.8 346.8 ;
      RECT  122.4 345.6 123.6 346.8 ;
      RECT  127.2 345.6 128.4 346.8 ;
      RECT  132.0 345.6 133.2 346.8 ;
      RECT  136.8 345.6 138.0 346.8 ;
      RECT  141.6 345.6 142.8 346.8 ;
      RECT  146.4 345.6 147.6 346.8 ;
      RECT  151.2 345.6 152.4 346.8 ;
      RECT  156.0 345.6 157.2 346.8 ;
      RECT  160.8 345.6 162.0 346.8 ;
      RECT  165.6 345.6 166.8 346.8 ;
      RECT  170.4 345.6 171.6 346.8 ;
      RECT  175.2 345.6 176.4 346.8 ;
      RECT  180.0 345.6 181.2 346.8 ;
      RECT  184.8 345.6 186.0 346.8 ;
      RECT  189.6 345.6 190.8 346.8 ;
      RECT  194.4 345.6 195.6 346.8 ;
      RECT  199.2 345.6 200.4 346.8 ;
      RECT  204.0 345.6 205.2 346.8 ;
      RECT  208.8 345.6 210.0 346.8 ;
      RECT  213.6 345.6 214.8 346.8 ;
      RECT  218.4 345.6 219.6 346.8 ;
      RECT  223.2 345.6 224.4 346.8 ;
      RECT  2.4 350.4 3.6 351.6 ;
      RECT  7.2 350.4 8.4 351.6 ;
      RECT  12.0 350.4 13.2 351.6 ;
      RECT  16.8 350.4 18.0 351.6 ;
      RECT  21.6 350.4 22.8 351.6 ;
      RECT  26.4 350.4 27.6 351.6 ;
      RECT  31.2 350.4 32.4 351.6 ;
      RECT  36.0 350.4 37.2 351.6 ;
      RECT  40.8 350.4 42.0 351.6 ;
      RECT  45.6 350.4 46.8 351.6 ;
      RECT  50.4 350.4 51.6 351.6 ;
      RECT  55.2 350.4 56.4 351.6 ;
      RECT  60.0 350.4 61.2 351.6 ;
      RECT  64.8 350.4 66.0 351.6 ;
      RECT  69.6 350.4 70.8 351.6 ;
      RECT  79.2 350.4 80.4 351.6 ;
      RECT  84.0 350.4 85.2 351.6 ;
      RECT  88.8 350.4 90.0 351.6 ;
      RECT  93.6 350.4 94.8 351.6 ;
      RECT  98.4 350.4 99.6 351.6 ;
      RECT  103.2 350.4 104.4 351.6 ;
      RECT  108.0 350.4 109.2 351.6 ;
      RECT  112.8 350.4 114.0 351.6 ;
      RECT  117.6 350.4 118.8 351.6 ;
      RECT  122.4 350.4 123.6 351.6 ;
      RECT  127.2 350.4 128.4 351.6 ;
      RECT  132.0 350.4 133.2 351.6 ;
      RECT  136.8 350.4 138.0 351.6 ;
      RECT  2.4 355.2 3.6 356.4 ;
      RECT  7.2 355.2 8.4 356.4 ;
      RECT  12.0 355.2 13.2 356.4 ;
      RECT  16.8 355.2 18.0 356.4 ;
      RECT  21.6 355.2 22.8 356.4 ;
      RECT  26.4 355.2 27.6 356.4 ;
      RECT  31.2 355.2 32.4 356.4 ;
      RECT  36.0 355.2 37.2 356.4 ;
      RECT  40.8 355.2 42.0 356.4 ;
      RECT  45.6 355.2 46.8 356.4 ;
      RECT  50.4 355.2 51.6 356.4 ;
      RECT  55.2 355.2 56.4 356.4 ;
      RECT  60.0 355.2 61.2 356.4 ;
      RECT  64.8 355.2 66.0 356.4 ;
      RECT  69.6 355.2 70.8 356.4 ;
      RECT  74.4 355.2 75.6 356.4 ;
      RECT  79.2 355.2 80.4 356.4 ;
      RECT  84.0 355.2 85.2 356.4 ;
      RECT  88.8 355.2 90.0 356.4 ;
      RECT  93.6 355.2 94.8 356.4 ;
      RECT  98.4 355.2 99.6 356.4 ;
      RECT  103.2 355.2 104.4 356.4 ;
      RECT  108.0 355.2 109.2 356.4 ;
      RECT  112.8 355.2 114.0 356.4 ;
      RECT  117.6 355.2 118.8 356.4 ;
      RECT  122.4 355.2 123.6 356.4 ;
      RECT  127.2 355.2 128.4 356.4 ;
      RECT  132.0 355.2 133.2 356.4 ;
      RECT  136.8 355.2 138.0 356.4 ;
      RECT  141.6 355.2 142.8 356.4 ;
      RECT  146.4 355.2 147.6 356.4 ;
      RECT  151.2 355.2 152.4 356.4 ;
      RECT  156.0 355.2 157.2 356.4 ;
      RECT  160.8 355.2 162.0 356.4 ;
      RECT  165.6 355.2 166.8 356.4 ;
      RECT  170.4 355.2 171.6 356.4 ;
      RECT  175.2 355.2 176.4 356.4 ;
      RECT  180.0 355.2 181.2 356.4 ;
      RECT  184.8 355.2 186.0 356.4 ;
      RECT  189.6 355.2 190.8 356.4 ;
      RECT  194.4 355.2 195.6 356.4 ;
      RECT  199.2 355.2 200.4 356.4 ;
      RECT  204.0 355.2 205.2 356.4 ;
      RECT  208.8 355.2 210.0 356.4 ;
      RECT  213.6 355.2 214.8 356.4 ;
      RECT  218.4 355.2 219.6 356.4 ;
      RECT  223.2 355.2 224.4 356.4 ;
      RECT  2.4 360.0 3.6 361.2 ;
      RECT  7.2 360.0 8.4 361.2 ;
      RECT  12.0 360.0 13.2 361.2 ;
      RECT  16.8 360.0 18.0 361.2 ;
      RECT  21.6 360.0 22.8 361.2 ;
      RECT  26.4 360.0 27.6 361.2 ;
      RECT  31.2 360.0 32.4 361.2 ;
      RECT  36.0 360.0 37.2 361.2 ;
      RECT  40.8 360.0 42.0 361.2 ;
      RECT  45.6 360.0 46.8 361.2 ;
      RECT  50.4 360.0 51.6 361.2 ;
      RECT  55.2 360.0 56.4 361.2 ;
      RECT  60.0 360.0 61.2 361.2 ;
      RECT  64.8 360.0 66.0 361.2 ;
      RECT  69.6 360.0 70.8 361.2 ;
      RECT  74.4 360.0 75.6 361.2 ;
      RECT  79.2 360.0 80.4 361.2 ;
      RECT  84.0 360.0 85.2 361.2 ;
      RECT  88.8 360.0 90.0 361.2 ;
      RECT  93.6 360.0 94.8 361.2 ;
      RECT  98.4 360.0 99.6 361.2 ;
      RECT  103.2 360.0 104.4 361.2 ;
      RECT  108.0 360.0 109.2 361.2 ;
      RECT  112.8 360.0 114.0 361.2 ;
      RECT  117.6 360.0 118.8 361.2 ;
      RECT  122.4 360.0 123.6 361.2 ;
      RECT  127.2 360.0 128.4 361.2 ;
      RECT  132.0 360.0 133.2 361.2 ;
      RECT  136.8 360.0 138.0 361.2 ;
      RECT  141.6 360.0 142.8 361.2 ;
      RECT  146.4 360.0 147.6 361.2 ;
      RECT  151.2 360.0 152.4 361.2 ;
      RECT  156.0 360.0 157.2 361.2 ;
      RECT  160.8 360.0 162.0 361.2 ;
      RECT  165.6 360.0 166.8 361.2 ;
      RECT  170.4 360.0 171.6 361.2 ;
      RECT  175.2 360.0 176.4 361.2 ;
      RECT  180.0 360.0 181.2 361.2 ;
      RECT  184.8 360.0 186.0 361.2 ;
      RECT  189.6 360.0 190.8 361.2 ;
      RECT  194.4 360.0 195.6 361.2 ;
      RECT  199.2 360.0 200.4 361.2 ;
      RECT  204.0 360.0 205.2 361.2 ;
      RECT  208.8 360.0 210.0 361.2 ;
      RECT  213.6 360.0 214.8 361.2 ;
      RECT  218.4 360.0 219.6 361.2 ;
      RECT  223.2 360.0 224.4 361.2 ;
      RECT  2.4 364.8 3.6 366.0 ;
      RECT  7.2 364.8 8.4 366.0 ;
      RECT  12.0 364.8 13.2 366.0 ;
      RECT  16.8 364.8 18.0 366.0 ;
      RECT  21.6 364.8 22.8 366.0 ;
      RECT  26.4 364.8 27.6 366.0 ;
      RECT  31.2 364.8 32.4 366.0 ;
      RECT  36.0 364.8 37.2 366.0 ;
      RECT  40.8 364.8 42.0 366.0 ;
      RECT  45.6 364.8 46.8 366.0 ;
      RECT  50.4 364.8 51.6 366.0 ;
      RECT  55.2 364.8 56.4 366.0 ;
      RECT  60.0 364.8 61.2 366.0 ;
      RECT  64.8 364.8 66.0 366.0 ;
      RECT  69.6 364.8 70.8 366.0 ;
      RECT  74.4 364.8 75.6 366.0 ;
      RECT  79.2 364.8 80.4 366.0 ;
      RECT  84.0 364.8 85.2 366.0 ;
      RECT  88.8 364.8 90.0 366.0 ;
      RECT  93.6 364.8 94.8 366.0 ;
      RECT  98.4 364.8 99.6 366.0 ;
      RECT  103.2 364.8 104.4 366.0 ;
      RECT  108.0 364.8 109.2 366.0 ;
      RECT  112.8 364.8 114.0 366.0 ;
      RECT  117.6 364.8 118.8 366.0 ;
      RECT  122.4 364.8 123.6 366.0 ;
      RECT  127.2 364.8 128.4 366.0 ;
      RECT  132.0 364.8 133.2 366.0 ;
      RECT  136.8 364.8 138.0 366.0 ;
      RECT  141.6 364.8 142.8 366.0 ;
      RECT  146.4 364.8 147.6 366.0 ;
      RECT  151.2 364.8 152.4 366.0 ;
      RECT  156.0 364.8 157.2 366.0 ;
      RECT  160.8 364.8 162.0 366.0 ;
      RECT  165.6 364.8 166.8 366.0 ;
      RECT  170.4 364.8 171.6 366.0 ;
      RECT  175.2 364.8 176.4 366.0 ;
      RECT  180.0 364.8 181.2 366.0 ;
      RECT  184.8 364.8 186.0 366.0 ;
      RECT  189.6 364.8 190.8 366.0 ;
      RECT  194.4 364.8 195.6 366.0 ;
      RECT  199.2 364.8 200.4 366.0 ;
      RECT  204.0 364.8 205.2 366.0 ;
      RECT  208.8 364.8 210.0 366.0 ;
      RECT  213.6 364.8 214.8 366.0 ;
      RECT  218.4 364.8 219.6 366.0 ;
      RECT  223.2 364.8 224.4 366.0 ;
      RECT  2.4 369.6 3.6 370.8 ;
      RECT  7.2 369.6 8.4 370.8 ;
      RECT  12.0 369.6 13.2 370.8 ;
      RECT  16.8 369.6 18.0 370.8 ;
      RECT  21.6 369.6 22.8 370.8 ;
      RECT  26.4 369.6 27.6 370.8 ;
      RECT  31.2 369.6 32.4 370.8 ;
      RECT  36.0 369.6 37.2 370.8 ;
      RECT  40.8 369.6 42.0 370.8 ;
      RECT  45.6 369.6 46.8 370.8 ;
      RECT  50.4 369.6 51.6 370.8 ;
      RECT  55.2 369.6 56.4 370.8 ;
      RECT  60.0 369.6 61.2 370.8 ;
      RECT  64.8 369.6 66.0 370.8 ;
      RECT  69.6 369.6 70.8 370.8 ;
      RECT  74.4 369.6 75.6 370.8 ;
      RECT  79.2 369.6 80.4 370.8 ;
      RECT  84.0 369.6 85.2 370.8 ;
      RECT  88.8 369.6 90.0 370.8 ;
      RECT  93.6 369.6 94.8 370.8 ;
      RECT  98.4 369.6 99.6 370.8 ;
      RECT  103.2 369.6 104.4 370.8 ;
      RECT  108.0 369.6 109.2 370.8 ;
      RECT  112.8 369.6 114.0 370.8 ;
      RECT  117.6 369.6 118.8 370.8 ;
      RECT  122.4 369.6 123.6 370.8 ;
      RECT  127.2 369.6 128.4 370.8 ;
      RECT  132.0 369.6 133.2 370.8 ;
      RECT  136.8 369.6 138.0 370.8 ;
      RECT  141.6 369.6 142.8 370.8 ;
      RECT  146.4 369.6 147.6 370.8 ;
      RECT  151.2 369.6 152.4 370.8 ;
      RECT  156.0 369.6 157.2 370.8 ;
      RECT  160.8 369.6 162.0 370.8 ;
      RECT  165.6 369.6 166.8 370.8 ;
      RECT  170.4 369.6 171.6 370.8 ;
      RECT  175.2 369.6 176.4 370.8 ;
      RECT  180.0 369.6 181.2 370.8 ;
      RECT  4.8 2.4 6.0 3.6 ;
      RECT  9.6 2.4 10.8 3.6 ;
      RECT  14.4 2.4 15.6 3.6 ;
      RECT  19.2 2.4 20.4 3.6 ;
      RECT  24.0 2.4 25.2 3.6 ;
      RECT  28.8 2.4 30.0 3.6 ;
      RECT  33.6 2.4 34.8 3.6 ;
      RECT  38.4 2.4 39.6 3.6 ;
      RECT  43.2 2.4 44.4 3.6 ;
      RECT  48.0 2.4 49.2 3.6 ;
      RECT  52.8 2.4 54.0 3.6 ;
      RECT  57.6 2.4 58.8 3.6 ;
      RECT  62.4 2.4 63.6 3.6 ;
      RECT  67.2 2.4 68.4 3.6 ;
      RECT  72.0 2.4 73.2 3.6 ;
      RECT  76.8 2.4 78.0 3.6 ;
      RECT  91.2 2.4 92.4 3.6 ;
      RECT  96.0 2.4 97.2 3.6 ;
      RECT  100.8 2.4 102.0 3.6 ;
      RECT  105.6 2.4 106.8 3.6 ;
      RECT  110.4 2.4 111.6 3.6 ;
      RECT  115.2 2.4 116.4 3.6 ;
      RECT  120.0 2.4 121.2 3.6 ;
      RECT  124.8 2.4 126.0 3.6 ;
      RECT  129.6 2.4 130.8 3.6 ;
      RECT  134.4 2.4 135.6 3.6 ;
      RECT  139.2 2.4 140.4 3.6 ;
      RECT  144.0 2.4 145.2 3.6 ;
      RECT  148.8 2.4 150.0 3.6 ;
      RECT  153.6 2.4 154.8 3.6 ;
      RECT  158.4 2.4 159.6 3.6 ;
      RECT  163.2 2.4 164.4 3.6 ;
      RECT  168.0 2.4 169.2 3.6 ;
      RECT  172.8 2.4 174.0 3.6 ;
      RECT  177.6 2.4 178.8 3.6 ;
      RECT  182.4 2.4 183.6 3.6 ;
      RECT  187.2 2.4 188.4 3.6 ;
      RECT  192.0 2.4 193.2 3.6 ;
      RECT  196.8 2.4 198.0 3.6 ;
      RECT  201.6 2.4 202.8 3.6 ;
      RECT  206.4 2.4 207.6 3.6 ;
      RECT  211.2 2.4 212.4 3.6 ;
      RECT  216.0 2.4 217.2 3.6 ;
      RECT  220.8 2.4 222.0 3.6 ;
      RECT  225.6 2.4 226.8 3.6 ;
      RECT  4.8 7.2 6.0 8.4 ;
      RECT  9.6 7.2 10.8 8.4 ;
      RECT  14.4 7.2 15.6 8.4 ;
      RECT  19.2 7.2 20.4 8.4 ;
      RECT  24.0 7.2 25.2 8.4 ;
      RECT  28.8 7.2 30.0 8.4 ;
      RECT  33.6 7.2 34.8 8.4 ;
      RECT  38.4 7.2 39.6 8.4 ;
      RECT  43.2 7.2 44.4 8.4 ;
      RECT  48.0 7.2 49.2 8.4 ;
      RECT  52.8 7.2 54.0 8.4 ;
      RECT  57.6 7.2 58.8 8.4 ;
      RECT  62.4 7.2 63.6 8.4 ;
      RECT  67.2 7.2 68.4 8.4 ;
      RECT  72.0 7.2 73.2 8.4 ;
      RECT  76.8 7.2 78.0 8.4 ;
      RECT  81.6 7.2 82.8 8.4 ;
      RECT  86.4 7.2 87.6 8.4 ;
      RECT  91.2 7.2 92.4 8.4 ;
      RECT  96.0 7.2 97.2 8.4 ;
      RECT  100.8 7.2 102.0 8.4 ;
      RECT  105.6 7.2 106.8 8.4 ;
      RECT  110.4 7.2 111.6 8.4 ;
      RECT  115.2 7.2 116.4 8.4 ;
      RECT  120.0 7.2 121.2 8.4 ;
      RECT  124.8 7.2 126.0 8.4 ;
      RECT  129.6 7.2 130.8 8.4 ;
      RECT  134.4 7.2 135.6 8.4 ;
      RECT  139.2 7.2 140.4 8.4 ;
      RECT  144.0 7.2 145.2 8.4 ;
      RECT  148.8 7.2 150.0 8.4 ;
      RECT  153.6 7.2 154.8 8.4 ;
      RECT  158.4 7.2 159.6 8.4 ;
      RECT  163.2 7.2 164.4 8.4 ;
      RECT  168.0 7.2 169.2 8.4 ;
      RECT  172.8 7.2 174.0 8.4 ;
      RECT  177.6 7.2 178.8 8.4 ;
      RECT  182.4 7.2 183.6 8.4 ;
      RECT  187.2 7.2 188.4 8.4 ;
      RECT  192.0 7.2 193.2 8.4 ;
      RECT  196.8 7.2 198.0 8.4 ;
      RECT  201.6 7.2 202.8 8.4 ;
      RECT  206.4 7.2 207.6 8.4 ;
      RECT  211.2 7.2 212.4 8.4 ;
      RECT  216.0 7.2 217.2 8.4 ;
      RECT  220.8 7.2 222.0 8.4 ;
      RECT  225.6 7.2 226.8 8.4 ;
      RECT  52.8 12.0 54.0 13.2 ;
      RECT  57.6 12.0 58.8 13.2 ;
      RECT  62.4 12.0 63.6 13.2 ;
      RECT  67.2 12.0 68.4 13.2 ;
      RECT  72.0 12.0 73.2 13.2 ;
      RECT  76.8 12.0 78.0 13.2 ;
      RECT  81.6 12.0 82.8 13.2 ;
      RECT  86.4 12.0 87.6 13.2 ;
      RECT  91.2 12.0 92.4 13.2 ;
      RECT  96.0 12.0 97.2 13.2 ;
      RECT  100.8 12.0 102.0 13.2 ;
      RECT  105.6 12.0 106.8 13.2 ;
      RECT  110.4 12.0 111.6 13.2 ;
      RECT  115.2 12.0 116.4 13.2 ;
      RECT  120.0 12.0 121.2 13.2 ;
      RECT  124.8 12.0 126.0 13.2 ;
      RECT  129.6 12.0 130.8 13.2 ;
      RECT  134.4 12.0 135.6 13.2 ;
      RECT  139.2 12.0 140.4 13.2 ;
      RECT  144.0 12.0 145.2 13.2 ;
      RECT  148.8 12.0 150.0 13.2 ;
      RECT  153.6 12.0 154.8 13.2 ;
      RECT  158.4 12.0 159.6 13.2 ;
      RECT  163.2 12.0 164.4 13.2 ;
      RECT  168.0 12.0 169.2 13.2 ;
      RECT  172.8 12.0 174.0 13.2 ;
      RECT  177.6 12.0 178.8 13.2 ;
      RECT  182.4 12.0 183.6 13.2 ;
      RECT  187.2 12.0 188.4 13.2 ;
      RECT  192.0 12.0 193.2 13.2 ;
      RECT  196.8 12.0 198.0 13.2 ;
      RECT  201.6 12.0 202.8 13.2 ;
      RECT  206.4 12.0 207.6 13.2 ;
      RECT  211.2 12.0 212.4 13.2 ;
      RECT  216.0 12.0 217.2 13.2 ;
      RECT  220.8 12.0 222.0 13.2 ;
      RECT  225.6 12.0 226.8 13.2 ;
      RECT  4.8 16.8 6.0 18.0 ;
      RECT  9.6 16.8 10.8 18.0 ;
      RECT  14.4 16.8 15.6 18.0 ;
      RECT  19.2 16.8 20.4 18.0 ;
      RECT  24.0 16.8 25.2 18.0 ;
      RECT  28.8 16.8 30.0 18.0 ;
      RECT  33.6 16.8 34.8 18.0 ;
      RECT  38.4 16.8 39.6 18.0 ;
      RECT  43.2 16.8 44.4 18.0 ;
      RECT  48.0 16.8 49.2 18.0 ;
      RECT  52.8 16.8 54.0 18.0 ;
      RECT  57.6 16.8 58.8 18.0 ;
      RECT  62.4 16.8 63.6 18.0 ;
      RECT  67.2 16.8 68.4 18.0 ;
      RECT  72.0 16.8 73.2 18.0 ;
      RECT  76.8 16.8 78.0 18.0 ;
      RECT  81.6 16.8 82.8 18.0 ;
      RECT  86.4 16.8 87.6 18.0 ;
      RECT  91.2 16.8 92.4 18.0 ;
      RECT  96.0 16.8 97.2 18.0 ;
      RECT  100.8 16.8 102.0 18.0 ;
      RECT  105.6 16.8 106.8 18.0 ;
      RECT  110.4 16.8 111.6 18.0 ;
      RECT  115.2 16.8 116.4 18.0 ;
      RECT  120.0 16.8 121.2 18.0 ;
      RECT  124.8 16.8 126.0 18.0 ;
      RECT  129.6 16.8 130.8 18.0 ;
      RECT  134.4 16.8 135.6 18.0 ;
      RECT  139.2 16.8 140.4 18.0 ;
      RECT  144.0 16.8 145.2 18.0 ;
      RECT  148.8 16.8 150.0 18.0 ;
      RECT  153.6 16.8 154.8 18.0 ;
      RECT  158.4 16.8 159.6 18.0 ;
      RECT  163.2 16.8 164.4 18.0 ;
      RECT  168.0 16.8 169.2 18.0 ;
      RECT  172.8 16.8 174.0 18.0 ;
      RECT  177.6 16.8 178.8 18.0 ;
      RECT  182.4 16.8 183.6 18.0 ;
      RECT  187.2 16.8 188.4 18.0 ;
      RECT  192.0 16.8 193.2 18.0 ;
      RECT  196.8 16.8 198.0 18.0 ;
      RECT  201.6 16.8 202.8 18.0 ;
      RECT  206.4 16.8 207.6 18.0 ;
      RECT  211.2 16.8 212.4 18.0 ;
      RECT  216.0 16.8 217.2 18.0 ;
      RECT  220.8 16.8 222.0 18.0 ;
      RECT  225.6 16.8 226.8 18.0 ;
      RECT  4.8 21.6 6.0 22.8 ;
      RECT  9.6 21.6 10.8 22.8 ;
      RECT  14.4 21.6 15.6 22.8 ;
      RECT  19.2 21.6 20.4 22.8 ;
      RECT  24.0 21.6 25.2 22.8 ;
      RECT  28.8 21.6 30.0 22.8 ;
      RECT  33.6 21.6 34.8 22.8 ;
      RECT  38.4 21.6 39.6 22.8 ;
      RECT  43.2 21.6 44.4 22.8 ;
      RECT  48.0 21.6 49.2 22.8 ;
      RECT  52.8 21.6 54.0 22.8 ;
      RECT  57.6 21.6 58.8 22.8 ;
      RECT  62.4 21.6 63.6 22.8 ;
      RECT  67.2 21.6 68.4 22.8 ;
      RECT  72.0 21.6 73.2 22.8 ;
      RECT  76.8 21.6 78.0 22.8 ;
      RECT  81.6 21.6 82.8 22.8 ;
      RECT  86.4 21.6 87.6 22.8 ;
      RECT  91.2 21.6 92.4 22.8 ;
      RECT  96.0 21.6 97.2 22.8 ;
      RECT  100.8 21.6 102.0 22.8 ;
      RECT  105.6 21.6 106.8 22.8 ;
      RECT  110.4 21.6 111.6 22.8 ;
      RECT  115.2 21.6 116.4 22.8 ;
      RECT  120.0 21.6 121.2 22.8 ;
      RECT  124.8 21.6 126.0 22.8 ;
      RECT  129.6 21.6 130.8 22.8 ;
      RECT  134.4 21.6 135.6 22.8 ;
      RECT  139.2 21.6 140.4 22.8 ;
      RECT  144.0 21.6 145.2 22.8 ;
      RECT  148.8 21.6 150.0 22.8 ;
      RECT  153.6 21.6 154.8 22.8 ;
      RECT  158.4 21.6 159.6 22.8 ;
      RECT  163.2 21.6 164.4 22.8 ;
      RECT  168.0 21.6 169.2 22.8 ;
      RECT  172.8 21.6 174.0 22.8 ;
      RECT  177.6 21.6 178.8 22.8 ;
      RECT  182.4 21.6 183.6 22.8 ;
      RECT  187.2 21.6 188.4 22.8 ;
      RECT  192.0 21.6 193.2 22.8 ;
      RECT  196.8 21.6 198.0 22.8 ;
      RECT  201.6 21.6 202.8 22.8 ;
      RECT  206.4 21.6 207.6 22.8 ;
      RECT  211.2 21.6 212.4 22.8 ;
      RECT  216.0 21.6 217.2 22.8 ;
      RECT  220.8 21.6 222.0 22.8 ;
      RECT  225.6 21.6 226.8 22.8 ;
      RECT  4.8 26.4 6.0 27.6 ;
      RECT  9.6 26.4 10.8 27.6 ;
      RECT  14.4 26.4 15.6 27.6 ;
      RECT  19.2 26.4 20.4 27.6 ;
      RECT  24.0 26.4 25.2 27.6 ;
      RECT  28.8 26.4 30.0 27.6 ;
      RECT  33.6 26.4 34.8 27.6 ;
      RECT  38.4 26.4 39.6 27.6 ;
      RECT  43.2 26.4 44.4 27.6 ;
      RECT  48.0 26.4 49.2 27.6 ;
      RECT  52.8 26.4 54.0 27.6 ;
      RECT  57.6 26.4 58.8 27.6 ;
      RECT  62.4 26.4 63.6 27.6 ;
      RECT  67.2 26.4 68.4 27.6 ;
      RECT  72.0 26.4 73.2 27.6 ;
      RECT  76.8 26.4 78.0 27.6 ;
      RECT  81.6 26.4 82.8 27.6 ;
      RECT  86.4 26.4 87.6 27.6 ;
      RECT  91.2 26.4 92.4 27.6 ;
      RECT  96.0 26.4 97.2 27.6 ;
      RECT  100.8 26.4 102.0 27.6 ;
      RECT  105.6 26.4 106.8 27.6 ;
      RECT  110.4 26.4 111.6 27.6 ;
      RECT  115.2 26.4 116.4 27.6 ;
      RECT  120.0 26.4 121.2 27.6 ;
      RECT  124.8 26.4 126.0 27.6 ;
      RECT  129.6 26.4 130.8 27.6 ;
      RECT  134.4 26.4 135.6 27.6 ;
      RECT  139.2 26.4 140.4 27.6 ;
      RECT  144.0 26.4 145.2 27.6 ;
      RECT  148.8 26.4 150.0 27.6 ;
      RECT  153.6 26.4 154.8 27.6 ;
      RECT  158.4 26.4 159.6 27.6 ;
      RECT  163.2 26.4 164.4 27.6 ;
      RECT  168.0 26.4 169.2 27.6 ;
      RECT  172.8 26.4 174.0 27.6 ;
      RECT  177.6 26.4 178.8 27.6 ;
      RECT  182.4 26.4 183.6 27.6 ;
      RECT  187.2 26.4 188.4 27.6 ;
      RECT  192.0 26.4 193.2 27.6 ;
      RECT  196.8 26.4 198.0 27.6 ;
      RECT  201.6 26.4 202.8 27.6 ;
      RECT  206.4 26.4 207.6 27.6 ;
      RECT  211.2 26.4 212.4 27.6 ;
      RECT  216.0 26.4 217.2 27.6 ;
      RECT  220.8 26.4 222.0 27.6 ;
      RECT  225.6 26.4 226.8 27.6 ;
      RECT  86.4 31.2 87.6 32.4 ;
      RECT  91.2 31.2 92.4 32.4 ;
      RECT  96.0 31.2 97.2 32.4 ;
      RECT  100.8 31.2 102.0 32.4 ;
      RECT  105.6 31.2 106.8 32.4 ;
      RECT  110.4 31.2 111.6 32.4 ;
      RECT  115.2 31.2 116.4 32.4 ;
      RECT  120.0 31.2 121.2 32.4 ;
      RECT  124.8 31.2 126.0 32.4 ;
      RECT  129.6 31.2 130.8 32.4 ;
      RECT  134.4 31.2 135.6 32.4 ;
      RECT  139.2 31.2 140.4 32.4 ;
      RECT  144.0 31.2 145.2 32.4 ;
      RECT  148.8 31.2 150.0 32.4 ;
      RECT  153.6 31.2 154.8 32.4 ;
      RECT  158.4 31.2 159.6 32.4 ;
      RECT  163.2 31.2 164.4 32.4 ;
      RECT  168.0 31.2 169.2 32.4 ;
      RECT  172.8 31.2 174.0 32.4 ;
      RECT  177.6 31.2 178.8 32.4 ;
      RECT  182.4 31.2 183.6 32.4 ;
      RECT  187.2 31.2 188.4 32.4 ;
      RECT  192.0 31.2 193.2 32.4 ;
      RECT  196.8 31.2 198.0 32.4 ;
      RECT  201.6 31.2 202.8 32.4 ;
      RECT  206.4 31.2 207.6 32.4 ;
      RECT  211.2 31.2 212.4 32.4 ;
      RECT  216.0 31.2 217.2 32.4 ;
      RECT  220.8 31.2 222.0 32.4 ;
      RECT  225.6 31.2 226.8 32.4 ;
      RECT  4.8 36.0 6.0 37.2 ;
      RECT  9.6 36.0 10.8 37.2 ;
      RECT  14.4 36.0 15.6 37.2 ;
      RECT  19.2 36.0 20.4 37.2 ;
      RECT  24.0 36.0 25.2 37.2 ;
      RECT  28.8 36.0 30.0 37.2 ;
      RECT  33.6 36.0 34.8 37.2 ;
      RECT  38.4 36.0 39.6 37.2 ;
      RECT  62.4 36.0 63.6 37.2 ;
      RECT  67.2 36.0 68.4 37.2 ;
      RECT  72.0 36.0 73.2 37.2 ;
      RECT  76.8 36.0 78.0 37.2 ;
      RECT  81.6 36.0 82.8 37.2 ;
      RECT  86.4 36.0 87.6 37.2 ;
      RECT  91.2 36.0 92.4 37.2 ;
      RECT  96.0 36.0 97.2 37.2 ;
      RECT  100.8 36.0 102.0 37.2 ;
      RECT  105.6 36.0 106.8 37.2 ;
      RECT  110.4 36.0 111.6 37.2 ;
      RECT  115.2 36.0 116.4 37.2 ;
      RECT  120.0 36.0 121.2 37.2 ;
      RECT  124.8 36.0 126.0 37.2 ;
      RECT  129.6 36.0 130.8 37.2 ;
      RECT  134.4 36.0 135.6 37.2 ;
      RECT  139.2 36.0 140.4 37.2 ;
      RECT  144.0 36.0 145.2 37.2 ;
      RECT  148.8 36.0 150.0 37.2 ;
      RECT  153.6 36.0 154.8 37.2 ;
      RECT  158.4 36.0 159.6 37.2 ;
      RECT  163.2 36.0 164.4 37.2 ;
      RECT  168.0 36.0 169.2 37.2 ;
      RECT  172.8 36.0 174.0 37.2 ;
      RECT  177.6 36.0 178.8 37.2 ;
      RECT  182.4 36.0 183.6 37.2 ;
      RECT  187.2 36.0 188.4 37.2 ;
      RECT  192.0 36.0 193.2 37.2 ;
      RECT  196.8 36.0 198.0 37.2 ;
      RECT  201.6 36.0 202.8 37.2 ;
      RECT  206.4 36.0 207.6 37.2 ;
      RECT  211.2 36.0 212.4 37.2 ;
      RECT  216.0 36.0 217.2 37.2 ;
      RECT  220.8 36.0 222.0 37.2 ;
      RECT  225.6 36.0 226.8 37.2 ;
      RECT  4.8 40.8 6.0 42.0 ;
      RECT  9.6 40.8 10.8 42.0 ;
      RECT  14.4 40.8 15.6 42.0 ;
      RECT  19.2 40.8 20.4 42.0 ;
      RECT  24.0 40.8 25.2 42.0 ;
      RECT  28.8 40.8 30.0 42.0 ;
      RECT  33.6 40.8 34.8 42.0 ;
      RECT  38.4 40.8 39.6 42.0 ;
      RECT  43.2 40.8 44.4 42.0 ;
      RECT  48.0 40.8 49.2 42.0 ;
      RECT  52.8 40.8 54.0 42.0 ;
      RECT  57.6 40.8 58.8 42.0 ;
      RECT  62.4 40.8 63.6 42.0 ;
      RECT  67.2 40.8 68.4 42.0 ;
      RECT  72.0 40.8 73.2 42.0 ;
      RECT  76.8 40.8 78.0 42.0 ;
      RECT  91.2 40.8 92.4 42.0 ;
      RECT  96.0 40.8 97.2 42.0 ;
      RECT  100.8 40.8 102.0 42.0 ;
      RECT  105.6 40.8 106.8 42.0 ;
      RECT  110.4 40.8 111.6 42.0 ;
      RECT  115.2 40.8 116.4 42.0 ;
      RECT  120.0 40.8 121.2 42.0 ;
      RECT  124.8 40.8 126.0 42.0 ;
      RECT  129.6 40.8 130.8 42.0 ;
      RECT  134.4 40.8 135.6 42.0 ;
      RECT  139.2 40.8 140.4 42.0 ;
      RECT  144.0 40.8 145.2 42.0 ;
      RECT  148.8 40.8 150.0 42.0 ;
      RECT  153.6 40.8 154.8 42.0 ;
      RECT  158.4 40.8 159.6 42.0 ;
      RECT  163.2 40.8 164.4 42.0 ;
      RECT  168.0 40.8 169.2 42.0 ;
      RECT  172.8 40.8 174.0 42.0 ;
      RECT  177.6 40.8 178.8 42.0 ;
      RECT  182.4 40.8 183.6 42.0 ;
      RECT  187.2 40.8 188.4 42.0 ;
      RECT  192.0 40.8 193.2 42.0 ;
      RECT  196.8 40.8 198.0 42.0 ;
      RECT  201.6 40.8 202.8 42.0 ;
      RECT  206.4 40.8 207.6 42.0 ;
      RECT  211.2 40.8 212.4 42.0 ;
      RECT  216.0 40.8 217.2 42.0 ;
      RECT  220.8 40.8 222.0 42.0 ;
      RECT  225.6 40.8 226.8 42.0 ;
      RECT  4.8 45.6 6.0 46.8 ;
      RECT  9.6 45.6 10.8 46.8 ;
      RECT  14.4 45.6 15.6 46.8 ;
      RECT  19.2 45.6 20.4 46.8 ;
      RECT  24.0 45.6 25.2 46.8 ;
      RECT  28.8 45.6 30.0 46.8 ;
      RECT  33.6 45.6 34.8 46.8 ;
      RECT  38.4 45.6 39.6 46.8 ;
      RECT  43.2 45.6 44.4 46.8 ;
      RECT  48.0 45.6 49.2 46.8 ;
      RECT  52.8 45.6 54.0 46.8 ;
      RECT  57.6 45.6 58.8 46.8 ;
      RECT  62.4 45.6 63.6 46.8 ;
      RECT  67.2 45.6 68.4 46.8 ;
      RECT  72.0 45.6 73.2 46.8 ;
      RECT  76.8 45.6 78.0 46.8 ;
      RECT  81.6 45.6 82.8 46.8 ;
      RECT  86.4 45.6 87.6 46.8 ;
      RECT  91.2 45.6 92.4 46.8 ;
      RECT  96.0 45.6 97.2 46.8 ;
      RECT  100.8 45.6 102.0 46.8 ;
      RECT  105.6 45.6 106.8 46.8 ;
      RECT  110.4 45.6 111.6 46.8 ;
      RECT  115.2 45.6 116.4 46.8 ;
      RECT  120.0 45.6 121.2 46.8 ;
      RECT  124.8 45.6 126.0 46.8 ;
      RECT  129.6 45.6 130.8 46.8 ;
      RECT  134.4 45.6 135.6 46.8 ;
      RECT  139.2 45.6 140.4 46.8 ;
      RECT  144.0 45.6 145.2 46.8 ;
      RECT  148.8 45.6 150.0 46.8 ;
      RECT  153.6 45.6 154.8 46.8 ;
      RECT  158.4 45.6 159.6 46.8 ;
      RECT  163.2 45.6 164.4 46.8 ;
      RECT  168.0 45.6 169.2 46.8 ;
      RECT  172.8 45.6 174.0 46.8 ;
      RECT  177.6 45.6 178.8 46.8 ;
      RECT  182.4 45.6 183.6 46.8 ;
      RECT  187.2 45.6 188.4 46.8 ;
      RECT  4.8 50.4 6.0 51.6 ;
      RECT  9.6 50.4 10.8 51.6 ;
      RECT  14.4 50.4 15.6 51.6 ;
      RECT  19.2 50.4 20.4 51.6 ;
      RECT  24.0 50.4 25.2 51.6 ;
      RECT  28.8 50.4 30.0 51.6 ;
      RECT  33.6 50.4 34.8 51.6 ;
      RECT  81.6 50.4 82.8 51.6 ;
      RECT  86.4 50.4 87.6 51.6 ;
      RECT  91.2 50.4 92.4 51.6 ;
      RECT  96.0 50.4 97.2 51.6 ;
      RECT  100.8 50.4 102.0 51.6 ;
      RECT  105.6 50.4 106.8 51.6 ;
      RECT  110.4 50.4 111.6 51.6 ;
      RECT  115.2 50.4 116.4 51.6 ;
      RECT  120.0 50.4 121.2 51.6 ;
      RECT  124.8 50.4 126.0 51.6 ;
      RECT  129.6 50.4 130.8 51.6 ;
      RECT  134.4 50.4 135.6 51.6 ;
      RECT  139.2 50.4 140.4 51.6 ;
      RECT  144.0 50.4 145.2 51.6 ;
      RECT  148.8 50.4 150.0 51.6 ;
      RECT  153.6 50.4 154.8 51.6 ;
      RECT  158.4 50.4 159.6 51.6 ;
      RECT  163.2 50.4 164.4 51.6 ;
      RECT  168.0 50.4 169.2 51.6 ;
      RECT  172.8 50.4 174.0 51.6 ;
      RECT  177.6 50.4 178.8 51.6 ;
      RECT  182.4 50.4 183.6 51.6 ;
      RECT  187.2 50.4 188.4 51.6 ;
      RECT  192.0 50.4 193.2 51.6 ;
      RECT  196.8 50.4 198.0 51.6 ;
      RECT  201.6 50.4 202.8 51.6 ;
      RECT  206.4 50.4 207.6 51.6 ;
      RECT  211.2 50.4 212.4 51.6 ;
      RECT  216.0 50.4 217.2 51.6 ;
      RECT  220.8 50.4 222.0 51.6 ;
      RECT  225.6 50.4 226.8 51.6 ;
      RECT  4.8 55.2 6.0 56.4 ;
      RECT  9.6 55.2 10.8 56.4 ;
      RECT  14.4 55.2 15.6 56.4 ;
      RECT  19.2 55.2 20.4 56.4 ;
      RECT  24.0 55.2 25.2 56.4 ;
      RECT  28.8 55.2 30.0 56.4 ;
      RECT  33.6 55.2 34.8 56.4 ;
      RECT  38.4 55.2 39.6 56.4 ;
      RECT  43.2 55.2 44.4 56.4 ;
      RECT  48.0 55.2 49.2 56.4 ;
      RECT  52.8 55.2 54.0 56.4 ;
      RECT  57.6 55.2 58.8 56.4 ;
      RECT  62.4 55.2 63.6 56.4 ;
      RECT  67.2 55.2 68.4 56.4 ;
      RECT  72.0 55.2 73.2 56.4 ;
      RECT  76.8 55.2 78.0 56.4 ;
      RECT  81.6 55.2 82.8 56.4 ;
      RECT  86.4 55.2 87.6 56.4 ;
      RECT  91.2 55.2 92.4 56.4 ;
      RECT  96.0 55.2 97.2 56.4 ;
      RECT  100.8 55.2 102.0 56.4 ;
      RECT  105.6 55.2 106.8 56.4 ;
      RECT  110.4 55.2 111.6 56.4 ;
      RECT  115.2 55.2 116.4 56.4 ;
      RECT  120.0 55.2 121.2 56.4 ;
      RECT  124.8 55.2 126.0 56.4 ;
      RECT  129.6 55.2 130.8 56.4 ;
      RECT  134.4 55.2 135.6 56.4 ;
      RECT  139.2 55.2 140.4 56.4 ;
      RECT  144.0 55.2 145.2 56.4 ;
      RECT  148.8 55.2 150.0 56.4 ;
      RECT  153.6 55.2 154.8 56.4 ;
      RECT  158.4 55.2 159.6 56.4 ;
      RECT  163.2 55.2 164.4 56.4 ;
      RECT  168.0 55.2 169.2 56.4 ;
      RECT  172.8 55.2 174.0 56.4 ;
      RECT  177.6 55.2 178.8 56.4 ;
      RECT  182.4 55.2 183.6 56.4 ;
      RECT  187.2 55.2 188.4 56.4 ;
      RECT  192.0 55.2 193.2 56.4 ;
      RECT  196.8 55.2 198.0 56.4 ;
      RECT  201.6 55.2 202.8 56.4 ;
      RECT  206.4 55.2 207.6 56.4 ;
      RECT  211.2 55.2 212.4 56.4 ;
      RECT  216.0 55.2 217.2 56.4 ;
      RECT  220.8 55.2 222.0 56.4 ;
      RECT  225.6 55.2 226.8 56.4 ;
      RECT  4.8 60.0 6.0 61.2 ;
      RECT  9.6 60.0 10.8 61.2 ;
      RECT  14.4 60.0 15.6 61.2 ;
      RECT  19.2 60.0 20.4 61.2 ;
      RECT  24.0 60.0 25.2 61.2 ;
      RECT  28.8 60.0 30.0 61.2 ;
      RECT  33.6 60.0 34.8 61.2 ;
      RECT  38.4 60.0 39.6 61.2 ;
      RECT  43.2 60.0 44.4 61.2 ;
      RECT  48.0 60.0 49.2 61.2 ;
      RECT  52.8 60.0 54.0 61.2 ;
      RECT  57.6 60.0 58.8 61.2 ;
      RECT  62.4 60.0 63.6 61.2 ;
      RECT  67.2 60.0 68.4 61.2 ;
      RECT  72.0 60.0 73.2 61.2 ;
      RECT  76.8 60.0 78.0 61.2 ;
      RECT  81.6 60.0 82.8 61.2 ;
      RECT  86.4 60.0 87.6 61.2 ;
      RECT  91.2 60.0 92.4 61.2 ;
      RECT  96.0 60.0 97.2 61.2 ;
      RECT  100.8 60.0 102.0 61.2 ;
      RECT  105.6 60.0 106.8 61.2 ;
      RECT  110.4 60.0 111.6 61.2 ;
      RECT  115.2 60.0 116.4 61.2 ;
      RECT  120.0 60.0 121.2 61.2 ;
      RECT  124.8 60.0 126.0 61.2 ;
      RECT  129.6 60.0 130.8 61.2 ;
      RECT  134.4 60.0 135.6 61.2 ;
      RECT  139.2 60.0 140.4 61.2 ;
      RECT  144.0 60.0 145.2 61.2 ;
      RECT  148.8 60.0 150.0 61.2 ;
      RECT  153.6 60.0 154.8 61.2 ;
      RECT  158.4 60.0 159.6 61.2 ;
      RECT  163.2 60.0 164.4 61.2 ;
      RECT  168.0 60.0 169.2 61.2 ;
      RECT  172.8 60.0 174.0 61.2 ;
      RECT  177.6 60.0 178.8 61.2 ;
      RECT  182.4 60.0 183.6 61.2 ;
      RECT  187.2 60.0 188.4 61.2 ;
      RECT  192.0 60.0 193.2 61.2 ;
      RECT  196.8 60.0 198.0 61.2 ;
      RECT  201.6 60.0 202.8 61.2 ;
      RECT  206.4 60.0 207.6 61.2 ;
      RECT  211.2 60.0 212.4 61.2 ;
      RECT  216.0 60.0 217.2 61.2 ;
      RECT  220.8 60.0 222.0 61.2 ;
      RECT  225.6 60.0 226.8 61.2 ;
      RECT  4.8 64.8 6.0 66.0 ;
      RECT  9.6 64.8 10.8 66.0 ;
      RECT  14.4 64.8 15.6 66.0 ;
      RECT  19.2 64.8 20.4 66.0 ;
      RECT  24.0 64.8 25.2 66.0 ;
      RECT  28.8 64.8 30.0 66.0 ;
      RECT  33.6 64.8 34.8 66.0 ;
      RECT  38.4 64.8 39.6 66.0 ;
      RECT  43.2 64.8 44.4 66.0 ;
      RECT  48.0 64.8 49.2 66.0 ;
      RECT  52.8 64.8 54.0 66.0 ;
      RECT  57.6 64.8 58.8 66.0 ;
      RECT  62.4 64.8 63.6 66.0 ;
      RECT  67.2 64.8 68.4 66.0 ;
      RECT  72.0 64.8 73.2 66.0 ;
      RECT  76.8 64.8 78.0 66.0 ;
      RECT  81.6 64.8 82.8 66.0 ;
      RECT  86.4 64.8 87.6 66.0 ;
      RECT  91.2 64.8 92.4 66.0 ;
      RECT  96.0 64.8 97.2 66.0 ;
      RECT  100.8 64.8 102.0 66.0 ;
      RECT  105.6 64.8 106.8 66.0 ;
      RECT  110.4 64.8 111.6 66.0 ;
      RECT  115.2 64.8 116.4 66.0 ;
      RECT  120.0 64.8 121.2 66.0 ;
      RECT  124.8 64.8 126.0 66.0 ;
      RECT  129.6 64.8 130.8 66.0 ;
      RECT  134.4 64.8 135.6 66.0 ;
      RECT  139.2 64.8 140.4 66.0 ;
      RECT  144.0 64.8 145.2 66.0 ;
      RECT  148.8 64.8 150.0 66.0 ;
      RECT  153.6 64.8 154.8 66.0 ;
      RECT  158.4 64.8 159.6 66.0 ;
      RECT  163.2 64.8 164.4 66.0 ;
      RECT  168.0 64.8 169.2 66.0 ;
      RECT  172.8 64.8 174.0 66.0 ;
      RECT  177.6 64.8 178.8 66.0 ;
      RECT  182.4 64.8 183.6 66.0 ;
      RECT  187.2 64.8 188.4 66.0 ;
      RECT  192.0 64.8 193.2 66.0 ;
      RECT  196.8 64.8 198.0 66.0 ;
      RECT  201.6 64.8 202.8 66.0 ;
      RECT  206.4 64.8 207.6 66.0 ;
      RECT  211.2 64.8 212.4 66.0 ;
      RECT  216.0 64.8 217.2 66.0 ;
      RECT  220.8 64.8 222.0 66.0 ;
      RECT  225.6 64.8 226.8 66.0 ;
      RECT  4.8 69.6 6.0 70.8 ;
      RECT  9.6 69.6 10.8 70.8 ;
      RECT  14.4 69.6 15.6 70.8 ;
      RECT  19.2 69.6 20.4 70.8 ;
      RECT  24.0 69.6 25.2 70.8 ;
      RECT  28.8 69.6 30.0 70.8 ;
      RECT  33.6 69.6 34.8 70.8 ;
      RECT  38.4 69.6 39.6 70.8 ;
      RECT  43.2 69.6 44.4 70.8 ;
      RECT  48.0 69.6 49.2 70.8 ;
      RECT  52.8 69.6 54.0 70.8 ;
      RECT  57.6 69.6 58.8 70.8 ;
      RECT  62.4 69.6 63.6 70.8 ;
      RECT  67.2 69.6 68.4 70.8 ;
      RECT  72.0 69.6 73.2 70.8 ;
      RECT  76.8 69.6 78.0 70.8 ;
      RECT  81.6 69.6 82.8 70.8 ;
      RECT  86.4 69.6 87.6 70.8 ;
      RECT  91.2 69.6 92.4 70.8 ;
      RECT  96.0 69.6 97.2 70.8 ;
      RECT  100.8 69.6 102.0 70.8 ;
      RECT  105.6 69.6 106.8 70.8 ;
      RECT  110.4 69.6 111.6 70.8 ;
      RECT  115.2 69.6 116.4 70.8 ;
      RECT  120.0 69.6 121.2 70.8 ;
      RECT  124.8 69.6 126.0 70.8 ;
      RECT  129.6 69.6 130.8 70.8 ;
      RECT  134.4 69.6 135.6 70.8 ;
      RECT  139.2 69.6 140.4 70.8 ;
      RECT  144.0 69.6 145.2 70.8 ;
      RECT  148.8 69.6 150.0 70.8 ;
      RECT  153.6 69.6 154.8 70.8 ;
      RECT  158.4 69.6 159.6 70.8 ;
      RECT  163.2 69.6 164.4 70.8 ;
      RECT  168.0 69.6 169.2 70.8 ;
      RECT  172.8 69.6 174.0 70.8 ;
      RECT  177.6 69.6 178.8 70.8 ;
      RECT  182.4 69.6 183.6 70.8 ;
      RECT  187.2 69.6 188.4 70.8 ;
      RECT  192.0 69.6 193.2 70.8 ;
      RECT  196.8 69.6 198.0 70.8 ;
      RECT  201.6 69.6 202.8 70.8 ;
      RECT  206.4 69.6 207.6 70.8 ;
      RECT  211.2 69.6 212.4 70.8 ;
      RECT  216.0 69.6 217.2 70.8 ;
      RECT  220.8 69.6 222.0 70.8 ;
      RECT  225.6 69.6 226.8 70.8 ;
      RECT  4.8 74.4 6.0 75.6 ;
      RECT  9.6 74.4 10.8 75.6 ;
      RECT  14.4 74.4 15.6 75.6 ;
      RECT  19.2 74.4 20.4 75.6 ;
      RECT  24.0 74.4 25.2 75.6 ;
      RECT  28.8 74.4 30.0 75.6 ;
      RECT  33.6 74.4 34.8 75.6 ;
      RECT  38.4 74.4 39.6 75.6 ;
      RECT  43.2 74.4 44.4 75.6 ;
      RECT  48.0 74.4 49.2 75.6 ;
      RECT  52.8 74.4 54.0 75.6 ;
      RECT  57.6 74.4 58.8 75.6 ;
      RECT  62.4 74.4 63.6 75.6 ;
      RECT  67.2 74.4 68.4 75.6 ;
      RECT  72.0 74.4 73.2 75.6 ;
      RECT  76.8 74.4 78.0 75.6 ;
      RECT  81.6 74.4 82.8 75.6 ;
      RECT  187.2 74.4 188.4 75.6 ;
      RECT  192.0 74.4 193.2 75.6 ;
      RECT  196.8 74.4 198.0 75.6 ;
      RECT  201.6 74.4 202.8 75.6 ;
      RECT  206.4 74.4 207.6 75.6 ;
      RECT  211.2 74.4 212.4 75.6 ;
      RECT  216.0 74.4 217.2 75.6 ;
      RECT  220.8 74.4 222.0 75.6 ;
      RECT  225.6 74.4 226.8 75.6 ;
      RECT  4.8 79.2 6.0 80.4 ;
      RECT  9.6 79.2 10.8 80.4 ;
      RECT  14.4 79.2 15.6 80.4 ;
      RECT  19.2 79.2 20.4 80.4 ;
      RECT  24.0 79.2 25.2 80.4 ;
      RECT  28.8 79.2 30.0 80.4 ;
      RECT  33.6 79.2 34.8 80.4 ;
      RECT  38.4 79.2 39.6 80.4 ;
      RECT  43.2 79.2 44.4 80.4 ;
      RECT  48.0 79.2 49.2 80.4 ;
      RECT  52.8 79.2 54.0 80.4 ;
      RECT  57.6 79.2 58.8 80.4 ;
      RECT  62.4 79.2 63.6 80.4 ;
      RECT  67.2 79.2 68.4 80.4 ;
      RECT  72.0 79.2 73.2 80.4 ;
      RECT  76.8 79.2 78.0 80.4 ;
      RECT  81.6 79.2 82.8 80.4 ;
      RECT  86.4 79.2 87.6 80.4 ;
      RECT  91.2 79.2 92.4 80.4 ;
      RECT  96.0 79.2 97.2 80.4 ;
      RECT  100.8 79.2 102.0 80.4 ;
      RECT  105.6 79.2 106.8 80.4 ;
      RECT  110.4 79.2 111.6 80.4 ;
      RECT  115.2 79.2 116.4 80.4 ;
      RECT  120.0 79.2 121.2 80.4 ;
      RECT  124.8 79.2 126.0 80.4 ;
      RECT  129.6 79.2 130.8 80.4 ;
      RECT  134.4 79.2 135.6 80.4 ;
      RECT  139.2 79.2 140.4 80.4 ;
      RECT  144.0 79.2 145.2 80.4 ;
      RECT  148.8 79.2 150.0 80.4 ;
      RECT  153.6 79.2 154.8 80.4 ;
      RECT  158.4 79.2 159.6 80.4 ;
      RECT  163.2 79.2 164.4 80.4 ;
      RECT  168.0 79.2 169.2 80.4 ;
      RECT  172.8 79.2 174.0 80.4 ;
      RECT  177.6 79.2 178.8 80.4 ;
      RECT  182.4 79.2 183.6 80.4 ;
      RECT  187.2 79.2 188.4 80.4 ;
      RECT  192.0 79.2 193.2 80.4 ;
      RECT  196.8 79.2 198.0 80.4 ;
      RECT  201.6 79.2 202.8 80.4 ;
      RECT  206.4 79.2 207.6 80.4 ;
      RECT  211.2 79.2 212.4 80.4 ;
      RECT  216.0 79.2 217.2 80.4 ;
      RECT  220.8 79.2 222.0 80.4 ;
      RECT  225.6 79.2 226.8 80.4 ;
      RECT  4.8 84.0 6.0 85.2 ;
      RECT  9.6 84.0 10.8 85.2 ;
      RECT  14.4 84.0 15.6 85.2 ;
      RECT  19.2 84.0 20.4 85.2 ;
      RECT  24.0 84.0 25.2 85.2 ;
      RECT  28.8 84.0 30.0 85.2 ;
      RECT  33.6 84.0 34.8 85.2 ;
      RECT  38.4 84.0 39.6 85.2 ;
      RECT  43.2 84.0 44.4 85.2 ;
      RECT  48.0 84.0 49.2 85.2 ;
      RECT  52.8 84.0 54.0 85.2 ;
      RECT  57.6 84.0 58.8 85.2 ;
      RECT  62.4 84.0 63.6 85.2 ;
      RECT  67.2 84.0 68.4 85.2 ;
      RECT  72.0 84.0 73.2 85.2 ;
      RECT  76.8 84.0 78.0 85.2 ;
      RECT  81.6 84.0 82.8 85.2 ;
      RECT  86.4 84.0 87.6 85.2 ;
      RECT  91.2 84.0 92.4 85.2 ;
      RECT  96.0 84.0 97.2 85.2 ;
      RECT  100.8 84.0 102.0 85.2 ;
      RECT  105.6 84.0 106.8 85.2 ;
      RECT  110.4 84.0 111.6 85.2 ;
      RECT  115.2 84.0 116.4 85.2 ;
      RECT  120.0 84.0 121.2 85.2 ;
      RECT  124.8 84.0 126.0 85.2 ;
      RECT  129.6 84.0 130.8 85.2 ;
      RECT  134.4 84.0 135.6 85.2 ;
      RECT  139.2 84.0 140.4 85.2 ;
      RECT  144.0 84.0 145.2 85.2 ;
      RECT  148.8 84.0 150.0 85.2 ;
      RECT  153.6 84.0 154.8 85.2 ;
      RECT  158.4 84.0 159.6 85.2 ;
      RECT  163.2 84.0 164.4 85.2 ;
      RECT  168.0 84.0 169.2 85.2 ;
      RECT  172.8 84.0 174.0 85.2 ;
      RECT  177.6 84.0 178.8 85.2 ;
      RECT  182.4 84.0 183.6 85.2 ;
      RECT  187.2 84.0 188.4 85.2 ;
      RECT  192.0 84.0 193.2 85.2 ;
      RECT  196.8 84.0 198.0 85.2 ;
      RECT  201.6 84.0 202.8 85.2 ;
      RECT  206.4 84.0 207.6 85.2 ;
      RECT  211.2 84.0 212.4 85.2 ;
      RECT  216.0 84.0 217.2 85.2 ;
      RECT  220.8 84.0 222.0 85.2 ;
      RECT  225.6 84.0 226.8 85.2 ;
      RECT  4.8 88.8 6.0 90.0 ;
      RECT  9.6 88.8 10.8 90.0 ;
      RECT  14.4 88.8 15.6 90.0 ;
      RECT  19.2 88.8 20.4 90.0 ;
      RECT  24.0 88.8 25.2 90.0 ;
      RECT  28.8 88.8 30.0 90.0 ;
      RECT  33.6 88.8 34.8 90.0 ;
      RECT  38.4 88.8 39.6 90.0 ;
      RECT  43.2 88.8 44.4 90.0 ;
      RECT  48.0 88.8 49.2 90.0 ;
      RECT  52.8 88.8 54.0 90.0 ;
      RECT  57.6 88.8 58.8 90.0 ;
      RECT  62.4 88.8 63.6 90.0 ;
      RECT  67.2 88.8 68.4 90.0 ;
      RECT  72.0 88.8 73.2 90.0 ;
      RECT  76.8 88.8 78.0 90.0 ;
      RECT  81.6 88.8 82.8 90.0 ;
      RECT  4.8 93.6 6.0 94.8 ;
      RECT  9.6 93.6 10.8 94.8 ;
      RECT  14.4 93.6 15.6 94.8 ;
      RECT  19.2 93.6 20.4 94.8 ;
      RECT  24.0 93.6 25.2 94.8 ;
      RECT  28.8 93.6 30.0 94.8 ;
      RECT  33.6 93.6 34.8 94.8 ;
      RECT  38.4 93.6 39.6 94.8 ;
      RECT  43.2 93.6 44.4 94.8 ;
      RECT  48.0 93.6 49.2 94.8 ;
      RECT  52.8 93.6 54.0 94.8 ;
      RECT  57.6 93.6 58.8 94.8 ;
      RECT  62.4 93.6 63.6 94.8 ;
      RECT  67.2 93.6 68.4 94.8 ;
      RECT  72.0 93.6 73.2 94.8 ;
      RECT  76.8 93.6 78.0 94.8 ;
      RECT  81.6 93.6 82.8 94.8 ;
      RECT  86.4 93.6 87.6 94.8 ;
      RECT  91.2 93.6 92.4 94.8 ;
      RECT  96.0 93.6 97.2 94.8 ;
      RECT  100.8 93.6 102.0 94.8 ;
      RECT  105.6 93.6 106.8 94.8 ;
      RECT  110.4 93.6 111.6 94.8 ;
      RECT  115.2 93.6 116.4 94.8 ;
      RECT  120.0 93.6 121.2 94.8 ;
      RECT  124.8 93.6 126.0 94.8 ;
      RECT  129.6 93.6 130.8 94.8 ;
      RECT  134.4 93.6 135.6 94.8 ;
      RECT  139.2 93.6 140.4 94.8 ;
      RECT  144.0 93.6 145.2 94.8 ;
      RECT  148.8 93.6 150.0 94.8 ;
      RECT  153.6 93.6 154.8 94.8 ;
      RECT  158.4 93.6 159.6 94.8 ;
      RECT  163.2 93.6 164.4 94.8 ;
      RECT  168.0 93.6 169.2 94.8 ;
      RECT  172.8 93.6 174.0 94.8 ;
      RECT  177.6 93.6 178.8 94.8 ;
      RECT  182.4 93.6 183.6 94.8 ;
      RECT  187.2 93.6 188.4 94.8 ;
      RECT  192.0 93.6 193.2 94.8 ;
      RECT  196.8 93.6 198.0 94.8 ;
      RECT  4.8 98.4 6.0 99.6 ;
      RECT  9.6 98.4 10.8 99.6 ;
      RECT  14.4 98.4 15.6 99.6 ;
      RECT  19.2 98.4 20.4 99.6 ;
      RECT  24.0 98.4 25.2 99.6 ;
      RECT  28.8 98.4 30.0 99.6 ;
      RECT  33.6 98.4 34.8 99.6 ;
      RECT  38.4 98.4 39.6 99.6 ;
      RECT  43.2 98.4 44.4 99.6 ;
      RECT  48.0 98.4 49.2 99.6 ;
      RECT  52.8 98.4 54.0 99.6 ;
      RECT  57.6 98.4 58.8 99.6 ;
      RECT  62.4 98.4 63.6 99.6 ;
      RECT  67.2 98.4 68.4 99.6 ;
      RECT  72.0 98.4 73.2 99.6 ;
      RECT  76.8 98.4 78.0 99.6 ;
      RECT  81.6 98.4 82.8 99.6 ;
      RECT  86.4 98.4 87.6 99.6 ;
      RECT  91.2 98.4 92.4 99.6 ;
      RECT  96.0 98.4 97.2 99.6 ;
      RECT  100.8 98.4 102.0 99.6 ;
      RECT  105.6 98.4 106.8 99.6 ;
      RECT  110.4 98.4 111.6 99.6 ;
      RECT  115.2 98.4 116.4 99.6 ;
      RECT  120.0 98.4 121.2 99.6 ;
      RECT  124.8 98.4 126.0 99.6 ;
      RECT  129.6 98.4 130.8 99.6 ;
      RECT  134.4 98.4 135.6 99.6 ;
      RECT  139.2 98.4 140.4 99.6 ;
      RECT  144.0 98.4 145.2 99.6 ;
      RECT  148.8 98.4 150.0 99.6 ;
      RECT  153.6 98.4 154.8 99.6 ;
      RECT  158.4 98.4 159.6 99.6 ;
      RECT  163.2 98.4 164.4 99.6 ;
      RECT  168.0 98.4 169.2 99.6 ;
      RECT  172.8 98.4 174.0 99.6 ;
      RECT  177.6 98.4 178.8 99.6 ;
      RECT  182.4 98.4 183.6 99.6 ;
      RECT  187.2 98.4 188.4 99.6 ;
      RECT  192.0 98.4 193.2 99.6 ;
      RECT  196.8 98.4 198.0 99.6 ;
      RECT  201.6 98.4 202.8 99.6 ;
      RECT  206.4 98.4 207.6 99.6 ;
      RECT  211.2 98.4 212.4 99.6 ;
      RECT  216.0 98.4 217.2 99.6 ;
      RECT  220.8 98.4 222.0 99.6 ;
      RECT  225.6 98.4 226.8 99.6 ;
      RECT  4.8 103.2 6.0 104.4 ;
      RECT  9.6 103.2 10.8 104.4 ;
      RECT  14.4 103.2 15.6 104.4 ;
      RECT  19.2 103.2 20.4 104.4 ;
      RECT  24.0 103.2 25.2 104.4 ;
      RECT  28.8 103.2 30.0 104.4 ;
      RECT  33.6 103.2 34.8 104.4 ;
      RECT  38.4 103.2 39.6 104.4 ;
      RECT  43.2 103.2 44.4 104.4 ;
      RECT  48.0 103.2 49.2 104.4 ;
      RECT  52.8 103.2 54.0 104.4 ;
      RECT  57.6 103.2 58.8 104.4 ;
      RECT  62.4 103.2 63.6 104.4 ;
      RECT  67.2 103.2 68.4 104.4 ;
      RECT  72.0 103.2 73.2 104.4 ;
      RECT  76.8 103.2 78.0 104.4 ;
      RECT  81.6 103.2 82.8 104.4 ;
      RECT  86.4 103.2 87.6 104.4 ;
      RECT  91.2 103.2 92.4 104.4 ;
      RECT  96.0 103.2 97.2 104.4 ;
      RECT  100.8 103.2 102.0 104.4 ;
      RECT  105.6 103.2 106.8 104.4 ;
      RECT  110.4 103.2 111.6 104.4 ;
      RECT  115.2 103.2 116.4 104.4 ;
      RECT  120.0 103.2 121.2 104.4 ;
      RECT  124.8 103.2 126.0 104.4 ;
      RECT  129.6 103.2 130.8 104.4 ;
      RECT  134.4 103.2 135.6 104.4 ;
      RECT  139.2 103.2 140.4 104.4 ;
      RECT  144.0 103.2 145.2 104.4 ;
      RECT  148.8 103.2 150.0 104.4 ;
      RECT  153.6 103.2 154.8 104.4 ;
      RECT  158.4 103.2 159.6 104.4 ;
      RECT  163.2 103.2 164.4 104.4 ;
      RECT  168.0 103.2 169.2 104.4 ;
      RECT  172.8 103.2 174.0 104.4 ;
      RECT  177.6 103.2 178.8 104.4 ;
      RECT  182.4 103.2 183.6 104.4 ;
      RECT  187.2 103.2 188.4 104.4 ;
      RECT  192.0 103.2 193.2 104.4 ;
      RECT  196.8 103.2 198.0 104.4 ;
      RECT  201.6 103.2 202.8 104.4 ;
      RECT  206.4 103.2 207.6 104.4 ;
      RECT  211.2 103.2 212.4 104.4 ;
      RECT  216.0 103.2 217.2 104.4 ;
      RECT  220.8 103.2 222.0 104.4 ;
      RECT  225.6 103.2 226.8 104.4 ;
      RECT  4.8 108.0 6.0 109.2 ;
      RECT  9.6 108.0 10.8 109.2 ;
      RECT  14.4 108.0 15.6 109.2 ;
      RECT  19.2 108.0 20.4 109.2 ;
      RECT  24.0 108.0 25.2 109.2 ;
      RECT  28.8 108.0 30.0 109.2 ;
      RECT  33.6 108.0 34.8 109.2 ;
      RECT  38.4 108.0 39.6 109.2 ;
      RECT  43.2 108.0 44.4 109.2 ;
      RECT  48.0 108.0 49.2 109.2 ;
      RECT  52.8 108.0 54.0 109.2 ;
      RECT  57.6 108.0 58.8 109.2 ;
      RECT  62.4 108.0 63.6 109.2 ;
      RECT  67.2 108.0 68.4 109.2 ;
      RECT  72.0 108.0 73.2 109.2 ;
      RECT  76.8 108.0 78.0 109.2 ;
      RECT  81.6 108.0 82.8 109.2 ;
      RECT  86.4 108.0 87.6 109.2 ;
      RECT  91.2 108.0 92.4 109.2 ;
      RECT  96.0 108.0 97.2 109.2 ;
      RECT  100.8 108.0 102.0 109.2 ;
      RECT  105.6 108.0 106.8 109.2 ;
      RECT  110.4 108.0 111.6 109.2 ;
      RECT  115.2 108.0 116.4 109.2 ;
      RECT  120.0 108.0 121.2 109.2 ;
      RECT  124.8 108.0 126.0 109.2 ;
      RECT  129.6 108.0 130.8 109.2 ;
      RECT  134.4 108.0 135.6 109.2 ;
      RECT  139.2 108.0 140.4 109.2 ;
      RECT  144.0 108.0 145.2 109.2 ;
      RECT  148.8 108.0 150.0 109.2 ;
      RECT  153.6 108.0 154.8 109.2 ;
      RECT  158.4 108.0 159.6 109.2 ;
      RECT  163.2 108.0 164.4 109.2 ;
      RECT  168.0 108.0 169.2 109.2 ;
      RECT  172.8 108.0 174.0 109.2 ;
      RECT  177.6 108.0 178.8 109.2 ;
      RECT  182.4 108.0 183.6 109.2 ;
      RECT  187.2 108.0 188.4 109.2 ;
      RECT  192.0 108.0 193.2 109.2 ;
      RECT  196.8 108.0 198.0 109.2 ;
      RECT  4.8 112.8 6.0 114.0 ;
      RECT  9.6 112.8 10.8 114.0 ;
      RECT  14.4 112.8 15.6 114.0 ;
      RECT  19.2 112.8 20.4 114.0 ;
      RECT  24.0 112.8 25.2 114.0 ;
      RECT  28.8 112.8 30.0 114.0 ;
      RECT  33.6 112.8 34.8 114.0 ;
      RECT  38.4 112.8 39.6 114.0 ;
      RECT  43.2 112.8 44.4 114.0 ;
      RECT  48.0 112.8 49.2 114.0 ;
      RECT  52.8 112.8 54.0 114.0 ;
      RECT  57.6 112.8 58.8 114.0 ;
      RECT  62.4 112.8 63.6 114.0 ;
      RECT  67.2 112.8 68.4 114.0 ;
      RECT  72.0 112.8 73.2 114.0 ;
      RECT  76.8 112.8 78.0 114.0 ;
      RECT  81.6 112.8 82.8 114.0 ;
      RECT  187.2 112.8 188.4 114.0 ;
      RECT  192.0 112.8 193.2 114.0 ;
      RECT  196.8 112.8 198.0 114.0 ;
      RECT  201.6 112.8 202.8 114.0 ;
      RECT  206.4 112.8 207.6 114.0 ;
      RECT  211.2 112.8 212.4 114.0 ;
      RECT  216.0 112.8 217.2 114.0 ;
      RECT  220.8 112.8 222.0 114.0 ;
      RECT  225.6 112.8 226.8 114.0 ;
      RECT  4.8 117.6 6.0 118.8 ;
      RECT  9.6 117.6 10.8 118.8 ;
      RECT  14.4 117.6 15.6 118.8 ;
      RECT  19.2 117.6 20.4 118.8 ;
      RECT  24.0 117.6 25.2 118.8 ;
      RECT  28.8 117.6 30.0 118.8 ;
      RECT  33.6 117.6 34.8 118.8 ;
      RECT  38.4 117.6 39.6 118.8 ;
      RECT  43.2 117.6 44.4 118.8 ;
      RECT  48.0 117.6 49.2 118.8 ;
      RECT  52.8 117.6 54.0 118.8 ;
      RECT  57.6 117.6 58.8 118.8 ;
      RECT  62.4 117.6 63.6 118.8 ;
      RECT  67.2 117.6 68.4 118.8 ;
      RECT  72.0 117.6 73.2 118.8 ;
      RECT  76.8 117.6 78.0 118.8 ;
      RECT  81.6 117.6 82.8 118.8 ;
      RECT  86.4 117.6 87.6 118.8 ;
      RECT  91.2 117.6 92.4 118.8 ;
      RECT  96.0 117.6 97.2 118.8 ;
      RECT  100.8 117.6 102.0 118.8 ;
      RECT  105.6 117.6 106.8 118.8 ;
      RECT  110.4 117.6 111.6 118.8 ;
      RECT  115.2 117.6 116.4 118.8 ;
      RECT  120.0 117.6 121.2 118.8 ;
      RECT  124.8 117.6 126.0 118.8 ;
      RECT  129.6 117.6 130.8 118.8 ;
      RECT  134.4 117.6 135.6 118.8 ;
      RECT  139.2 117.6 140.4 118.8 ;
      RECT  144.0 117.6 145.2 118.8 ;
      RECT  148.8 117.6 150.0 118.8 ;
      RECT  153.6 117.6 154.8 118.8 ;
      RECT  158.4 117.6 159.6 118.8 ;
      RECT  163.2 117.6 164.4 118.8 ;
      RECT  168.0 117.6 169.2 118.8 ;
      RECT  172.8 117.6 174.0 118.8 ;
      RECT  177.6 117.6 178.8 118.8 ;
      RECT  182.4 117.6 183.6 118.8 ;
      RECT  187.2 117.6 188.4 118.8 ;
      RECT  192.0 117.6 193.2 118.8 ;
      RECT  196.8 117.6 198.0 118.8 ;
      RECT  201.6 117.6 202.8 118.8 ;
      RECT  206.4 117.6 207.6 118.8 ;
      RECT  211.2 117.6 212.4 118.8 ;
      RECT  216.0 117.6 217.2 118.8 ;
      RECT  220.8 117.6 222.0 118.8 ;
      RECT  225.6 117.6 226.8 118.8 ;
      RECT  4.8 122.4 6.0 123.6 ;
      RECT  9.6 122.4 10.8 123.6 ;
      RECT  14.4 122.4 15.6 123.6 ;
      RECT  19.2 122.4 20.4 123.6 ;
      RECT  24.0 122.4 25.2 123.6 ;
      RECT  28.8 122.4 30.0 123.6 ;
      RECT  33.6 122.4 34.8 123.6 ;
      RECT  38.4 122.4 39.6 123.6 ;
      RECT  43.2 122.4 44.4 123.6 ;
      RECT  48.0 122.4 49.2 123.6 ;
      RECT  52.8 122.4 54.0 123.6 ;
      RECT  57.6 122.4 58.8 123.6 ;
      RECT  62.4 122.4 63.6 123.6 ;
      RECT  67.2 122.4 68.4 123.6 ;
      RECT  72.0 122.4 73.2 123.6 ;
      RECT  76.8 122.4 78.0 123.6 ;
      RECT  91.2 122.4 92.4 123.6 ;
      RECT  96.0 122.4 97.2 123.6 ;
      RECT  100.8 122.4 102.0 123.6 ;
      RECT  105.6 122.4 106.8 123.6 ;
      RECT  110.4 122.4 111.6 123.6 ;
      RECT  115.2 122.4 116.4 123.6 ;
      RECT  120.0 122.4 121.2 123.6 ;
      RECT  124.8 122.4 126.0 123.6 ;
      RECT  129.6 122.4 130.8 123.6 ;
      RECT  134.4 122.4 135.6 123.6 ;
      RECT  139.2 122.4 140.4 123.6 ;
      RECT  144.0 122.4 145.2 123.6 ;
      RECT  148.8 122.4 150.0 123.6 ;
      RECT  153.6 122.4 154.8 123.6 ;
      RECT  158.4 122.4 159.6 123.6 ;
      RECT  163.2 122.4 164.4 123.6 ;
      RECT  168.0 122.4 169.2 123.6 ;
      RECT  172.8 122.4 174.0 123.6 ;
      RECT  177.6 122.4 178.8 123.6 ;
      RECT  182.4 122.4 183.6 123.6 ;
      RECT  187.2 122.4 188.4 123.6 ;
      RECT  192.0 122.4 193.2 123.6 ;
      RECT  196.8 122.4 198.0 123.6 ;
      RECT  201.6 122.4 202.8 123.6 ;
      RECT  206.4 122.4 207.6 123.6 ;
      RECT  211.2 122.4 212.4 123.6 ;
      RECT  216.0 122.4 217.2 123.6 ;
      RECT  220.8 122.4 222.0 123.6 ;
      RECT  225.6 122.4 226.8 123.6 ;
      RECT  4.8 127.2 6.0 128.4 ;
      RECT  9.6 127.2 10.8 128.4 ;
      RECT  14.4 127.2 15.6 128.4 ;
      RECT  19.2 127.2 20.4 128.4 ;
      RECT  24.0 127.2 25.2 128.4 ;
      RECT  28.8 127.2 30.0 128.4 ;
      RECT  33.6 127.2 34.8 128.4 ;
      RECT  38.4 127.2 39.6 128.4 ;
      RECT  43.2 127.2 44.4 128.4 ;
      RECT  48.0 127.2 49.2 128.4 ;
      RECT  52.8 127.2 54.0 128.4 ;
      RECT  57.6 127.2 58.8 128.4 ;
      RECT  62.4 127.2 63.6 128.4 ;
      RECT  67.2 127.2 68.4 128.4 ;
      RECT  72.0 127.2 73.2 128.4 ;
      RECT  76.8 127.2 78.0 128.4 ;
      RECT  81.6 127.2 82.8 128.4 ;
      RECT  86.4 127.2 87.6 128.4 ;
      RECT  91.2 127.2 92.4 128.4 ;
      RECT  96.0 127.2 97.2 128.4 ;
      RECT  100.8 127.2 102.0 128.4 ;
      RECT  105.6 127.2 106.8 128.4 ;
      RECT  110.4 127.2 111.6 128.4 ;
      RECT  115.2 127.2 116.4 128.4 ;
      RECT  120.0 127.2 121.2 128.4 ;
      RECT  124.8 127.2 126.0 128.4 ;
      RECT  129.6 127.2 130.8 128.4 ;
      RECT  134.4 127.2 135.6 128.4 ;
      RECT  139.2 127.2 140.4 128.4 ;
      RECT  144.0 127.2 145.2 128.4 ;
      RECT  148.8 127.2 150.0 128.4 ;
      RECT  153.6 127.2 154.8 128.4 ;
      RECT  158.4 127.2 159.6 128.4 ;
      RECT  163.2 127.2 164.4 128.4 ;
      RECT  168.0 127.2 169.2 128.4 ;
      RECT  172.8 127.2 174.0 128.4 ;
      RECT  177.6 127.2 178.8 128.4 ;
      RECT  182.4 127.2 183.6 128.4 ;
      RECT  187.2 127.2 188.4 128.4 ;
      RECT  192.0 127.2 193.2 128.4 ;
      RECT  196.8 127.2 198.0 128.4 ;
      RECT  201.6 127.2 202.8 128.4 ;
      RECT  206.4 127.2 207.6 128.4 ;
      RECT  211.2 127.2 212.4 128.4 ;
      RECT  216.0 127.2 217.2 128.4 ;
      RECT  220.8 127.2 222.0 128.4 ;
      RECT  225.6 127.2 226.8 128.4 ;
      RECT  4.8 132.0 6.0 133.2 ;
      RECT  9.6 132.0 10.8 133.2 ;
      RECT  14.4 132.0 15.6 133.2 ;
      RECT  19.2 132.0 20.4 133.2 ;
      RECT  24.0 132.0 25.2 133.2 ;
      RECT  28.8 132.0 30.0 133.2 ;
      RECT  57.6 132.0 58.8 133.2 ;
      RECT  62.4 132.0 63.6 133.2 ;
      RECT  67.2 132.0 68.4 133.2 ;
      RECT  72.0 132.0 73.2 133.2 ;
      RECT  76.8 132.0 78.0 133.2 ;
      RECT  81.6 132.0 82.8 133.2 ;
      RECT  86.4 132.0 87.6 133.2 ;
      RECT  91.2 132.0 92.4 133.2 ;
      RECT  96.0 132.0 97.2 133.2 ;
      RECT  100.8 132.0 102.0 133.2 ;
      RECT  105.6 132.0 106.8 133.2 ;
      RECT  110.4 132.0 111.6 133.2 ;
      RECT  115.2 132.0 116.4 133.2 ;
      RECT  120.0 132.0 121.2 133.2 ;
      RECT  124.8 132.0 126.0 133.2 ;
      RECT  129.6 132.0 130.8 133.2 ;
      RECT  134.4 132.0 135.6 133.2 ;
      RECT  139.2 132.0 140.4 133.2 ;
      RECT  144.0 132.0 145.2 133.2 ;
      RECT  148.8 132.0 150.0 133.2 ;
      RECT  153.6 132.0 154.8 133.2 ;
      RECT  158.4 132.0 159.6 133.2 ;
      RECT  163.2 132.0 164.4 133.2 ;
      RECT  168.0 132.0 169.2 133.2 ;
      RECT  172.8 132.0 174.0 133.2 ;
      RECT  177.6 132.0 178.8 133.2 ;
      RECT  182.4 132.0 183.6 133.2 ;
      RECT  187.2 132.0 188.4 133.2 ;
      RECT  192.0 132.0 193.2 133.2 ;
      RECT  196.8 132.0 198.0 133.2 ;
      RECT  201.6 132.0 202.8 133.2 ;
      RECT  206.4 132.0 207.6 133.2 ;
      RECT  211.2 132.0 212.4 133.2 ;
      RECT  216.0 132.0 217.2 133.2 ;
      RECT  220.8 132.0 222.0 133.2 ;
      RECT  225.6 132.0 226.8 133.2 ;
      RECT  4.8 136.8 6.0 138.0 ;
      RECT  9.6 136.8 10.8 138.0 ;
      RECT  14.4 136.8 15.6 138.0 ;
      RECT  19.2 136.8 20.4 138.0 ;
      RECT  24.0 136.8 25.2 138.0 ;
      RECT  28.8 136.8 30.0 138.0 ;
      RECT  33.6 136.8 34.8 138.0 ;
      RECT  38.4 136.8 39.6 138.0 ;
      RECT  43.2 136.8 44.4 138.0 ;
      RECT  48.0 136.8 49.2 138.0 ;
      RECT  52.8 136.8 54.0 138.0 ;
      RECT  57.6 136.8 58.8 138.0 ;
      RECT  62.4 136.8 63.6 138.0 ;
      RECT  67.2 136.8 68.4 138.0 ;
      RECT  72.0 136.8 73.2 138.0 ;
      RECT  76.8 136.8 78.0 138.0 ;
      RECT  81.6 136.8 82.8 138.0 ;
      RECT  86.4 136.8 87.6 138.0 ;
      RECT  91.2 136.8 92.4 138.0 ;
      RECT  96.0 136.8 97.2 138.0 ;
      RECT  100.8 136.8 102.0 138.0 ;
      RECT  105.6 136.8 106.8 138.0 ;
      RECT  110.4 136.8 111.6 138.0 ;
      RECT  115.2 136.8 116.4 138.0 ;
      RECT  120.0 136.8 121.2 138.0 ;
      RECT  124.8 136.8 126.0 138.0 ;
      RECT  129.6 136.8 130.8 138.0 ;
      RECT  134.4 136.8 135.6 138.0 ;
      RECT  139.2 136.8 140.4 138.0 ;
      RECT  144.0 136.8 145.2 138.0 ;
      RECT  148.8 136.8 150.0 138.0 ;
      RECT  153.6 136.8 154.8 138.0 ;
      RECT  158.4 136.8 159.6 138.0 ;
      RECT  163.2 136.8 164.4 138.0 ;
      RECT  168.0 136.8 169.2 138.0 ;
      RECT  172.8 136.8 174.0 138.0 ;
      RECT  177.6 136.8 178.8 138.0 ;
      RECT  182.4 136.8 183.6 138.0 ;
      RECT  187.2 136.8 188.4 138.0 ;
      RECT  192.0 136.8 193.2 138.0 ;
      RECT  196.8 136.8 198.0 138.0 ;
      RECT  201.6 136.8 202.8 138.0 ;
      RECT  206.4 136.8 207.6 138.0 ;
      RECT  211.2 136.8 212.4 138.0 ;
      RECT  216.0 136.8 217.2 138.0 ;
      RECT  220.8 136.8 222.0 138.0 ;
      RECT  225.6 136.8 226.8 138.0 ;
      RECT  4.8 141.6 6.0 142.8 ;
      RECT  9.6 141.6 10.8 142.8 ;
      RECT  14.4 141.6 15.6 142.8 ;
      RECT  19.2 141.6 20.4 142.8 ;
      RECT  24.0 141.6 25.2 142.8 ;
      RECT  28.8 141.6 30.0 142.8 ;
      RECT  33.6 141.6 34.8 142.8 ;
      RECT  38.4 141.6 39.6 142.8 ;
      RECT  43.2 141.6 44.4 142.8 ;
      RECT  48.0 141.6 49.2 142.8 ;
      RECT  52.8 141.6 54.0 142.8 ;
      RECT  57.6 141.6 58.8 142.8 ;
      RECT  62.4 141.6 63.6 142.8 ;
      RECT  67.2 141.6 68.4 142.8 ;
      RECT  72.0 141.6 73.2 142.8 ;
      RECT  76.8 141.6 78.0 142.8 ;
      RECT  81.6 141.6 82.8 142.8 ;
      RECT  86.4 141.6 87.6 142.8 ;
      RECT  91.2 141.6 92.4 142.8 ;
      RECT  96.0 141.6 97.2 142.8 ;
      RECT  100.8 141.6 102.0 142.8 ;
      RECT  105.6 141.6 106.8 142.8 ;
      RECT  110.4 141.6 111.6 142.8 ;
      RECT  115.2 141.6 116.4 142.8 ;
      RECT  120.0 141.6 121.2 142.8 ;
      RECT  124.8 141.6 126.0 142.8 ;
      RECT  129.6 141.6 130.8 142.8 ;
      RECT  134.4 141.6 135.6 142.8 ;
      RECT  139.2 141.6 140.4 142.8 ;
      RECT  144.0 141.6 145.2 142.8 ;
      RECT  148.8 141.6 150.0 142.8 ;
      RECT  153.6 141.6 154.8 142.8 ;
      RECT  158.4 141.6 159.6 142.8 ;
      RECT  163.2 141.6 164.4 142.8 ;
      RECT  168.0 141.6 169.2 142.8 ;
      RECT  172.8 141.6 174.0 142.8 ;
      RECT  177.6 141.6 178.8 142.8 ;
      RECT  182.4 141.6 183.6 142.8 ;
      RECT  187.2 141.6 188.4 142.8 ;
      RECT  192.0 141.6 193.2 142.8 ;
      RECT  196.8 141.6 198.0 142.8 ;
      RECT  201.6 141.6 202.8 142.8 ;
      RECT  206.4 141.6 207.6 142.8 ;
      RECT  211.2 141.6 212.4 142.8 ;
      RECT  216.0 141.6 217.2 142.8 ;
      RECT  220.8 141.6 222.0 142.8 ;
      RECT  225.6 141.6 226.8 142.8 ;
      RECT  4.8 146.4 6.0 147.6 ;
      RECT  9.6 146.4 10.8 147.6 ;
      RECT  14.4 146.4 15.6 147.6 ;
      RECT  19.2 146.4 20.4 147.6 ;
      RECT  24.0 146.4 25.2 147.6 ;
      RECT  28.8 146.4 30.0 147.6 ;
      RECT  33.6 146.4 34.8 147.6 ;
      RECT  38.4 146.4 39.6 147.6 ;
      RECT  43.2 146.4 44.4 147.6 ;
      RECT  48.0 146.4 49.2 147.6 ;
      RECT  52.8 146.4 54.0 147.6 ;
      RECT  57.6 146.4 58.8 147.6 ;
      RECT  62.4 146.4 63.6 147.6 ;
      RECT  67.2 146.4 68.4 147.6 ;
      RECT  72.0 146.4 73.2 147.6 ;
      RECT  76.8 146.4 78.0 147.6 ;
      RECT  81.6 146.4 82.8 147.6 ;
      RECT  86.4 146.4 87.6 147.6 ;
      RECT  91.2 146.4 92.4 147.6 ;
      RECT  96.0 146.4 97.2 147.6 ;
      RECT  100.8 146.4 102.0 147.6 ;
      RECT  105.6 146.4 106.8 147.6 ;
      RECT  110.4 146.4 111.6 147.6 ;
      RECT  115.2 146.4 116.4 147.6 ;
      RECT  120.0 146.4 121.2 147.6 ;
      RECT  124.8 146.4 126.0 147.6 ;
      RECT  129.6 146.4 130.8 147.6 ;
      RECT  134.4 146.4 135.6 147.6 ;
      RECT  139.2 146.4 140.4 147.6 ;
      RECT  144.0 146.4 145.2 147.6 ;
      RECT  148.8 146.4 150.0 147.6 ;
      RECT  153.6 146.4 154.8 147.6 ;
      RECT  158.4 146.4 159.6 147.6 ;
      RECT  163.2 146.4 164.4 147.6 ;
      RECT  168.0 146.4 169.2 147.6 ;
      RECT  172.8 146.4 174.0 147.6 ;
      RECT  177.6 146.4 178.8 147.6 ;
      RECT  182.4 146.4 183.6 147.6 ;
      RECT  187.2 146.4 188.4 147.6 ;
      RECT  192.0 146.4 193.2 147.6 ;
      RECT  196.8 146.4 198.0 147.6 ;
      RECT  4.8 151.2 6.0 152.4 ;
      RECT  9.6 151.2 10.8 152.4 ;
      RECT  14.4 151.2 15.6 152.4 ;
      RECT  19.2 151.2 20.4 152.4 ;
      RECT  24.0 151.2 25.2 152.4 ;
      RECT  28.8 151.2 30.0 152.4 ;
      RECT  33.6 151.2 34.8 152.4 ;
      RECT  38.4 151.2 39.6 152.4 ;
      RECT  43.2 151.2 44.4 152.4 ;
      RECT  48.0 151.2 49.2 152.4 ;
      RECT  52.8 151.2 54.0 152.4 ;
      RECT  57.6 151.2 58.8 152.4 ;
      RECT  62.4 151.2 63.6 152.4 ;
      RECT  67.2 151.2 68.4 152.4 ;
      RECT  72.0 151.2 73.2 152.4 ;
      RECT  76.8 151.2 78.0 152.4 ;
      RECT  81.6 151.2 82.8 152.4 ;
      RECT  187.2 151.2 188.4 152.4 ;
      RECT  192.0 151.2 193.2 152.4 ;
      RECT  196.8 151.2 198.0 152.4 ;
      RECT  201.6 151.2 202.8 152.4 ;
      RECT  206.4 151.2 207.6 152.4 ;
      RECT  211.2 151.2 212.4 152.4 ;
      RECT  216.0 151.2 217.2 152.4 ;
      RECT  220.8 151.2 222.0 152.4 ;
      RECT  225.6 151.2 226.8 152.4 ;
      RECT  4.8 156.0 6.0 157.2 ;
      RECT  9.6 156.0 10.8 157.2 ;
      RECT  14.4 156.0 15.6 157.2 ;
      RECT  19.2 156.0 20.4 157.2 ;
      RECT  24.0 156.0 25.2 157.2 ;
      RECT  28.8 156.0 30.0 157.2 ;
      RECT  33.6 156.0 34.8 157.2 ;
      RECT  38.4 156.0 39.6 157.2 ;
      RECT  43.2 156.0 44.4 157.2 ;
      RECT  48.0 156.0 49.2 157.2 ;
      RECT  52.8 156.0 54.0 157.2 ;
      RECT  57.6 156.0 58.8 157.2 ;
      RECT  62.4 156.0 63.6 157.2 ;
      RECT  67.2 156.0 68.4 157.2 ;
      RECT  72.0 156.0 73.2 157.2 ;
      RECT  76.8 156.0 78.0 157.2 ;
      RECT  81.6 156.0 82.8 157.2 ;
      RECT  86.4 156.0 87.6 157.2 ;
      RECT  91.2 156.0 92.4 157.2 ;
      RECT  96.0 156.0 97.2 157.2 ;
      RECT  100.8 156.0 102.0 157.2 ;
      RECT  105.6 156.0 106.8 157.2 ;
      RECT  110.4 156.0 111.6 157.2 ;
      RECT  115.2 156.0 116.4 157.2 ;
      RECT  120.0 156.0 121.2 157.2 ;
      RECT  124.8 156.0 126.0 157.2 ;
      RECT  129.6 156.0 130.8 157.2 ;
      RECT  134.4 156.0 135.6 157.2 ;
      RECT  139.2 156.0 140.4 157.2 ;
      RECT  144.0 156.0 145.2 157.2 ;
      RECT  148.8 156.0 150.0 157.2 ;
      RECT  153.6 156.0 154.8 157.2 ;
      RECT  158.4 156.0 159.6 157.2 ;
      RECT  163.2 156.0 164.4 157.2 ;
      RECT  168.0 156.0 169.2 157.2 ;
      RECT  172.8 156.0 174.0 157.2 ;
      RECT  177.6 156.0 178.8 157.2 ;
      RECT  182.4 156.0 183.6 157.2 ;
      RECT  187.2 156.0 188.4 157.2 ;
      RECT  192.0 156.0 193.2 157.2 ;
      RECT  196.8 156.0 198.0 157.2 ;
      RECT  201.6 156.0 202.8 157.2 ;
      RECT  206.4 156.0 207.6 157.2 ;
      RECT  211.2 156.0 212.4 157.2 ;
      RECT  216.0 156.0 217.2 157.2 ;
      RECT  220.8 156.0 222.0 157.2 ;
      RECT  225.6 156.0 226.8 157.2 ;
      RECT  4.8 160.8 6.0 162.0 ;
      RECT  9.6 160.8 10.8 162.0 ;
      RECT  14.4 160.8 15.6 162.0 ;
      RECT  19.2 160.8 20.4 162.0 ;
      RECT  24.0 160.8 25.2 162.0 ;
      RECT  28.8 160.8 30.0 162.0 ;
      RECT  33.6 160.8 34.8 162.0 ;
      RECT  38.4 160.8 39.6 162.0 ;
      RECT  43.2 160.8 44.4 162.0 ;
      RECT  48.0 160.8 49.2 162.0 ;
      RECT  52.8 160.8 54.0 162.0 ;
      RECT  57.6 160.8 58.8 162.0 ;
      RECT  62.4 160.8 63.6 162.0 ;
      RECT  67.2 160.8 68.4 162.0 ;
      RECT  72.0 160.8 73.2 162.0 ;
      RECT  76.8 160.8 78.0 162.0 ;
      RECT  91.2 160.8 92.4 162.0 ;
      RECT  96.0 160.8 97.2 162.0 ;
      RECT  100.8 160.8 102.0 162.0 ;
      RECT  105.6 160.8 106.8 162.0 ;
      RECT  110.4 160.8 111.6 162.0 ;
      RECT  115.2 160.8 116.4 162.0 ;
      RECT  120.0 160.8 121.2 162.0 ;
      RECT  124.8 160.8 126.0 162.0 ;
      RECT  129.6 160.8 130.8 162.0 ;
      RECT  134.4 160.8 135.6 162.0 ;
      RECT  139.2 160.8 140.4 162.0 ;
      RECT  144.0 160.8 145.2 162.0 ;
      RECT  148.8 160.8 150.0 162.0 ;
      RECT  153.6 160.8 154.8 162.0 ;
      RECT  158.4 160.8 159.6 162.0 ;
      RECT  163.2 160.8 164.4 162.0 ;
      RECT  168.0 160.8 169.2 162.0 ;
      RECT  172.8 160.8 174.0 162.0 ;
      RECT  177.6 160.8 178.8 162.0 ;
      RECT  182.4 160.8 183.6 162.0 ;
      RECT  187.2 160.8 188.4 162.0 ;
      RECT  192.0 160.8 193.2 162.0 ;
      RECT  196.8 160.8 198.0 162.0 ;
      RECT  201.6 160.8 202.8 162.0 ;
      RECT  206.4 160.8 207.6 162.0 ;
      RECT  211.2 160.8 212.4 162.0 ;
      RECT  216.0 160.8 217.2 162.0 ;
      RECT  220.8 160.8 222.0 162.0 ;
      RECT  225.6 160.8 226.8 162.0 ;
      RECT  201.6 165.6 202.8 166.8 ;
      RECT  206.4 165.6 207.6 166.8 ;
      RECT  211.2 165.6 212.4 166.8 ;
      RECT  216.0 165.6 217.2 166.8 ;
      RECT  220.8 165.6 222.0 166.8 ;
      RECT  225.6 165.6 226.8 166.8 ;
      RECT  33.6 170.4 34.8 171.6 ;
      RECT  38.4 170.4 39.6 171.6 ;
      RECT  43.2 170.4 44.4 171.6 ;
      RECT  48.0 170.4 49.2 171.6 ;
      RECT  52.8 170.4 54.0 171.6 ;
      RECT  57.6 170.4 58.8 171.6 ;
      RECT  62.4 170.4 63.6 171.6 ;
      RECT  67.2 170.4 68.4 171.6 ;
      RECT  72.0 170.4 73.2 171.6 ;
      RECT  76.8 170.4 78.0 171.6 ;
      RECT  81.6 170.4 82.8 171.6 ;
      RECT  86.4 170.4 87.6 171.6 ;
      RECT  91.2 170.4 92.4 171.6 ;
      RECT  96.0 170.4 97.2 171.6 ;
      RECT  100.8 170.4 102.0 171.6 ;
      RECT  105.6 170.4 106.8 171.6 ;
      RECT  110.4 170.4 111.6 171.6 ;
      RECT  115.2 170.4 116.4 171.6 ;
      RECT  120.0 170.4 121.2 171.6 ;
      RECT  124.8 170.4 126.0 171.6 ;
      RECT  129.6 170.4 130.8 171.6 ;
      RECT  134.4 170.4 135.6 171.6 ;
      RECT  139.2 170.4 140.4 171.6 ;
      RECT  144.0 170.4 145.2 171.6 ;
      RECT  148.8 170.4 150.0 171.6 ;
      RECT  153.6 170.4 154.8 171.6 ;
      RECT  158.4 170.4 159.6 171.6 ;
      RECT  163.2 170.4 164.4 171.6 ;
      RECT  168.0 170.4 169.2 171.6 ;
      RECT  172.8 170.4 174.0 171.6 ;
      RECT  177.6 170.4 178.8 171.6 ;
      RECT  182.4 170.4 183.6 171.6 ;
      RECT  187.2 170.4 188.4 171.6 ;
      RECT  192.0 170.4 193.2 171.6 ;
      RECT  196.8 170.4 198.0 171.6 ;
      RECT  201.6 170.4 202.8 171.6 ;
      RECT  206.4 170.4 207.6 171.6 ;
      RECT  211.2 170.4 212.4 171.6 ;
      RECT  216.0 170.4 217.2 171.6 ;
      RECT  220.8 170.4 222.0 171.6 ;
      RECT  225.6 170.4 226.8 171.6 ;
      RECT  4.8 175.2 6.0 176.4 ;
      RECT  9.6 175.2 10.8 176.4 ;
      RECT  14.4 175.2 15.6 176.4 ;
      RECT  19.2 175.2 20.4 176.4 ;
      RECT  24.0 175.2 25.2 176.4 ;
      RECT  28.8 175.2 30.0 176.4 ;
      RECT  33.6 175.2 34.8 176.4 ;
      RECT  38.4 175.2 39.6 176.4 ;
      RECT  43.2 175.2 44.4 176.4 ;
      RECT  48.0 175.2 49.2 176.4 ;
      RECT  52.8 175.2 54.0 176.4 ;
      RECT  57.6 175.2 58.8 176.4 ;
      RECT  62.4 175.2 63.6 176.4 ;
      RECT  67.2 175.2 68.4 176.4 ;
      RECT  72.0 175.2 73.2 176.4 ;
      RECT  76.8 175.2 78.0 176.4 ;
      RECT  81.6 175.2 82.8 176.4 ;
      RECT  86.4 175.2 87.6 176.4 ;
      RECT  91.2 175.2 92.4 176.4 ;
      RECT  96.0 175.2 97.2 176.4 ;
      RECT  100.8 175.2 102.0 176.4 ;
      RECT  105.6 175.2 106.8 176.4 ;
      RECT  110.4 175.2 111.6 176.4 ;
      RECT  115.2 175.2 116.4 176.4 ;
      RECT  120.0 175.2 121.2 176.4 ;
      RECT  124.8 175.2 126.0 176.4 ;
      RECT  129.6 175.2 130.8 176.4 ;
      RECT  134.4 175.2 135.6 176.4 ;
      RECT  139.2 175.2 140.4 176.4 ;
      RECT  144.0 175.2 145.2 176.4 ;
      RECT  148.8 175.2 150.0 176.4 ;
      RECT  153.6 175.2 154.8 176.4 ;
      RECT  158.4 175.2 159.6 176.4 ;
      RECT  163.2 175.2 164.4 176.4 ;
      RECT  168.0 175.2 169.2 176.4 ;
      RECT  172.8 175.2 174.0 176.4 ;
      RECT  177.6 175.2 178.8 176.4 ;
      RECT  182.4 175.2 183.6 176.4 ;
      RECT  187.2 175.2 188.4 176.4 ;
      RECT  192.0 175.2 193.2 176.4 ;
      RECT  196.8 175.2 198.0 176.4 ;
      RECT  201.6 175.2 202.8 176.4 ;
      RECT  206.4 175.2 207.6 176.4 ;
      RECT  211.2 175.2 212.4 176.4 ;
      RECT  216.0 175.2 217.2 176.4 ;
      RECT  220.8 175.2 222.0 176.4 ;
      RECT  225.6 175.2 226.8 176.4 ;
      RECT  33.6 180.0 34.8 181.2 ;
      RECT  38.4 180.0 39.6 181.2 ;
      RECT  43.2 180.0 44.4 181.2 ;
      RECT  48.0 180.0 49.2 181.2 ;
      RECT  52.8 180.0 54.0 181.2 ;
      RECT  57.6 180.0 58.8 181.2 ;
      RECT  62.4 180.0 63.6 181.2 ;
      RECT  67.2 180.0 68.4 181.2 ;
      RECT  72.0 180.0 73.2 181.2 ;
      RECT  76.8 180.0 78.0 181.2 ;
      RECT  81.6 180.0 82.8 181.2 ;
      RECT  86.4 180.0 87.6 181.2 ;
      RECT  91.2 180.0 92.4 181.2 ;
      RECT  96.0 180.0 97.2 181.2 ;
      RECT  100.8 180.0 102.0 181.2 ;
      RECT  105.6 180.0 106.8 181.2 ;
      RECT  110.4 180.0 111.6 181.2 ;
      RECT  115.2 180.0 116.4 181.2 ;
      RECT  120.0 180.0 121.2 181.2 ;
      RECT  124.8 180.0 126.0 181.2 ;
      RECT  129.6 180.0 130.8 181.2 ;
      RECT  134.4 180.0 135.6 181.2 ;
      RECT  139.2 180.0 140.4 181.2 ;
      RECT  144.0 180.0 145.2 181.2 ;
      RECT  148.8 180.0 150.0 181.2 ;
      RECT  153.6 180.0 154.8 181.2 ;
      RECT  158.4 180.0 159.6 181.2 ;
      RECT  163.2 180.0 164.4 181.2 ;
      RECT  168.0 180.0 169.2 181.2 ;
      RECT  172.8 180.0 174.0 181.2 ;
      RECT  177.6 180.0 178.8 181.2 ;
      RECT  24.0 184.8 25.2 186.0 ;
      RECT  28.8 184.8 30.0 186.0 ;
      RECT  33.6 184.8 34.8 186.0 ;
      RECT  38.4 184.8 39.6 186.0 ;
      RECT  43.2 184.8 44.4 186.0 ;
      RECT  48.0 184.8 49.2 186.0 ;
      RECT  52.8 184.8 54.0 186.0 ;
      RECT  57.6 184.8 58.8 186.0 ;
      RECT  62.4 184.8 63.6 186.0 ;
      RECT  67.2 184.8 68.4 186.0 ;
      RECT  72.0 184.8 73.2 186.0 ;
      RECT  76.8 184.8 78.0 186.0 ;
      RECT  81.6 184.8 82.8 186.0 ;
      RECT  86.4 184.8 87.6 186.0 ;
      RECT  91.2 184.8 92.4 186.0 ;
      RECT  96.0 184.8 97.2 186.0 ;
      RECT  100.8 184.8 102.0 186.0 ;
      RECT  105.6 184.8 106.8 186.0 ;
      RECT  110.4 184.8 111.6 186.0 ;
      RECT  115.2 184.8 116.4 186.0 ;
      RECT  120.0 184.8 121.2 186.0 ;
      RECT  124.8 184.8 126.0 186.0 ;
      RECT  129.6 184.8 130.8 186.0 ;
      RECT  134.4 184.8 135.6 186.0 ;
      RECT  139.2 184.8 140.4 186.0 ;
      RECT  144.0 184.8 145.2 186.0 ;
      RECT  148.8 184.8 150.0 186.0 ;
      RECT  153.6 184.8 154.8 186.0 ;
      RECT  158.4 184.8 159.6 186.0 ;
      RECT  163.2 184.8 164.4 186.0 ;
      RECT  168.0 184.8 169.2 186.0 ;
      RECT  172.8 184.8 174.0 186.0 ;
      RECT  177.6 184.8 178.8 186.0 ;
      RECT  182.4 184.8 183.6 186.0 ;
      RECT  187.2 184.8 188.4 186.0 ;
      RECT  192.0 184.8 193.2 186.0 ;
      RECT  196.8 184.8 198.0 186.0 ;
      RECT  201.6 184.8 202.8 186.0 ;
      RECT  206.4 184.8 207.6 186.0 ;
      RECT  211.2 184.8 212.4 186.0 ;
      RECT  216.0 184.8 217.2 186.0 ;
      RECT  220.8 184.8 222.0 186.0 ;
      RECT  225.6 184.8 226.8 186.0 ;
      RECT  33.6 189.6 34.8 190.8 ;
      RECT  38.4 189.6 39.6 190.8 ;
      RECT  43.2 189.6 44.4 190.8 ;
      RECT  48.0 189.6 49.2 190.8 ;
      RECT  52.8 189.6 54.0 190.8 ;
      RECT  57.6 189.6 58.8 190.8 ;
      RECT  62.4 189.6 63.6 190.8 ;
      RECT  67.2 189.6 68.4 190.8 ;
      RECT  72.0 189.6 73.2 190.8 ;
      RECT  76.8 189.6 78.0 190.8 ;
      RECT  81.6 189.6 82.8 190.8 ;
      RECT  86.4 189.6 87.6 190.8 ;
      RECT  91.2 189.6 92.4 190.8 ;
      RECT  96.0 189.6 97.2 190.8 ;
      RECT  100.8 189.6 102.0 190.8 ;
      RECT  105.6 189.6 106.8 190.8 ;
      RECT  110.4 189.6 111.6 190.8 ;
      RECT  115.2 189.6 116.4 190.8 ;
      RECT  120.0 189.6 121.2 190.8 ;
      RECT  124.8 189.6 126.0 190.8 ;
      RECT  129.6 189.6 130.8 190.8 ;
      RECT  134.4 189.6 135.6 190.8 ;
      RECT  139.2 189.6 140.4 190.8 ;
      RECT  144.0 189.6 145.2 190.8 ;
      RECT  148.8 189.6 150.0 190.8 ;
      RECT  153.6 189.6 154.8 190.8 ;
      RECT  158.4 189.6 159.6 190.8 ;
      RECT  163.2 189.6 164.4 190.8 ;
      RECT  168.0 189.6 169.2 190.8 ;
      RECT  172.8 189.6 174.0 190.8 ;
      RECT  177.6 189.6 178.8 190.8 ;
      RECT  4.8 194.4 6.0 195.6 ;
      RECT  9.6 194.4 10.8 195.6 ;
      RECT  14.4 194.4 15.6 195.6 ;
      RECT  19.2 194.4 20.4 195.6 ;
      RECT  24.0 194.4 25.2 195.6 ;
      RECT  28.8 194.4 30.0 195.6 ;
      RECT  33.6 194.4 34.8 195.6 ;
      RECT  38.4 194.4 39.6 195.6 ;
      RECT  43.2 194.4 44.4 195.6 ;
      RECT  48.0 194.4 49.2 195.6 ;
      RECT  52.8 194.4 54.0 195.6 ;
      RECT  57.6 194.4 58.8 195.6 ;
      RECT  62.4 194.4 63.6 195.6 ;
      RECT  67.2 194.4 68.4 195.6 ;
      RECT  72.0 194.4 73.2 195.6 ;
      RECT  76.8 194.4 78.0 195.6 ;
      RECT  81.6 194.4 82.8 195.6 ;
      RECT  86.4 194.4 87.6 195.6 ;
      RECT  91.2 194.4 92.4 195.6 ;
      RECT  96.0 194.4 97.2 195.6 ;
      RECT  177.6 194.4 178.8 195.6 ;
      RECT  182.4 194.4 183.6 195.6 ;
      RECT  187.2 194.4 188.4 195.6 ;
      RECT  192.0 194.4 193.2 195.6 ;
      RECT  196.8 194.4 198.0 195.6 ;
      RECT  201.6 194.4 202.8 195.6 ;
      RECT  206.4 194.4 207.6 195.6 ;
      RECT  211.2 194.4 212.4 195.6 ;
      RECT  216.0 194.4 217.2 195.6 ;
      RECT  220.8 194.4 222.0 195.6 ;
      RECT  225.6 194.4 226.8 195.6 ;
      RECT  33.6 199.2 34.8 200.4 ;
      RECT  38.4 199.2 39.6 200.4 ;
      RECT  43.2 199.2 44.4 200.4 ;
      RECT  48.0 199.2 49.2 200.4 ;
      RECT  52.8 199.2 54.0 200.4 ;
      RECT  57.6 199.2 58.8 200.4 ;
      RECT  62.4 199.2 63.6 200.4 ;
      RECT  67.2 199.2 68.4 200.4 ;
      RECT  72.0 199.2 73.2 200.4 ;
      RECT  76.8 199.2 78.0 200.4 ;
      RECT  81.6 199.2 82.8 200.4 ;
      RECT  86.4 199.2 87.6 200.4 ;
      RECT  91.2 199.2 92.4 200.4 ;
      RECT  96.0 199.2 97.2 200.4 ;
      RECT  100.8 199.2 102.0 200.4 ;
      RECT  105.6 199.2 106.8 200.4 ;
      RECT  110.4 199.2 111.6 200.4 ;
      RECT  115.2 199.2 116.4 200.4 ;
      RECT  120.0 199.2 121.2 200.4 ;
      RECT  124.8 199.2 126.0 200.4 ;
      RECT  129.6 199.2 130.8 200.4 ;
      RECT  134.4 199.2 135.6 200.4 ;
      RECT  139.2 199.2 140.4 200.4 ;
      RECT  144.0 199.2 145.2 200.4 ;
      RECT  148.8 199.2 150.0 200.4 ;
      RECT  153.6 199.2 154.8 200.4 ;
      RECT  158.4 199.2 159.6 200.4 ;
      RECT  163.2 199.2 164.4 200.4 ;
      RECT  168.0 199.2 169.2 200.4 ;
      RECT  172.8 199.2 174.0 200.4 ;
      RECT  177.6 199.2 178.8 200.4 ;
      RECT  24.0 204.0 25.2 205.2 ;
      RECT  28.8 204.0 30.0 205.2 ;
      RECT  33.6 204.0 34.8 205.2 ;
      RECT  38.4 204.0 39.6 205.2 ;
      RECT  43.2 204.0 44.4 205.2 ;
      RECT  48.0 204.0 49.2 205.2 ;
      RECT  52.8 204.0 54.0 205.2 ;
      RECT  57.6 204.0 58.8 205.2 ;
      RECT  62.4 204.0 63.6 205.2 ;
      RECT  67.2 204.0 68.4 205.2 ;
      RECT  72.0 204.0 73.2 205.2 ;
      RECT  76.8 204.0 78.0 205.2 ;
      RECT  81.6 204.0 82.8 205.2 ;
      RECT  139.2 204.0 140.4 205.2 ;
      RECT  144.0 204.0 145.2 205.2 ;
      RECT  148.8 204.0 150.0 205.2 ;
      RECT  153.6 204.0 154.8 205.2 ;
      RECT  158.4 204.0 159.6 205.2 ;
      RECT  163.2 204.0 164.4 205.2 ;
      RECT  168.0 204.0 169.2 205.2 ;
      RECT  172.8 204.0 174.0 205.2 ;
      RECT  177.6 204.0 178.8 205.2 ;
      RECT  182.4 204.0 183.6 205.2 ;
      RECT  187.2 204.0 188.4 205.2 ;
      RECT  192.0 204.0 193.2 205.2 ;
      RECT  196.8 204.0 198.0 205.2 ;
      RECT  201.6 204.0 202.8 205.2 ;
      RECT  206.4 204.0 207.6 205.2 ;
      RECT  211.2 204.0 212.4 205.2 ;
      RECT  216.0 204.0 217.2 205.2 ;
      RECT  220.8 204.0 222.0 205.2 ;
      RECT  225.6 204.0 226.8 205.2 ;
      RECT  4.8 208.8 6.0 210.0 ;
      RECT  9.6 208.8 10.8 210.0 ;
      RECT  14.4 208.8 15.6 210.0 ;
      RECT  19.2 208.8 20.4 210.0 ;
      RECT  24.0 208.8 25.2 210.0 ;
      RECT  28.8 208.8 30.0 210.0 ;
      RECT  33.6 208.8 34.8 210.0 ;
      RECT  38.4 208.8 39.6 210.0 ;
      RECT  43.2 208.8 44.4 210.0 ;
      RECT  48.0 208.8 49.2 210.0 ;
      RECT  52.8 208.8 54.0 210.0 ;
      RECT  57.6 208.8 58.8 210.0 ;
      RECT  62.4 208.8 63.6 210.0 ;
      RECT  67.2 208.8 68.4 210.0 ;
      RECT  72.0 208.8 73.2 210.0 ;
      RECT  76.8 208.8 78.0 210.0 ;
      RECT  81.6 208.8 82.8 210.0 ;
      RECT  86.4 208.8 87.6 210.0 ;
      RECT  91.2 208.8 92.4 210.0 ;
      RECT  96.0 208.8 97.2 210.0 ;
      RECT  100.8 208.8 102.0 210.0 ;
      RECT  105.6 208.8 106.8 210.0 ;
      RECT  110.4 208.8 111.6 210.0 ;
      RECT  115.2 208.8 116.4 210.0 ;
      RECT  120.0 208.8 121.2 210.0 ;
      RECT  124.8 208.8 126.0 210.0 ;
      RECT  129.6 208.8 130.8 210.0 ;
      RECT  134.4 208.8 135.6 210.0 ;
      RECT  139.2 208.8 140.4 210.0 ;
      RECT  144.0 208.8 145.2 210.0 ;
      RECT  148.8 208.8 150.0 210.0 ;
      RECT  153.6 208.8 154.8 210.0 ;
      RECT  158.4 208.8 159.6 210.0 ;
      RECT  163.2 208.8 164.4 210.0 ;
      RECT  168.0 208.8 169.2 210.0 ;
      RECT  172.8 208.8 174.0 210.0 ;
      RECT  177.6 208.8 178.8 210.0 ;
      RECT  4.8 213.6 6.0 214.8 ;
      RECT  9.6 213.6 10.8 214.8 ;
      RECT  14.4 213.6 15.6 214.8 ;
      RECT  19.2 213.6 20.4 214.8 ;
      RECT  24.0 213.6 25.2 214.8 ;
      RECT  28.8 213.6 30.0 214.8 ;
      RECT  33.6 213.6 34.8 214.8 ;
      RECT  38.4 213.6 39.6 214.8 ;
      RECT  43.2 213.6 44.4 214.8 ;
      RECT  48.0 213.6 49.2 214.8 ;
      RECT  52.8 213.6 54.0 214.8 ;
      RECT  57.6 213.6 58.8 214.8 ;
      RECT  62.4 213.6 63.6 214.8 ;
      RECT  67.2 213.6 68.4 214.8 ;
      RECT  72.0 213.6 73.2 214.8 ;
      RECT  76.8 213.6 78.0 214.8 ;
      RECT  81.6 213.6 82.8 214.8 ;
      RECT  86.4 213.6 87.6 214.8 ;
      RECT  91.2 213.6 92.4 214.8 ;
      RECT  96.0 213.6 97.2 214.8 ;
      RECT  177.6 213.6 178.8 214.8 ;
      RECT  182.4 213.6 183.6 214.8 ;
      RECT  187.2 213.6 188.4 214.8 ;
      RECT  192.0 213.6 193.2 214.8 ;
      RECT  196.8 213.6 198.0 214.8 ;
      RECT  201.6 213.6 202.8 214.8 ;
      RECT  206.4 213.6 207.6 214.8 ;
      RECT  211.2 213.6 212.4 214.8 ;
      RECT  216.0 213.6 217.2 214.8 ;
      RECT  220.8 213.6 222.0 214.8 ;
      RECT  225.6 213.6 226.8 214.8 ;
      RECT  4.8 218.4 6.0 219.6 ;
      RECT  9.6 218.4 10.8 219.6 ;
      RECT  14.4 218.4 15.6 219.6 ;
      RECT  19.2 218.4 20.4 219.6 ;
      RECT  24.0 218.4 25.2 219.6 ;
      RECT  28.8 218.4 30.0 219.6 ;
      RECT  33.6 218.4 34.8 219.6 ;
      RECT  38.4 218.4 39.6 219.6 ;
      RECT  43.2 218.4 44.4 219.6 ;
      RECT  48.0 218.4 49.2 219.6 ;
      RECT  52.8 218.4 54.0 219.6 ;
      RECT  57.6 218.4 58.8 219.6 ;
      RECT  62.4 218.4 63.6 219.6 ;
      RECT  67.2 218.4 68.4 219.6 ;
      RECT  72.0 218.4 73.2 219.6 ;
      RECT  76.8 218.4 78.0 219.6 ;
      RECT  81.6 218.4 82.8 219.6 ;
      RECT  86.4 218.4 87.6 219.6 ;
      RECT  91.2 218.4 92.4 219.6 ;
      RECT  96.0 218.4 97.2 219.6 ;
      RECT  100.8 218.4 102.0 219.6 ;
      RECT  105.6 218.4 106.8 219.6 ;
      RECT  110.4 218.4 111.6 219.6 ;
      RECT  115.2 218.4 116.4 219.6 ;
      RECT  120.0 218.4 121.2 219.6 ;
      RECT  124.8 218.4 126.0 219.6 ;
      RECT  129.6 218.4 130.8 219.6 ;
      RECT  134.4 218.4 135.6 219.6 ;
      RECT  139.2 218.4 140.4 219.6 ;
      RECT  144.0 218.4 145.2 219.6 ;
      RECT  148.8 218.4 150.0 219.6 ;
      RECT  153.6 218.4 154.8 219.6 ;
      RECT  158.4 218.4 159.6 219.6 ;
      RECT  163.2 218.4 164.4 219.6 ;
      RECT  168.0 218.4 169.2 219.6 ;
      RECT  172.8 218.4 174.0 219.6 ;
      RECT  177.6 218.4 178.8 219.6 ;
      RECT  33.6 223.2 34.8 224.4 ;
      RECT  38.4 223.2 39.6 224.4 ;
      RECT  43.2 223.2 44.4 224.4 ;
      RECT  48.0 223.2 49.2 224.4 ;
      RECT  52.8 223.2 54.0 224.4 ;
      RECT  57.6 223.2 58.8 224.4 ;
      RECT  62.4 223.2 63.6 224.4 ;
      RECT  67.2 223.2 68.4 224.4 ;
      RECT  72.0 223.2 73.2 224.4 ;
      RECT  76.8 223.2 78.0 224.4 ;
      RECT  81.6 223.2 82.8 224.4 ;
      RECT  86.4 223.2 87.6 224.4 ;
      RECT  91.2 223.2 92.4 224.4 ;
      RECT  96.0 223.2 97.2 224.4 ;
      RECT  100.8 223.2 102.0 224.4 ;
      RECT  105.6 223.2 106.8 224.4 ;
      RECT  110.4 223.2 111.6 224.4 ;
      RECT  115.2 223.2 116.4 224.4 ;
      RECT  120.0 223.2 121.2 224.4 ;
      RECT  139.2 223.2 140.4 224.4 ;
      RECT  144.0 223.2 145.2 224.4 ;
      RECT  148.8 223.2 150.0 224.4 ;
      RECT  153.6 223.2 154.8 224.4 ;
      RECT  158.4 223.2 159.6 224.4 ;
      RECT  163.2 223.2 164.4 224.4 ;
      RECT  168.0 223.2 169.2 224.4 ;
      RECT  172.8 223.2 174.0 224.4 ;
      RECT  177.6 223.2 178.8 224.4 ;
      RECT  182.4 223.2 183.6 224.4 ;
      RECT  187.2 223.2 188.4 224.4 ;
      RECT  192.0 223.2 193.2 224.4 ;
      RECT  196.8 223.2 198.0 224.4 ;
      RECT  201.6 223.2 202.8 224.4 ;
      RECT  206.4 223.2 207.6 224.4 ;
      RECT  211.2 223.2 212.4 224.4 ;
      RECT  216.0 223.2 217.2 224.4 ;
      RECT  220.8 223.2 222.0 224.4 ;
      RECT  225.6 223.2 226.8 224.4 ;
      RECT  24.0 228.0 25.2 229.2 ;
      RECT  28.8 228.0 30.0 229.2 ;
      RECT  33.6 228.0 34.8 229.2 ;
      RECT  38.4 228.0 39.6 229.2 ;
      RECT  43.2 228.0 44.4 229.2 ;
      RECT  48.0 228.0 49.2 229.2 ;
      RECT  52.8 228.0 54.0 229.2 ;
      RECT  57.6 228.0 58.8 229.2 ;
      RECT  62.4 228.0 63.6 229.2 ;
      RECT  67.2 228.0 68.4 229.2 ;
      RECT  72.0 228.0 73.2 229.2 ;
      RECT  76.8 228.0 78.0 229.2 ;
      RECT  81.6 228.0 82.8 229.2 ;
      RECT  86.4 228.0 87.6 229.2 ;
      RECT  91.2 228.0 92.4 229.2 ;
      RECT  96.0 228.0 97.2 229.2 ;
      RECT  100.8 228.0 102.0 229.2 ;
      RECT  105.6 228.0 106.8 229.2 ;
      RECT  110.4 228.0 111.6 229.2 ;
      RECT  115.2 228.0 116.4 229.2 ;
      RECT  120.0 228.0 121.2 229.2 ;
      RECT  124.8 228.0 126.0 229.2 ;
      RECT  129.6 228.0 130.8 229.2 ;
      RECT  134.4 228.0 135.6 229.2 ;
      RECT  139.2 228.0 140.4 229.2 ;
      RECT  144.0 228.0 145.2 229.2 ;
      RECT  148.8 228.0 150.0 229.2 ;
      RECT  153.6 228.0 154.8 229.2 ;
      RECT  158.4 228.0 159.6 229.2 ;
      RECT  163.2 228.0 164.4 229.2 ;
      RECT  168.0 228.0 169.2 229.2 ;
      RECT  172.8 228.0 174.0 229.2 ;
      RECT  177.6 228.0 178.8 229.2 ;
      RECT  33.6 232.8 34.8 234.0 ;
      RECT  38.4 232.8 39.6 234.0 ;
      RECT  43.2 232.8 44.4 234.0 ;
      RECT  48.0 232.8 49.2 234.0 ;
      RECT  52.8 232.8 54.0 234.0 ;
      RECT  57.6 232.8 58.8 234.0 ;
      RECT  62.4 232.8 63.6 234.0 ;
      RECT  67.2 232.8 68.4 234.0 ;
      RECT  72.0 232.8 73.2 234.0 ;
      RECT  76.8 232.8 78.0 234.0 ;
      RECT  81.6 232.8 82.8 234.0 ;
      RECT  86.4 232.8 87.6 234.0 ;
      RECT  91.2 232.8 92.4 234.0 ;
      RECT  96.0 232.8 97.2 234.0 ;
      RECT  100.8 232.8 102.0 234.0 ;
      RECT  105.6 232.8 106.8 234.0 ;
      RECT  110.4 232.8 111.6 234.0 ;
      RECT  115.2 232.8 116.4 234.0 ;
      RECT  120.0 232.8 121.2 234.0 ;
      RECT  124.8 232.8 126.0 234.0 ;
      RECT  129.6 232.8 130.8 234.0 ;
      RECT  134.4 232.8 135.6 234.0 ;
      RECT  139.2 232.8 140.4 234.0 ;
      RECT  144.0 232.8 145.2 234.0 ;
      RECT  148.8 232.8 150.0 234.0 ;
      RECT  153.6 232.8 154.8 234.0 ;
      RECT  158.4 232.8 159.6 234.0 ;
      RECT  163.2 232.8 164.4 234.0 ;
      RECT  168.0 232.8 169.2 234.0 ;
      RECT  172.8 232.8 174.0 234.0 ;
      RECT  177.6 232.8 178.8 234.0 ;
      RECT  182.4 232.8 183.6 234.0 ;
      RECT  187.2 232.8 188.4 234.0 ;
      RECT  192.0 232.8 193.2 234.0 ;
      RECT  196.8 232.8 198.0 234.0 ;
      RECT  201.6 232.8 202.8 234.0 ;
      RECT  206.4 232.8 207.6 234.0 ;
      RECT  211.2 232.8 212.4 234.0 ;
      RECT  216.0 232.8 217.2 234.0 ;
      RECT  220.8 232.8 222.0 234.0 ;
      RECT  225.6 232.8 226.8 234.0 ;
      RECT  4.8 237.6 6.0 238.8 ;
      RECT  9.6 237.6 10.8 238.8 ;
      RECT  14.4 237.6 15.6 238.8 ;
      RECT  19.2 237.6 20.4 238.8 ;
      RECT  24.0 237.6 25.2 238.8 ;
      RECT  28.8 237.6 30.0 238.8 ;
      RECT  33.6 237.6 34.8 238.8 ;
      RECT  38.4 237.6 39.6 238.8 ;
      RECT  43.2 237.6 44.4 238.8 ;
      RECT  48.0 237.6 49.2 238.8 ;
      RECT  52.8 237.6 54.0 238.8 ;
      RECT  57.6 237.6 58.8 238.8 ;
      RECT  62.4 237.6 63.6 238.8 ;
      RECT  67.2 237.6 68.4 238.8 ;
      RECT  72.0 237.6 73.2 238.8 ;
      RECT  76.8 237.6 78.0 238.8 ;
      RECT  81.6 237.6 82.8 238.8 ;
      RECT  86.4 237.6 87.6 238.8 ;
      RECT  91.2 237.6 92.4 238.8 ;
      RECT  96.0 237.6 97.2 238.8 ;
      RECT  177.6 237.6 178.8 238.8 ;
      RECT  182.4 237.6 183.6 238.8 ;
      RECT  187.2 237.6 188.4 238.8 ;
      RECT  192.0 237.6 193.2 238.8 ;
      RECT  196.8 237.6 198.0 238.8 ;
      RECT  201.6 237.6 202.8 238.8 ;
      RECT  206.4 237.6 207.6 238.8 ;
      RECT  211.2 237.6 212.4 238.8 ;
      RECT  216.0 237.6 217.2 238.8 ;
      RECT  220.8 237.6 222.0 238.8 ;
      RECT  225.6 237.6 226.8 238.8 ;
      RECT  33.6 242.4 34.8 243.6 ;
      RECT  38.4 242.4 39.6 243.6 ;
      RECT  43.2 242.4 44.4 243.6 ;
      RECT  48.0 242.4 49.2 243.6 ;
      RECT  52.8 242.4 54.0 243.6 ;
      RECT  57.6 242.4 58.8 243.6 ;
      RECT  62.4 242.4 63.6 243.6 ;
      RECT  67.2 242.4 68.4 243.6 ;
      RECT  72.0 242.4 73.2 243.6 ;
      RECT  76.8 242.4 78.0 243.6 ;
      RECT  81.6 242.4 82.8 243.6 ;
      RECT  86.4 242.4 87.6 243.6 ;
      RECT  91.2 242.4 92.4 243.6 ;
      RECT  96.0 242.4 97.2 243.6 ;
      RECT  100.8 242.4 102.0 243.6 ;
      RECT  105.6 242.4 106.8 243.6 ;
      RECT  110.4 242.4 111.6 243.6 ;
      RECT  115.2 242.4 116.4 243.6 ;
      RECT  120.0 242.4 121.2 243.6 ;
      RECT  124.8 242.4 126.0 243.6 ;
      RECT  129.6 242.4 130.8 243.6 ;
      RECT  134.4 242.4 135.6 243.6 ;
      RECT  139.2 242.4 140.4 243.6 ;
      RECT  144.0 242.4 145.2 243.6 ;
      RECT  148.8 242.4 150.0 243.6 ;
      RECT  153.6 242.4 154.8 243.6 ;
      RECT  158.4 242.4 159.6 243.6 ;
      RECT  163.2 242.4 164.4 243.6 ;
      RECT  168.0 242.4 169.2 243.6 ;
      RECT  172.8 242.4 174.0 243.6 ;
      RECT  177.6 242.4 178.8 243.6 ;
      RECT  24.0 247.2 25.2 248.4 ;
      RECT  28.8 247.2 30.0 248.4 ;
      RECT  33.6 247.2 34.8 248.4 ;
      RECT  38.4 247.2 39.6 248.4 ;
      RECT  43.2 247.2 44.4 248.4 ;
      RECT  48.0 247.2 49.2 248.4 ;
      RECT  52.8 247.2 54.0 248.4 ;
      RECT  57.6 247.2 58.8 248.4 ;
      RECT  62.4 247.2 63.6 248.4 ;
      RECT  67.2 247.2 68.4 248.4 ;
      RECT  72.0 247.2 73.2 248.4 ;
      RECT  76.8 247.2 78.0 248.4 ;
      RECT  81.6 247.2 82.8 248.4 ;
      RECT  86.4 247.2 87.6 248.4 ;
      RECT  144.0 247.2 145.2 248.4 ;
      RECT  148.8 247.2 150.0 248.4 ;
      RECT  153.6 247.2 154.8 248.4 ;
      RECT  158.4 247.2 159.6 248.4 ;
      RECT  163.2 247.2 164.4 248.4 ;
      RECT  168.0 247.2 169.2 248.4 ;
      RECT  172.8 247.2 174.0 248.4 ;
      RECT  177.6 247.2 178.8 248.4 ;
      RECT  182.4 247.2 183.6 248.4 ;
      RECT  187.2 247.2 188.4 248.4 ;
      RECT  192.0 247.2 193.2 248.4 ;
      RECT  196.8 247.2 198.0 248.4 ;
      RECT  201.6 247.2 202.8 248.4 ;
      RECT  206.4 247.2 207.6 248.4 ;
      RECT  211.2 247.2 212.4 248.4 ;
      RECT  216.0 247.2 217.2 248.4 ;
      RECT  220.8 247.2 222.0 248.4 ;
      RECT  225.6 247.2 226.8 248.4 ;
      RECT  33.6 252.0 34.8 253.2 ;
      RECT  38.4 252.0 39.6 253.2 ;
      RECT  43.2 252.0 44.4 253.2 ;
      RECT  48.0 252.0 49.2 253.2 ;
      RECT  52.8 252.0 54.0 253.2 ;
      RECT  57.6 252.0 58.8 253.2 ;
      RECT  62.4 252.0 63.6 253.2 ;
      RECT  67.2 252.0 68.4 253.2 ;
      RECT  72.0 252.0 73.2 253.2 ;
      RECT  76.8 252.0 78.0 253.2 ;
      RECT  81.6 252.0 82.8 253.2 ;
      RECT  86.4 252.0 87.6 253.2 ;
      RECT  91.2 252.0 92.4 253.2 ;
      RECT  96.0 252.0 97.2 253.2 ;
      RECT  100.8 252.0 102.0 253.2 ;
      RECT  105.6 252.0 106.8 253.2 ;
      RECT  110.4 252.0 111.6 253.2 ;
      RECT  115.2 252.0 116.4 253.2 ;
      RECT  120.0 252.0 121.2 253.2 ;
      RECT  124.8 252.0 126.0 253.2 ;
      RECT  129.6 252.0 130.8 253.2 ;
      RECT  134.4 252.0 135.6 253.2 ;
      RECT  139.2 252.0 140.4 253.2 ;
      RECT  144.0 252.0 145.2 253.2 ;
      RECT  148.8 252.0 150.0 253.2 ;
      RECT  153.6 252.0 154.8 253.2 ;
      RECT  158.4 252.0 159.6 253.2 ;
      RECT  163.2 252.0 164.4 253.2 ;
      RECT  168.0 252.0 169.2 253.2 ;
      RECT  172.8 252.0 174.0 253.2 ;
      RECT  177.6 252.0 178.8 253.2 ;
      RECT  4.8 256.8 6.0 258.0 ;
      RECT  9.6 256.8 10.8 258.0 ;
      RECT  14.4 256.8 15.6 258.0 ;
      RECT  19.2 256.8 20.4 258.0 ;
      RECT  24.0 256.8 25.2 258.0 ;
      RECT  28.8 256.8 30.0 258.0 ;
      RECT  33.6 256.8 34.8 258.0 ;
      RECT  38.4 256.8 39.6 258.0 ;
      RECT  43.2 256.8 44.4 258.0 ;
      RECT  48.0 256.8 49.2 258.0 ;
      RECT  52.8 256.8 54.0 258.0 ;
      RECT  57.6 256.8 58.8 258.0 ;
      RECT  62.4 256.8 63.6 258.0 ;
      RECT  67.2 256.8 68.4 258.0 ;
      RECT  72.0 256.8 73.2 258.0 ;
      RECT  76.8 256.8 78.0 258.0 ;
      RECT  81.6 256.8 82.8 258.0 ;
      RECT  86.4 256.8 87.6 258.0 ;
      RECT  177.6 256.8 178.8 258.0 ;
      RECT  182.4 256.8 183.6 258.0 ;
      RECT  187.2 256.8 188.4 258.0 ;
      RECT  192.0 256.8 193.2 258.0 ;
      RECT  196.8 256.8 198.0 258.0 ;
      RECT  201.6 256.8 202.8 258.0 ;
      RECT  206.4 256.8 207.6 258.0 ;
      RECT  211.2 256.8 212.4 258.0 ;
      RECT  216.0 256.8 217.2 258.0 ;
      RECT  220.8 256.8 222.0 258.0 ;
      RECT  225.6 256.8 226.8 258.0 ;
      RECT  4.8 261.6 6.0 262.8 ;
      RECT  9.6 261.6 10.8 262.8 ;
      RECT  14.4 261.6 15.6 262.8 ;
      RECT  19.2 261.6 20.4 262.8 ;
      RECT  24.0 261.6 25.2 262.8 ;
      RECT  28.8 261.6 30.0 262.8 ;
      RECT  33.6 261.6 34.8 262.8 ;
      RECT  38.4 261.6 39.6 262.8 ;
      RECT  43.2 261.6 44.4 262.8 ;
      RECT  48.0 261.6 49.2 262.8 ;
      RECT  52.8 261.6 54.0 262.8 ;
      RECT  57.6 261.6 58.8 262.8 ;
      RECT  62.4 261.6 63.6 262.8 ;
      RECT  67.2 261.6 68.4 262.8 ;
      RECT  72.0 261.6 73.2 262.8 ;
      RECT  76.8 261.6 78.0 262.8 ;
      RECT  81.6 261.6 82.8 262.8 ;
      RECT  86.4 261.6 87.6 262.8 ;
      RECT  91.2 261.6 92.4 262.8 ;
      RECT  96.0 261.6 97.2 262.8 ;
      RECT  100.8 261.6 102.0 262.8 ;
      RECT  105.6 261.6 106.8 262.8 ;
      RECT  110.4 261.6 111.6 262.8 ;
      RECT  115.2 261.6 116.4 262.8 ;
      RECT  120.0 261.6 121.2 262.8 ;
      RECT  124.8 261.6 126.0 262.8 ;
      RECT  129.6 261.6 130.8 262.8 ;
      RECT  134.4 261.6 135.6 262.8 ;
      RECT  139.2 261.6 140.4 262.8 ;
      RECT  144.0 261.6 145.2 262.8 ;
      RECT  148.8 261.6 150.0 262.8 ;
      RECT  153.6 261.6 154.8 262.8 ;
      RECT  158.4 261.6 159.6 262.8 ;
      RECT  163.2 261.6 164.4 262.8 ;
      RECT  168.0 261.6 169.2 262.8 ;
      RECT  172.8 261.6 174.0 262.8 ;
      RECT  177.6 261.6 178.8 262.8 ;
      RECT  4.8 266.4 6.0 267.6 ;
      RECT  9.6 266.4 10.8 267.6 ;
      RECT  14.4 266.4 15.6 267.6 ;
      RECT  19.2 266.4 20.4 267.6 ;
      RECT  24.0 266.4 25.2 267.6 ;
      RECT  28.8 266.4 30.0 267.6 ;
      RECT  33.6 266.4 34.8 267.6 ;
      RECT  38.4 266.4 39.6 267.6 ;
      RECT  43.2 266.4 44.4 267.6 ;
      RECT  48.0 266.4 49.2 267.6 ;
      RECT  52.8 266.4 54.0 267.6 ;
      RECT  57.6 266.4 58.8 267.6 ;
      RECT  62.4 266.4 63.6 267.6 ;
      RECT  67.2 266.4 68.4 267.6 ;
      RECT  72.0 266.4 73.2 267.6 ;
      RECT  76.8 266.4 78.0 267.6 ;
      RECT  81.6 266.4 82.8 267.6 ;
      RECT  86.4 266.4 87.6 267.6 ;
      RECT  91.2 266.4 92.4 267.6 ;
      RECT  96.0 266.4 97.2 267.6 ;
      RECT  100.8 266.4 102.0 267.6 ;
      RECT  105.6 266.4 106.8 267.6 ;
      RECT  110.4 266.4 111.6 267.6 ;
      RECT  115.2 266.4 116.4 267.6 ;
      RECT  120.0 266.4 121.2 267.6 ;
      RECT  144.0 266.4 145.2 267.6 ;
      RECT  148.8 266.4 150.0 267.6 ;
      RECT  153.6 266.4 154.8 267.6 ;
      RECT  158.4 266.4 159.6 267.6 ;
      RECT  163.2 266.4 164.4 267.6 ;
      RECT  168.0 266.4 169.2 267.6 ;
      RECT  172.8 266.4 174.0 267.6 ;
      RECT  177.6 266.4 178.8 267.6 ;
      RECT  182.4 266.4 183.6 267.6 ;
      RECT  187.2 266.4 188.4 267.6 ;
      RECT  192.0 266.4 193.2 267.6 ;
      RECT  196.8 266.4 198.0 267.6 ;
      RECT  201.6 266.4 202.8 267.6 ;
      RECT  206.4 266.4 207.6 267.6 ;
      RECT  211.2 266.4 212.4 267.6 ;
      RECT  216.0 266.4 217.2 267.6 ;
      RECT  220.8 266.4 222.0 267.6 ;
      RECT  225.6 266.4 226.8 267.6 ;
      RECT  4.8 271.2 6.0 272.4 ;
      RECT  9.6 271.2 10.8 272.4 ;
      RECT  14.4 271.2 15.6 272.4 ;
      RECT  19.2 271.2 20.4 272.4 ;
      RECT  24.0 271.2 25.2 272.4 ;
      RECT  28.8 271.2 30.0 272.4 ;
      RECT  33.6 271.2 34.8 272.4 ;
      RECT  38.4 271.2 39.6 272.4 ;
      RECT  43.2 271.2 44.4 272.4 ;
      RECT  48.0 271.2 49.2 272.4 ;
      RECT  52.8 271.2 54.0 272.4 ;
      RECT  57.6 271.2 58.8 272.4 ;
      RECT  62.4 271.2 63.6 272.4 ;
      RECT  67.2 271.2 68.4 272.4 ;
      RECT  72.0 271.2 73.2 272.4 ;
      RECT  76.8 271.2 78.0 272.4 ;
      RECT  81.6 271.2 82.8 272.4 ;
      RECT  86.4 271.2 87.6 272.4 ;
      RECT  91.2 271.2 92.4 272.4 ;
      RECT  96.0 271.2 97.2 272.4 ;
      RECT  100.8 271.2 102.0 272.4 ;
      RECT  105.6 271.2 106.8 272.4 ;
      RECT  110.4 271.2 111.6 272.4 ;
      RECT  115.2 271.2 116.4 272.4 ;
      RECT  120.0 271.2 121.2 272.4 ;
      RECT  124.8 271.2 126.0 272.4 ;
      RECT  129.6 271.2 130.8 272.4 ;
      RECT  134.4 271.2 135.6 272.4 ;
      RECT  139.2 271.2 140.4 272.4 ;
      RECT  144.0 271.2 145.2 272.4 ;
      RECT  148.8 271.2 150.0 272.4 ;
      RECT  153.6 271.2 154.8 272.4 ;
      RECT  158.4 271.2 159.6 272.4 ;
      RECT  163.2 271.2 164.4 272.4 ;
      RECT  168.0 271.2 169.2 272.4 ;
      RECT  172.8 271.2 174.0 272.4 ;
      RECT  177.6 271.2 178.8 272.4 ;
      RECT  4.8 276.0 6.0 277.2 ;
      RECT  9.6 276.0 10.8 277.2 ;
      RECT  14.4 276.0 15.6 277.2 ;
      RECT  19.2 276.0 20.4 277.2 ;
      RECT  24.0 276.0 25.2 277.2 ;
      RECT  28.8 276.0 30.0 277.2 ;
      RECT  33.6 276.0 34.8 277.2 ;
      RECT  38.4 276.0 39.6 277.2 ;
      RECT  43.2 276.0 44.4 277.2 ;
      RECT  48.0 276.0 49.2 277.2 ;
      RECT  52.8 276.0 54.0 277.2 ;
      RECT  57.6 276.0 58.8 277.2 ;
      RECT  62.4 276.0 63.6 277.2 ;
      RECT  67.2 276.0 68.4 277.2 ;
      RECT  72.0 276.0 73.2 277.2 ;
      RECT  76.8 276.0 78.0 277.2 ;
      RECT  81.6 276.0 82.8 277.2 ;
      RECT  86.4 276.0 87.6 277.2 ;
      RECT  91.2 276.0 92.4 277.2 ;
      RECT  96.0 276.0 97.2 277.2 ;
      RECT  177.6 276.0 178.8 277.2 ;
      RECT  182.4 276.0 183.6 277.2 ;
      RECT  187.2 276.0 188.4 277.2 ;
      RECT  192.0 276.0 193.2 277.2 ;
      RECT  196.8 276.0 198.0 277.2 ;
      RECT  201.6 276.0 202.8 277.2 ;
      RECT  206.4 276.0 207.6 277.2 ;
      RECT  211.2 276.0 212.4 277.2 ;
      RECT  216.0 276.0 217.2 277.2 ;
      RECT  220.8 276.0 222.0 277.2 ;
      RECT  225.6 276.0 226.8 277.2 ;
      RECT  4.8 280.8 6.0 282.0 ;
      RECT  9.6 280.8 10.8 282.0 ;
      RECT  14.4 280.8 15.6 282.0 ;
      RECT  19.2 280.8 20.4 282.0 ;
      RECT  24.0 280.8 25.2 282.0 ;
      RECT  28.8 280.8 30.0 282.0 ;
      RECT  33.6 280.8 34.8 282.0 ;
      RECT  38.4 280.8 39.6 282.0 ;
      RECT  43.2 280.8 44.4 282.0 ;
      RECT  48.0 280.8 49.2 282.0 ;
      RECT  52.8 280.8 54.0 282.0 ;
      RECT  57.6 280.8 58.8 282.0 ;
      RECT  62.4 280.8 63.6 282.0 ;
      RECT  67.2 280.8 68.4 282.0 ;
      RECT  72.0 280.8 73.2 282.0 ;
      RECT  76.8 280.8 78.0 282.0 ;
      RECT  81.6 280.8 82.8 282.0 ;
      RECT  86.4 280.8 87.6 282.0 ;
      RECT  91.2 280.8 92.4 282.0 ;
      RECT  96.0 280.8 97.2 282.0 ;
      RECT  100.8 280.8 102.0 282.0 ;
      RECT  105.6 280.8 106.8 282.0 ;
      RECT  110.4 280.8 111.6 282.0 ;
      RECT  115.2 280.8 116.4 282.0 ;
      RECT  120.0 280.8 121.2 282.0 ;
      RECT  124.8 280.8 126.0 282.0 ;
      RECT  129.6 280.8 130.8 282.0 ;
      RECT  134.4 280.8 135.6 282.0 ;
      RECT  139.2 280.8 140.4 282.0 ;
      RECT  144.0 280.8 145.2 282.0 ;
      RECT  148.8 280.8 150.0 282.0 ;
      RECT  153.6 280.8 154.8 282.0 ;
      RECT  158.4 280.8 159.6 282.0 ;
      RECT  163.2 280.8 164.4 282.0 ;
      RECT  168.0 280.8 169.2 282.0 ;
      RECT  172.8 280.8 174.0 282.0 ;
      RECT  177.6 280.8 178.8 282.0 ;
      RECT  4.8 285.6 6.0 286.8 ;
      RECT  9.6 285.6 10.8 286.8 ;
      RECT  14.4 285.6 15.6 286.8 ;
      RECT  19.2 285.6 20.4 286.8 ;
      RECT  24.0 285.6 25.2 286.8 ;
      RECT  28.8 285.6 30.0 286.8 ;
      RECT  33.6 285.6 34.8 286.8 ;
      RECT  38.4 285.6 39.6 286.8 ;
      RECT  43.2 285.6 44.4 286.8 ;
      RECT  48.0 285.6 49.2 286.8 ;
      RECT  52.8 285.6 54.0 286.8 ;
      RECT  57.6 285.6 58.8 286.8 ;
      RECT  62.4 285.6 63.6 286.8 ;
      RECT  67.2 285.6 68.4 286.8 ;
      RECT  72.0 285.6 73.2 286.8 ;
      RECT  76.8 285.6 78.0 286.8 ;
      RECT  81.6 285.6 82.8 286.8 ;
      RECT  86.4 285.6 87.6 286.8 ;
      RECT  91.2 285.6 92.4 286.8 ;
      RECT  96.0 285.6 97.2 286.8 ;
      RECT  100.8 285.6 102.0 286.8 ;
      RECT  105.6 285.6 106.8 286.8 ;
      RECT  110.4 285.6 111.6 286.8 ;
      RECT  115.2 285.6 116.4 286.8 ;
      RECT  120.0 285.6 121.2 286.8 ;
      RECT  124.8 285.6 126.0 286.8 ;
      RECT  129.6 285.6 130.8 286.8 ;
      RECT  134.4 285.6 135.6 286.8 ;
      RECT  139.2 285.6 140.4 286.8 ;
      RECT  144.0 285.6 145.2 286.8 ;
      RECT  148.8 285.6 150.0 286.8 ;
      RECT  153.6 285.6 154.8 286.8 ;
      RECT  158.4 285.6 159.6 286.8 ;
      RECT  163.2 285.6 164.4 286.8 ;
      RECT  168.0 285.6 169.2 286.8 ;
      RECT  172.8 285.6 174.0 286.8 ;
      RECT  177.6 285.6 178.8 286.8 ;
      RECT  182.4 285.6 183.6 286.8 ;
      RECT  187.2 285.6 188.4 286.8 ;
      RECT  192.0 285.6 193.2 286.8 ;
      RECT  196.8 285.6 198.0 286.8 ;
      RECT  201.6 285.6 202.8 286.8 ;
      RECT  206.4 285.6 207.6 286.8 ;
      RECT  211.2 285.6 212.4 286.8 ;
      RECT  216.0 285.6 217.2 286.8 ;
      RECT  220.8 285.6 222.0 286.8 ;
      RECT  225.6 285.6 226.8 286.8 ;
      RECT  4.8 290.4 6.0 291.6 ;
      RECT  9.6 290.4 10.8 291.6 ;
      RECT  14.4 290.4 15.6 291.6 ;
      RECT  19.2 290.4 20.4 291.6 ;
      RECT  24.0 290.4 25.2 291.6 ;
      RECT  28.8 290.4 30.0 291.6 ;
      RECT  33.6 290.4 34.8 291.6 ;
      RECT  38.4 290.4 39.6 291.6 ;
      RECT  43.2 290.4 44.4 291.6 ;
      RECT  48.0 290.4 49.2 291.6 ;
      RECT  52.8 290.4 54.0 291.6 ;
      RECT  57.6 290.4 58.8 291.6 ;
      RECT  62.4 290.4 63.6 291.6 ;
      RECT  67.2 290.4 68.4 291.6 ;
      RECT  81.6 290.4 82.8 291.6 ;
      RECT  86.4 290.4 87.6 291.6 ;
      RECT  91.2 290.4 92.4 291.6 ;
      RECT  96.0 290.4 97.2 291.6 ;
      RECT  100.8 290.4 102.0 291.6 ;
      RECT  105.6 290.4 106.8 291.6 ;
      RECT  110.4 290.4 111.6 291.6 ;
      RECT  115.2 290.4 116.4 291.6 ;
      RECT  120.0 290.4 121.2 291.6 ;
      RECT  124.8 290.4 126.0 291.6 ;
      RECT  129.6 290.4 130.8 291.6 ;
      RECT  134.4 290.4 135.6 291.6 ;
      RECT  139.2 290.4 140.4 291.6 ;
      RECT  144.0 290.4 145.2 291.6 ;
      RECT  148.8 290.4 150.0 291.6 ;
      RECT  153.6 290.4 154.8 291.6 ;
      RECT  158.4 290.4 159.6 291.6 ;
      RECT  163.2 290.4 164.4 291.6 ;
      RECT  168.0 290.4 169.2 291.6 ;
      RECT  172.8 290.4 174.0 291.6 ;
      RECT  177.6 290.4 178.8 291.6 ;
      RECT  4.8 295.2 6.0 296.4 ;
      RECT  9.6 295.2 10.8 296.4 ;
      RECT  14.4 295.2 15.6 296.4 ;
      RECT  19.2 295.2 20.4 296.4 ;
      RECT  24.0 295.2 25.2 296.4 ;
      RECT  28.8 295.2 30.0 296.4 ;
      RECT  33.6 295.2 34.8 296.4 ;
      RECT  38.4 295.2 39.6 296.4 ;
      RECT  43.2 295.2 44.4 296.4 ;
      RECT  48.0 295.2 49.2 296.4 ;
      RECT  52.8 295.2 54.0 296.4 ;
      RECT  57.6 295.2 58.8 296.4 ;
      RECT  62.4 295.2 63.6 296.4 ;
      RECT  67.2 295.2 68.4 296.4 ;
      RECT  72.0 295.2 73.2 296.4 ;
      RECT  76.8 295.2 78.0 296.4 ;
      RECT  81.6 295.2 82.8 296.4 ;
      RECT  86.4 295.2 87.6 296.4 ;
      RECT  91.2 295.2 92.4 296.4 ;
      RECT  96.0 295.2 97.2 296.4 ;
      RECT  100.8 295.2 102.0 296.4 ;
      RECT  105.6 295.2 106.8 296.4 ;
      RECT  110.4 295.2 111.6 296.4 ;
      RECT  115.2 295.2 116.4 296.4 ;
      RECT  120.0 295.2 121.2 296.4 ;
      RECT  124.8 295.2 126.0 296.4 ;
      RECT  129.6 295.2 130.8 296.4 ;
      RECT  134.4 295.2 135.6 296.4 ;
      RECT  139.2 295.2 140.4 296.4 ;
      RECT  144.0 295.2 145.2 296.4 ;
      RECT  148.8 295.2 150.0 296.4 ;
      RECT  153.6 295.2 154.8 296.4 ;
      RECT  158.4 295.2 159.6 296.4 ;
      RECT  163.2 295.2 164.4 296.4 ;
      RECT  168.0 295.2 169.2 296.4 ;
      RECT  172.8 295.2 174.0 296.4 ;
      RECT  177.6 295.2 178.8 296.4 ;
      RECT  182.4 295.2 183.6 296.4 ;
      RECT  187.2 295.2 188.4 296.4 ;
      RECT  192.0 295.2 193.2 296.4 ;
      RECT  196.8 295.2 198.0 296.4 ;
      RECT  201.6 295.2 202.8 296.4 ;
      RECT  206.4 295.2 207.6 296.4 ;
      RECT  211.2 295.2 212.4 296.4 ;
      RECT  216.0 295.2 217.2 296.4 ;
      RECT  220.8 295.2 222.0 296.4 ;
      RECT  225.6 295.2 226.8 296.4 ;
      RECT  4.8 300.0 6.0 301.2 ;
      RECT  9.6 300.0 10.8 301.2 ;
      RECT  14.4 300.0 15.6 301.2 ;
      RECT  19.2 300.0 20.4 301.2 ;
      RECT  24.0 300.0 25.2 301.2 ;
      RECT  28.8 300.0 30.0 301.2 ;
      RECT  33.6 300.0 34.8 301.2 ;
      RECT  38.4 300.0 39.6 301.2 ;
      RECT  43.2 300.0 44.4 301.2 ;
      RECT  48.0 300.0 49.2 301.2 ;
      RECT  52.8 300.0 54.0 301.2 ;
      RECT  57.6 300.0 58.8 301.2 ;
      RECT  62.4 300.0 63.6 301.2 ;
      RECT  67.2 300.0 68.4 301.2 ;
      RECT  72.0 300.0 73.2 301.2 ;
      RECT  76.8 300.0 78.0 301.2 ;
      RECT  81.6 300.0 82.8 301.2 ;
      RECT  86.4 300.0 87.6 301.2 ;
      RECT  91.2 300.0 92.4 301.2 ;
      RECT  96.0 300.0 97.2 301.2 ;
      RECT  100.8 300.0 102.0 301.2 ;
      RECT  105.6 300.0 106.8 301.2 ;
      RECT  110.4 300.0 111.6 301.2 ;
      RECT  115.2 300.0 116.4 301.2 ;
      RECT  120.0 300.0 121.2 301.2 ;
      RECT  124.8 300.0 126.0 301.2 ;
      RECT  129.6 300.0 130.8 301.2 ;
      RECT  134.4 300.0 135.6 301.2 ;
      RECT  139.2 300.0 140.4 301.2 ;
      RECT  177.6 300.0 178.8 301.2 ;
      RECT  182.4 300.0 183.6 301.2 ;
      RECT  187.2 300.0 188.4 301.2 ;
      RECT  192.0 300.0 193.2 301.2 ;
      RECT  196.8 300.0 198.0 301.2 ;
      RECT  201.6 300.0 202.8 301.2 ;
      RECT  206.4 300.0 207.6 301.2 ;
      RECT  211.2 300.0 212.4 301.2 ;
      RECT  216.0 300.0 217.2 301.2 ;
      RECT  220.8 300.0 222.0 301.2 ;
      RECT  225.6 300.0 226.8 301.2 ;
      RECT  4.8 304.8 6.0 306.0 ;
      RECT  9.6 304.8 10.8 306.0 ;
      RECT  14.4 304.8 15.6 306.0 ;
      RECT  19.2 304.8 20.4 306.0 ;
      RECT  24.0 304.8 25.2 306.0 ;
      RECT  28.8 304.8 30.0 306.0 ;
      RECT  33.6 304.8 34.8 306.0 ;
      RECT  38.4 304.8 39.6 306.0 ;
      RECT  43.2 304.8 44.4 306.0 ;
      RECT  48.0 304.8 49.2 306.0 ;
      RECT  52.8 304.8 54.0 306.0 ;
      RECT  57.6 304.8 58.8 306.0 ;
      RECT  62.4 304.8 63.6 306.0 ;
      RECT  67.2 304.8 68.4 306.0 ;
      RECT  72.0 304.8 73.2 306.0 ;
      RECT  76.8 304.8 78.0 306.0 ;
      RECT  81.6 304.8 82.8 306.0 ;
      RECT  86.4 304.8 87.6 306.0 ;
      RECT  91.2 304.8 92.4 306.0 ;
      RECT  96.0 304.8 97.2 306.0 ;
      RECT  100.8 304.8 102.0 306.0 ;
      RECT  105.6 304.8 106.8 306.0 ;
      RECT  110.4 304.8 111.6 306.0 ;
      RECT  115.2 304.8 116.4 306.0 ;
      RECT  120.0 304.8 121.2 306.0 ;
      RECT  124.8 304.8 126.0 306.0 ;
      RECT  129.6 304.8 130.8 306.0 ;
      RECT  134.4 304.8 135.6 306.0 ;
      RECT  139.2 304.8 140.4 306.0 ;
      RECT  144.0 304.8 145.2 306.0 ;
      RECT  148.8 304.8 150.0 306.0 ;
      RECT  153.6 304.8 154.8 306.0 ;
      RECT  158.4 304.8 159.6 306.0 ;
      RECT  163.2 304.8 164.4 306.0 ;
      RECT  168.0 304.8 169.2 306.0 ;
      RECT  172.8 304.8 174.0 306.0 ;
      RECT  177.6 304.8 178.8 306.0 ;
      RECT  4.8 309.6 6.0 310.8 ;
      RECT  9.6 309.6 10.8 310.8 ;
      RECT  14.4 309.6 15.6 310.8 ;
      RECT  19.2 309.6 20.4 310.8 ;
      RECT  24.0 309.6 25.2 310.8 ;
      RECT  28.8 309.6 30.0 310.8 ;
      RECT  33.6 309.6 34.8 310.8 ;
      RECT  38.4 309.6 39.6 310.8 ;
      RECT  43.2 309.6 44.4 310.8 ;
      RECT  48.0 309.6 49.2 310.8 ;
      RECT  52.8 309.6 54.0 310.8 ;
      RECT  57.6 309.6 58.8 310.8 ;
      RECT  62.4 309.6 63.6 310.8 ;
      RECT  67.2 309.6 68.4 310.8 ;
      RECT  72.0 309.6 73.2 310.8 ;
      RECT  76.8 309.6 78.0 310.8 ;
      RECT  81.6 309.6 82.8 310.8 ;
      RECT  86.4 309.6 87.6 310.8 ;
      RECT  91.2 309.6 92.4 310.8 ;
      RECT  96.0 309.6 97.2 310.8 ;
      RECT  100.8 309.6 102.0 310.8 ;
      RECT  105.6 309.6 106.8 310.8 ;
      RECT  110.4 309.6 111.6 310.8 ;
      RECT  115.2 309.6 116.4 310.8 ;
      RECT  120.0 309.6 121.2 310.8 ;
      RECT  124.8 309.6 126.0 310.8 ;
      RECT  129.6 309.6 130.8 310.8 ;
      RECT  134.4 309.6 135.6 310.8 ;
      RECT  139.2 309.6 140.4 310.8 ;
      RECT  144.0 309.6 145.2 310.8 ;
      RECT  148.8 309.6 150.0 310.8 ;
      RECT  153.6 309.6 154.8 310.8 ;
      RECT  158.4 309.6 159.6 310.8 ;
      RECT  163.2 309.6 164.4 310.8 ;
      RECT  168.0 309.6 169.2 310.8 ;
      RECT  172.8 309.6 174.0 310.8 ;
      RECT  177.6 309.6 178.8 310.8 ;
      RECT  182.4 309.6 183.6 310.8 ;
      RECT  187.2 309.6 188.4 310.8 ;
      RECT  192.0 309.6 193.2 310.8 ;
      RECT  196.8 309.6 198.0 310.8 ;
      RECT  201.6 309.6 202.8 310.8 ;
      RECT  206.4 309.6 207.6 310.8 ;
      RECT  211.2 309.6 212.4 310.8 ;
      RECT  216.0 309.6 217.2 310.8 ;
      RECT  220.8 309.6 222.0 310.8 ;
      RECT  225.6 309.6 226.8 310.8 ;
      RECT  4.8 314.4 6.0 315.6 ;
      RECT  9.6 314.4 10.8 315.6 ;
      RECT  14.4 314.4 15.6 315.6 ;
      RECT  19.2 314.4 20.4 315.6 ;
      RECT  24.0 314.4 25.2 315.6 ;
      RECT  28.8 314.4 30.0 315.6 ;
      RECT  33.6 314.4 34.8 315.6 ;
      RECT  38.4 314.4 39.6 315.6 ;
      RECT  43.2 314.4 44.4 315.6 ;
      RECT  48.0 314.4 49.2 315.6 ;
      RECT  52.8 314.4 54.0 315.6 ;
      RECT  57.6 314.4 58.8 315.6 ;
      RECT  62.4 314.4 63.6 315.6 ;
      RECT  67.2 314.4 68.4 315.6 ;
      RECT  72.0 314.4 73.2 315.6 ;
      RECT  76.8 314.4 78.0 315.6 ;
      RECT  81.6 314.4 82.8 315.6 ;
      RECT  86.4 314.4 87.6 315.6 ;
      RECT  91.2 314.4 92.4 315.6 ;
      RECT  96.0 314.4 97.2 315.6 ;
      RECT  100.8 314.4 102.0 315.6 ;
      RECT  105.6 314.4 106.8 315.6 ;
      RECT  110.4 314.4 111.6 315.6 ;
      RECT  115.2 314.4 116.4 315.6 ;
      RECT  120.0 314.4 121.2 315.6 ;
      RECT  124.8 314.4 126.0 315.6 ;
      RECT  129.6 314.4 130.8 315.6 ;
      RECT  134.4 314.4 135.6 315.6 ;
      RECT  139.2 314.4 140.4 315.6 ;
      RECT  144.0 314.4 145.2 315.6 ;
      RECT  148.8 314.4 150.0 315.6 ;
      RECT  153.6 314.4 154.8 315.6 ;
      RECT  158.4 314.4 159.6 315.6 ;
      RECT  163.2 314.4 164.4 315.6 ;
      RECT  168.0 314.4 169.2 315.6 ;
      RECT  172.8 314.4 174.0 315.6 ;
      RECT  177.6 314.4 178.8 315.6 ;
      RECT  4.8 319.2 6.0 320.4 ;
      RECT  9.6 319.2 10.8 320.4 ;
      RECT  14.4 319.2 15.6 320.4 ;
      RECT  19.2 319.2 20.4 320.4 ;
      RECT  24.0 319.2 25.2 320.4 ;
      RECT  28.8 319.2 30.0 320.4 ;
      RECT  33.6 319.2 34.8 320.4 ;
      RECT  38.4 319.2 39.6 320.4 ;
      RECT  43.2 319.2 44.4 320.4 ;
      RECT  48.0 319.2 49.2 320.4 ;
      RECT  52.8 319.2 54.0 320.4 ;
      RECT  57.6 319.2 58.8 320.4 ;
      RECT  62.4 319.2 63.6 320.4 ;
      RECT  67.2 319.2 68.4 320.4 ;
      RECT  72.0 319.2 73.2 320.4 ;
      RECT  76.8 319.2 78.0 320.4 ;
      RECT  81.6 319.2 82.8 320.4 ;
      RECT  86.4 319.2 87.6 320.4 ;
      RECT  91.2 319.2 92.4 320.4 ;
      RECT  96.0 319.2 97.2 320.4 ;
      RECT  100.8 319.2 102.0 320.4 ;
      RECT  105.6 319.2 106.8 320.4 ;
      RECT  110.4 319.2 111.6 320.4 ;
      RECT  115.2 319.2 116.4 320.4 ;
      RECT  120.0 319.2 121.2 320.4 ;
      RECT  124.8 319.2 126.0 320.4 ;
      RECT  129.6 319.2 130.8 320.4 ;
      RECT  134.4 319.2 135.6 320.4 ;
      RECT  139.2 319.2 140.4 320.4 ;
      RECT  177.6 319.2 178.8 320.4 ;
      RECT  182.4 319.2 183.6 320.4 ;
      RECT  187.2 319.2 188.4 320.4 ;
      RECT  192.0 319.2 193.2 320.4 ;
      RECT  196.8 319.2 198.0 320.4 ;
      RECT  201.6 319.2 202.8 320.4 ;
      RECT  206.4 319.2 207.6 320.4 ;
      RECT  211.2 319.2 212.4 320.4 ;
      RECT  216.0 319.2 217.2 320.4 ;
      RECT  220.8 319.2 222.0 320.4 ;
      RECT  225.6 319.2 226.8 320.4 ;
      RECT  4.8 324.0 6.0 325.2 ;
      RECT  9.6 324.0 10.8 325.2 ;
      RECT  14.4 324.0 15.6 325.2 ;
      RECT  19.2 324.0 20.4 325.2 ;
      RECT  24.0 324.0 25.2 325.2 ;
      RECT  28.8 324.0 30.0 325.2 ;
      RECT  33.6 324.0 34.8 325.2 ;
      RECT  38.4 324.0 39.6 325.2 ;
      RECT  43.2 324.0 44.4 325.2 ;
      RECT  48.0 324.0 49.2 325.2 ;
      RECT  52.8 324.0 54.0 325.2 ;
      RECT  57.6 324.0 58.8 325.2 ;
      RECT  62.4 324.0 63.6 325.2 ;
      RECT  67.2 324.0 68.4 325.2 ;
      RECT  72.0 324.0 73.2 325.2 ;
      RECT  76.8 324.0 78.0 325.2 ;
      RECT  96.0 324.0 97.2 325.2 ;
      RECT  100.8 324.0 102.0 325.2 ;
      RECT  105.6 324.0 106.8 325.2 ;
      RECT  110.4 324.0 111.6 325.2 ;
      RECT  115.2 324.0 116.4 325.2 ;
      RECT  120.0 324.0 121.2 325.2 ;
      RECT  124.8 324.0 126.0 325.2 ;
      RECT  129.6 324.0 130.8 325.2 ;
      RECT  134.4 324.0 135.6 325.2 ;
      RECT  139.2 324.0 140.4 325.2 ;
      RECT  144.0 324.0 145.2 325.2 ;
      RECT  148.8 324.0 150.0 325.2 ;
      RECT  153.6 324.0 154.8 325.2 ;
      RECT  158.4 324.0 159.6 325.2 ;
      RECT  163.2 324.0 164.4 325.2 ;
      RECT  168.0 324.0 169.2 325.2 ;
      RECT  172.8 324.0 174.0 325.2 ;
      RECT  177.6 324.0 178.8 325.2 ;
      RECT  4.8 328.8 6.0 330.0 ;
      RECT  9.6 328.8 10.8 330.0 ;
      RECT  14.4 328.8 15.6 330.0 ;
      RECT  19.2 328.8 20.4 330.0 ;
      RECT  24.0 328.8 25.2 330.0 ;
      RECT  28.8 328.8 30.0 330.0 ;
      RECT  33.6 328.8 34.8 330.0 ;
      RECT  38.4 328.8 39.6 330.0 ;
      RECT  43.2 328.8 44.4 330.0 ;
      RECT  48.0 328.8 49.2 330.0 ;
      RECT  52.8 328.8 54.0 330.0 ;
      RECT  57.6 328.8 58.8 330.0 ;
      RECT  62.4 328.8 63.6 330.0 ;
      RECT  67.2 328.8 68.4 330.0 ;
      RECT  72.0 328.8 73.2 330.0 ;
      RECT  76.8 328.8 78.0 330.0 ;
      RECT  81.6 328.8 82.8 330.0 ;
      RECT  86.4 328.8 87.6 330.0 ;
      RECT  91.2 328.8 92.4 330.0 ;
      RECT  96.0 328.8 97.2 330.0 ;
      RECT  100.8 328.8 102.0 330.0 ;
      RECT  105.6 328.8 106.8 330.0 ;
      RECT  110.4 328.8 111.6 330.0 ;
      RECT  115.2 328.8 116.4 330.0 ;
      RECT  120.0 328.8 121.2 330.0 ;
      RECT  124.8 328.8 126.0 330.0 ;
      RECT  129.6 328.8 130.8 330.0 ;
      RECT  134.4 328.8 135.6 330.0 ;
      RECT  139.2 328.8 140.4 330.0 ;
      RECT  144.0 328.8 145.2 330.0 ;
      RECT  148.8 328.8 150.0 330.0 ;
      RECT  153.6 328.8 154.8 330.0 ;
      RECT  158.4 328.8 159.6 330.0 ;
      RECT  163.2 328.8 164.4 330.0 ;
      RECT  168.0 328.8 169.2 330.0 ;
      RECT  172.8 328.8 174.0 330.0 ;
      RECT  177.6 328.8 178.8 330.0 ;
      RECT  182.4 328.8 183.6 330.0 ;
      RECT  187.2 328.8 188.4 330.0 ;
      RECT  192.0 328.8 193.2 330.0 ;
      RECT  196.8 328.8 198.0 330.0 ;
      RECT  201.6 328.8 202.8 330.0 ;
      RECT  206.4 328.8 207.6 330.0 ;
      RECT  211.2 328.8 212.4 330.0 ;
      RECT  216.0 328.8 217.2 330.0 ;
      RECT  220.8 328.8 222.0 330.0 ;
      RECT  225.6 328.8 226.8 330.0 ;
      RECT  4.8 333.6 6.0 334.8 ;
      RECT  9.6 333.6 10.8 334.8 ;
      RECT  14.4 333.6 15.6 334.8 ;
      RECT  19.2 333.6 20.4 334.8 ;
      RECT  24.0 333.6 25.2 334.8 ;
      RECT  28.8 333.6 30.0 334.8 ;
      RECT  33.6 333.6 34.8 334.8 ;
      RECT  38.4 333.6 39.6 334.8 ;
      RECT  43.2 333.6 44.4 334.8 ;
      RECT  48.0 333.6 49.2 334.8 ;
      RECT  52.8 333.6 54.0 334.8 ;
      RECT  57.6 333.6 58.8 334.8 ;
      RECT  62.4 333.6 63.6 334.8 ;
      RECT  67.2 333.6 68.4 334.8 ;
      RECT  81.6 333.6 82.8 334.8 ;
      RECT  86.4 333.6 87.6 334.8 ;
      RECT  91.2 333.6 92.4 334.8 ;
      RECT  96.0 333.6 97.2 334.8 ;
      RECT  100.8 333.6 102.0 334.8 ;
      RECT  105.6 333.6 106.8 334.8 ;
      RECT  110.4 333.6 111.6 334.8 ;
      RECT  115.2 333.6 116.4 334.8 ;
      RECT  120.0 333.6 121.2 334.8 ;
      RECT  124.8 333.6 126.0 334.8 ;
      RECT  129.6 333.6 130.8 334.8 ;
      RECT  134.4 333.6 135.6 334.8 ;
      RECT  139.2 333.6 140.4 334.8 ;
      RECT  144.0 333.6 145.2 334.8 ;
      RECT  148.8 333.6 150.0 334.8 ;
      RECT  153.6 333.6 154.8 334.8 ;
      RECT  158.4 333.6 159.6 334.8 ;
      RECT  163.2 333.6 164.4 334.8 ;
      RECT  168.0 333.6 169.2 334.8 ;
      RECT  172.8 333.6 174.0 334.8 ;
      RECT  177.6 333.6 178.8 334.8 ;
      RECT  4.8 338.4 6.0 339.6 ;
      RECT  9.6 338.4 10.8 339.6 ;
      RECT  14.4 338.4 15.6 339.6 ;
      RECT  19.2 338.4 20.4 339.6 ;
      RECT  24.0 338.4 25.2 339.6 ;
      RECT  28.8 338.4 30.0 339.6 ;
      RECT  33.6 338.4 34.8 339.6 ;
      RECT  38.4 338.4 39.6 339.6 ;
      RECT  43.2 338.4 44.4 339.6 ;
      RECT  48.0 338.4 49.2 339.6 ;
      RECT  52.8 338.4 54.0 339.6 ;
      RECT  57.6 338.4 58.8 339.6 ;
      RECT  62.4 338.4 63.6 339.6 ;
      RECT  67.2 338.4 68.4 339.6 ;
      RECT  72.0 338.4 73.2 339.6 ;
      RECT  76.8 338.4 78.0 339.6 ;
      RECT  81.6 338.4 82.8 339.6 ;
      RECT  86.4 338.4 87.6 339.6 ;
      RECT  91.2 338.4 92.4 339.6 ;
      RECT  96.0 338.4 97.2 339.6 ;
      RECT  100.8 338.4 102.0 339.6 ;
      RECT  105.6 338.4 106.8 339.6 ;
      RECT  110.4 338.4 111.6 339.6 ;
      RECT  115.2 338.4 116.4 339.6 ;
      RECT  120.0 338.4 121.2 339.6 ;
      RECT  124.8 338.4 126.0 339.6 ;
      RECT  129.6 338.4 130.8 339.6 ;
      RECT  134.4 338.4 135.6 339.6 ;
      RECT  139.2 338.4 140.4 339.6 ;
      RECT  177.6 338.4 178.8 339.6 ;
      RECT  182.4 338.4 183.6 339.6 ;
      RECT  187.2 338.4 188.4 339.6 ;
      RECT  192.0 338.4 193.2 339.6 ;
      RECT  196.8 338.4 198.0 339.6 ;
      RECT  201.6 338.4 202.8 339.6 ;
      RECT  206.4 338.4 207.6 339.6 ;
      RECT  211.2 338.4 212.4 339.6 ;
      RECT  216.0 338.4 217.2 339.6 ;
      RECT  220.8 338.4 222.0 339.6 ;
      RECT  225.6 338.4 226.8 339.6 ;
      RECT  4.8 343.2 6.0 344.4 ;
      RECT  9.6 343.2 10.8 344.4 ;
      RECT  14.4 343.2 15.6 344.4 ;
      RECT  19.2 343.2 20.4 344.4 ;
      RECT  24.0 343.2 25.2 344.4 ;
      RECT  28.8 343.2 30.0 344.4 ;
      RECT  33.6 343.2 34.8 344.4 ;
      RECT  38.4 343.2 39.6 344.4 ;
      RECT  43.2 343.2 44.4 344.4 ;
      RECT  48.0 343.2 49.2 344.4 ;
      RECT  52.8 343.2 54.0 344.4 ;
      RECT  57.6 343.2 58.8 344.4 ;
      RECT  62.4 343.2 63.6 344.4 ;
      RECT  67.2 343.2 68.4 344.4 ;
      RECT  72.0 343.2 73.2 344.4 ;
      RECT  76.8 343.2 78.0 344.4 ;
      RECT  100.8 343.2 102.0 344.4 ;
      RECT  105.6 343.2 106.8 344.4 ;
      RECT  110.4 343.2 111.6 344.4 ;
      RECT  115.2 343.2 116.4 344.4 ;
      RECT  120.0 343.2 121.2 344.4 ;
      RECT  124.8 343.2 126.0 344.4 ;
      RECT  129.6 343.2 130.8 344.4 ;
      RECT  134.4 343.2 135.6 344.4 ;
      RECT  139.2 343.2 140.4 344.4 ;
      RECT  144.0 343.2 145.2 344.4 ;
      RECT  148.8 343.2 150.0 344.4 ;
      RECT  153.6 343.2 154.8 344.4 ;
      RECT  158.4 343.2 159.6 344.4 ;
      RECT  163.2 343.2 164.4 344.4 ;
      RECT  168.0 343.2 169.2 344.4 ;
      RECT  172.8 343.2 174.0 344.4 ;
      RECT  177.6 343.2 178.8 344.4 ;
      RECT  4.8 348.0 6.0 349.2 ;
      RECT  9.6 348.0 10.8 349.2 ;
      RECT  14.4 348.0 15.6 349.2 ;
      RECT  19.2 348.0 20.4 349.2 ;
      RECT  24.0 348.0 25.2 349.2 ;
      RECT  28.8 348.0 30.0 349.2 ;
      RECT  33.6 348.0 34.8 349.2 ;
      RECT  38.4 348.0 39.6 349.2 ;
      RECT  43.2 348.0 44.4 349.2 ;
      RECT  48.0 348.0 49.2 349.2 ;
      RECT  52.8 348.0 54.0 349.2 ;
      RECT  57.6 348.0 58.8 349.2 ;
      RECT  62.4 348.0 63.6 349.2 ;
      RECT  67.2 348.0 68.4 349.2 ;
      RECT  72.0 348.0 73.2 349.2 ;
      RECT  76.8 348.0 78.0 349.2 ;
      RECT  81.6 348.0 82.8 349.2 ;
      RECT  86.4 348.0 87.6 349.2 ;
      RECT  91.2 348.0 92.4 349.2 ;
      RECT  96.0 348.0 97.2 349.2 ;
      RECT  100.8 348.0 102.0 349.2 ;
      RECT  105.6 348.0 106.8 349.2 ;
      RECT  110.4 348.0 111.6 349.2 ;
      RECT  115.2 348.0 116.4 349.2 ;
      RECT  120.0 348.0 121.2 349.2 ;
      RECT  124.8 348.0 126.0 349.2 ;
      RECT  129.6 348.0 130.8 349.2 ;
      RECT  134.4 348.0 135.6 349.2 ;
      RECT  139.2 348.0 140.4 349.2 ;
      RECT  144.0 348.0 145.2 349.2 ;
      RECT  148.8 348.0 150.0 349.2 ;
      RECT  153.6 348.0 154.8 349.2 ;
      RECT  158.4 348.0 159.6 349.2 ;
      RECT  163.2 348.0 164.4 349.2 ;
      RECT  168.0 348.0 169.2 349.2 ;
      RECT  172.8 348.0 174.0 349.2 ;
      RECT  177.6 348.0 178.8 349.2 ;
      RECT  182.4 348.0 183.6 349.2 ;
      RECT  187.2 348.0 188.4 349.2 ;
      RECT  192.0 348.0 193.2 349.2 ;
      RECT  196.8 348.0 198.0 349.2 ;
      RECT  201.6 348.0 202.8 349.2 ;
      RECT  206.4 348.0 207.6 349.2 ;
      RECT  211.2 348.0 212.4 349.2 ;
      RECT  216.0 348.0 217.2 349.2 ;
      RECT  220.8 348.0 222.0 349.2 ;
      RECT  225.6 348.0 226.8 349.2 ;
      RECT  4.8 352.8 6.0 354.0 ;
      RECT  9.6 352.8 10.8 354.0 ;
      RECT  14.4 352.8 15.6 354.0 ;
      RECT  19.2 352.8 20.4 354.0 ;
      RECT  24.0 352.8 25.2 354.0 ;
      RECT  28.8 352.8 30.0 354.0 ;
      RECT  33.6 352.8 34.8 354.0 ;
      RECT  38.4 352.8 39.6 354.0 ;
      RECT  43.2 352.8 44.4 354.0 ;
      RECT  48.0 352.8 49.2 354.0 ;
      RECT  52.8 352.8 54.0 354.0 ;
      RECT  57.6 352.8 58.8 354.0 ;
      RECT  62.4 352.8 63.6 354.0 ;
      RECT  67.2 352.8 68.4 354.0 ;
      RECT  72.0 352.8 73.2 354.0 ;
      RECT  76.8 352.8 78.0 354.0 ;
      RECT  81.6 352.8 82.8 354.0 ;
      RECT  86.4 352.8 87.6 354.0 ;
      RECT  91.2 352.8 92.4 354.0 ;
      RECT  96.0 352.8 97.2 354.0 ;
      RECT  100.8 352.8 102.0 354.0 ;
      RECT  105.6 352.8 106.8 354.0 ;
      RECT  110.4 352.8 111.6 354.0 ;
      RECT  115.2 352.8 116.4 354.0 ;
      RECT  120.0 352.8 121.2 354.0 ;
      RECT  124.8 352.8 126.0 354.0 ;
      RECT  129.6 352.8 130.8 354.0 ;
      RECT  134.4 352.8 135.6 354.0 ;
      RECT  139.2 352.8 140.4 354.0 ;
      RECT  144.0 352.8 145.2 354.0 ;
      RECT  148.8 352.8 150.0 354.0 ;
      RECT  153.6 352.8 154.8 354.0 ;
      RECT  158.4 352.8 159.6 354.0 ;
      RECT  163.2 352.8 164.4 354.0 ;
      RECT  168.0 352.8 169.2 354.0 ;
      RECT  172.8 352.8 174.0 354.0 ;
      RECT  177.6 352.8 178.8 354.0 ;
      RECT  4.8 357.6 6.0 358.8 ;
      RECT  9.6 357.6 10.8 358.8 ;
      RECT  14.4 357.6 15.6 358.8 ;
      RECT  19.2 357.6 20.4 358.8 ;
      RECT  24.0 357.6 25.2 358.8 ;
      RECT  28.8 357.6 30.0 358.8 ;
      RECT  33.6 357.6 34.8 358.8 ;
      RECT  38.4 357.6 39.6 358.8 ;
      RECT  43.2 357.6 44.4 358.8 ;
      RECT  48.0 357.6 49.2 358.8 ;
      RECT  52.8 357.6 54.0 358.8 ;
      RECT  57.6 357.6 58.8 358.8 ;
      RECT  62.4 357.6 63.6 358.8 ;
      RECT  67.2 357.6 68.4 358.8 ;
      RECT  72.0 357.6 73.2 358.8 ;
      RECT  76.8 357.6 78.0 358.8 ;
      RECT  81.6 357.6 82.8 358.8 ;
      RECT  86.4 357.6 87.6 358.8 ;
      RECT  91.2 357.6 92.4 358.8 ;
      RECT  96.0 357.6 97.2 358.8 ;
      RECT  100.8 357.6 102.0 358.8 ;
      RECT  105.6 357.6 106.8 358.8 ;
      RECT  110.4 357.6 111.6 358.8 ;
      RECT  115.2 357.6 116.4 358.8 ;
      RECT  120.0 357.6 121.2 358.8 ;
      RECT  124.8 357.6 126.0 358.8 ;
      RECT  129.6 357.6 130.8 358.8 ;
      RECT  134.4 357.6 135.6 358.8 ;
      RECT  139.2 357.6 140.4 358.8 ;
      RECT  144.0 357.6 145.2 358.8 ;
      RECT  148.8 357.6 150.0 358.8 ;
      RECT  153.6 357.6 154.8 358.8 ;
      RECT  158.4 357.6 159.6 358.8 ;
      RECT  163.2 357.6 164.4 358.8 ;
      RECT  168.0 357.6 169.2 358.8 ;
      RECT  172.8 357.6 174.0 358.8 ;
      RECT  177.6 357.6 178.8 358.8 ;
      RECT  182.4 357.6 183.6 358.8 ;
      RECT  187.2 357.6 188.4 358.8 ;
      RECT  192.0 357.6 193.2 358.8 ;
      RECT  196.8 357.6 198.0 358.8 ;
      RECT  201.6 357.6 202.8 358.8 ;
      RECT  206.4 357.6 207.6 358.8 ;
      RECT  211.2 357.6 212.4 358.8 ;
      RECT  216.0 357.6 217.2 358.8 ;
      RECT  220.8 357.6 222.0 358.8 ;
      RECT  225.6 357.6 226.8 358.8 ;
      RECT  4.8 362.4 6.0 363.6 ;
      RECT  9.6 362.4 10.8 363.6 ;
      RECT  14.4 362.4 15.6 363.6 ;
      RECT  19.2 362.4 20.4 363.6 ;
      RECT  24.0 362.4 25.2 363.6 ;
      RECT  28.8 362.4 30.0 363.6 ;
      RECT  33.6 362.4 34.8 363.6 ;
      RECT  38.4 362.4 39.6 363.6 ;
      RECT  43.2 362.4 44.4 363.6 ;
      RECT  48.0 362.4 49.2 363.6 ;
      RECT  52.8 362.4 54.0 363.6 ;
      RECT  57.6 362.4 58.8 363.6 ;
      RECT  62.4 362.4 63.6 363.6 ;
      RECT  67.2 362.4 68.4 363.6 ;
      RECT  72.0 362.4 73.2 363.6 ;
      RECT  76.8 362.4 78.0 363.6 ;
      RECT  100.8 362.4 102.0 363.6 ;
      RECT  105.6 362.4 106.8 363.6 ;
      RECT  110.4 362.4 111.6 363.6 ;
      RECT  115.2 362.4 116.4 363.6 ;
      RECT  120.0 362.4 121.2 363.6 ;
      RECT  124.8 362.4 126.0 363.6 ;
      RECT  129.6 362.4 130.8 363.6 ;
      RECT  134.4 362.4 135.6 363.6 ;
      RECT  139.2 362.4 140.4 363.6 ;
      RECT  177.6 362.4 178.8 363.6 ;
      RECT  182.4 362.4 183.6 363.6 ;
      RECT  187.2 362.4 188.4 363.6 ;
      RECT  192.0 362.4 193.2 363.6 ;
      RECT  196.8 362.4 198.0 363.6 ;
      RECT  201.6 362.4 202.8 363.6 ;
      RECT  206.4 362.4 207.6 363.6 ;
      RECT  211.2 362.4 212.4 363.6 ;
      RECT  216.0 362.4 217.2 363.6 ;
      RECT  220.8 362.4 222.0 363.6 ;
      RECT  225.6 362.4 226.8 363.6 ;
      RECT  4.8 367.2 6.0 368.4 ;
      RECT  9.6 367.2 10.8 368.4 ;
      RECT  14.4 367.2 15.6 368.4 ;
      RECT  19.2 367.2 20.4 368.4 ;
      RECT  24.0 367.2 25.2 368.4 ;
      RECT  28.8 367.2 30.0 368.4 ;
      RECT  33.6 367.2 34.8 368.4 ;
      RECT  38.4 367.2 39.6 368.4 ;
      RECT  43.2 367.2 44.4 368.4 ;
      RECT  48.0 367.2 49.2 368.4 ;
      RECT  52.8 367.2 54.0 368.4 ;
      RECT  57.6 367.2 58.8 368.4 ;
      RECT  62.4 367.2 63.6 368.4 ;
      RECT  67.2 367.2 68.4 368.4 ;
      RECT  72.0 367.2 73.2 368.4 ;
      RECT  76.8 367.2 78.0 368.4 ;
      RECT  81.6 367.2 82.8 368.4 ;
      RECT  86.4 367.2 87.6 368.4 ;
      RECT  91.2 367.2 92.4 368.4 ;
      RECT  96.0 367.2 97.2 368.4 ;
      RECT  100.8 367.2 102.0 368.4 ;
      RECT  105.6 367.2 106.8 368.4 ;
      RECT  110.4 367.2 111.6 368.4 ;
      RECT  115.2 367.2 116.4 368.4 ;
      RECT  120.0 367.2 121.2 368.4 ;
      RECT  124.8 367.2 126.0 368.4 ;
      RECT  129.6 367.2 130.8 368.4 ;
      RECT  134.4 367.2 135.6 368.4 ;
      RECT  139.2 367.2 140.4 368.4 ;
      RECT  144.0 367.2 145.2 368.4 ;
      RECT  148.8 367.2 150.0 368.4 ;
      RECT  153.6 367.2 154.8 368.4 ;
      RECT  158.4 367.2 159.6 368.4 ;
      RECT  163.2 367.2 164.4 368.4 ;
      RECT  168.0 367.2 169.2 368.4 ;
      RECT  172.8 367.2 174.0 368.4 ;
      RECT  177.6 367.2 178.8 368.4 ;
      RECT  105.6 247.2 106.8 248.4 ;
      RECT  105.6 204.0 106.8 205.2 ;
      RECT  187.2 369.6 188.4 370.8 ;
      RECT  196.8 369.6 198.0 370.8 ;
      RECT  201.6 369.6 202.8 370.8 ;
      RECT  211.2 369.6 212.4 370.8 ;
      RECT  216.0 369.6 217.2 370.8 ;
   END
   END    sram_2_16_scn4m_subm
END    LIBRARY
