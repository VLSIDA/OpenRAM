magic
tech sky130A
magscale 1 2
timestamp 1591909763
<< nwell >>
rect -8 676 1176 1467
<< nmos >>
rect 81 102 111 302
rect 167 102 197 302
rect 239 102 269 302
rect 359 102 389 302
rect 431 102 461 302
rect 517 102 547 302
rect 589 102 619 302
rect 709 102 739 302
rect 781 102 811 302
rect 867 102 897 302
rect 1057 102 1087 302
<< pmos >>
rect 81 712 111 1312
rect 167 712 197 1312
rect 239 712 269 1312
rect 359 712 389 1312
rect 431 712 461 1312
rect 517 712 547 1312
rect 589 712 619 1312
rect 709 712 739 1312
rect 781 712 811 1312
rect 867 712 897 1312
rect 1057 712 1087 1312
<< ndiff >>
rect 28 254 81 302
rect 28 118 36 254
rect 70 118 81 254
rect 28 102 81 118
rect 111 254 167 302
rect 111 118 122 254
rect 156 118 167 254
rect 111 102 167 118
rect 197 102 239 302
rect 269 254 359 302
rect 269 118 280 254
rect 348 118 359 254
rect 269 102 359 118
rect 389 102 431 302
rect 461 254 517 302
rect 461 118 472 254
rect 506 118 517 254
rect 461 102 517 118
rect 547 102 589 302
rect 619 254 709 302
rect 619 118 630 254
rect 698 118 709 254
rect 619 102 709 118
rect 739 102 781 302
rect 811 254 867 302
rect 811 118 822 254
rect 856 118 867 254
rect 811 102 867 118
rect 897 254 950 302
rect 897 118 908 254
rect 942 118 950 254
rect 897 102 950 118
rect 1004 254 1057 302
rect 1004 118 1012 254
rect 1046 118 1057 254
rect 1004 102 1057 118
rect 1087 254 1140 302
rect 1087 118 1098 254
rect 1132 118 1140 254
rect 1087 102 1140 118
<< pdiff >>
rect 28 1296 81 1312
rect 28 820 36 1296
rect 70 820 81 1296
rect 28 712 81 820
rect 111 1296 167 1312
rect 111 820 122 1296
rect 156 820 167 1296
rect 111 712 167 820
rect 197 712 239 1312
rect 269 1296 359 1312
rect 269 820 280 1296
rect 348 820 359 1296
rect 269 712 359 820
rect 389 712 431 1312
rect 461 1296 517 1312
rect 461 820 472 1296
rect 506 820 517 1296
rect 461 712 517 820
rect 547 712 589 1312
rect 619 1296 709 1312
rect 619 820 630 1296
rect 698 820 709 1296
rect 619 712 709 820
rect 739 712 781 1312
rect 811 1296 867 1312
rect 811 820 822 1296
rect 856 820 867 1296
rect 811 712 867 820
rect 897 1296 950 1312
rect 897 820 908 1296
rect 942 820 950 1296
rect 897 712 950 820
rect 1004 1296 1057 1312
rect 1004 820 1012 1296
rect 1046 820 1057 1296
rect 1004 712 1057 820
rect 1087 1296 1140 1312
rect 1087 820 1098 1296
rect 1132 820 1140 1296
rect 1087 712 1140 820
<< ndiffc >>
rect 36 118 70 254
rect 122 118 156 254
rect 280 118 348 254
rect 472 118 506 254
rect 630 118 698 254
rect 822 118 856 254
rect 908 118 942 254
rect 1012 118 1046 254
rect 1098 118 1132 254
<< pdiffc >>
rect 36 820 70 1296
rect 122 820 156 1296
rect 280 820 348 1296
rect 472 820 506 1296
rect 630 820 698 1296
rect 822 820 856 1296
rect 908 820 942 1296
rect 1012 820 1046 1296
rect 1098 820 1132 1296
<< psubdiff >>
rect 28 -17 52 17
rect 86 -17 110 17
rect 164 -17 188 17
rect 222 -17 246 17
rect 300 -17 324 17
rect 358 -17 382 17
rect 436 -17 460 17
rect 494 -17 518 17
rect 572 -17 596 17
rect 630 -17 654 17
rect 708 -17 732 17
rect 766 -17 790 17
rect 844 -17 868 17
rect 902 -17 926 17
rect 980 -17 1004 17
rect 1038 -17 1062 17
<< nsubdiff >>
rect 28 1397 52 1431
rect 86 1397 110 1431
rect 164 1397 188 1431
rect 222 1397 246 1431
rect 300 1397 324 1431
rect 358 1397 382 1431
rect 436 1397 460 1431
rect 494 1397 518 1431
rect 572 1397 596 1431
rect 630 1397 654 1431
rect 708 1397 732 1431
rect 766 1397 790 1431
rect 844 1397 868 1431
rect 902 1397 926 1431
rect 980 1397 1004 1431
rect 1038 1397 1062 1431
<< psubdiffcont >>
rect 52 -17 86 17
rect 188 -17 222 17
rect 324 -17 358 17
rect 460 -17 494 17
rect 596 -17 630 17
rect 732 -17 766 17
rect 868 -17 902 17
rect 1004 -17 1038 17
<< nsubdiffcont >>
rect 52 1397 86 1431
rect 188 1397 222 1431
rect 324 1397 358 1431
rect 460 1397 494 1431
rect 596 1397 630 1431
rect 732 1397 766 1431
rect 868 1397 902 1431
rect 1004 1397 1038 1431
<< poly >>
rect 81 1312 111 1338
rect 167 1312 197 1338
rect 239 1312 269 1338
rect 359 1312 389 1338
rect 431 1312 461 1338
rect 517 1312 547 1338
rect 589 1312 619 1338
rect 709 1312 739 1338
rect 781 1312 811 1338
rect 867 1312 897 1338
rect 1057 1312 1087 1338
rect 81 697 111 712
rect 70 677 111 697
rect 47 667 111 677
rect 47 661 101 667
rect 47 627 57 661
rect 91 627 101 661
rect 47 611 101 627
rect 71 447 101 611
rect 167 597 197 712
rect 239 672 269 712
rect 239 656 293 672
rect 239 622 249 656
rect 283 622 293 656
rect 239 606 293 622
rect 143 581 197 597
rect 143 547 153 581
rect 187 547 197 581
rect 143 531 197 547
rect 359 531 389 712
rect 431 667 461 712
rect 517 667 547 712
rect 431 657 547 667
rect 431 623 472 657
rect 506 623 547 657
rect 431 613 547 623
rect 589 531 619 712
rect 709 672 739 712
rect 685 656 739 672
rect 685 622 695 656
rect 729 622 739 656
rect 685 606 739 622
rect 781 597 811 712
rect 867 677 897 712
rect 867 661 938 677
rect 867 647 894 661
rect 878 627 894 647
rect 928 627 938 661
rect 878 611 938 627
rect 781 581 835 597
rect 781 547 791 581
rect 825 547 835 581
rect 781 531 835 547
rect 71 417 111 447
rect 81 302 111 417
rect 167 302 197 531
rect 239 501 739 531
rect 239 302 269 501
rect 685 467 695 501
rect 729 467 739 501
rect 685 451 739 467
rect 335 421 389 437
rect 335 387 345 421
rect 379 387 389 421
rect 335 371 389 387
rect 359 302 389 371
rect 431 421 547 431
rect 431 387 472 421
rect 506 387 547 421
rect 431 377 547 387
rect 431 302 461 377
rect 517 302 547 377
rect 589 421 643 437
rect 589 387 599 421
rect 633 387 643 421
rect 589 371 643 387
rect 589 302 619 371
rect 709 302 739 451
rect 781 302 811 531
rect 878 481 908 611
rect 1057 517 1087 712
rect 867 371 908 481
rect 1033 501 1087 517
rect 1033 467 1043 501
rect 1077 467 1087 501
rect 1033 451 1087 467
rect 867 302 897 371
rect 1057 302 1087 451
rect 81 76 111 102
rect 167 76 197 102
rect 239 76 269 102
rect 359 76 389 102
rect 431 76 461 102
rect 517 76 547 102
rect 589 76 619 102
rect 709 76 739 102
rect 781 76 811 102
rect 867 76 897 102
rect 1057 76 1087 102
<< polycont >>
rect 57 627 91 661
rect 249 622 283 656
rect 153 547 187 581
rect 472 623 506 657
rect 695 622 729 656
rect 894 627 928 661
rect 791 547 825 581
rect 695 467 729 501
rect 345 387 379 421
rect 472 387 506 421
rect 599 387 633 421
rect 1043 467 1077 501
<< locali >>
rect 0 1431 1168 1432
rect 0 1397 52 1431
rect 86 1397 188 1431
rect 222 1397 324 1431
rect 358 1397 460 1431
rect 494 1397 596 1431
rect 630 1397 732 1431
rect 766 1397 868 1431
rect 902 1397 1004 1431
rect 1038 1397 1168 1431
rect 0 1396 1168 1397
rect 36 1296 70 1312
rect 122 1296 156 1396
rect 122 804 156 820
rect 280 1296 348 1312
rect 280 804 297 820
rect 331 804 348 820
rect 472 1296 506 1396
rect 472 804 506 820
rect 630 1296 698 1312
rect 630 804 647 820
rect 681 804 698 820
rect 822 1296 856 1396
rect 822 804 856 820
rect 908 1296 942 1312
rect 1012 1296 1046 1396
rect 1012 804 1046 820
rect 1098 1296 1132 1312
rect 41 707 379 741
rect 413 707 1132 741
rect 41 627 57 661
rect 91 627 113 661
rect 249 656 283 707
rect 456 623 472 657
rect 506 623 522 657
rect 249 606 283 622
rect 137 547 153 581
rect 187 547 203 581
rect 472 566 506 623
rect 239 532 506 566
rect 239 501 273 532
rect 70 467 273 501
rect 472 421 506 532
rect 599 421 633 707
rect 695 656 729 707
rect 894 661 928 707
rect 878 627 894 661
rect 928 627 944 661
rect 695 606 729 622
rect 1098 581 1132 618
rect 775 547 791 581
rect 825 547 1132 581
rect 679 467 695 501
rect 729 467 908 501
rect 1012 467 1020 501
rect 1077 467 1093 501
rect 328 387 345 421
rect 456 387 472 421
rect 506 387 522 421
rect 583 387 599 421
rect 633 387 649 421
rect 1012 341 1046 467
rect 647 307 1046 341
rect 647 270 681 307
rect 36 261 70 270
rect 36 102 70 118
rect 122 254 156 270
rect 122 20 156 118
rect 280 261 348 270
rect 280 254 297 261
rect 331 254 348 261
rect 280 102 348 118
rect 472 254 506 270
rect 472 20 506 118
rect 630 261 698 270
rect 630 254 647 261
rect 681 254 698 261
rect 630 102 698 118
rect 822 254 856 270
rect 822 20 856 118
rect 908 261 942 271
rect 908 102 942 118
rect 1012 254 1046 270
rect 1012 20 1046 118
rect 1098 261 1132 271
rect 1098 102 1132 118
rect 0 17 1168 20
rect 0 -17 52 17
rect 86 -17 188 17
rect 222 -17 324 17
rect 358 -17 460 17
rect 494 -17 596 17
rect 630 -17 732 17
rect 766 -17 868 17
rect 902 -17 1004 17
rect 1038 -17 1168 17
rect 0 -20 1168 -17
<< viali >>
rect 36 820 70 821
rect 36 787 70 820
rect 297 820 331 821
rect 297 787 331 820
rect 647 820 681 821
rect 647 787 681 820
rect 908 820 942 821
rect 908 787 942 820
rect 1098 820 1132 821
rect 1098 787 1132 820
rect 379 707 413 741
rect 113 627 147 661
rect 153 547 187 581
rect 36 467 70 501
rect 1098 618 1132 652
rect 908 467 942 501
rect 1020 467 1043 501
rect 1043 467 1054 501
rect 379 387 413 421
rect 36 254 70 261
rect 36 227 70 254
rect 297 254 331 261
rect 297 227 331 254
rect 647 254 681 261
rect 647 227 681 254
rect 908 254 942 261
rect 908 227 942 254
rect 1098 254 1132 261
rect 1098 227 1132 254
<< metal1 >>
rect 24 821 82 827
rect 24 787 36 821
rect 70 787 82 821
rect 24 781 82 787
rect 285 821 343 827
rect 285 787 297 821
rect 331 787 343 821
rect 285 781 343 787
rect 635 821 693 827
rect 635 787 647 821
rect 681 787 693 821
rect 635 781 693 787
rect 896 821 954 827
rect 896 787 908 821
rect 942 787 954 821
rect 896 781 954 787
rect 1086 821 1144 827
rect 1086 787 1098 821
rect 1132 787 1144 821
rect 1086 781 1144 787
rect 36 507 70 781
rect 101 661 159 667
rect 297 661 331 781
rect 369 750 423 756
rect 367 701 369 747
rect 423 701 425 747
rect 369 692 423 698
rect 101 627 113 661
rect 147 627 331 661
rect 101 621 159 627
rect 137 538 143 590
rect 197 538 203 590
rect 24 501 82 507
rect 24 467 36 501
rect 70 467 82 501
rect 24 461 82 467
rect 36 267 70 461
rect 297 267 331 627
rect 379 436 413 692
rect 369 427 423 436
rect 367 421 425 427
rect 367 387 379 421
rect 413 387 425 421
rect 367 381 425 387
rect 369 372 423 381
rect 647 267 681 781
rect 908 507 942 781
rect 1098 661 1132 781
rect 1082 609 1088 661
rect 1142 609 1148 661
rect 896 501 954 507
rect 896 467 908 501
rect 942 467 954 501
rect 896 461 954 467
rect 908 267 942 461
rect 1004 458 1010 510
rect 1064 458 1070 510
rect 1098 267 1132 609
rect 24 261 82 267
rect 24 227 36 261
rect 70 227 82 261
rect 24 221 82 227
rect 285 261 343 267
rect 285 227 297 261
rect 331 227 343 261
rect 285 221 343 227
rect 635 261 693 267
rect 635 227 647 261
rect 681 227 693 261
rect 635 221 693 227
rect 896 261 954 267
rect 896 227 908 261
rect 942 227 954 261
rect 896 221 954 227
rect 1086 261 1144 267
rect 1086 227 1098 261
rect 1132 227 1144 261
rect 1086 221 1144 227
<< via1 >>
rect 369 741 423 750
rect 369 707 379 741
rect 379 707 413 741
rect 413 707 423 741
rect 369 698 423 707
rect 143 581 197 590
rect 143 547 153 581
rect 153 547 187 581
rect 187 547 197 581
rect 143 538 197 547
rect 1088 652 1142 661
rect 1088 618 1098 652
rect 1098 618 1132 652
rect 1132 618 1142 652
rect 1088 609 1142 618
rect 1010 501 1064 510
rect 1010 467 1020 501
rect 1020 467 1054 501
rect 1054 467 1064 501
rect 1010 458 1064 467
<< metal2 >>
rect 369 750 423 756
rect 369 692 423 698
rect 1082 609 1088 661
rect 1142 609 1148 661
rect 137 538 143 590
rect 197 538 203 590
rect 1004 458 1010 510
rect 1064 458 1070 510
<< labels >>
rlabel metal2 1146 659 1146 659 1 Q
rlabel metal2 419 753 419 753 1 clk
rlabel metal2 1007 504 1007 504 1 ON
rlabel metal2 139 586 139 586 1 D
rlabel locali 544 0 544 0 1 gnd
rlabel locali 548 1416 548 1416 1 vdd
<< properties >>
string FIXED_BBOX 0 0 1168 1414
string BBOX_FIXED 0 0 1168 1414
<< end >>
