VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_2_16_1_freepdk45
   CLASS BLOCK ;
   SIZE 23.88 BY 46.6 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  12.7725 1.0375 12.85 1.1725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  15.6325 1.0375 15.71 1.1725 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  7.0525 37.7375 7.13 37.8725 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  7.0525 40.4775 7.13 40.6125 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  7.0525 42.6875 7.13 42.8225 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  7.0525 45.4275 7.13 45.5625 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  0.245 1.0375 0.3225 1.1725 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  0.245 3.7775 0.3225 3.9125 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  6.155 1.1575 6.225 1.2275 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal2 ;
         RECT  21.375 12.825 21.445 13.2225 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal2 ;
         RECT  22.08 12.825 22.15 13.2225 ;
      END
   END dout0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  21.655 45.5475 21.79 45.6825 ;
         LAYER metal3 ;
         RECT  8.12 39.1125 8.255 39.2475 ;
         LAYER metal3 ;
         RECT  -0.0675 2.4125 0.0675 2.5475 ;
         LAYER metal3 ;
         RECT  23.065 24.0275 23.2 24.1625 ;
         LAYER metal3 ;
         RECT  20.95 45.5475 21.085 45.6825 ;
         LAYER metal3 ;
         RECT  2.125 36.3725 2.26 36.5075 ;
         LAYER metal3 ;
         RECT  18.6925 34.7875 18.8275 34.9225 ;
         LAYER metal3 ;
         RECT  9.46 17.2575 9.595 17.3925 ;
         LAYER metal3 ;
         RECT  8.12 44.0525 8.255 44.1875 ;
         LAYER metal3 ;
         RECT  23.065 40.1675 23.2 40.3025 ;
         LAYER metal3 ;
         RECT  17.1025 29.4075 17.2375 29.5425 ;
         LAYER metal3 ;
         RECT  21.0075 19.3325 21.0775 19.4675 ;
         LAYER metal3 ;
         RECT  18.6925 37.4775 18.8275 37.6125 ;
         LAYER metal3 ;
         RECT  17.1025 40.1675 17.2375 40.3025 ;
         LAYER metal3 ;
         RECT  0.75 32.7325 0.885 32.8675 ;
         LAYER metal3 ;
         RECT  17.915 21.3375 18.05 21.4725 ;
         LAYER metal3 ;
         RECT  18.6925 26.7175 18.8275 26.8525 ;
         LAYER metal3 ;
         RECT  23.065 34.7875 23.2 34.9225 ;
         LAYER metal3 ;
         RECT  18.6925 40.1675 18.8275 40.3025 ;
         LAYER metal3 ;
         RECT  2.125 32.7325 2.26 32.8675 ;
         LAYER metal3 ;
         RECT  16.7 2.4025 16.835 2.5375 ;
         LAYER metal3 ;
         RECT  9.46 2.4075 9.595 2.5425 ;
         LAYER metal3 ;
         RECT  23.065 26.7175 23.2 26.8525 ;
         LAYER metal3 ;
         RECT  22.3975 13.2925 22.4675 13.4275 ;
         LAYER metal3 ;
         RECT  11.0325 26.7175 11.1675 26.8525 ;
         LAYER metal3 ;
         RECT  20.245 29.4075 20.38 29.5425 ;
         LAYER metal3 ;
         RECT  20.245 37.4775 20.38 37.6125 ;
         LAYER metal3 ;
         RECT  11.0325 32.0975 11.1675 32.2325 ;
         LAYER metal3 ;
         RECT  21.7125 19.3325 21.7825 19.4675 ;
         LAYER metal3 ;
         RECT  20.245 40.1675 20.38 40.3025 ;
         LAYER metal3 ;
         RECT  17.1025 24.0275 17.2375 24.1625 ;
         LAYER metal3 ;
         RECT  12.56 32.0975 12.695 32.2325 ;
         LAYER metal3 ;
         RECT  22.2175 8.5075 22.2875 8.6425 ;
         LAYER metal3 ;
         RECT  21.6925 13.2925 21.7625 13.4275 ;
         LAYER metal3 ;
         RECT  -0.0675 2.4025 0.0675 2.5375 ;
         LAYER metal3 ;
         RECT  2.125 29.0925 2.26 29.2275 ;
         LAYER metal3 ;
         RECT  17.1025 26.7175 17.2375 26.8525 ;
         LAYER metal3 ;
         RECT  12.56 34.7875 12.695 34.9225 ;
         LAYER metal3 ;
         RECT  23.065 45.5475 23.2 45.6825 ;
         LAYER metal3 ;
         RECT  20.245 32.0975 20.38 32.2325 ;
         LAYER metal3 ;
         RECT  13.84 2.4025 13.975 2.5375 ;
         LAYER metal3 ;
         RECT  22.36 45.5475 22.495 45.6825 ;
         LAYER metal3 ;
         RECT  20.245 34.7875 20.38 34.9225 ;
         LAYER metal3 ;
         RECT  20.245 21.3375 20.38 21.4725 ;
         LAYER metal3 ;
         RECT  2.125 21.8125 2.26 21.9475 ;
         LAYER metal3 ;
         RECT  17.1025 42.8575 17.2375 42.9925 ;
         LAYER metal3 ;
         RECT  20.245 42.8575 20.38 42.9925 ;
         LAYER metal3 ;
         RECT  18.6925 24.0275 18.8275 24.1625 ;
         LAYER metal3 ;
         RECT  8.12 44.0625 8.255 44.1975 ;
         LAYER metal3 ;
         RECT  18.6925 42.8575 18.8275 42.9925 ;
         LAYER metal3 ;
         RECT  20.95 21.3375 21.085 21.4725 ;
         LAYER metal3 ;
         RECT  22.4175 19.3325 22.4875 19.4675 ;
         LAYER metal3 ;
         RECT  17.1025 37.4775 17.2375 37.6125 ;
         LAYER metal3 ;
         RECT  23.065 42.8575 23.2 42.9925 ;
         LAYER metal3 ;
         RECT  21.655 21.3375 21.79 21.4725 ;
         LAYER metal3 ;
         RECT  18.6925 32.0975 18.8275 32.2325 ;
         LAYER metal3 ;
         RECT  20.245 45.5475 20.38 45.6825 ;
         LAYER metal3 ;
         RECT  17.1025 34.7875 17.2375 34.9225 ;
         LAYER metal3 ;
         RECT  2.125 25.4525 2.26 25.5875 ;
         LAYER metal3 ;
         RECT  8.12 39.1025 8.255 39.2375 ;
         LAYER metal3 ;
         RECT  23.065 37.4775 23.2 37.6125 ;
         LAYER metal3 ;
         RECT  0.75 29.0925 0.885 29.2275 ;
         LAYER metal3 ;
         RECT  20.245 24.0275 20.38 24.1625 ;
         LAYER metal3 ;
         RECT  9.46 12.3075 9.595 12.4425 ;
         LAYER metal3 ;
         RECT  11.0325 24.0275 11.1675 24.1625 ;
         LAYER metal3 ;
         RECT  23.065 21.3375 23.2 21.4725 ;
         LAYER metal3 ;
         RECT  23.065 29.4075 23.2 29.5425 ;
         LAYER metal3 ;
         RECT  9.46 7.3575 9.595 7.4925 ;
         LAYER metal3 ;
         RECT  0.75 21.8125 0.885 21.9475 ;
         LAYER metal3 ;
         RECT  0.75 25.4525 0.885 25.5875 ;
         LAYER metal3 ;
         RECT  22.36 21.3375 22.495 21.4725 ;
         LAYER metal3 ;
         RECT  11.0325 34.7875 11.1675 34.9225 ;
         LAYER metal3 ;
         RECT  17.1025 32.0975 17.2375 32.2325 ;
         LAYER metal3 ;
         RECT  12.56 24.0275 12.695 24.1625 ;
         LAYER metal3 ;
         RECT  18.6925 29.4075 18.8275 29.5425 ;
         LAYER metal3 ;
         RECT  21.5125 8.5075 21.5825 8.6425 ;
         LAYER metal3 ;
         RECT  12.56 26.7175 12.695 26.8525 ;
         LAYER metal3 ;
         RECT  20.245 26.7175 20.38 26.8525 ;
         LAYER metal3 ;
         RECT  0.75 36.3725 0.885 36.5075 ;
         LAYER metal3 ;
         RECT  23.065 32.0975 23.2 32.2325 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  17.1025 22.6825 17.2375 22.8175 ;
         LAYER metal3 ;
         RECT  18.6925 33.4425 18.8275 33.5775 ;
         LAYER metal3 ;
         RECT  20.6025 44.2025 20.7375 44.3375 ;
         LAYER metal3 ;
         RECT  18.6925 44.2025 18.8275 44.3375 ;
         LAYER metal3 ;
         RECT  22.7175 30.7525 22.8525 30.8875 ;
         LAYER metal3 ;
         RECT  22.75 17.3275 22.82 17.4625 ;
         LAYER metal3 ;
         RECT  22.045 10.5575 22.115 10.6925 ;
         LAYER metal3 ;
         RECT  21.3075 44.2025 21.4425 44.3375 ;
         LAYER metal3 ;
         RECT  22.7175 36.1325 22.8525 36.2675 ;
         LAYER metal3 ;
         RECT  19.8975 30.7525 20.0325 30.8875 ;
         LAYER metal3 ;
         RECT  18.6925 30.7525 18.8275 30.8875 ;
         LAYER metal3 ;
         RECT  21.3075 19.9925 21.4425 20.1275 ;
         LAYER metal3 ;
         RECT  19.8975 44.2025 20.0325 44.3375 ;
         LAYER metal3 ;
         RECT  19.8975 38.8225 20.0325 38.9575 ;
         LAYER metal3 ;
         RECT  9.46 -0.0675 9.595 0.0675 ;
         LAYER metal3 ;
         RECT  9.46 9.8325 9.595 9.9675 ;
         LAYER metal3 ;
         RECT  19.8975 41.5125 20.0325 41.6475 ;
         LAYER metal3 ;
         RECT  19.8975 25.3725 20.0325 25.5075 ;
         LAYER metal3 ;
         RECT  23.6175 20.165 23.7525 20.235 ;
         LAYER metal3 ;
         RECT  19.8975 19.9925 20.0325 20.1275 ;
         LAYER metal3 ;
         RECT  17.1025 33.4425 17.2375 33.5775 ;
         LAYER metal3 ;
         RECT  17.1025 44.2025 17.2375 44.3375 ;
         LAYER metal3 ;
         RECT  22.0125 19.9925 22.1475 20.1275 ;
         LAYER metal3 ;
         RECT  18.6925 22.6825 18.8275 22.8175 ;
         LAYER metal3 ;
         RECT  22.0125 44.2025 22.1475 44.3375 ;
         LAYER metal3 ;
         RECT  13.89 -0.0675 14.025 0.0675 ;
         LAYER metal3 ;
         RECT  19.8975 36.1325 20.0325 36.2675 ;
         LAYER metal3 ;
         RECT  17.1025 41.5125 17.2375 41.6475 ;
         LAYER metal3 ;
         RECT  0.75 30.9125 0.885 31.0475 ;
         LAYER metal3 ;
         RECT  22.7175 28.0625 22.8525 28.1975 ;
         LAYER metal3 ;
         RECT  18.6925 28.0625 18.8275 28.1975 ;
         LAYER metal3 ;
         RECT  0.75 19.9925 0.885 20.1275 ;
         LAYER metal3 ;
         RECT  11.0325 25.3725 11.1675 25.5075 ;
         LAYER metal3 ;
         RECT  12.56 28.0625 12.695 28.1975 ;
         LAYER metal3 ;
         RECT  17.1025 38.8225 17.2375 38.9575 ;
         LAYER metal3 ;
         RECT  9.46 19.7325 9.595 19.8675 ;
         LAYER metal3 ;
         RECT  23.6175 44.375 23.7525 44.445 ;
         LAYER metal3 ;
         RECT  9.46 14.7825 9.595 14.9175 ;
         LAYER metal3 ;
         RECT  0.75 34.5525 0.885 34.6875 ;
         LAYER metal3 ;
         RECT  12.56 22.6825 12.695 22.8175 ;
         LAYER metal3 ;
         RECT  17.1025 28.0625 17.2375 28.1975 ;
         LAYER metal3 ;
         RECT  19.8975 22.6825 20.0325 22.8175 ;
         LAYER metal3 ;
         RECT  12.56 30.7525 12.695 30.8875 ;
         LAYER metal3 ;
         RECT  21.34 10.5575 21.41 10.6925 ;
         LAYER metal3 ;
         RECT  22.7175 33.4425 22.8525 33.5775 ;
         LAYER metal3 ;
         RECT  12.56 33.4425 12.695 33.5775 ;
         LAYER metal3 ;
         RECT  22.7175 19.9925 22.8525 20.1275 ;
         LAYER metal3 ;
         RECT  22.7175 41.5125 22.8525 41.6475 ;
         LAYER metal3 ;
         RECT  16.75 -0.0675 16.885 0.0675 ;
         LAYER metal3 ;
         RECT  11.0325 22.6825 11.1675 22.8175 ;
         LAYER metal3 ;
         RECT  19.8975 28.0625 20.0325 28.1975 ;
         LAYER metal3 ;
         RECT  2.125 19.9925 2.26 20.1275 ;
         LAYER metal3 ;
         RECT  17.1025 30.7525 17.2375 30.8875 ;
         LAYER metal3 ;
         RECT  18.6925 38.8225 18.8275 38.9575 ;
         LAYER metal3 ;
         RECT  12.56 36.1325 12.695 36.2675 ;
         LAYER metal3 ;
         RECT  17.1025 36.1325 17.2375 36.2675 ;
         LAYER metal3 ;
         RECT  11.0325 28.0625 11.1675 28.1975 ;
         LAYER metal3 ;
         RECT  11.0325 36.1325 11.1675 36.2675 ;
         LAYER metal3 ;
         RECT  19.7025 44.375 19.8375 44.445 ;
         LAYER metal3 ;
         RECT  18.6925 25.3725 18.8275 25.5075 ;
         LAYER metal3 ;
         RECT  8.17 41.5825 8.305 41.7175 ;
         LAYER metal3 ;
         RECT  20.6025 19.9925 20.7375 20.1275 ;
         LAYER metal3 ;
         RECT  0.75 23.6325 0.885 23.7675 ;
         LAYER metal3 ;
         RECT  2.125 34.5525 2.26 34.6875 ;
         LAYER metal3 ;
         RECT  22.7175 38.8225 22.8525 38.9575 ;
         LAYER metal3 ;
         RECT  18.6925 36.1325 18.8275 36.2675 ;
         LAYER metal3 ;
         RECT  -0.0675 -0.0675 0.0675 0.0675 ;
         LAYER metal3 ;
         RECT  8.17 36.6325 8.305 36.7675 ;
         LAYER metal3 ;
         RECT  2.125 23.6325 2.26 23.7675 ;
         LAYER metal3 ;
         RECT  -0.0675 4.8825 0.0675 5.0175 ;
         LAYER metal3 ;
         RECT  18.6925 41.5125 18.8275 41.6475 ;
         LAYER metal3 ;
         RECT  0.75 27.2725 0.885 27.4075 ;
         LAYER metal3 ;
         RECT  11.0325 33.4425 11.1675 33.5775 ;
         LAYER metal3 ;
         RECT  22.045 17.3275 22.115 17.4625 ;
         LAYER metal3 ;
         RECT  22.7175 22.6825 22.8525 22.8175 ;
         LAYER metal3 ;
         RECT  19.7025 20.165 19.8375 20.235 ;
         LAYER metal3 ;
         RECT  17.1025 25.3725 17.2375 25.5075 ;
         LAYER metal3 ;
         RECT  8.17 46.5325 8.305 46.6675 ;
         LAYER metal3 ;
         RECT  2.125 30.9125 2.26 31.0475 ;
         LAYER metal3 ;
         RECT  12.56 25.3725 12.695 25.5075 ;
         LAYER metal3 ;
         RECT  11.0325 30.7525 11.1675 30.8875 ;
         LAYER metal3 ;
         RECT  19.8975 33.4425 20.0325 33.5775 ;
         LAYER metal3 ;
         RECT  22.7175 25.3725 22.8525 25.5075 ;
         LAYER metal3 ;
         RECT  9.46 4.8825 9.595 5.0175 ;
         LAYER metal3 ;
         RECT  2.125 27.2725 2.26 27.4075 ;
         LAYER metal3 ;
         RECT  22.7175 44.2025 22.8525 44.3375 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  21.53 23.3975 21.595 23.5325 ;
      RECT  22.045 23.3975 22.115 23.5325 ;
      RECT  21.425 23.2325 21.595 23.2975 ;
      RECT  21.285 22.8575 22.17 22.9225 ;
      RECT  21.34 23.8625 21.41 24.0625 ;
      RECT  22.045 23.8625 22.11 23.9975 ;
      RECT  21.5975 23.0075 21.6625 23.1425 ;
      RECT  21.78 23.0075 21.845 23.1425 ;
      RECT  22.045 23.3975 22.11 23.5325 ;
      RECT  22.0125 22.7175 22.1475 22.7825 ;
      RECT  21.7725 23.5975 21.9075 23.6625 ;
      RECT  21.995 22.86 22.0475 22.9225 ;
      RECT  21.5475 23.7475 21.6825 23.8125 ;
      RECT  21.425 23.0075 21.495 23.2975 ;
      RECT  21.53 23.2325 21.595 23.9725 ;
      RECT  22.045 23.8625 22.115 24.0625 ;
      RECT  21.965 23.0075 22.03 23.1425 ;
      RECT  21.29 22.86 21.3425 22.9225 ;
      RECT  21.285 24.0625 22.17 24.1275 ;
      RECT  21.3425 23.5 21.4075 23.635 ;
      RECT  21.66 22.7175 21.795 22.7825 ;
      RECT  21.965 23.0075 22.035 23.2975 ;
      RECT  21.6425 22.8575 21.7775 22.9225 ;
      RECT  21.345 23.8625 21.41 23.9975 ;
      RECT  21.86 23.2325 22.035 23.2975 ;
      RECT  21.86 23.8625 21.925 23.9975 ;
      RECT  21.285 22.7175 22.17 22.7825 ;
      RECT  22.0475 23.5 22.1125 23.635 ;
      RECT  21.34 23.3975 21.41 23.5325 ;
      RECT  21.61 23.0075 21.675 23.1425 ;
      RECT  21.86 23.3975 21.925 23.5325 ;
      RECT  21.7925 23.0075 21.8575 23.1425 ;
      RECT  21.345 23.3975 21.41 23.5325 ;
      RECT  21.53 23.8625 21.595 23.9975 ;
      RECT  21.86 23.2325 21.925 23.8625 ;
      RECT  21.3075 22.7175 21.4425 22.7825 ;
      RECT  21.425 23.0075 21.49 23.1425 ;
      RECT  21.53 24.7925 21.595 24.6575 ;
      RECT  22.045 24.7925 22.115 24.6575 ;
      RECT  21.425 24.9575 21.595 24.8925 ;
      RECT  21.285 25.3325 22.17 25.2675 ;
      RECT  21.34 24.3275 21.41 24.1275 ;
      RECT  22.045 24.3275 22.11 24.1925 ;
      RECT  21.5975 25.1825 21.6625 25.0475 ;
      RECT  21.78 25.1825 21.845 25.0475 ;
      RECT  22.045 24.7925 22.11 24.6575 ;
      RECT  22.0125 25.4725 22.1475 25.4075 ;
      RECT  21.7725 24.5925 21.9075 24.5275 ;
      RECT  21.995 25.33 22.0475 25.2675 ;
      RECT  21.5475 24.4425 21.6825 24.3775 ;
      RECT  21.425 25.1825 21.495 24.8925 ;
      RECT  21.53 24.9575 21.595 24.2175 ;
      RECT  22.045 24.3275 22.115 24.1275 ;
      RECT  21.965 25.1825 22.03 25.0475 ;
      RECT  21.29 25.33 21.3425 25.2675 ;
      RECT  21.285 24.1275 22.17 24.0625 ;
      RECT  21.3425 24.69 21.4075 24.555 ;
      RECT  21.66 25.4725 21.795 25.4075 ;
      RECT  21.965 25.1825 22.035 24.8925 ;
      RECT  21.6425 25.3325 21.7775 25.2675 ;
      RECT  21.345 24.3275 21.41 24.1925 ;
      RECT  21.86 24.9575 22.035 24.8925 ;
      RECT  21.86 24.3275 21.925 24.1925 ;
      RECT  21.285 25.4725 22.17 25.4075 ;
      RECT  22.0475 24.69 22.1125 24.555 ;
      RECT  21.34 24.7925 21.41 24.6575 ;
      RECT  21.61 25.1825 21.675 25.0475 ;
      RECT  21.86 24.7925 21.925 24.6575 ;
      RECT  21.7925 25.1825 21.8575 25.0475 ;
      RECT  21.345 24.7925 21.41 24.6575 ;
      RECT  21.53 24.3275 21.595 24.1925 ;
      RECT  21.86 24.9575 21.925 24.3275 ;
      RECT  21.3075 25.4725 21.4425 25.4075 ;
      RECT  21.425 25.1825 21.49 25.0475 ;
      RECT  21.53 26.0875 21.595 26.2225 ;
      RECT  22.045 26.0875 22.115 26.2225 ;
      RECT  21.425 25.9225 21.595 25.9875 ;
      RECT  21.285 25.5475 22.17 25.6125 ;
      RECT  21.34 26.5525 21.41 26.7525 ;
      RECT  22.045 26.5525 22.11 26.6875 ;
      RECT  21.5975 25.6975 21.6625 25.8325 ;
      RECT  21.78 25.6975 21.845 25.8325 ;
      RECT  22.045 26.0875 22.11 26.2225 ;
      RECT  22.0125 25.4075 22.1475 25.4725 ;
      RECT  21.7725 26.2875 21.9075 26.3525 ;
      RECT  21.995 25.55 22.0475 25.6125 ;
      RECT  21.5475 26.4375 21.6825 26.5025 ;
      RECT  21.425 25.6975 21.495 25.9875 ;
      RECT  21.53 25.9225 21.595 26.6625 ;
      RECT  22.045 26.5525 22.115 26.7525 ;
      RECT  21.965 25.6975 22.03 25.8325 ;
      RECT  21.29 25.55 21.3425 25.6125 ;
      RECT  21.285 26.7525 22.17 26.8175 ;
      RECT  21.3425 26.19 21.4075 26.325 ;
      RECT  21.66 25.4075 21.795 25.4725 ;
      RECT  21.965 25.6975 22.035 25.9875 ;
      RECT  21.6425 25.5475 21.7775 25.6125 ;
      RECT  21.345 26.5525 21.41 26.6875 ;
      RECT  21.86 25.9225 22.035 25.9875 ;
      RECT  21.86 26.5525 21.925 26.6875 ;
      RECT  21.285 25.4075 22.17 25.4725 ;
      RECT  22.0475 26.19 22.1125 26.325 ;
      RECT  21.34 26.0875 21.41 26.2225 ;
      RECT  21.61 25.6975 21.675 25.8325 ;
      RECT  21.86 26.0875 21.925 26.2225 ;
      RECT  21.7925 25.6975 21.8575 25.8325 ;
      RECT  21.345 26.0875 21.41 26.2225 ;
      RECT  21.53 26.5525 21.595 26.6875 ;
      RECT  21.86 25.9225 21.925 26.5525 ;
      RECT  21.3075 25.4075 21.4425 25.4725 ;
      RECT  21.425 25.6975 21.49 25.8325 ;
      RECT  21.53 27.4825 21.595 27.3475 ;
      RECT  22.045 27.4825 22.115 27.3475 ;
      RECT  21.425 27.6475 21.595 27.5825 ;
      RECT  21.285 28.0225 22.17 27.9575 ;
      RECT  21.34 27.0175 21.41 26.8175 ;
      RECT  22.045 27.0175 22.11 26.8825 ;
      RECT  21.5975 27.8725 21.6625 27.7375 ;
      RECT  21.78 27.8725 21.845 27.7375 ;
      RECT  22.045 27.4825 22.11 27.3475 ;
      RECT  22.0125 28.1625 22.1475 28.0975 ;
      RECT  21.7725 27.2825 21.9075 27.2175 ;
      RECT  21.995 28.02 22.0475 27.9575 ;
      RECT  21.5475 27.1325 21.6825 27.0675 ;
      RECT  21.425 27.8725 21.495 27.5825 ;
      RECT  21.53 27.6475 21.595 26.9075 ;
      RECT  22.045 27.0175 22.115 26.8175 ;
      RECT  21.965 27.8725 22.03 27.7375 ;
      RECT  21.29 28.02 21.3425 27.9575 ;
      RECT  21.285 26.8175 22.17 26.7525 ;
      RECT  21.3425 27.38 21.4075 27.245 ;
      RECT  21.66 28.1625 21.795 28.0975 ;
      RECT  21.965 27.8725 22.035 27.5825 ;
      RECT  21.6425 28.0225 21.7775 27.9575 ;
      RECT  21.345 27.0175 21.41 26.8825 ;
      RECT  21.86 27.6475 22.035 27.5825 ;
      RECT  21.86 27.0175 21.925 26.8825 ;
      RECT  21.285 28.1625 22.17 28.0975 ;
      RECT  22.0475 27.38 22.1125 27.245 ;
      RECT  21.34 27.4825 21.41 27.3475 ;
      RECT  21.61 27.8725 21.675 27.7375 ;
      RECT  21.86 27.4825 21.925 27.3475 ;
      RECT  21.7925 27.8725 21.8575 27.7375 ;
      RECT  21.345 27.4825 21.41 27.3475 ;
      RECT  21.53 27.0175 21.595 26.8825 ;
      RECT  21.86 27.6475 21.925 27.0175 ;
      RECT  21.3075 28.1625 21.4425 28.0975 ;
      RECT  21.425 27.8725 21.49 27.7375 ;
      RECT  21.53 28.7775 21.595 28.9125 ;
      RECT  22.045 28.7775 22.115 28.9125 ;
      RECT  21.425 28.6125 21.595 28.6775 ;
      RECT  21.285 28.2375 22.17 28.3025 ;
      RECT  21.34 29.2425 21.41 29.4425 ;
      RECT  22.045 29.2425 22.11 29.3775 ;
      RECT  21.5975 28.3875 21.6625 28.5225 ;
      RECT  21.78 28.3875 21.845 28.5225 ;
      RECT  22.045 28.7775 22.11 28.9125 ;
      RECT  22.0125 28.0975 22.1475 28.1625 ;
      RECT  21.7725 28.9775 21.9075 29.0425 ;
      RECT  21.995 28.24 22.0475 28.3025 ;
      RECT  21.5475 29.1275 21.6825 29.1925 ;
      RECT  21.425 28.3875 21.495 28.6775 ;
      RECT  21.53 28.6125 21.595 29.3525 ;
      RECT  22.045 29.2425 22.115 29.4425 ;
      RECT  21.965 28.3875 22.03 28.5225 ;
      RECT  21.29 28.24 21.3425 28.3025 ;
      RECT  21.285 29.4425 22.17 29.5075 ;
      RECT  21.3425 28.88 21.4075 29.015 ;
      RECT  21.66 28.0975 21.795 28.1625 ;
      RECT  21.965 28.3875 22.035 28.6775 ;
      RECT  21.6425 28.2375 21.7775 28.3025 ;
      RECT  21.345 29.2425 21.41 29.3775 ;
      RECT  21.86 28.6125 22.035 28.6775 ;
      RECT  21.86 29.2425 21.925 29.3775 ;
      RECT  21.285 28.0975 22.17 28.1625 ;
      RECT  22.0475 28.88 22.1125 29.015 ;
      RECT  21.34 28.7775 21.41 28.9125 ;
      RECT  21.61 28.3875 21.675 28.5225 ;
      RECT  21.86 28.7775 21.925 28.9125 ;
      RECT  21.7925 28.3875 21.8575 28.5225 ;
      RECT  21.345 28.7775 21.41 28.9125 ;
      RECT  21.53 29.2425 21.595 29.3775 ;
      RECT  21.86 28.6125 21.925 29.2425 ;
      RECT  21.3075 28.0975 21.4425 28.1625 ;
      RECT  21.425 28.3875 21.49 28.5225 ;
      RECT  21.53 30.1725 21.595 30.0375 ;
      RECT  22.045 30.1725 22.115 30.0375 ;
      RECT  21.425 30.3375 21.595 30.2725 ;
      RECT  21.285 30.7125 22.17 30.6475 ;
      RECT  21.34 29.7075 21.41 29.5075 ;
      RECT  22.045 29.7075 22.11 29.5725 ;
      RECT  21.5975 30.5625 21.6625 30.4275 ;
      RECT  21.78 30.5625 21.845 30.4275 ;
      RECT  22.045 30.1725 22.11 30.0375 ;
      RECT  22.0125 30.8525 22.1475 30.7875 ;
      RECT  21.7725 29.9725 21.9075 29.9075 ;
      RECT  21.995 30.71 22.0475 30.6475 ;
      RECT  21.5475 29.8225 21.6825 29.7575 ;
      RECT  21.425 30.5625 21.495 30.2725 ;
      RECT  21.53 30.3375 21.595 29.5975 ;
      RECT  22.045 29.7075 22.115 29.5075 ;
      RECT  21.965 30.5625 22.03 30.4275 ;
      RECT  21.29 30.71 21.3425 30.6475 ;
      RECT  21.285 29.5075 22.17 29.4425 ;
      RECT  21.3425 30.07 21.4075 29.935 ;
      RECT  21.66 30.8525 21.795 30.7875 ;
      RECT  21.965 30.5625 22.035 30.2725 ;
      RECT  21.6425 30.7125 21.7775 30.6475 ;
      RECT  21.345 29.7075 21.41 29.5725 ;
      RECT  21.86 30.3375 22.035 30.2725 ;
      RECT  21.86 29.7075 21.925 29.5725 ;
      RECT  21.285 30.8525 22.17 30.7875 ;
      RECT  22.0475 30.07 22.1125 29.935 ;
      RECT  21.34 30.1725 21.41 30.0375 ;
      RECT  21.61 30.5625 21.675 30.4275 ;
      RECT  21.86 30.1725 21.925 30.0375 ;
      RECT  21.7925 30.5625 21.8575 30.4275 ;
      RECT  21.345 30.1725 21.41 30.0375 ;
      RECT  21.53 29.7075 21.595 29.5725 ;
      RECT  21.86 30.3375 21.925 29.7075 ;
      RECT  21.3075 30.8525 21.4425 30.7875 ;
      RECT  21.425 30.5625 21.49 30.4275 ;
      RECT  21.53 31.4675 21.595 31.6025 ;
      RECT  22.045 31.4675 22.115 31.6025 ;
      RECT  21.425 31.3025 21.595 31.3675 ;
      RECT  21.285 30.9275 22.17 30.9925 ;
      RECT  21.34 31.9325 21.41 32.1325 ;
      RECT  22.045 31.9325 22.11 32.0675 ;
      RECT  21.5975 31.0775 21.6625 31.2125 ;
      RECT  21.78 31.0775 21.845 31.2125 ;
      RECT  22.045 31.4675 22.11 31.6025 ;
      RECT  22.0125 30.7875 22.1475 30.8525 ;
      RECT  21.7725 31.6675 21.9075 31.7325 ;
      RECT  21.995 30.93 22.0475 30.9925 ;
      RECT  21.5475 31.8175 21.6825 31.8825 ;
      RECT  21.425 31.0775 21.495 31.3675 ;
      RECT  21.53 31.3025 21.595 32.0425 ;
      RECT  22.045 31.9325 22.115 32.1325 ;
      RECT  21.965 31.0775 22.03 31.2125 ;
      RECT  21.29 30.93 21.3425 30.9925 ;
      RECT  21.285 32.1325 22.17 32.1975 ;
      RECT  21.3425 31.57 21.4075 31.705 ;
      RECT  21.66 30.7875 21.795 30.8525 ;
      RECT  21.965 31.0775 22.035 31.3675 ;
      RECT  21.6425 30.9275 21.7775 30.9925 ;
      RECT  21.345 31.9325 21.41 32.0675 ;
      RECT  21.86 31.3025 22.035 31.3675 ;
      RECT  21.86 31.9325 21.925 32.0675 ;
      RECT  21.285 30.7875 22.17 30.8525 ;
      RECT  22.0475 31.57 22.1125 31.705 ;
      RECT  21.34 31.4675 21.41 31.6025 ;
      RECT  21.61 31.0775 21.675 31.2125 ;
      RECT  21.86 31.4675 21.925 31.6025 ;
      RECT  21.7925 31.0775 21.8575 31.2125 ;
      RECT  21.345 31.4675 21.41 31.6025 ;
      RECT  21.53 31.9325 21.595 32.0675 ;
      RECT  21.86 31.3025 21.925 31.9325 ;
      RECT  21.3075 30.7875 21.4425 30.8525 ;
      RECT  21.425 31.0775 21.49 31.2125 ;
      RECT  21.53 32.8625 21.595 32.7275 ;
      RECT  22.045 32.8625 22.115 32.7275 ;
      RECT  21.425 33.0275 21.595 32.9625 ;
      RECT  21.285 33.4025 22.17 33.3375 ;
      RECT  21.34 32.3975 21.41 32.1975 ;
      RECT  22.045 32.3975 22.11 32.2625 ;
      RECT  21.5975 33.2525 21.6625 33.1175 ;
      RECT  21.78 33.2525 21.845 33.1175 ;
      RECT  22.045 32.8625 22.11 32.7275 ;
      RECT  22.0125 33.5425 22.1475 33.4775 ;
      RECT  21.7725 32.6625 21.9075 32.5975 ;
      RECT  21.995 33.4 22.0475 33.3375 ;
      RECT  21.5475 32.5125 21.6825 32.4475 ;
      RECT  21.425 33.2525 21.495 32.9625 ;
      RECT  21.53 33.0275 21.595 32.2875 ;
      RECT  22.045 32.3975 22.115 32.1975 ;
      RECT  21.965 33.2525 22.03 33.1175 ;
      RECT  21.29 33.4 21.3425 33.3375 ;
      RECT  21.285 32.1975 22.17 32.1325 ;
      RECT  21.3425 32.76 21.4075 32.625 ;
      RECT  21.66 33.5425 21.795 33.4775 ;
      RECT  21.965 33.2525 22.035 32.9625 ;
      RECT  21.6425 33.4025 21.7775 33.3375 ;
      RECT  21.345 32.3975 21.41 32.2625 ;
      RECT  21.86 33.0275 22.035 32.9625 ;
      RECT  21.86 32.3975 21.925 32.2625 ;
      RECT  21.285 33.5425 22.17 33.4775 ;
      RECT  22.0475 32.76 22.1125 32.625 ;
      RECT  21.34 32.8625 21.41 32.7275 ;
      RECT  21.61 33.2525 21.675 33.1175 ;
      RECT  21.86 32.8625 21.925 32.7275 ;
      RECT  21.7925 33.2525 21.8575 33.1175 ;
      RECT  21.345 32.8625 21.41 32.7275 ;
      RECT  21.53 32.3975 21.595 32.2625 ;
      RECT  21.86 33.0275 21.925 32.3975 ;
      RECT  21.3075 33.5425 21.4425 33.4775 ;
      RECT  21.425 33.2525 21.49 33.1175 ;
      RECT  21.53 34.1575 21.595 34.2925 ;
      RECT  22.045 34.1575 22.115 34.2925 ;
      RECT  21.425 33.9925 21.595 34.0575 ;
      RECT  21.285 33.6175 22.17 33.6825 ;
      RECT  21.34 34.6225 21.41 34.8225 ;
      RECT  22.045 34.6225 22.11 34.7575 ;
      RECT  21.5975 33.7675 21.6625 33.9025 ;
      RECT  21.78 33.7675 21.845 33.9025 ;
      RECT  22.045 34.1575 22.11 34.2925 ;
      RECT  22.0125 33.4775 22.1475 33.5425 ;
      RECT  21.7725 34.3575 21.9075 34.4225 ;
      RECT  21.995 33.62 22.0475 33.6825 ;
      RECT  21.5475 34.5075 21.6825 34.5725 ;
      RECT  21.425 33.7675 21.495 34.0575 ;
      RECT  21.53 33.9925 21.595 34.7325 ;
      RECT  22.045 34.6225 22.115 34.8225 ;
      RECT  21.965 33.7675 22.03 33.9025 ;
      RECT  21.29 33.62 21.3425 33.6825 ;
      RECT  21.285 34.8225 22.17 34.8875 ;
      RECT  21.3425 34.26 21.4075 34.395 ;
      RECT  21.66 33.4775 21.795 33.5425 ;
      RECT  21.965 33.7675 22.035 34.0575 ;
      RECT  21.6425 33.6175 21.7775 33.6825 ;
      RECT  21.345 34.6225 21.41 34.7575 ;
      RECT  21.86 33.9925 22.035 34.0575 ;
      RECT  21.86 34.6225 21.925 34.7575 ;
      RECT  21.285 33.4775 22.17 33.5425 ;
      RECT  22.0475 34.26 22.1125 34.395 ;
      RECT  21.34 34.1575 21.41 34.2925 ;
      RECT  21.61 33.7675 21.675 33.9025 ;
      RECT  21.86 34.1575 21.925 34.2925 ;
      RECT  21.7925 33.7675 21.8575 33.9025 ;
      RECT  21.345 34.1575 21.41 34.2925 ;
      RECT  21.53 34.6225 21.595 34.7575 ;
      RECT  21.86 33.9925 21.925 34.6225 ;
      RECT  21.3075 33.4775 21.4425 33.5425 ;
      RECT  21.425 33.7675 21.49 33.9025 ;
      RECT  21.53 35.5525 21.595 35.4175 ;
      RECT  22.045 35.5525 22.115 35.4175 ;
      RECT  21.425 35.7175 21.595 35.6525 ;
      RECT  21.285 36.0925 22.17 36.0275 ;
      RECT  21.34 35.0875 21.41 34.8875 ;
      RECT  22.045 35.0875 22.11 34.9525 ;
      RECT  21.5975 35.9425 21.6625 35.8075 ;
      RECT  21.78 35.9425 21.845 35.8075 ;
      RECT  22.045 35.5525 22.11 35.4175 ;
      RECT  22.0125 36.2325 22.1475 36.1675 ;
      RECT  21.7725 35.3525 21.9075 35.2875 ;
      RECT  21.995 36.09 22.0475 36.0275 ;
      RECT  21.5475 35.2025 21.6825 35.1375 ;
      RECT  21.425 35.9425 21.495 35.6525 ;
      RECT  21.53 35.7175 21.595 34.9775 ;
      RECT  22.045 35.0875 22.115 34.8875 ;
      RECT  21.965 35.9425 22.03 35.8075 ;
      RECT  21.29 36.09 21.3425 36.0275 ;
      RECT  21.285 34.8875 22.17 34.8225 ;
      RECT  21.3425 35.45 21.4075 35.315 ;
      RECT  21.66 36.2325 21.795 36.1675 ;
      RECT  21.965 35.9425 22.035 35.6525 ;
      RECT  21.6425 36.0925 21.7775 36.0275 ;
      RECT  21.345 35.0875 21.41 34.9525 ;
      RECT  21.86 35.7175 22.035 35.6525 ;
      RECT  21.86 35.0875 21.925 34.9525 ;
      RECT  21.285 36.2325 22.17 36.1675 ;
      RECT  22.0475 35.45 22.1125 35.315 ;
      RECT  21.34 35.5525 21.41 35.4175 ;
      RECT  21.61 35.9425 21.675 35.8075 ;
      RECT  21.86 35.5525 21.925 35.4175 ;
      RECT  21.7925 35.9425 21.8575 35.8075 ;
      RECT  21.345 35.5525 21.41 35.4175 ;
      RECT  21.53 35.0875 21.595 34.9525 ;
      RECT  21.86 35.7175 21.925 35.0875 ;
      RECT  21.3075 36.2325 21.4425 36.1675 ;
      RECT  21.425 35.9425 21.49 35.8075 ;
      RECT  21.53 36.8475 21.595 36.9825 ;
      RECT  22.045 36.8475 22.115 36.9825 ;
      RECT  21.425 36.6825 21.595 36.7475 ;
      RECT  21.285 36.3075 22.17 36.3725 ;
      RECT  21.34 37.3125 21.41 37.5125 ;
      RECT  22.045 37.3125 22.11 37.4475 ;
      RECT  21.5975 36.4575 21.6625 36.5925 ;
      RECT  21.78 36.4575 21.845 36.5925 ;
      RECT  22.045 36.8475 22.11 36.9825 ;
      RECT  22.0125 36.1675 22.1475 36.2325 ;
      RECT  21.7725 37.0475 21.9075 37.1125 ;
      RECT  21.995 36.31 22.0475 36.3725 ;
      RECT  21.5475 37.1975 21.6825 37.2625 ;
      RECT  21.425 36.4575 21.495 36.7475 ;
      RECT  21.53 36.6825 21.595 37.4225 ;
      RECT  22.045 37.3125 22.115 37.5125 ;
      RECT  21.965 36.4575 22.03 36.5925 ;
      RECT  21.29 36.31 21.3425 36.3725 ;
      RECT  21.285 37.5125 22.17 37.5775 ;
      RECT  21.3425 36.95 21.4075 37.085 ;
      RECT  21.66 36.1675 21.795 36.2325 ;
      RECT  21.965 36.4575 22.035 36.7475 ;
      RECT  21.6425 36.3075 21.7775 36.3725 ;
      RECT  21.345 37.3125 21.41 37.4475 ;
      RECT  21.86 36.6825 22.035 36.7475 ;
      RECT  21.86 37.3125 21.925 37.4475 ;
      RECT  21.285 36.1675 22.17 36.2325 ;
      RECT  22.0475 36.95 22.1125 37.085 ;
      RECT  21.34 36.8475 21.41 36.9825 ;
      RECT  21.61 36.4575 21.675 36.5925 ;
      RECT  21.86 36.8475 21.925 36.9825 ;
      RECT  21.7925 36.4575 21.8575 36.5925 ;
      RECT  21.345 36.8475 21.41 36.9825 ;
      RECT  21.53 37.3125 21.595 37.4475 ;
      RECT  21.86 36.6825 21.925 37.3125 ;
      RECT  21.3075 36.1675 21.4425 36.2325 ;
      RECT  21.425 36.4575 21.49 36.5925 ;
      RECT  21.53 38.2425 21.595 38.1075 ;
      RECT  22.045 38.2425 22.115 38.1075 ;
      RECT  21.425 38.4075 21.595 38.3425 ;
      RECT  21.285 38.7825 22.17 38.7175 ;
      RECT  21.34 37.7775 21.41 37.5775 ;
      RECT  22.045 37.7775 22.11 37.6425 ;
      RECT  21.5975 38.6325 21.6625 38.4975 ;
      RECT  21.78 38.6325 21.845 38.4975 ;
      RECT  22.045 38.2425 22.11 38.1075 ;
      RECT  22.0125 38.9225 22.1475 38.8575 ;
      RECT  21.7725 38.0425 21.9075 37.9775 ;
      RECT  21.995 38.78 22.0475 38.7175 ;
      RECT  21.5475 37.8925 21.6825 37.8275 ;
      RECT  21.425 38.6325 21.495 38.3425 ;
      RECT  21.53 38.4075 21.595 37.6675 ;
      RECT  22.045 37.7775 22.115 37.5775 ;
      RECT  21.965 38.6325 22.03 38.4975 ;
      RECT  21.29 38.78 21.3425 38.7175 ;
      RECT  21.285 37.5775 22.17 37.5125 ;
      RECT  21.3425 38.14 21.4075 38.005 ;
      RECT  21.66 38.9225 21.795 38.8575 ;
      RECT  21.965 38.6325 22.035 38.3425 ;
      RECT  21.6425 38.7825 21.7775 38.7175 ;
      RECT  21.345 37.7775 21.41 37.6425 ;
      RECT  21.86 38.4075 22.035 38.3425 ;
      RECT  21.86 37.7775 21.925 37.6425 ;
      RECT  21.285 38.9225 22.17 38.8575 ;
      RECT  22.0475 38.14 22.1125 38.005 ;
      RECT  21.34 38.2425 21.41 38.1075 ;
      RECT  21.61 38.6325 21.675 38.4975 ;
      RECT  21.86 38.2425 21.925 38.1075 ;
      RECT  21.7925 38.6325 21.8575 38.4975 ;
      RECT  21.345 38.2425 21.41 38.1075 ;
      RECT  21.53 37.7775 21.595 37.6425 ;
      RECT  21.86 38.4075 21.925 37.7775 ;
      RECT  21.3075 38.9225 21.4425 38.8575 ;
      RECT  21.425 38.6325 21.49 38.4975 ;
      RECT  21.53 39.5375 21.595 39.6725 ;
      RECT  22.045 39.5375 22.115 39.6725 ;
      RECT  21.425 39.3725 21.595 39.4375 ;
      RECT  21.285 38.9975 22.17 39.0625 ;
      RECT  21.34 40.0025 21.41 40.2025 ;
      RECT  22.045 40.0025 22.11 40.1375 ;
      RECT  21.5975 39.1475 21.6625 39.2825 ;
      RECT  21.78 39.1475 21.845 39.2825 ;
      RECT  22.045 39.5375 22.11 39.6725 ;
      RECT  22.0125 38.8575 22.1475 38.9225 ;
      RECT  21.7725 39.7375 21.9075 39.8025 ;
      RECT  21.995 39.0 22.0475 39.0625 ;
      RECT  21.5475 39.8875 21.6825 39.9525 ;
      RECT  21.425 39.1475 21.495 39.4375 ;
      RECT  21.53 39.3725 21.595 40.1125 ;
      RECT  22.045 40.0025 22.115 40.2025 ;
      RECT  21.965 39.1475 22.03 39.2825 ;
      RECT  21.29 39.0 21.3425 39.0625 ;
      RECT  21.285 40.2025 22.17 40.2675 ;
      RECT  21.3425 39.64 21.4075 39.775 ;
      RECT  21.66 38.8575 21.795 38.9225 ;
      RECT  21.965 39.1475 22.035 39.4375 ;
      RECT  21.6425 38.9975 21.7775 39.0625 ;
      RECT  21.345 40.0025 21.41 40.1375 ;
      RECT  21.86 39.3725 22.035 39.4375 ;
      RECT  21.86 40.0025 21.925 40.1375 ;
      RECT  21.285 38.8575 22.17 38.9225 ;
      RECT  22.0475 39.64 22.1125 39.775 ;
      RECT  21.34 39.5375 21.41 39.6725 ;
      RECT  21.61 39.1475 21.675 39.2825 ;
      RECT  21.86 39.5375 21.925 39.6725 ;
      RECT  21.7925 39.1475 21.8575 39.2825 ;
      RECT  21.345 39.5375 21.41 39.6725 ;
      RECT  21.53 40.0025 21.595 40.1375 ;
      RECT  21.86 39.3725 21.925 40.0025 ;
      RECT  21.3075 38.8575 21.4425 38.9225 ;
      RECT  21.425 39.1475 21.49 39.2825 ;
      RECT  21.53 40.9325 21.595 40.7975 ;
      RECT  22.045 40.9325 22.115 40.7975 ;
      RECT  21.425 41.0975 21.595 41.0325 ;
      RECT  21.285 41.4725 22.17 41.4075 ;
      RECT  21.34 40.4675 21.41 40.2675 ;
      RECT  22.045 40.4675 22.11 40.3325 ;
      RECT  21.5975 41.3225 21.6625 41.1875 ;
      RECT  21.78 41.3225 21.845 41.1875 ;
      RECT  22.045 40.9325 22.11 40.7975 ;
      RECT  22.0125 41.6125 22.1475 41.5475 ;
      RECT  21.7725 40.7325 21.9075 40.6675 ;
      RECT  21.995 41.47 22.0475 41.4075 ;
      RECT  21.5475 40.5825 21.6825 40.5175 ;
      RECT  21.425 41.3225 21.495 41.0325 ;
      RECT  21.53 41.0975 21.595 40.3575 ;
      RECT  22.045 40.4675 22.115 40.2675 ;
      RECT  21.965 41.3225 22.03 41.1875 ;
      RECT  21.29 41.47 21.3425 41.4075 ;
      RECT  21.285 40.2675 22.17 40.2025 ;
      RECT  21.3425 40.83 21.4075 40.695 ;
      RECT  21.66 41.6125 21.795 41.5475 ;
      RECT  21.965 41.3225 22.035 41.0325 ;
      RECT  21.6425 41.4725 21.7775 41.4075 ;
      RECT  21.345 40.4675 21.41 40.3325 ;
      RECT  21.86 41.0975 22.035 41.0325 ;
      RECT  21.86 40.4675 21.925 40.3325 ;
      RECT  21.285 41.6125 22.17 41.5475 ;
      RECT  22.0475 40.83 22.1125 40.695 ;
      RECT  21.34 40.9325 21.41 40.7975 ;
      RECT  21.61 41.3225 21.675 41.1875 ;
      RECT  21.86 40.9325 21.925 40.7975 ;
      RECT  21.7925 41.3225 21.8575 41.1875 ;
      RECT  21.345 40.9325 21.41 40.7975 ;
      RECT  21.53 40.4675 21.595 40.3325 ;
      RECT  21.86 41.0975 21.925 40.4675 ;
      RECT  21.3075 41.6125 21.4425 41.5475 ;
      RECT  21.425 41.3225 21.49 41.1875 ;
      RECT  21.53 42.2275 21.595 42.3625 ;
      RECT  22.045 42.2275 22.115 42.3625 ;
      RECT  21.425 42.0625 21.595 42.1275 ;
      RECT  21.285 41.6875 22.17 41.7525 ;
      RECT  21.34 42.6925 21.41 42.8925 ;
      RECT  22.045 42.6925 22.11 42.8275 ;
      RECT  21.5975 41.8375 21.6625 41.9725 ;
      RECT  21.78 41.8375 21.845 41.9725 ;
      RECT  22.045 42.2275 22.11 42.3625 ;
      RECT  22.0125 41.5475 22.1475 41.6125 ;
      RECT  21.7725 42.4275 21.9075 42.4925 ;
      RECT  21.995 41.69 22.0475 41.7525 ;
      RECT  21.5475 42.5775 21.6825 42.6425 ;
      RECT  21.425 41.8375 21.495 42.1275 ;
      RECT  21.53 42.0625 21.595 42.8025 ;
      RECT  22.045 42.6925 22.115 42.8925 ;
      RECT  21.965 41.8375 22.03 41.9725 ;
      RECT  21.29 41.69 21.3425 41.7525 ;
      RECT  21.285 42.8925 22.17 42.9575 ;
      RECT  21.3425 42.33 21.4075 42.465 ;
      RECT  21.66 41.5475 21.795 41.6125 ;
      RECT  21.965 41.8375 22.035 42.1275 ;
      RECT  21.6425 41.6875 21.7775 41.7525 ;
      RECT  21.345 42.6925 21.41 42.8275 ;
      RECT  21.86 42.0625 22.035 42.1275 ;
      RECT  21.86 42.6925 21.925 42.8275 ;
      RECT  21.285 41.5475 22.17 41.6125 ;
      RECT  22.0475 42.33 22.1125 42.465 ;
      RECT  21.34 42.2275 21.41 42.3625 ;
      RECT  21.61 41.8375 21.675 41.9725 ;
      RECT  21.86 42.2275 21.925 42.3625 ;
      RECT  21.7925 41.8375 21.8575 41.9725 ;
      RECT  21.345 42.2275 21.41 42.3625 ;
      RECT  21.53 42.6925 21.595 42.8275 ;
      RECT  21.86 42.0625 21.925 42.6925 ;
      RECT  21.3075 41.5475 21.4425 41.6125 ;
      RECT  21.425 41.8375 21.49 41.9725 ;
      RECT  21.53 43.6225 21.595 43.4875 ;
      RECT  22.045 43.6225 22.115 43.4875 ;
      RECT  21.425 43.7875 21.595 43.7225 ;
      RECT  21.285 44.1625 22.17 44.0975 ;
      RECT  21.34 43.1575 21.41 42.9575 ;
      RECT  22.045 43.1575 22.11 43.0225 ;
      RECT  21.5975 44.0125 21.6625 43.8775 ;
      RECT  21.78 44.0125 21.845 43.8775 ;
      RECT  22.045 43.6225 22.11 43.4875 ;
      RECT  22.0125 44.3025 22.1475 44.2375 ;
      RECT  21.7725 43.4225 21.9075 43.3575 ;
      RECT  21.995 44.16 22.0475 44.0975 ;
      RECT  21.5475 43.2725 21.6825 43.2075 ;
      RECT  21.425 44.0125 21.495 43.7225 ;
      RECT  21.53 43.7875 21.595 43.0475 ;
      RECT  22.045 43.1575 22.115 42.9575 ;
      RECT  21.965 44.0125 22.03 43.8775 ;
      RECT  21.29 44.16 21.3425 44.0975 ;
      RECT  21.285 42.9575 22.17 42.8925 ;
      RECT  21.3425 43.52 21.4075 43.385 ;
      RECT  21.66 44.3025 21.795 44.2375 ;
      RECT  21.965 44.0125 22.035 43.7225 ;
      RECT  21.6425 44.1625 21.7775 44.0975 ;
      RECT  21.345 43.1575 21.41 43.0225 ;
      RECT  21.86 43.7875 22.035 43.7225 ;
      RECT  21.86 43.1575 21.925 43.0225 ;
      RECT  21.285 44.3025 22.17 44.2375 ;
      RECT  22.0475 43.52 22.1125 43.385 ;
      RECT  21.34 43.6225 21.41 43.4875 ;
      RECT  21.61 44.0125 21.675 43.8775 ;
      RECT  21.86 43.6225 21.925 43.4875 ;
      RECT  21.7925 44.0125 21.8575 43.8775 ;
      RECT  21.345 43.6225 21.41 43.4875 ;
      RECT  21.53 43.1575 21.595 43.0225 ;
      RECT  21.86 43.7875 21.925 43.1575 ;
      RECT  21.3075 44.3025 21.4425 44.2375 ;
      RECT  21.425 44.0125 21.49 43.8775 ;
      RECT  22.235 23.3975 22.3 23.5325 ;
      RECT  22.75 23.3975 22.82 23.5325 ;
      RECT  22.13 23.2325 22.3 23.2975 ;
      RECT  21.99 22.8575 22.875 22.9225 ;
      RECT  22.045 23.8625 22.115 24.0625 ;
      RECT  22.75 23.8625 22.815 23.9975 ;
      RECT  22.3025 23.0075 22.3675 23.1425 ;
      RECT  22.485 23.0075 22.55 23.1425 ;
      RECT  22.75 23.3975 22.815 23.5325 ;
      RECT  22.7175 22.7175 22.8525 22.7825 ;
      RECT  22.4775 23.5975 22.6125 23.6625 ;
      RECT  22.7 22.86 22.7525 22.9225 ;
      RECT  22.2525 23.7475 22.3875 23.8125 ;
      RECT  22.13 23.0075 22.2 23.2975 ;
      RECT  22.235 23.2325 22.3 23.9725 ;
      RECT  22.75 23.8625 22.82 24.0625 ;
      RECT  22.67 23.0075 22.735 23.1425 ;
      RECT  21.995 22.86 22.0475 22.9225 ;
      RECT  21.99 24.0625 22.875 24.1275 ;
      RECT  22.0475 23.5 22.1125 23.635 ;
      RECT  22.365 22.7175 22.5 22.7825 ;
      RECT  22.67 23.0075 22.74 23.2975 ;
      RECT  22.3475 22.8575 22.4825 22.9225 ;
      RECT  22.05 23.8625 22.115 23.9975 ;
      RECT  22.565 23.2325 22.74 23.2975 ;
      RECT  22.565 23.8625 22.63 23.9975 ;
      RECT  21.99 22.7175 22.875 22.7825 ;
      RECT  22.7525 23.5 22.8175 23.635 ;
      RECT  22.045 23.3975 22.115 23.5325 ;
      RECT  22.315 23.0075 22.38 23.1425 ;
      RECT  22.565 23.3975 22.63 23.5325 ;
      RECT  22.4975 23.0075 22.5625 23.1425 ;
      RECT  22.05 23.3975 22.115 23.5325 ;
      RECT  22.235 23.8625 22.3 23.9975 ;
      RECT  22.565 23.2325 22.63 23.8625 ;
      RECT  22.0125 22.7175 22.1475 22.7825 ;
      RECT  22.13 23.0075 22.195 23.1425 ;
      RECT  22.235 24.7925 22.3 24.6575 ;
      RECT  22.75 24.7925 22.82 24.6575 ;
      RECT  22.13 24.9575 22.3 24.8925 ;
      RECT  21.99 25.3325 22.875 25.2675 ;
      RECT  22.045 24.3275 22.115 24.1275 ;
      RECT  22.75 24.3275 22.815 24.1925 ;
      RECT  22.3025 25.1825 22.3675 25.0475 ;
      RECT  22.485 25.1825 22.55 25.0475 ;
      RECT  22.75 24.7925 22.815 24.6575 ;
      RECT  22.7175 25.4725 22.8525 25.4075 ;
      RECT  22.4775 24.5925 22.6125 24.5275 ;
      RECT  22.7 25.33 22.7525 25.2675 ;
      RECT  22.2525 24.4425 22.3875 24.3775 ;
      RECT  22.13 25.1825 22.2 24.8925 ;
      RECT  22.235 24.9575 22.3 24.2175 ;
      RECT  22.75 24.3275 22.82 24.1275 ;
      RECT  22.67 25.1825 22.735 25.0475 ;
      RECT  21.995 25.33 22.0475 25.2675 ;
      RECT  21.99 24.1275 22.875 24.0625 ;
      RECT  22.0475 24.69 22.1125 24.555 ;
      RECT  22.365 25.4725 22.5 25.4075 ;
      RECT  22.67 25.1825 22.74 24.8925 ;
      RECT  22.3475 25.3325 22.4825 25.2675 ;
      RECT  22.05 24.3275 22.115 24.1925 ;
      RECT  22.565 24.9575 22.74 24.8925 ;
      RECT  22.565 24.3275 22.63 24.1925 ;
      RECT  21.99 25.4725 22.875 25.4075 ;
      RECT  22.7525 24.69 22.8175 24.555 ;
      RECT  22.045 24.7925 22.115 24.6575 ;
      RECT  22.315 25.1825 22.38 25.0475 ;
      RECT  22.565 24.7925 22.63 24.6575 ;
      RECT  22.4975 25.1825 22.5625 25.0475 ;
      RECT  22.05 24.7925 22.115 24.6575 ;
      RECT  22.235 24.3275 22.3 24.1925 ;
      RECT  22.565 24.9575 22.63 24.3275 ;
      RECT  22.0125 25.4725 22.1475 25.4075 ;
      RECT  22.13 25.1825 22.195 25.0475 ;
      RECT  22.235 26.0875 22.3 26.2225 ;
      RECT  22.75 26.0875 22.82 26.2225 ;
      RECT  22.13 25.9225 22.3 25.9875 ;
      RECT  21.99 25.5475 22.875 25.6125 ;
      RECT  22.045 26.5525 22.115 26.7525 ;
      RECT  22.75 26.5525 22.815 26.6875 ;
      RECT  22.3025 25.6975 22.3675 25.8325 ;
      RECT  22.485 25.6975 22.55 25.8325 ;
      RECT  22.75 26.0875 22.815 26.2225 ;
      RECT  22.7175 25.4075 22.8525 25.4725 ;
      RECT  22.4775 26.2875 22.6125 26.3525 ;
      RECT  22.7 25.55 22.7525 25.6125 ;
      RECT  22.2525 26.4375 22.3875 26.5025 ;
      RECT  22.13 25.6975 22.2 25.9875 ;
      RECT  22.235 25.9225 22.3 26.6625 ;
      RECT  22.75 26.5525 22.82 26.7525 ;
      RECT  22.67 25.6975 22.735 25.8325 ;
      RECT  21.995 25.55 22.0475 25.6125 ;
      RECT  21.99 26.7525 22.875 26.8175 ;
      RECT  22.0475 26.19 22.1125 26.325 ;
      RECT  22.365 25.4075 22.5 25.4725 ;
      RECT  22.67 25.6975 22.74 25.9875 ;
      RECT  22.3475 25.5475 22.4825 25.6125 ;
      RECT  22.05 26.5525 22.115 26.6875 ;
      RECT  22.565 25.9225 22.74 25.9875 ;
      RECT  22.565 26.5525 22.63 26.6875 ;
      RECT  21.99 25.4075 22.875 25.4725 ;
      RECT  22.7525 26.19 22.8175 26.325 ;
      RECT  22.045 26.0875 22.115 26.2225 ;
      RECT  22.315 25.6975 22.38 25.8325 ;
      RECT  22.565 26.0875 22.63 26.2225 ;
      RECT  22.4975 25.6975 22.5625 25.8325 ;
      RECT  22.05 26.0875 22.115 26.2225 ;
      RECT  22.235 26.5525 22.3 26.6875 ;
      RECT  22.565 25.9225 22.63 26.5525 ;
      RECT  22.0125 25.4075 22.1475 25.4725 ;
      RECT  22.13 25.6975 22.195 25.8325 ;
      RECT  22.235 27.4825 22.3 27.3475 ;
      RECT  22.75 27.4825 22.82 27.3475 ;
      RECT  22.13 27.6475 22.3 27.5825 ;
      RECT  21.99 28.0225 22.875 27.9575 ;
      RECT  22.045 27.0175 22.115 26.8175 ;
      RECT  22.75 27.0175 22.815 26.8825 ;
      RECT  22.3025 27.8725 22.3675 27.7375 ;
      RECT  22.485 27.8725 22.55 27.7375 ;
      RECT  22.75 27.4825 22.815 27.3475 ;
      RECT  22.7175 28.1625 22.8525 28.0975 ;
      RECT  22.4775 27.2825 22.6125 27.2175 ;
      RECT  22.7 28.02 22.7525 27.9575 ;
      RECT  22.2525 27.1325 22.3875 27.0675 ;
      RECT  22.13 27.8725 22.2 27.5825 ;
      RECT  22.235 27.6475 22.3 26.9075 ;
      RECT  22.75 27.0175 22.82 26.8175 ;
      RECT  22.67 27.8725 22.735 27.7375 ;
      RECT  21.995 28.02 22.0475 27.9575 ;
      RECT  21.99 26.8175 22.875 26.7525 ;
      RECT  22.0475 27.38 22.1125 27.245 ;
      RECT  22.365 28.1625 22.5 28.0975 ;
      RECT  22.67 27.8725 22.74 27.5825 ;
      RECT  22.3475 28.0225 22.4825 27.9575 ;
      RECT  22.05 27.0175 22.115 26.8825 ;
      RECT  22.565 27.6475 22.74 27.5825 ;
      RECT  22.565 27.0175 22.63 26.8825 ;
      RECT  21.99 28.1625 22.875 28.0975 ;
      RECT  22.7525 27.38 22.8175 27.245 ;
      RECT  22.045 27.4825 22.115 27.3475 ;
      RECT  22.315 27.8725 22.38 27.7375 ;
      RECT  22.565 27.4825 22.63 27.3475 ;
      RECT  22.4975 27.8725 22.5625 27.7375 ;
      RECT  22.05 27.4825 22.115 27.3475 ;
      RECT  22.235 27.0175 22.3 26.8825 ;
      RECT  22.565 27.6475 22.63 27.0175 ;
      RECT  22.0125 28.1625 22.1475 28.0975 ;
      RECT  22.13 27.8725 22.195 27.7375 ;
      RECT  22.235 28.7775 22.3 28.9125 ;
      RECT  22.75 28.7775 22.82 28.9125 ;
      RECT  22.13 28.6125 22.3 28.6775 ;
      RECT  21.99 28.2375 22.875 28.3025 ;
      RECT  22.045 29.2425 22.115 29.4425 ;
      RECT  22.75 29.2425 22.815 29.3775 ;
      RECT  22.3025 28.3875 22.3675 28.5225 ;
      RECT  22.485 28.3875 22.55 28.5225 ;
      RECT  22.75 28.7775 22.815 28.9125 ;
      RECT  22.7175 28.0975 22.8525 28.1625 ;
      RECT  22.4775 28.9775 22.6125 29.0425 ;
      RECT  22.7 28.24 22.7525 28.3025 ;
      RECT  22.2525 29.1275 22.3875 29.1925 ;
      RECT  22.13 28.3875 22.2 28.6775 ;
      RECT  22.235 28.6125 22.3 29.3525 ;
      RECT  22.75 29.2425 22.82 29.4425 ;
      RECT  22.67 28.3875 22.735 28.5225 ;
      RECT  21.995 28.24 22.0475 28.3025 ;
      RECT  21.99 29.4425 22.875 29.5075 ;
      RECT  22.0475 28.88 22.1125 29.015 ;
      RECT  22.365 28.0975 22.5 28.1625 ;
      RECT  22.67 28.3875 22.74 28.6775 ;
      RECT  22.3475 28.2375 22.4825 28.3025 ;
      RECT  22.05 29.2425 22.115 29.3775 ;
      RECT  22.565 28.6125 22.74 28.6775 ;
      RECT  22.565 29.2425 22.63 29.3775 ;
      RECT  21.99 28.0975 22.875 28.1625 ;
      RECT  22.7525 28.88 22.8175 29.015 ;
      RECT  22.045 28.7775 22.115 28.9125 ;
      RECT  22.315 28.3875 22.38 28.5225 ;
      RECT  22.565 28.7775 22.63 28.9125 ;
      RECT  22.4975 28.3875 22.5625 28.5225 ;
      RECT  22.05 28.7775 22.115 28.9125 ;
      RECT  22.235 29.2425 22.3 29.3775 ;
      RECT  22.565 28.6125 22.63 29.2425 ;
      RECT  22.0125 28.0975 22.1475 28.1625 ;
      RECT  22.13 28.3875 22.195 28.5225 ;
      RECT  22.235 30.1725 22.3 30.0375 ;
      RECT  22.75 30.1725 22.82 30.0375 ;
      RECT  22.13 30.3375 22.3 30.2725 ;
      RECT  21.99 30.7125 22.875 30.6475 ;
      RECT  22.045 29.7075 22.115 29.5075 ;
      RECT  22.75 29.7075 22.815 29.5725 ;
      RECT  22.3025 30.5625 22.3675 30.4275 ;
      RECT  22.485 30.5625 22.55 30.4275 ;
      RECT  22.75 30.1725 22.815 30.0375 ;
      RECT  22.7175 30.8525 22.8525 30.7875 ;
      RECT  22.4775 29.9725 22.6125 29.9075 ;
      RECT  22.7 30.71 22.7525 30.6475 ;
      RECT  22.2525 29.8225 22.3875 29.7575 ;
      RECT  22.13 30.5625 22.2 30.2725 ;
      RECT  22.235 30.3375 22.3 29.5975 ;
      RECT  22.75 29.7075 22.82 29.5075 ;
      RECT  22.67 30.5625 22.735 30.4275 ;
      RECT  21.995 30.71 22.0475 30.6475 ;
      RECT  21.99 29.5075 22.875 29.4425 ;
      RECT  22.0475 30.07 22.1125 29.935 ;
      RECT  22.365 30.8525 22.5 30.7875 ;
      RECT  22.67 30.5625 22.74 30.2725 ;
      RECT  22.3475 30.7125 22.4825 30.6475 ;
      RECT  22.05 29.7075 22.115 29.5725 ;
      RECT  22.565 30.3375 22.74 30.2725 ;
      RECT  22.565 29.7075 22.63 29.5725 ;
      RECT  21.99 30.8525 22.875 30.7875 ;
      RECT  22.7525 30.07 22.8175 29.935 ;
      RECT  22.045 30.1725 22.115 30.0375 ;
      RECT  22.315 30.5625 22.38 30.4275 ;
      RECT  22.565 30.1725 22.63 30.0375 ;
      RECT  22.4975 30.5625 22.5625 30.4275 ;
      RECT  22.05 30.1725 22.115 30.0375 ;
      RECT  22.235 29.7075 22.3 29.5725 ;
      RECT  22.565 30.3375 22.63 29.7075 ;
      RECT  22.0125 30.8525 22.1475 30.7875 ;
      RECT  22.13 30.5625 22.195 30.4275 ;
      RECT  22.235 31.4675 22.3 31.6025 ;
      RECT  22.75 31.4675 22.82 31.6025 ;
      RECT  22.13 31.3025 22.3 31.3675 ;
      RECT  21.99 30.9275 22.875 30.9925 ;
      RECT  22.045 31.9325 22.115 32.1325 ;
      RECT  22.75 31.9325 22.815 32.0675 ;
      RECT  22.3025 31.0775 22.3675 31.2125 ;
      RECT  22.485 31.0775 22.55 31.2125 ;
      RECT  22.75 31.4675 22.815 31.6025 ;
      RECT  22.7175 30.7875 22.8525 30.8525 ;
      RECT  22.4775 31.6675 22.6125 31.7325 ;
      RECT  22.7 30.93 22.7525 30.9925 ;
      RECT  22.2525 31.8175 22.3875 31.8825 ;
      RECT  22.13 31.0775 22.2 31.3675 ;
      RECT  22.235 31.3025 22.3 32.0425 ;
      RECT  22.75 31.9325 22.82 32.1325 ;
      RECT  22.67 31.0775 22.735 31.2125 ;
      RECT  21.995 30.93 22.0475 30.9925 ;
      RECT  21.99 32.1325 22.875 32.1975 ;
      RECT  22.0475 31.57 22.1125 31.705 ;
      RECT  22.365 30.7875 22.5 30.8525 ;
      RECT  22.67 31.0775 22.74 31.3675 ;
      RECT  22.3475 30.9275 22.4825 30.9925 ;
      RECT  22.05 31.9325 22.115 32.0675 ;
      RECT  22.565 31.3025 22.74 31.3675 ;
      RECT  22.565 31.9325 22.63 32.0675 ;
      RECT  21.99 30.7875 22.875 30.8525 ;
      RECT  22.7525 31.57 22.8175 31.705 ;
      RECT  22.045 31.4675 22.115 31.6025 ;
      RECT  22.315 31.0775 22.38 31.2125 ;
      RECT  22.565 31.4675 22.63 31.6025 ;
      RECT  22.4975 31.0775 22.5625 31.2125 ;
      RECT  22.05 31.4675 22.115 31.6025 ;
      RECT  22.235 31.9325 22.3 32.0675 ;
      RECT  22.565 31.3025 22.63 31.9325 ;
      RECT  22.0125 30.7875 22.1475 30.8525 ;
      RECT  22.13 31.0775 22.195 31.2125 ;
      RECT  22.235 32.8625 22.3 32.7275 ;
      RECT  22.75 32.8625 22.82 32.7275 ;
      RECT  22.13 33.0275 22.3 32.9625 ;
      RECT  21.99 33.4025 22.875 33.3375 ;
      RECT  22.045 32.3975 22.115 32.1975 ;
      RECT  22.75 32.3975 22.815 32.2625 ;
      RECT  22.3025 33.2525 22.3675 33.1175 ;
      RECT  22.485 33.2525 22.55 33.1175 ;
      RECT  22.75 32.8625 22.815 32.7275 ;
      RECT  22.7175 33.5425 22.8525 33.4775 ;
      RECT  22.4775 32.6625 22.6125 32.5975 ;
      RECT  22.7 33.4 22.7525 33.3375 ;
      RECT  22.2525 32.5125 22.3875 32.4475 ;
      RECT  22.13 33.2525 22.2 32.9625 ;
      RECT  22.235 33.0275 22.3 32.2875 ;
      RECT  22.75 32.3975 22.82 32.1975 ;
      RECT  22.67 33.2525 22.735 33.1175 ;
      RECT  21.995 33.4 22.0475 33.3375 ;
      RECT  21.99 32.1975 22.875 32.1325 ;
      RECT  22.0475 32.76 22.1125 32.625 ;
      RECT  22.365 33.5425 22.5 33.4775 ;
      RECT  22.67 33.2525 22.74 32.9625 ;
      RECT  22.3475 33.4025 22.4825 33.3375 ;
      RECT  22.05 32.3975 22.115 32.2625 ;
      RECT  22.565 33.0275 22.74 32.9625 ;
      RECT  22.565 32.3975 22.63 32.2625 ;
      RECT  21.99 33.5425 22.875 33.4775 ;
      RECT  22.7525 32.76 22.8175 32.625 ;
      RECT  22.045 32.8625 22.115 32.7275 ;
      RECT  22.315 33.2525 22.38 33.1175 ;
      RECT  22.565 32.8625 22.63 32.7275 ;
      RECT  22.4975 33.2525 22.5625 33.1175 ;
      RECT  22.05 32.8625 22.115 32.7275 ;
      RECT  22.235 32.3975 22.3 32.2625 ;
      RECT  22.565 33.0275 22.63 32.3975 ;
      RECT  22.0125 33.5425 22.1475 33.4775 ;
      RECT  22.13 33.2525 22.195 33.1175 ;
      RECT  22.235 34.1575 22.3 34.2925 ;
      RECT  22.75 34.1575 22.82 34.2925 ;
      RECT  22.13 33.9925 22.3 34.0575 ;
      RECT  21.99 33.6175 22.875 33.6825 ;
      RECT  22.045 34.6225 22.115 34.8225 ;
      RECT  22.75 34.6225 22.815 34.7575 ;
      RECT  22.3025 33.7675 22.3675 33.9025 ;
      RECT  22.485 33.7675 22.55 33.9025 ;
      RECT  22.75 34.1575 22.815 34.2925 ;
      RECT  22.7175 33.4775 22.8525 33.5425 ;
      RECT  22.4775 34.3575 22.6125 34.4225 ;
      RECT  22.7 33.62 22.7525 33.6825 ;
      RECT  22.2525 34.5075 22.3875 34.5725 ;
      RECT  22.13 33.7675 22.2 34.0575 ;
      RECT  22.235 33.9925 22.3 34.7325 ;
      RECT  22.75 34.6225 22.82 34.8225 ;
      RECT  22.67 33.7675 22.735 33.9025 ;
      RECT  21.995 33.62 22.0475 33.6825 ;
      RECT  21.99 34.8225 22.875 34.8875 ;
      RECT  22.0475 34.26 22.1125 34.395 ;
      RECT  22.365 33.4775 22.5 33.5425 ;
      RECT  22.67 33.7675 22.74 34.0575 ;
      RECT  22.3475 33.6175 22.4825 33.6825 ;
      RECT  22.05 34.6225 22.115 34.7575 ;
      RECT  22.565 33.9925 22.74 34.0575 ;
      RECT  22.565 34.6225 22.63 34.7575 ;
      RECT  21.99 33.4775 22.875 33.5425 ;
      RECT  22.7525 34.26 22.8175 34.395 ;
      RECT  22.045 34.1575 22.115 34.2925 ;
      RECT  22.315 33.7675 22.38 33.9025 ;
      RECT  22.565 34.1575 22.63 34.2925 ;
      RECT  22.4975 33.7675 22.5625 33.9025 ;
      RECT  22.05 34.1575 22.115 34.2925 ;
      RECT  22.235 34.6225 22.3 34.7575 ;
      RECT  22.565 33.9925 22.63 34.6225 ;
      RECT  22.0125 33.4775 22.1475 33.5425 ;
      RECT  22.13 33.7675 22.195 33.9025 ;
      RECT  22.235 35.5525 22.3 35.4175 ;
      RECT  22.75 35.5525 22.82 35.4175 ;
      RECT  22.13 35.7175 22.3 35.6525 ;
      RECT  21.99 36.0925 22.875 36.0275 ;
      RECT  22.045 35.0875 22.115 34.8875 ;
      RECT  22.75 35.0875 22.815 34.9525 ;
      RECT  22.3025 35.9425 22.3675 35.8075 ;
      RECT  22.485 35.9425 22.55 35.8075 ;
      RECT  22.75 35.5525 22.815 35.4175 ;
      RECT  22.7175 36.2325 22.8525 36.1675 ;
      RECT  22.4775 35.3525 22.6125 35.2875 ;
      RECT  22.7 36.09 22.7525 36.0275 ;
      RECT  22.2525 35.2025 22.3875 35.1375 ;
      RECT  22.13 35.9425 22.2 35.6525 ;
      RECT  22.235 35.7175 22.3 34.9775 ;
      RECT  22.75 35.0875 22.82 34.8875 ;
      RECT  22.67 35.9425 22.735 35.8075 ;
      RECT  21.995 36.09 22.0475 36.0275 ;
      RECT  21.99 34.8875 22.875 34.8225 ;
      RECT  22.0475 35.45 22.1125 35.315 ;
      RECT  22.365 36.2325 22.5 36.1675 ;
      RECT  22.67 35.9425 22.74 35.6525 ;
      RECT  22.3475 36.0925 22.4825 36.0275 ;
      RECT  22.05 35.0875 22.115 34.9525 ;
      RECT  22.565 35.7175 22.74 35.6525 ;
      RECT  22.565 35.0875 22.63 34.9525 ;
      RECT  21.99 36.2325 22.875 36.1675 ;
      RECT  22.7525 35.45 22.8175 35.315 ;
      RECT  22.045 35.5525 22.115 35.4175 ;
      RECT  22.315 35.9425 22.38 35.8075 ;
      RECT  22.565 35.5525 22.63 35.4175 ;
      RECT  22.4975 35.9425 22.5625 35.8075 ;
      RECT  22.05 35.5525 22.115 35.4175 ;
      RECT  22.235 35.0875 22.3 34.9525 ;
      RECT  22.565 35.7175 22.63 35.0875 ;
      RECT  22.0125 36.2325 22.1475 36.1675 ;
      RECT  22.13 35.9425 22.195 35.8075 ;
      RECT  22.235 36.8475 22.3 36.9825 ;
      RECT  22.75 36.8475 22.82 36.9825 ;
      RECT  22.13 36.6825 22.3 36.7475 ;
      RECT  21.99 36.3075 22.875 36.3725 ;
      RECT  22.045 37.3125 22.115 37.5125 ;
      RECT  22.75 37.3125 22.815 37.4475 ;
      RECT  22.3025 36.4575 22.3675 36.5925 ;
      RECT  22.485 36.4575 22.55 36.5925 ;
      RECT  22.75 36.8475 22.815 36.9825 ;
      RECT  22.7175 36.1675 22.8525 36.2325 ;
      RECT  22.4775 37.0475 22.6125 37.1125 ;
      RECT  22.7 36.31 22.7525 36.3725 ;
      RECT  22.2525 37.1975 22.3875 37.2625 ;
      RECT  22.13 36.4575 22.2 36.7475 ;
      RECT  22.235 36.6825 22.3 37.4225 ;
      RECT  22.75 37.3125 22.82 37.5125 ;
      RECT  22.67 36.4575 22.735 36.5925 ;
      RECT  21.995 36.31 22.0475 36.3725 ;
      RECT  21.99 37.5125 22.875 37.5775 ;
      RECT  22.0475 36.95 22.1125 37.085 ;
      RECT  22.365 36.1675 22.5 36.2325 ;
      RECT  22.67 36.4575 22.74 36.7475 ;
      RECT  22.3475 36.3075 22.4825 36.3725 ;
      RECT  22.05 37.3125 22.115 37.4475 ;
      RECT  22.565 36.6825 22.74 36.7475 ;
      RECT  22.565 37.3125 22.63 37.4475 ;
      RECT  21.99 36.1675 22.875 36.2325 ;
      RECT  22.7525 36.95 22.8175 37.085 ;
      RECT  22.045 36.8475 22.115 36.9825 ;
      RECT  22.315 36.4575 22.38 36.5925 ;
      RECT  22.565 36.8475 22.63 36.9825 ;
      RECT  22.4975 36.4575 22.5625 36.5925 ;
      RECT  22.05 36.8475 22.115 36.9825 ;
      RECT  22.235 37.3125 22.3 37.4475 ;
      RECT  22.565 36.6825 22.63 37.3125 ;
      RECT  22.0125 36.1675 22.1475 36.2325 ;
      RECT  22.13 36.4575 22.195 36.5925 ;
      RECT  22.235 38.2425 22.3 38.1075 ;
      RECT  22.75 38.2425 22.82 38.1075 ;
      RECT  22.13 38.4075 22.3 38.3425 ;
      RECT  21.99 38.7825 22.875 38.7175 ;
      RECT  22.045 37.7775 22.115 37.5775 ;
      RECT  22.75 37.7775 22.815 37.6425 ;
      RECT  22.3025 38.6325 22.3675 38.4975 ;
      RECT  22.485 38.6325 22.55 38.4975 ;
      RECT  22.75 38.2425 22.815 38.1075 ;
      RECT  22.7175 38.9225 22.8525 38.8575 ;
      RECT  22.4775 38.0425 22.6125 37.9775 ;
      RECT  22.7 38.78 22.7525 38.7175 ;
      RECT  22.2525 37.8925 22.3875 37.8275 ;
      RECT  22.13 38.6325 22.2 38.3425 ;
      RECT  22.235 38.4075 22.3 37.6675 ;
      RECT  22.75 37.7775 22.82 37.5775 ;
      RECT  22.67 38.6325 22.735 38.4975 ;
      RECT  21.995 38.78 22.0475 38.7175 ;
      RECT  21.99 37.5775 22.875 37.5125 ;
      RECT  22.0475 38.14 22.1125 38.005 ;
      RECT  22.365 38.9225 22.5 38.8575 ;
      RECT  22.67 38.6325 22.74 38.3425 ;
      RECT  22.3475 38.7825 22.4825 38.7175 ;
      RECT  22.05 37.7775 22.115 37.6425 ;
      RECT  22.565 38.4075 22.74 38.3425 ;
      RECT  22.565 37.7775 22.63 37.6425 ;
      RECT  21.99 38.9225 22.875 38.8575 ;
      RECT  22.7525 38.14 22.8175 38.005 ;
      RECT  22.045 38.2425 22.115 38.1075 ;
      RECT  22.315 38.6325 22.38 38.4975 ;
      RECT  22.565 38.2425 22.63 38.1075 ;
      RECT  22.4975 38.6325 22.5625 38.4975 ;
      RECT  22.05 38.2425 22.115 38.1075 ;
      RECT  22.235 37.7775 22.3 37.6425 ;
      RECT  22.565 38.4075 22.63 37.7775 ;
      RECT  22.0125 38.9225 22.1475 38.8575 ;
      RECT  22.13 38.6325 22.195 38.4975 ;
      RECT  22.235 39.5375 22.3 39.6725 ;
      RECT  22.75 39.5375 22.82 39.6725 ;
      RECT  22.13 39.3725 22.3 39.4375 ;
      RECT  21.99 38.9975 22.875 39.0625 ;
      RECT  22.045 40.0025 22.115 40.2025 ;
      RECT  22.75 40.0025 22.815 40.1375 ;
      RECT  22.3025 39.1475 22.3675 39.2825 ;
      RECT  22.485 39.1475 22.55 39.2825 ;
      RECT  22.75 39.5375 22.815 39.6725 ;
      RECT  22.7175 38.8575 22.8525 38.9225 ;
      RECT  22.4775 39.7375 22.6125 39.8025 ;
      RECT  22.7 39.0 22.7525 39.0625 ;
      RECT  22.2525 39.8875 22.3875 39.9525 ;
      RECT  22.13 39.1475 22.2 39.4375 ;
      RECT  22.235 39.3725 22.3 40.1125 ;
      RECT  22.75 40.0025 22.82 40.2025 ;
      RECT  22.67 39.1475 22.735 39.2825 ;
      RECT  21.995 39.0 22.0475 39.0625 ;
      RECT  21.99 40.2025 22.875 40.2675 ;
      RECT  22.0475 39.64 22.1125 39.775 ;
      RECT  22.365 38.8575 22.5 38.9225 ;
      RECT  22.67 39.1475 22.74 39.4375 ;
      RECT  22.3475 38.9975 22.4825 39.0625 ;
      RECT  22.05 40.0025 22.115 40.1375 ;
      RECT  22.565 39.3725 22.74 39.4375 ;
      RECT  22.565 40.0025 22.63 40.1375 ;
      RECT  21.99 38.8575 22.875 38.9225 ;
      RECT  22.7525 39.64 22.8175 39.775 ;
      RECT  22.045 39.5375 22.115 39.6725 ;
      RECT  22.315 39.1475 22.38 39.2825 ;
      RECT  22.565 39.5375 22.63 39.6725 ;
      RECT  22.4975 39.1475 22.5625 39.2825 ;
      RECT  22.05 39.5375 22.115 39.6725 ;
      RECT  22.235 40.0025 22.3 40.1375 ;
      RECT  22.565 39.3725 22.63 40.0025 ;
      RECT  22.0125 38.8575 22.1475 38.9225 ;
      RECT  22.13 39.1475 22.195 39.2825 ;
      RECT  22.235 40.9325 22.3 40.7975 ;
      RECT  22.75 40.9325 22.82 40.7975 ;
      RECT  22.13 41.0975 22.3 41.0325 ;
      RECT  21.99 41.4725 22.875 41.4075 ;
      RECT  22.045 40.4675 22.115 40.2675 ;
      RECT  22.75 40.4675 22.815 40.3325 ;
      RECT  22.3025 41.3225 22.3675 41.1875 ;
      RECT  22.485 41.3225 22.55 41.1875 ;
      RECT  22.75 40.9325 22.815 40.7975 ;
      RECT  22.7175 41.6125 22.8525 41.5475 ;
      RECT  22.4775 40.7325 22.6125 40.6675 ;
      RECT  22.7 41.47 22.7525 41.4075 ;
      RECT  22.2525 40.5825 22.3875 40.5175 ;
      RECT  22.13 41.3225 22.2 41.0325 ;
      RECT  22.235 41.0975 22.3 40.3575 ;
      RECT  22.75 40.4675 22.82 40.2675 ;
      RECT  22.67 41.3225 22.735 41.1875 ;
      RECT  21.995 41.47 22.0475 41.4075 ;
      RECT  21.99 40.2675 22.875 40.2025 ;
      RECT  22.0475 40.83 22.1125 40.695 ;
      RECT  22.365 41.6125 22.5 41.5475 ;
      RECT  22.67 41.3225 22.74 41.0325 ;
      RECT  22.3475 41.4725 22.4825 41.4075 ;
      RECT  22.05 40.4675 22.115 40.3325 ;
      RECT  22.565 41.0975 22.74 41.0325 ;
      RECT  22.565 40.4675 22.63 40.3325 ;
      RECT  21.99 41.6125 22.875 41.5475 ;
      RECT  22.7525 40.83 22.8175 40.695 ;
      RECT  22.045 40.9325 22.115 40.7975 ;
      RECT  22.315 41.3225 22.38 41.1875 ;
      RECT  22.565 40.9325 22.63 40.7975 ;
      RECT  22.4975 41.3225 22.5625 41.1875 ;
      RECT  22.05 40.9325 22.115 40.7975 ;
      RECT  22.235 40.4675 22.3 40.3325 ;
      RECT  22.565 41.0975 22.63 40.4675 ;
      RECT  22.0125 41.6125 22.1475 41.5475 ;
      RECT  22.13 41.3225 22.195 41.1875 ;
      RECT  22.235 42.2275 22.3 42.3625 ;
      RECT  22.75 42.2275 22.82 42.3625 ;
      RECT  22.13 42.0625 22.3 42.1275 ;
      RECT  21.99 41.6875 22.875 41.7525 ;
      RECT  22.045 42.6925 22.115 42.8925 ;
      RECT  22.75 42.6925 22.815 42.8275 ;
      RECT  22.3025 41.8375 22.3675 41.9725 ;
      RECT  22.485 41.8375 22.55 41.9725 ;
      RECT  22.75 42.2275 22.815 42.3625 ;
      RECT  22.7175 41.5475 22.8525 41.6125 ;
      RECT  22.4775 42.4275 22.6125 42.4925 ;
      RECT  22.7 41.69 22.7525 41.7525 ;
      RECT  22.2525 42.5775 22.3875 42.6425 ;
      RECT  22.13 41.8375 22.2 42.1275 ;
      RECT  22.235 42.0625 22.3 42.8025 ;
      RECT  22.75 42.6925 22.82 42.8925 ;
      RECT  22.67 41.8375 22.735 41.9725 ;
      RECT  21.995 41.69 22.0475 41.7525 ;
      RECT  21.99 42.8925 22.875 42.9575 ;
      RECT  22.0475 42.33 22.1125 42.465 ;
      RECT  22.365 41.5475 22.5 41.6125 ;
      RECT  22.67 41.8375 22.74 42.1275 ;
      RECT  22.3475 41.6875 22.4825 41.7525 ;
      RECT  22.05 42.6925 22.115 42.8275 ;
      RECT  22.565 42.0625 22.74 42.1275 ;
      RECT  22.565 42.6925 22.63 42.8275 ;
      RECT  21.99 41.5475 22.875 41.6125 ;
      RECT  22.7525 42.33 22.8175 42.465 ;
      RECT  22.045 42.2275 22.115 42.3625 ;
      RECT  22.315 41.8375 22.38 41.9725 ;
      RECT  22.565 42.2275 22.63 42.3625 ;
      RECT  22.4975 41.8375 22.5625 41.9725 ;
      RECT  22.05 42.2275 22.115 42.3625 ;
      RECT  22.235 42.6925 22.3 42.8275 ;
      RECT  22.565 42.0625 22.63 42.6925 ;
      RECT  22.0125 41.5475 22.1475 41.6125 ;
      RECT  22.13 41.8375 22.195 41.9725 ;
      RECT  22.235 43.6225 22.3 43.4875 ;
      RECT  22.75 43.6225 22.82 43.4875 ;
      RECT  22.13 43.7875 22.3 43.7225 ;
      RECT  21.99 44.1625 22.875 44.0975 ;
      RECT  22.045 43.1575 22.115 42.9575 ;
      RECT  22.75 43.1575 22.815 43.0225 ;
      RECT  22.3025 44.0125 22.3675 43.8775 ;
      RECT  22.485 44.0125 22.55 43.8775 ;
      RECT  22.75 43.6225 22.815 43.4875 ;
      RECT  22.7175 44.3025 22.8525 44.2375 ;
      RECT  22.4775 43.4225 22.6125 43.3575 ;
      RECT  22.7 44.16 22.7525 44.0975 ;
      RECT  22.2525 43.2725 22.3875 43.2075 ;
      RECT  22.13 44.0125 22.2 43.7225 ;
      RECT  22.235 43.7875 22.3 43.0475 ;
      RECT  22.75 43.1575 22.82 42.9575 ;
      RECT  22.67 44.0125 22.735 43.8775 ;
      RECT  21.995 44.16 22.0475 44.0975 ;
      RECT  21.99 42.9575 22.875 42.8925 ;
      RECT  22.0475 43.52 22.1125 43.385 ;
      RECT  22.365 44.3025 22.5 44.2375 ;
      RECT  22.67 44.0125 22.74 43.7225 ;
      RECT  22.3475 44.1625 22.4825 44.0975 ;
      RECT  22.05 43.1575 22.115 43.0225 ;
      RECT  22.565 43.7875 22.74 43.7225 ;
      RECT  22.565 43.1575 22.63 43.0225 ;
      RECT  21.99 44.3025 22.875 44.2375 ;
      RECT  22.7525 43.52 22.8175 43.385 ;
      RECT  22.045 43.6225 22.115 43.4875 ;
      RECT  22.315 44.0125 22.38 43.8775 ;
      RECT  22.565 43.6225 22.63 43.4875 ;
      RECT  22.4975 44.0125 22.5625 43.8775 ;
      RECT  22.05 43.6225 22.115 43.4875 ;
      RECT  22.235 43.1575 22.3 43.0225 ;
      RECT  22.565 43.7875 22.63 43.1575 ;
      RECT  22.0125 44.3025 22.1475 44.2375 ;
      RECT  22.13 44.0125 22.195 43.8775 ;
      RECT  21.375 22.8575 22.785 22.9225 ;
      RECT  21.375 25.2675 22.785 25.3325 ;
      RECT  21.375 25.5475 22.785 25.6125 ;
      RECT  21.375 27.9575 22.785 28.0225 ;
      RECT  21.375 28.2375 22.785 28.3025 ;
      RECT  21.375 30.6475 22.785 30.7125 ;
      RECT  21.375 30.9275 22.785 30.9925 ;
      RECT  21.375 33.3375 22.785 33.4025 ;
      RECT  21.375 33.6175 22.785 33.6825 ;
      RECT  21.375 36.0275 22.785 36.0925 ;
      RECT  21.375 36.3075 22.785 36.3725 ;
      RECT  21.375 38.7175 22.785 38.7825 ;
      RECT  21.375 38.9975 22.785 39.0625 ;
      RECT  21.375 41.4075 22.785 41.4725 ;
      RECT  21.375 41.6875 22.785 41.7525 ;
      RECT  21.375 44.0975 22.785 44.1625 ;
      RECT  20.825 20.7075 20.89 20.8425 ;
      RECT  21.34 20.7075 21.41 20.8425 ;
      RECT  20.72 20.5425 20.89 20.6075 ;
      RECT  20.58 20.1675 21.465 20.2325 ;
      RECT  20.635 21.1725 20.705 21.3725 ;
      RECT  21.34 21.1725 21.405 21.3075 ;
      RECT  20.8925 20.3175 20.9575 20.4525 ;
      RECT  21.075 20.3175 21.14 20.4525 ;
      RECT  21.34 20.7075 21.405 20.8425 ;
      RECT  21.3075 20.0275 21.4425 20.0925 ;
      RECT  21.0675 20.9075 21.2025 20.9725 ;
      RECT  21.29 20.17 21.3425 20.2325 ;
      RECT  20.8425 21.0575 20.9775 21.1225 ;
      RECT  20.72 20.3175 20.79 20.6075 ;
      RECT  20.825 20.5425 20.89 21.2825 ;
      RECT  21.34 21.1725 21.41 21.3725 ;
      RECT  21.26 20.3175 21.325 20.4525 ;
      RECT  20.585 20.17 20.6375 20.2325 ;
      RECT  20.58 21.3725 21.465 21.4375 ;
      RECT  20.6375 20.81 20.7025 20.945 ;
      RECT  20.955 20.0275 21.09 20.0925 ;
      RECT  21.26 20.3175 21.33 20.6075 ;
      RECT  20.9375 20.1675 21.0725 20.2325 ;
      RECT  20.64 21.1725 20.705 21.3075 ;
      RECT  21.155 20.5425 21.33 20.6075 ;
      RECT  21.155 21.1725 21.22 21.3075 ;
      RECT  20.58 20.0275 21.465 20.0925 ;
      RECT  21.3425 20.81 21.4075 20.945 ;
      RECT  20.635 20.7075 20.705 20.8425 ;
      RECT  20.905 20.3175 20.97 20.4525 ;
      RECT  21.155 20.7075 21.22 20.8425 ;
      RECT  21.0875 20.3175 21.1525 20.4525 ;
      RECT  20.64 20.7075 20.705 20.8425 ;
      RECT  20.825 21.1725 20.89 21.3075 ;
      RECT  21.155 20.5425 21.22 21.1725 ;
      RECT  20.6025 20.0275 20.7375 20.0925 ;
      RECT  20.72 20.3175 20.785 20.4525 ;
      RECT  20.825 22.1025 20.89 21.9675 ;
      RECT  20.72 22.2675 20.89 22.2025 ;
      RECT  21.34 22.1025 21.41 21.9675 ;
      RECT  20.58 22.6425 21.465 22.5775 ;
      RECT  20.635 21.6375 20.705 21.4375 ;
      RECT  21.34 21.6375 21.405 21.5025 ;
      RECT  20.8925 22.4925 20.9575 22.3575 ;
      RECT  21.075 22.4925 21.14 22.3575 ;
      RECT  21.34 22.1025 21.405 21.9675 ;
      RECT  21.3075 22.7825 21.4425 22.7175 ;
      RECT  21.0675 21.9025 21.2025 21.8375 ;
      RECT  21.29 22.64 21.3425 22.5775 ;
      RECT  20.8425 21.7525 20.9775 21.6875 ;
      RECT  20.72 22.4925 20.79 22.2025 ;
      RECT  20.825 22.2675 20.89 21.5275 ;
      RECT  21.34 21.6375 21.41 21.4375 ;
      RECT  20.585 22.64 20.6375 22.5775 ;
      RECT  20.58 21.4375 21.465 21.3725 ;
      RECT  21.26 22.4925 21.325 22.3575 ;
      RECT  20.6375 22.0 20.7025 21.865 ;
      RECT  21.26 22.4925 21.33 22.2025 ;
      RECT  20.955 22.7825 21.09 22.7175 ;
      RECT  20.9375 22.6425 21.0725 22.5775 ;
      RECT  21.155 22.2675 21.33 22.2025 ;
      RECT  20.64 21.6375 20.705 21.5025 ;
      RECT  20.58 22.7825 21.465 22.7175 ;
      RECT  21.3425 22.0 21.4075 21.865 ;
      RECT  20.635 22.1025 20.705 21.9675 ;
      RECT  20.905 22.4925 20.97 22.3575 ;
      RECT  21.155 22.1025 21.22 21.9675 ;
      RECT  21.0875 22.4925 21.1525 22.3575 ;
      RECT  20.64 22.1025 20.705 21.9675 ;
      RECT  21.155 21.6375 21.22 21.425 ;
      RECT  20.825 21.6375 20.89 21.5025 ;
      RECT  21.155 22.2675 21.22 21.6375 ;
      RECT  20.6025 22.7825 20.7375 22.7175 ;
      RECT  20.72 22.4925 20.785 22.3575 ;
      RECT  20.825 23.3975 20.89 23.5325 ;
      RECT  20.72 23.2325 20.89 23.2975 ;
      RECT  21.34 23.3975 21.41 23.5325 ;
      RECT  20.58 22.8575 21.465 22.9225 ;
      RECT  20.635 23.8625 20.705 24.0625 ;
      RECT  21.34 23.8625 21.405 23.9975 ;
      RECT  20.8925 23.0075 20.9575 23.1425 ;
      RECT  21.075 23.0075 21.14 23.1425 ;
      RECT  21.34 23.3975 21.405 23.5325 ;
      RECT  21.3075 22.7175 21.4425 22.7825 ;
      RECT  21.0675 23.5975 21.2025 23.6625 ;
      RECT  21.29 22.86 21.3425 22.9225 ;
      RECT  20.8425 23.7475 20.9775 23.8125 ;
      RECT  20.72 23.0075 20.79 23.2975 ;
      RECT  20.825 23.2325 20.89 23.9725 ;
      RECT  21.34 23.8625 21.41 24.0625 ;
      RECT  20.585 22.86 20.6375 22.9225 ;
      RECT  20.58 24.0625 21.465 24.1275 ;
      RECT  21.26 23.0075 21.325 23.1425 ;
      RECT  20.6375 23.5 20.7025 23.635 ;
      RECT  21.26 23.0075 21.33 23.2975 ;
      RECT  20.955 22.7175 21.09 22.7825 ;
      RECT  20.9375 22.8575 21.0725 22.9225 ;
      RECT  21.155 23.2325 21.33 23.2975 ;
      RECT  20.64 23.8625 20.705 23.9975 ;
      RECT  20.58 22.7175 21.465 22.7825 ;
      RECT  21.3425 23.5 21.4075 23.635 ;
      RECT  20.635 23.3975 20.705 23.5325 ;
      RECT  20.905 23.0075 20.97 23.1425 ;
      RECT  21.155 23.3975 21.22 23.5325 ;
      RECT  21.0875 23.0075 21.1525 23.1425 ;
      RECT  20.64 23.3975 20.705 23.5325 ;
      RECT  21.155 23.8625 21.22 24.075 ;
      RECT  20.825 23.8625 20.89 23.9975 ;
      RECT  21.155 23.2325 21.22 23.8625 ;
      RECT  20.6025 22.7175 20.7375 22.7825 ;
      RECT  20.72 23.0075 20.785 23.1425 ;
      RECT  20.825 24.7925 20.89 24.6575 ;
      RECT  20.72 24.9575 20.89 24.8925 ;
      RECT  21.34 24.7925 21.41 24.6575 ;
      RECT  20.58 25.3325 21.465 25.2675 ;
      RECT  20.635 24.3275 20.705 24.1275 ;
      RECT  21.34 24.3275 21.405 24.1925 ;
      RECT  20.8925 25.1825 20.9575 25.0475 ;
      RECT  21.075 25.1825 21.14 25.0475 ;
      RECT  21.34 24.7925 21.405 24.6575 ;
      RECT  21.3075 25.4725 21.4425 25.4075 ;
      RECT  21.0675 24.5925 21.2025 24.5275 ;
      RECT  21.29 25.33 21.3425 25.2675 ;
      RECT  20.8425 24.4425 20.9775 24.3775 ;
      RECT  20.72 25.1825 20.79 24.8925 ;
      RECT  20.825 24.9575 20.89 24.2175 ;
      RECT  21.34 24.3275 21.41 24.1275 ;
      RECT  20.585 25.33 20.6375 25.2675 ;
      RECT  20.58 24.1275 21.465 24.0625 ;
      RECT  21.26 25.1825 21.325 25.0475 ;
      RECT  20.6375 24.69 20.7025 24.555 ;
      RECT  21.26 25.1825 21.33 24.8925 ;
      RECT  20.955 25.4725 21.09 25.4075 ;
      RECT  20.9375 25.3325 21.0725 25.2675 ;
      RECT  21.155 24.9575 21.33 24.8925 ;
      RECT  20.64 24.3275 20.705 24.1925 ;
      RECT  20.58 25.4725 21.465 25.4075 ;
      RECT  21.3425 24.69 21.4075 24.555 ;
      RECT  20.635 24.7925 20.705 24.6575 ;
      RECT  20.905 25.1825 20.97 25.0475 ;
      RECT  21.155 24.7925 21.22 24.6575 ;
      RECT  21.0875 25.1825 21.1525 25.0475 ;
      RECT  20.64 24.7925 20.705 24.6575 ;
      RECT  21.155 24.3275 21.22 24.115 ;
      RECT  20.825 24.3275 20.89 24.1925 ;
      RECT  21.155 24.9575 21.22 24.3275 ;
      RECT  20.6025 25.4725 20.7375 25.4075 ;
      RECT  20.72 25.1825 20.785 25.0475 ;
      RECT  20.825 26.0875 20.89 26.2225 ;
      RECT  20.72 25.9225 20.89 25.9875 ;
      RECT  21.34 26.0875 21.41 26.2225 ;
      RECT  20.58 25.5475 21.465 25.6125 ;
      RECT  20.635 26.5525 20.705 26.7525 ;
      RECT  21.34 26.5525 21.405 26.6875 ;
      RECT  20.8925 25.6975 20.9575 25.8325 ;
      RECT  21.075 25.6975 21.14 25.8325 ;
      RECT  21.34 26.0875 21.405 26.2225 ;
      RECT  21.3075 25.4075 21.4425 25.4725 ;
      RECT  21.0675 26.2875 21.2025 26.3525 ;
      RECT  21.29 25.55 21.3425 25.6125 ;
      RECT  20.8425 26.4375 20.9775 26.5025 ;
      RECT  20.72 25.6975 20.79 25.9875 ;
      RECT  20.825 25.9225 20.89 26.6625 ;
      RECT  21.34 26.5525 21.41 26.7525 ;
      RECT  20.585 25.55 20.6375 25.6125 ;
      RECT  20.58 26.7525 21.465 26.8175 ;
      RECT  21.26 25.6975 21.325 25.8325 ;
      RECT  20.6375 26.19 20.7025 26.325 ;
      RECT  21.26 25.6975 21.33 25.9875 ;
      RECT  20.955 25.4075 21.09 25.4725 ;
      RECT  20.9375 25.5475 21.0725 25.6125 ;
      RECT  21.155 25.9225 21.33 25.9875 ;
      RECT  20.64 26.5525 20.705 26.6875 ;
      RECT  20.58 25.4075 21.465 25.4725 ;
      RECT  21.3425 26.19 21.4075 26.325 ;
      RECT  20.635 26.0875 20.705 26.2225 ;
      RECT  20.905 25.6975 20.97 25.8325 ;
      RECT  21.155 26.0875 21.22 26.2225 ;
      RECT  21.0875 25.6975 21.1525 25.8325 ;
      RECT  20.64 26.0875 20.705 26.2225 ;
      RECT  21.155 26.5525 21.22 26.765 ;
      RECT  20.825 26.5525 20.89 26.6875 ;
      RECT  21.155 25.9225 21.22 26.5525 ;
      RECT  20.6025 25.4075 20.7375 25.4725 ;
      RECT  20.72 25.6975 20.785 25.8325 ;
      RECT  20.825 27.4825 20.89 27.3475 ;
      RECT  20.72 27.6475 20.89 27.5825 ;
      RECT  21.34 27.4825 21.41 27.3475 ;
      RECT  20.58 28.0225 21.465 27.9575 ;
      RECT  20.635 27.0175 20.705 26.8175 ;
      RECT  21.34 27.0175 21.405 26.8825 ;
      RECT  20.8925 27.8725 20.9575 27.7375 ;
      RECT  21.075 27.8725 21.14 27.7375 ;
      RECT  21.34 27.4825 21.405 27.3475 ;
      RECT  21.3075 28.1625 21.4425 28.0975 ;
      RECT  21.0675 27.2825 21.2025 27.2175 ;
      RECT  21.29 28.02 21.3425 27.9575 ;
      RECT  20.8425 27.1325 20.9775 27.0675 ;
      RECT  20.72 27.8725 20.79 27.5825 ;
      RECT  20.825 27.6475 20.89 26.9075 ;
      RECT  21.34 27.0175 21.41 26.8175 ;
      RECT  20.585 28.02 20.6375 27.9575 ;
      RECT  20.58 26.8175 21.465 26.7525 ;
      RECT  21.26 27.8725 21.325 27.7375 ;
      RECT  20.6375 27.38 20.7025 27.245 ;
      RECT  21.26 27.8725 21.33 27.5825 ;
      RECT  20.955 28.1625 21.09 28.0975 ;
      RECT  20.9375 28.0225 21.0725 27.9575 ;
      RECT  21.155 27.6475 21.33 27.5825 ;
      RECT  20.64 27.0175 20.705 26.8825 ;
      RECT  20.58 28.1625 21.465 28.0975 ;
      RECT  21.3425 27.38 21.4075 27.245 ;
      RECT  20.635 27.4825 20.705 27.3475 ;
      RECT  20.905 27.8725 20.97 27.7375 ;
      RECT  21.155 27.4825 21.22 27.3475 ;
      RECT  21.0875 27.8725 21.1525 27.7375 ;
      RECT  20.64 27.4825 20.705 27.3475 ;
      RECT  21.155 27.0175 21.22 26.805 ;
      RECT  20.825 27.0175 20.89 26.8825 ;
      RECT  21.155 27.6475 21.22 27.0175 ;
      RECT  20.6025 28.1625 20.7375 28.0975 ;
      RECT  20.72 27.8725 20.785 27.7375 ;
      RECT  20.825 28.7775 20.89 28.9125 ;
      RECT  20.72 28.6125 20.89 28.6775 ;
      RECT  21.34 28.7775 21.41 28.9125 ;
      RECT  20.58 28.2375 21.465 28.3025 ;
      RECT  20.635 29.2425 20.705 29.4425 ;
      RECT  21.34 29.2425 21.405 29.3775 ;
      RECT  20.8925 28.3875 20.9575 28.5225 ;
      RECT  21.075 28.3875 21.14 28.5225 ;
      RECT  21.34 28.7775 21.405 28.9125 ;
      RECT  21.3075 28.0975 21.4425 28.1625 ;
      RECT  21.0675 28.9775 21.2025 29.0425 ;
      RECT  21.29 28.24 21.3425 28.3025 ;
      RECT  20.8425 29.1275 20.9775 29.1925 ;
      RECT  20.72 28.3875 20.79 28.6775 ;
      RECT  20.825 28.6125 20.89 29.3525 ;
      RECT  21.34 29.2425 21.41 29.4425 ;
      RECT  20.585 28.24 20.6375 28.3025 ;
      RECT  20.58 29.4425 21.465 29.5075 ;
      RECT  21.26 28.3875 21.325 28.5225 ;
      RECT  20.6375 28.88 20.7025 29.015 ;
      RECT  21.26 28.3875 21.33 28.6775 ;
      RECT  20.955 28.0975 21.09 28.1625 ;
      RECT  20.9375 28.2375 21.0725 28.3025 ;
      RECT  21.155 28.6125 21.33 28.6775 ;
      RECT  20.64 29.2425 20.705 29.3775 ;
      RECT  20.58 28.0975 21.465 28.1625 ;
      RECT  21.3425 28.88 21.4075 29.015 ;
      RECT  20.635 28.7775 20.705 28.9125 ;
      RECT  20.905 28.3875 20.97 28.5225 ;
      RECT  21.155 28.7775 21.22 28.9125 ;
      RECT  21.0875 28.3875 21.1525 28.5225 ;
      RECT  20.64 28.7775 20.705 28.9125 ;
      RECT  21.155 29.2425 21.22 29.455 ;
      RECT  20.825 29.2425 20.89 29.3775 ;
      RECT  21.155 28.6125 21.22 29.2425 ;
      RECT  20.6025 28.0975 20.7375 28.1625 ;
      RECT  20.72 28.3875 20.785 28.5225 ;
      RECT  20.825 30.1725 20.89 30.0375 ;
      RECT  20.72 30.3375 20.89 30.2725 ;
      RECT  21.34 30.1725 21.41 30.0375 ;
      RECT  20.58 30.7125 21.465 30.6475 ;
      RECT  20.635 29.7075 20.705 29.5075 ;
      RECT  21.34 29.7075 21.405 29.5725 ;
      RECT  20.8925 30.5625 20.9575 30.4275 ;
      RECT  21.075 30.5625 21.14 30.4275 ;
      RECT  21.34 30.1725 21.405 30.0375 ;
      RECT  21.3075 30.8525 21.4425 30.7875 ;
      RECT  21.0675 29.9725 21.2025 29.9075 ;
      RECT  21.29 30.71 21.3425 30.6475 ;
      RECT  20.8425 29.8225 20.9775 29.7575 ;
      RECT  20.72 30.5625 20.79 30.2725 ;
      RECT  20.825 30.3375 20.89 29.5975 ;
      RECT  21.34 29.7075 21.41 29.5075 ;
      RECT  20.585 30.71 20.6375 30.6475 ;
      RECT  20.58 29.5075 21.465 29.4425 ;
      RECT  21.26 30.5625 21.325 30.4275 ;
      RECT  20.6375 30.07 20.7025 29.935 ;
      RECT  21.26 30.5625 21.33 30.2725 ;
      RECT  20.955 30.8525 21.09 30.7875 ;
      RECT  20.9375 30.7125 21.0725 30.6475 ;
      RECT  21.155 30.3375 21.33 30.2725 ;
      RECT  20.64 29.7075 20.705 29.5725 ;
      RECT  20.58 30.8525 21.465 30.7875 ;
      RECT  21.3425 30.07 21.4075 29.935 ;
      RECT  20.635 30.1725 20.705 30.0375 ;
      RECT  20.905 30.5625 20.97 30.4275 ;
      RECT  21.155 30.1725 21.22 30.0375 ;
      RECT  21.0875 30.5625 21.1525 30.4275 ;
      RECT  20.64 30.1725 20.705 30.0375 ;
      RECT  21.155 29.7075 21.22 29.495 ;
      RECT  20.825 29.7075 20.89 29.5725 ;
      RECT  21.155 30.3375 21.22 29.7075 ;
      RECT  20.6025 30.8525 20.7375 30.7875 ;
      RECT  20.72 30.5625 20.785 30.4275 ;
      RECT  20.825 31.4675 20.89 31.6025 ;
      RECT  20.72 31.3025 20.89 31.3675 ;
      RECT  21.34 31.4675 21.41 31.6025 ;
      RECT  20.58 30.9275 21.465 30.9925 ;
      RECT  20.635 31.9325 20.705 32.1325 ;
      RECT  21.34 31.9325 21.405 32.0675 ;
      RECT  20.8925 31.0775 20.9575 31.2125 ;
      RECT  21.075 31.0775 21.14 31.2125 ;
      RECT  21.34 31.4675 21.405 31.6025 ;
      RECT  21.3075 30.7875 21.4425 30.8525 ;
      RECT  21.0675 31.6675 21.2025 31.7325 ;
      RECT  21.29 30.93 21.3425 30.9925 ;
      RECT  20.8425 31.8175 20.9775 31.8825 ;
      RECT  20.72 31.0775 20.79 31.3675 ;
      RECT  20.825 31.3025 20.89 32.0425 ;
      RECT  21.34 31.9325 21.41 32.1325 ;
      RECT  20.585 30.93 20.6375 30.9925 ;
      RECT  20.58 32.1325 21.465 32.1975 ;
      RECT  21.26 31.0775 21.325 31.2125 ;
      RECT  20.6375 31.57 20.7025 31.705 ;
      RECT  21.26 31.0775 21.33 31.3675 ;
      RECT  20.955 30.7875 21.09 30.8525 ;
      RECT  20.9375 30.9275 21.0725 30.9925 ;
      RECT  21.155 31.3025 21.33 31.3675 ;
      RECT  20.64 31.9325 20.705 32.0675 ;
      RECT  20.58 30.7875 21.465 30.8525 ;
      RECT  21.3425 31.57 21.4075 31.705 ;
      RECT  20.635 31.4675 20.705 31.6025 ;
      RECT  20.905 31.0775 20.97 31.2125 ;
      RECT  21.155 31.4675 21.22 31.6025 ;
      RECT  21.0875 31.0775 21.1525 31.2125 ;
      RECT  20.64 31.4675 20.705 31.6025 ;
      RECT  21.155 31.9325 21.22 32.145 ;
      RECT  20.825 31.9325 20.89 32.0675 ;
      RECT  21.155 31.3025 21.22 31.9325 ;
      RECT  20.6025 30.7875 20.7375 30.8525 ;
      RECT  20.72 31.0775 20.785 31.2125 ;
      RECT  20.825 32.8625 20.89 32.7275 ;
      RECT  20.72 33.0275 20.89 32.9625 ;
      RECT  21.34 32.8625 21.41 32.7275 ;
      RECT  20.58 33.4025 21.465 33.3375 ;
      RECT  20.635 32.3975 20.705 32.1975 ;
      RECT  21.34 32.3975 21.405 32.2625 ;
      RECT  20.8925 33.2525 20.9575 33.1175 ;
      RECT  21.075 33.2525 21.14 33.1175 ;
      RECT  21.34 32.8625 21.405 32.7275 ;
      RECT  21.3075 33.5425 21.4425 33.4775 ;
      RECT  21.0675 32.6625 21.2025 32.5975 ;
      RECT  21.29 33.4 21.3425 33.3375 ;
      RECT  20.8425 32.5125 20.9775 32.4475 ;
      RECT  20.72 33.2525 20.79 32.9625 ;
      RECT  20.825 33.0275 20.89 32.2875 ;
      RECT  21.34 32.3975 21.41 32.1975 ;
      RECT  20.585 33.4 20.6375 33.3375 ;
      RECT  20.58 32.1975 21.465 32.1325 ;
      RECT  21.26 33.2525 21.325 33.1175 ;
      RECT  20.6375 32.76 20.7025 32.625 ;
      RECT  21.26 33.2525 21.33 32.9625 ;
      RECT  20.955 33.5425 21.09 33.4775 ;
      RECT  20.9375 33.4025 21.0725 33.3375 ;
      RECT  21.155 33.0275 21.33 32.9625 ;
      RECT  20.64 32.3975 20.705 32.2625 ;
      RECT  20.58 33.5425 21.465 33.4775 ;
      RECT  21.3425 32.76 21.4075 32.625 ;
      RECT  20.635 32.8625 20.705 32.7275 ;
      RECT  20.905 33.2525 20.97 33.1175 ;
      RECT  21.155 32.8625 21.22 32.7275 ;
      RECT  21.0875 33.2525 21.1525 33.1175 ;
      RECT  20.64 32.8625 20.705 32.7275 ;
      RECT  21.155 32.3975 21.22 32.185 ;
      RECT  20.825 32.3975 20.89 32.2625 ;
      RECT  21.155 33.0275 21.22 32.3975 ;
      RECT  20.6025 33.5425 20.7375 33.4775 ;
      RECT  20.72 33.2525 20.785 33.1175 ;
      RECT  20.825 34.1575 20.89 34.2925 ;
      RECT  20.72 33.9925 20.89 34.0575 ;
      RECT  21.34 34.1575 21.41 34.2925 ;
      RECT  20.58 33.6175 21.465 33.6825 ;
      RECT  20.635 34.6225 20.705 34.8225 ;
      RECT  21.34 34.6225 21.405 34.7575 ;
      RECT  20.8925 33.7675 20.9575 33.9025 ;
      RECT  21.075 33.7675 21.14 33.9025 ;
      RECT  21.34 34.1575 21.405 34.2925 ;
      RECT  21.3075 33.4775 21.4425 33.5425 ;
      RECT  21.0675 34.3575 21.2025 34.4225 ;
      RECT  21.29 33.62 21.3425 33.6825 ;
      RECT  20.8425 34.5075 20.9775 34.5725 ;
      RECT  20.72 33.7675 20.79 34.0575 ;
      RECT  20.825 33.9925 20.89 34.7325 ;
      RECT  21.34 34.6225 21.41 34.8225 ;
      RECT  20.585 33.62 20.6375 33.6825 ;
      RECT  20.58 34.8225 21.465 34.8875 ;
      RECT  21.26 33.7675 21.325 33.9025 ;
      RECT  20.6375 34.26 20.7025 34.395 ;
      RECT  21.26 33.7675 21.33 34.0575 ;
      RECT  20.955 33.4775 21.09 33.5425 ;
      RECT  20.9375 33.6175 21.0725 33.6825 ;
      RECT  21.155 33.9925 21.33 34.0575 ;
      RECT  20.64 34.6225 20.705 34.7575 ;
      RECT  20.58 33.4775 21.465 33.5425 ;
      RECT  21.3425 34.26 21.4075 34.395 ;
      RECT  20.635 34.1575 20.705 34.2925 ;
      RECT  20.905 33.7675 20.97 33.9025 ;
      RECT  21.155 34.1575 21.22 34.2925 ;
      RECT  21.0875 33.7675 21.1525 33.9025 ;
      RECT  20.64 34.1575 20.705 34.2925 ;
      RECT  21.155 34.6225 21.22 34.835 ;
      RECT  20.825 34.6225 20.89 34.7575 ;
      RECT  21.155 33.9925 21.22 34.6225 ;
      RECT  20.6025 33.4775 20.7375 33.5425 ;
      RECT  20.72 33.7675 20.785 33.9025 ;
      RECT  20.825 35.5525 20.89 35.4175 ;
      RECT  20.72 35.7175 20.89 35.6525 ;
      RECT  21.34 35.5525 21.41 35.4175 ;
      RECT  20.58 36.0925 21.465 36.0275 ;
      RECT  20.635 35.0875 20.705 34.8875 ;
      RECT  21.34 35.0875 21.405 34.9525 ;
      RECT  20.8925 35.9425 20.9575 35.8075 ;
      RECT  21.075 35.9425 21.14 35.8075 ;
      RECT  21.34 35.5525 21.405 35.4175 ;
      RECT  21.3075 36.2325 21.4425 36.1675 ;
      RECT  21.0675 35.3525 21.2025 35.2875 ;
      RECT  21.29 36.09 21.3425 36.0275 ;
      RECT  20.8425 35.2025 20.9775 35.1375 ;
      RECT  20.72 35.9425 20.79 35.6525 ;
      RECT  20.825 35.7175 20.89 34.9775 ;
      RECT  21.34 35.0875 21.41 34.8875 ;
      RECT  20.585 36.09 20.6375 36.0275 ;
      RECT  20.58 34.8875 21.465 34.8225 ;
      RECT  21.26 35.9425 21.325 35.8075 ;
      RECT  20.6375 35.45 20.7025 35.315 ;
      RECT  21.26 35.9425 21.33 35.6525 ;
      RECT  20.955 36.2325 21.09 36.1675 ;
      RECT  20.9375 36.0925 21.0725 36.0275 ;
      RECT  21.155 35.7175 21.33 35.6525 ;
      RECT  20.64 35.0875 20.705 34.9525 ;
      RECT  20.58 36.2325 21.465 36.1675 ;
      RECT  21.3425 35.45 21.4075 35.315 ;
      RECT  20.635 35.5525 20.705 35.4175 ;
      RECT  20.905 35.9425 20.97 35.8075 ;
      RECT  21.155 35.5525 21.22 35.4175 ;
      RECT  21.0875 35.9425 21.1525 35.8075 ;
      RECT  20.64 35.5525 20.705 35.4175 ;
      RECT  21.155 35.0875 21.22 34.875 ;
      RECT  20.825 35.0875 20.89 34.9525 ;
      RECT  21.155 35.7175 21.22 35.0875 ;
      RECT  20.6025 36.2325 20.7375 36.1675 ;
      RECT  20.72 35.9425 20.785 35.8075 ;
      RECT  20.825 36.8475 20.89 36.9825 ;
      RECT  20.72 36.6825 20.89 36.7475 ;
      RECT  21.34 36.8475 21.41 36.9825 ;
      RECT  20.58 36.3075 21.465 36.3725 ;
      RECT  20.635 37.3125 20.705 37.5125 ;
      RECT  21.34 37.3125 21.405 37.4475 ;
      RECT  20.8925 36.4575 20.9575 36.5925 ;
      RECT  21.075 36.4575 21.14 36.5925 ;
      RECT  21.34 36.8475 21.405 36.9825 ;
      RECT  21.3075 36.1675 21.4425 36.2325 ;
      RECT  21.0675 37.0475 21.2025 37.1125 ;
      RECT  21.29 36.31 21.3425 36.3725 ;
      RECT  20.8425 37.1975 20.9775 37.2625 ;
      RECT  20.72 36.4575 20.79 36.7475 ;
      RECT  20.825 36.6825 20.89 37.4225 ;
      RECT  21.34 37.3125 21.41 37.5125 ;
      RECT  20.585 36.31 20.6375 36.3725 ;
      RECT  20.58 37.5125 21.465 37.5775 ;
      RECT  21.26 36.4575 21.325 36.5925 ;
      RECT  20.6375 36.95 20.7025 37.085 ;
      RECT  21.26 36.4575 21.33 36.7475 ;
      RECT  20.955 36.1675 21.09 36.2325 ;
      RECT  20.9375 36.3075 21.0725 36.3725 ;
      RECT  21.155 36.6825 21.33 36.7475 ;
      RECT  20.64 37.3125 20.705 37.4475 ;
      RECT  20.58 36.1675 21.465 36.2325 ;
      RECT  21.3425 36.95 21.4075 37.085 ;
      RECT  20.635 36.8475 20.705 36.9825 ;
      RECT  20.905 36.4575 20.97 36.5925 ;
      RECT  21.155 36.8475 21.22 36.9825 ;
      RECT  21.0875 36.4575 21.1525 36.5925 ;
      RECT  20.64 36.8475 20.705 36.9825 ;
      RECT  21.155 37.3125 21.22 37.525 ;
      RECT  20.825 37.3125 20.89 37.4475 ;
      RECT  21.155 36.6825 21.22 37.3125 ;
      RECT  20.6025 36.1675 20.7375 36.2325 ;
      RECT  20.72 36.4575 20.785 36.5925 ;
      RECT  20.825 38.2425 20.89 38.1075 ;
      RECT  20.72 38.4075 20.89 38.3425 ;
      RECT  21.34 38.2425 21.41 38.1075 ;
      RECT  20.58 38.7825 21.465 38.7175 ;
      RECT  20.635 37.7775 20.705 37.5775 ;
      RECT  21.34 37.7775 21.405 37.6425 ;
      RECT  20.8925 38.6325 20.9575 38.4975 ;
      RECT  21.075 38.6325 21.14 38.4975 ;
      RECT  21.34 38.2425 21.405 38.1075 ;
      RECT  21.3075 38.9225 21.4425 38.8575 ;
      RECT  21.0675 38.0425 21.2025 37.9775 ;
      RECT  21.29 38.78 21.3425 38.7175 ;
      RECT  20.8425 37.8925 20.9775 37.8275 ;
      RECT  20.72 38.6325 20.79 38.3425 ;
      RECT  20.825 38.4075 20.89 37.6675 ;
      RECT  21.34 37.7775 21.41 37.5775 ;
      RECT  20.585 38.78 20.6375 38.7175 ;
      RECT  20.58 37.5775 21.465 37.5125 ;
      RECT  21.26 38.6325 21.325 38.4975 ;
      RECT  20.6375 38.14 20.7025 38.005 ;
      RECT  21.26 38.6325 21.33 38.3425 ;
      RECT  20.955 38.9225 21.09 38.8575 ;
      RECT  20.9375 38.7825 21.0725 38.7175 ;
      RECT  21.155 38.4075 21.33 38.3425 ;
      RECT  20.64 37.7775 20.705 37.6425 ;
      RECT  20.58 38.9225 21.465 38.8575 ;
      RECT  21.3425 38.14 21.4075 38.005 ;
      RECT  20.635 38.2425 20.705 38.1075 ;
      RECT  20.905 38.6325 20.97 38.4975 ;
      RECT  21.155 38.2425 21.22 38.1075 ;
      RECT  21.0875 38.6325 21.1525 38.4975 ;
      RECT  20.64 38.2425 20.705 38.1075 ;
      RECT  21.155 37.7775 21.22 37.565 ;
      RECT  20.825 37.7775 20.89 37.6425 ;
      RECT  21.155 38.4075 21.22 37.7775 ;
      RECT  20.6025 38.9225 20.7375 38.8575 ;
      RECT  20.72 38.6325 20.785 38.4975 ;
      RECT  20.825 39.5375 20.89 39.6725 ;
      RECT  20.72 39.3725 20.89 39.4375 ;
      RECT  21.34 39.5375 21.41 39.6725 ;
      RECT  20.58 38.9975 21.465 39.0625 ;
      RECT  20.635 40.0025 20.705 40.2025 ;
      RECT  21.34 40.0025 21.405 40.1375 ;
      RECT  20.8925 39.1475 20.9575 39.2825 ;
      RECT  21.075 39.1475 21.14 39.2825 ;
      RECT  21.34 39.5375 21.405 39.6725 ;
      RECT  21.3075 38.8575 21.4425 38.9225 ;
      RECT  21.0675 39.7375 21.2025 39.8025 ;
      RECT  21.29 39.0 21.3425 39.0625 ;
      RECT  20.8425 39.8875 20.9775 39.9525 ;
      RECT  20.72 39.1475 20.79 39.4375 ;
      RECT  20.825 39.3725 20.89 40.1125 ;
      RECT  21.34 40.0025 21.41 40.2025 ;
      RECT  20.585 39.0 20.6375 39.0625 ;
      RECT  20.58 40.2025 21.465 40.2675 ;
      RECT  21.26 39.1475 21.325 39.2825 ;
      RECT  20.6375 39.64 20.7025 39.775 ;
      RECT  21.26 39.1475 21.33 39.4375 ;
      RECT  20.955 38.8575 21.09 38.9225 ;
      RECT  20.9375 38.9975 21.0725 39.0625 ;
      RECT  21.155 39.3725 21.33 39.4375 ;
      RECT  20.64 40.0025 20.705 40.1375 ;
      RECT  20.58 38.8575 21.465 38.9225 ;
      RECT  21.3425 39.64 21.4075 39.775 ;
      RECT  20.635 39.5375 20.705 39.6725 ;
      RECT  20.905 39.1475 20.97 39.2825 ;
      RECT  21.155 39.5375 21.22 39.6725 ;
      RECT  21.0875 39.1475 21.1525 39.2825 ;
      RECT  20.64 39.5375 20.705 39.6725 ;
      RECT  21.155 40.0025 21.22 40.215 ;
      RECT  20.825 40.0025 20.89 40.1375 ;
      RECT  21.155 39.3725 21.22 40.0025 ;
      RECT  20.6025 38.8575 20.7375 38.9225 ;
      RECT  20.72 39.1475 20.785 39.2825 ;
      RECT  20.825 40.9325 20.89 40.7975 ;
      RECT  20.72 41.0975 20.89 41.0325 ;
      RECT  21.34 40.9325 21.41 40.7975 ;
      RECT  20.58 41.4725 21.465 41.4075 ;
      RECT  20.635 40.4675 20.705 40.2675 ;
      RECT  21.34 40.4675 21.405 40.3325 ;
      RECT  20.8925 41.3225 20.9575 41.1875 ;
      RECT  21.075 41.3225 21.14 41.1875 ;
      RECT  21.34 40.9325 21.405 40.7975 ;
      RECT  21.3075 41.6125 21.4425 41.5475 ;
      RECT  21.0675 40.7325 21.2025 40.6675 ;
      RECT  21.29 41.47 21.3425 41.4075 ;
      RECT  20.8425 40.5825 20.9775 40.5175 ;
      RECT  20.72 41.3225 20.79 41.0325 ;
      RECT  20.825 41.0975 20.89 40.3575 ;
      RECT  21.34 40.4675 21.41 40.2675 ;
      RECT  20.585 41.47 20.6375 41.4075 ;
      RECT  20.58 40.2675 21.465 40.2025 ;
      RECT  21.26 41.3225 21.325 41.1875 ;
      RECT  20.6375 40.83 20.7025 40.695 ;
      RECT  21.26 41.3225 21.33 41.0325 ;
      RECT  20.955 41.6125 21.09 41.5475 ;
      RECT  20.9375 41.4725 21.0725 41.4075 ;
      RECT  21.155 41.0975 21.33 41.0325 ;
      RECT  20.64 40.4675 20.705 40.3325 ;
      RECT  20.58 41.6125 21.465 41.5475 ;
      RECT  21.3425 40.83 21.4075 40.695 ;
      RECT  20.635 40.9325 20.705 40.7975 ;
      RECT  20.905 41.3225 20.97 41.1875 ;
      RECT  21.155 40.9325 21.22 40.7975 ;
      RECT  21.0875 41.3225 21.1525 41.1875 ;
      RECT  20.64 40.9325 20.705 40.7975 ;
      RECT  21.155 40.4675 21.22 40.255 ;
      RECT  20.825 40.4675 20.89 40.3325 ;
      RECT  21.155 41.0975 21.22 40.4675 ;
      RECT  20.6025 41.6125 20.7375 41.5475 ;
      RECT  20.72 41.3225 20.785 41.1875 ;
      RECT  20.825 42.2275 20.89 42.3625 ;
      RECT  20.72 42.0625 20.89 42.1275 ;
      RECT  21.34 42.2275 21.41 42.3625 ;
      RECT  20.58 41.6875 21.465 41.7525 ;
      RECT  20.635 42.6925 20.705 42.8925 ;
      RECT  21.34 42.6925 21.405 42.8275 ;
      RECT  20.8925 41.8375 20.9575 41.9725 ;
      RECT  21.075 41.8375 21.14 41.9725 ;
      RECT  21.34 42.2275 21.405 42.3625 ;
      RECT  21.3075 41.5475 21.4425 41.6125 ;
      RECT  21.0675 42.4275 21.2025 42.4925 ;
      RECT  21.29 41.69 21.3425 41.7525 ;
      RECT  20.8425 42.5775 20.9775 42.6425 ;
      RECT  20.72 41.8375 20.79 42.1275 ;
      RECT  20.825 42.0625 20.89 42.8025 ;
      RECT  21.34 42.6925 21.41 42.8925 ;
      RECT  20.585 41.69 20.6375 41.7525 ;
      RECT  20.58 42.8925 21.465 42.9575 ;
      RECT  21.26 41.8375 21.325 41.9725 ;
      RECT  20.6375 42.33 20.7025 42.465 ;
      RECT  21.26 41.8375 21.33 42.1275 ;
      RECT  20.955 41.5475 21.09 41.6125 ;
      RECT  20.9375 41.6875 21.0725 41.7525 ;
      RECT  21.155 42.0625 21.33 42.1275 ;
      RECT  20.64 42.6925 20.705 42.8275 ;
      RECT  20.58 41.5475 21.465 41.6125 ;
      RECT  21.3425 42.33 21.4075 42.465 ;
      RECT  20.635 42.2275 20.705 42.3625 ;
      RECT  20.905 41.8375 20.97 41.9725 ;
      RECT  21.155 42.2275 21.22 42.3625 ;
      RECT  21.0875 41.8375 21.1525 41.9725 ;
      RECT  20.64 42.2275 20.705 42.3625 ;
      RECT  21.155 42.6925 21.22 42.905 ;
      RECT  20.825 42.6925 20.89 42.8275 ;
      RECT  21.155 42.0625 21.22 42.6925 ;
      RECT  20.6025 41.5475 20.7375 41.6125 ;
      RECT  20.72 41.8375 20.785 41.9725 ;
      RECT  20.825 43.6225 20.89 43.4875 ;
      RECT  20.72 43.7875 20.89 43.7225 ;
      RECT  21.34 43.6225 21.41 43.4875 ;
      RECT  20.58 44.1625 21.465 44.0975 ;
      RECT  20.635 43.1575 20.705 42.9575 ;
      RECT  21.34 43.1575 21.405 43.0225 ;
      RECT  20.8925 44.0125 20.9575 43.8775 ;
      RECT  21.075 44.0125 21.14 43.8775 ;
      RECT  21.34 43.6225 21.405 43.4875 ;
      RECT  21.3075 44.3025 21.4425 44.2375 ;
      RECT  21.0675 43.4225 21.2025 43.3575 ;
      RECT  21.29 44.16 21.3425 44.0975 ;
      RECT  20.8425 43.2725 20.9775 43.2075 ;
      RECT  20.72 44.0125 20.79 43.7225 ;
      RECT  20.825 43.7875 20.89 43.0475 ;
      RECT  21.34 43.1575 21.41 42.9575 ;
      RECT  20.585 44.16 20.6375 44.0975 ;
      RECT  20.58 42.9575 21.465 42.8925 ;
      RECT  21.26 44.0125 21.325 43.8775 ;
      RECT  20.6375 43.52 20.7025 43.385 ;
      RECT  21.26 44.0125 21.33 43.7225 ;
      RECT  20.955 44.3025 21.09 44.2375 ;
      RECT  20.9375 44.1625 21.0725 44.0975 ;
      RECT  21.155 43.7875 21.33 43.7225 ;
      RECT  20.64 43.1575 20.705 43.0225 ;
      RECT  20.58 44.3025 21.465 44.2375 ;
      RECT  21.3425 43.52 21.4075 43.385 ;
      RECT  20.635 43.6225 20.705 43.4875 ;
      RECT  20.905 44.0125 20.97 43.8775 ;
      RECT  21.155 43.6225 21.22 43.4875 ;
      RECT  21.0875 44.0125 21.1525 43.8775 ;
      RECT  20.64 43.6225 20.705 43.4875 ;
      RECT  21.155 43.1575 21.22 42.945 ;
      RECT  20.825 43.1575 20.89 43.0225 ;
      RECT  21.155 43.7875 21.22 43.1575 ;
      RECT  20.6025 44.3025 20.7375 44.2375 ;
      RECT  20.72 44.0125 20.785 43.8775 ;
      RECT  20.825 44.9175 20.89 45.0525 ;
      RECT  21.34 44.9175 21.41 45.0525 ;
      RECT  20.72 44.7525 20.89 44.8175 ;
      RECT  20.58 44.3775 21.465 44.4425 ;
      RECT  20.635 45.3825 20.705 45.5825 ;
      RECT  21.34 45.3825 21.405 45.5175 ;
      RECT  20.8925 44.5275 20.9575 44.6625 ;
      RECT  21.075 44.5275 21.14 44.6625 ;
      RECT  21.34 44.9175 21.405 45.0525 ;
      RECT  21.3075 44.2375 21.4425 44.3025 ;
      RECT  21.0675 45.1175 21.2025 45.1825 ;
      RECT  21.29 44.38 21.3425 44.4425 ;
      RECT  20.8425 45.2675 20.9775 45.3325 ;
      RECT  20.72 44.5275 20.79 44.8175 ;
      RECT  20.825 44.7525 20.89 45.4925 ;
      RECT  21.34 45.3825 21.41 45.5825 ;
      RECT  21.26 44.5275 21.325 44.6625 ;
      RECT  20.585 44.38 20.6375 44.4425 ;
      RECT  20.58 45.5825 21.465 45.6475 ;
      RECT  20.6375 45.02 20.7025 45.155 ;
      RECT  20.955 44.2375 21.09 44.3025 ;
      RECT  21.26 44.5275 21.33 44.8175 ;
      RECT  20.9375 44.3775 21.0725 44.4425 ;
      RECT  20.64 45.3825 20.705 45.5175 ;
      RECT  21.155 44.7525 21.33 44.8175 ;
      RECT  21.155 45.3825 21.22 45.5175 ;
      RECT  20.58 44.2375 21.465 44.3025 ;
      RECT  21.3425 45.02 21.4075 45.155 ;
      RECT  20.635 44.9175 20.705 45.0525 ;
      RECT  20.905 44.5275 20.97 44.6625 ;
      RECT  21.155 44.9175 21.22 45.0525 ;
      RECT  21.0875 44.5275 21.1525 44.6625 ;
      RECT  20.64 44.9175 20.705 45.0525 ;
      RECT  20.825 45.3825 20.89 45.5175 ;
      RECT  21.155 44.7525 21.22 45.3825 ;
      RECT  20.6025 44.2375 20.7375 44.3025 ;
      RECT  20.72 44.5275 20.785 44.6625 ;
      RECT  20.67 20.1675 21.375 20.2325 ;
      RECT  20.67 22.5775 21.375 22.6425 ;
      RECT  20.67 22.8575 21.375 22.9225 ;
      RECT  20.67 25.2675 21.375 25.3325 ;
      RECT  20.67 25.5475 21.375 25.6125 ;
      RECT  20.67 27.9575 21.375 28.0225 ;
      RECT  20.67 28.2375 21.375 28.3025 ;
      RECT  20.67 30.6475 21.375 30.7125 ;
      RECT  20.67 30.9275 21.375 30.9925 ;
      RECT  20.67 33.3375 21.375 33.4025 ;
      RECT  20.67 33.6175 21.375 33.6825 ;
      RECT  20.67 36.0275 21.375 36.0925 ;
      RECT  20.67 36.3075 21.375 36.3725 ;
      RECT  20.67 38.7175 21.375 38.7825 ;
      RECT  20.67 38.9975 21.375 39.0625 ;
      RECT  20.67 41.4075 21.375 41.4725 ;
      RECT  20.67 41.6875 21.375 41.7525 ;
      RECT  20.67 44.0975 21.375 44.1625 ;
      RECT  20.67 44.3775 21.375 44.4425 ;
      RECT  21.53 22.1025 21.595 21.9675 ;
      RECT  22.045 22.1025 22.115 21.9675 ;
      RECT  21.425 22.2675 21.595 22.2025 ;
      RECT  21.285 22.6425 22.17 22.5775 ;
      RECT  21.34 21.6375 21.41 21.4375 ;
      RECT  22.045 21.6375 22.11 21.5025 ;
      RECT  21.5975 22.4925 21.6625 22.3575 ;
      RECT  21.78 22.4925 21.845 22.3575 ;
      RECT  22.045 22.1025 22.11 21.9675 ;
      RECT  22.0125 22.7825 22.1475 22.7175 ;
      RECT  21.7725 21.9025 21.9075 21.8375 ;
      RECT  21.995 22.64 22.0475 22.5775 ;
      RECT  21.5475 21.7525 21.6825 21.6875 ;
      RECT  21.425 22.4925 21.495 22.2025 ;
      RECT  21.53 22.2675 21.595 21.5275 ;
      RECT  22.045 21.6375 22.115 21.4375 ;
      RECT  21.965 22.4925 22.03 22.3575 ;
      RECT  21.29 22.64 21.3425 22.5775 ;
      RECT  21.285 21.4375 22.17 21.3725 ;
      RECT  21.3425 22.0 21.4075 21.865 ;
      RECT  21.66 22.7825 21.795 22.7175 ;
      RECT  21.965 22.4925 22.035 22.2025 ;
      RECT  21.6425 22.6425 21.7775 22.5775 ;
      RECT  21.345 21.6375 21.41 21.5025 ;
      RECT  21.86 22.2675 22.035 22.2025 ;
      RECT  21.86 21.6375 21.925 21.5025 ;
      RECT  21.285 22.7825 22.17 22.7175 ;
      RECT  22.0475 22.0 22.1125 21.865 ;
      RECT  21.34 22.1025 21.41 21.9675 ;
      RECT  21.61 22.4925 21.675 22.3575 ;
      RECT  21.86 22.1025 21.925 21.9675 ;
      RECT  21.7925 22.4925 21.8575 22.3575 ;
      RECT  21.345 22.1025 21.41 21.9675 ;
      RECT  21.53 21.6375 21.595 21.5025 ;
      RECT  21.86 22.2675 21.925 21.6375 ;
      RECT  21.3075 22.7825 21.4425 22.7175 ;
      RECT  21.425 22.4925 21.49 22.3575 ;
      RECT  22.235 22.1025 22.3 21.9675 ;
      RECT  22.75 22.1025 22.82 21.9675 ;
      RECT  22.13 22.2675 22.3 22.2025 ;
      RECT  21.99 22.6425 22.875 22.5775 ;
      RECT  22.045 21.6375 22.115 21.4375 ;
      RECT  22.75 21.6375 22.815 21.5025 ;
      RECT  22.3025 22.4925 22.3675 22.3575 ;
      RECT  22.485 22.4925 22.55 22.3575 ;
      RECT  22.75 22.1025 22.815 21.9675 ;
      RECT  22.7175 22.7825 22.8525 22.7175 ;
      RECT  22.4775 21.9025 22.6125 21.8375 ;
      RECT  22.7 22.64 22.7525 22.5775 ;
      RECT  22.2525 21.7525 22.3875 21.6875 ;
      RECT  22.13 22.4925 22.2 22.2025 ;
      RECT  22.235 22.2675 22.3 21.5275 ;
      RECT  22.75 21.6375 22.82 21.4375 ;
      RECT  22.67 22.4925 22.735 22.3575 ;
      RECT  21.995 22.64 22.0475 22.5775 ;
      RECT  21.99 21.4375 22.875 21.3725 ;
      RECT  22.0475 22.0 22.1125 21.865 ;
      RECT  22.365 22.7825 22.5 22.7175 ;
      RECT  22.67 22.4925 22.74 22.2025 ;
      RECT  22.3475 22.6425 22.4825 22.5775 ;
      RECT  22.05 21.6375 22.115 21.5025 ;
      RECT  22.565 22.2675 22.74 22.2025 ;
      RECT  22.565 21.6375 22.63 21.5025 ;
      RECT  21.99 22.7825 22.875 22.7175 ;
      RECT  22.7525 22.0 22.8175 21.865 ;
      RECT  22.045 22.1025 22.115 21.9675 ;
      RECT  22.315 22.4925 22.38 22.3575 ;
      RECT  22.565 22.1025 22.63 21.9675 ;
      RECT  22.4975 22.4925 22.5625 22.3575 ;
      RECT  22.05 22.1025 22.115 21.9675 ;
      RECT  22.235 21.6375 22.3 21.5025 ;
      RECT  22.565 22.2675 22.63 21.6375 ;
      RECT  22.0125 22.7825 22.1475 22.7175 ;
      RECT  22.13 22.4925 22.195 22.3575 ;
      RECT  21.375 22.6425 22.785 22.5775 ;
      RECT  21.53 20.7075 21.595 20.8425 ;
      RECT  22.045 20.7075 22.115 20.8425 ;
      RECT  21.425 20.5425 21.595 20.6075 ;
      RECT  21.285 20.1675 22.17 20.2325 ;
      RECT  21.34 21.1725 21.41 21.3725 ;
      RECT  22.045 21.1725 22.11 21.3075 ;
      RECT  21.5975 20.3175 21.6625 20.4525 ;
      RECT  21.78 20.3175 21.845 20.4525 ;
      RECT  22.045 20.7075 22.11 20.8425 ;
      RECT  22.0125 20.0275 22.1475 20.0925 ;
      RECT  21.7725 20.9075 21.9075 20.9725 ;
      RECT  21.995 20.17 22.0475 20.2325 ;
      RECT  21.5475 21.0575 21.6825 21.1225 ;
      RECT  21.425 20.3175 21.495 20.6075 ;
      RECT  21.53 20.5425 21.595 21.2825 ;
      RECT  22.045 21.1725 22.115 21.3725 ;
      RECT  21.965 20.3175 22.03 20.4525 ;
      RECT  21.29 20.17 21.3425 20.2325 ;
      RECT  21.285 21.3725 22.17 21.4375 ;
      RECT  21.3425 20.81 21.4075 20.945 ;
      RECT  21.66 20.0275 21.795 20.0925 ;
      RECT  21.965 20.3175 22.035 20.6075 ;
      RECT  21.6425 20.1675 21.7775 20.2325 ;
      RECT  21.345 21.1725 21.41 21.3075 ;
      RECT  21.86 20.5425 22.035 20.6075 ;
      RECT  21.86 21.1725 21.925 21.3075 ;
      RECT  21.285 20.0275 22.17 20.0925 ;
      RECT  22.0475 20.81 22.1125 20.945 ;
      RECT  21.34 20.7075 21.41 20.8425 ;
      RECT  21.61 20.3175 21.675 20.4525 ;
      RECT  21.86 20.7075 21.925 20.8425 ;
      RECT  21.7925 20.3175 21.8575 20.4525 ;
      RECT  21.345 20.7075 21.41 20.8425 ;
      RECT  21.53 21.1725 21.595 21.3075 ;
      RECT  21.86 20.5425 21.925 21.1725 ;
      RECT  21.3075 20.0275 21.4425 20.0925 ;
      RECT  21.425 20.3175 21.49 20.4525 ;
      RECT  22.235 20.7075 22.3 20.8425 ;
      RECT  22.75 20.7075 22.82 20.8425 ;
      RECT  22.13 20.5425 22.3 20.6075 ;
      RECT  21.99 20.1675 22.875 20.2325 ;
      RECT  22.045 21.1725 22.115 21.3725 ;
      RECT  22.75 21.1725 22.815 21.3075 ;
      RECT  22.3025 20.3175 22.3675 20.4525 ;
      RECT  22.485 20.3175 22.55 20.4525 ;
      RECT  22.75 20.7075 22.815 20.8425 ;
      RECT  22.7175 20.0275 22.8525 20.0925 ;
      RECT  22.4775 20.9075 22.6125 20.9725 ;
      RECT  22.7 20.17 22.7525 20.2325 ;
      RECT  22.2525 21.0575 22.3875 21.1225 ;
      RECT  22.13 20.3175 22.2 20.6075 ;
      RECT  22.235 20.5425 22.3 21.2825 ;
      RECT  22.75 21.1725 22.82 21.3725 ;
      RECT  22.67 20.3175 22.735 20.4525 ;
      RECT  21.995 20.17 22.0475 20.2325 ;
      RECT  21.99 21.3725 22.875 21.4375 ;
      RECT  22.0475 20.81 22.1125 20.945 ;
      RECT  22.365 20.0275 22.5 20.0925 ;
      RECT  22.67 20.3175 22.74 20.6075 ;
      RECT  22.3475 20.1675 22.4825 20.2325 ;
      RECT  22.05 21.1725 22.115 21.3075 ;
      RECT  22.565 20.5425 22.74 20.6075 ;
      RECT  22.565 21.1725 22.63 21.3075 ;
      RECT  21.99 20.0275 22.875 20.0925 ;
      RECT  22.7525 20.81 22.8175 20.945 ;
      RECT  22.045 20.7075 22.115 20.8425 ;
      RECT  22.315 20.3175 22.38 20.4525 ;
      RECT  22.565 20.7075 22.63 20.8425 ;
      RECT  22.4975 20.3175 22.5625 20.4525 ;
      RECT  22.05 20.7075 22.115 20.8425 ;
      RECT  22.235 21.1725 22.3 21.3075 ;
      RECT  22.565 20.5425 22.63 21.1725 ;
      RECT  22.0125 20.0275 22.1475 20.0925 ;
      RECT  22.13 20.3175 22.195 20.4525 ;
      RECT  21.375 20.1675 22.785 20.2325 ;
      RECT  21.53 44.9175 21.595 45.0525 ;
      RECT  22.045 44.9175 22.115 45.0525 ;
      RECT  21.425 44.7525 21.595 44.8175 ;
      RECT  21.285 44.3775 22.17 44.4425 ;
      RECT  21.34 45.3825 21.41 45.5825 ;
      RECT  22.045 45.3825 22.11 45.5175 ;
      RECT  21.5975 44.5275 21.6625 44.6625 ;
      RECT  21.78 44.5275 21.845 44.6625 ;
      RECT  22.045 44.9175 22.11 45.0525 ;
      RECT  22.0125 44.2375 22.1475 44.3025 ;
      RECT  21.7725 45.1175 21.9075 45.1825 ;
      RECT  21.995 44.38 22.0475 44.4425 ;
      RECT  21.5475 45.2675 21.6825 45.3325 ;
      RECT  21.425 44.5275 21.495 44.8175 ;
      RECT  21.53 44.7525 21.595 45.4925 ;
      RECT  22.045 45.3825 22.115 45.5825 ;
      RECT  21.965 44.5275 22.03 44.6625 ;
      RECT  21.29 44.38 21.3425 44.4425 ;
      RECT  21.285 45.5825 22.17 45.6475 ;
      RECT  21.3425 45.02 21.4075 45.155 ;
      RECT  21.66 44.2375 21.795 44.3025 ;
      RECT  21.965 44.5275 22.035 44.8175 ;
      RECT  21.6425 44.3775 21.7775 44.4425 ;
      RECT  21.345 45.3825 21.41 45.5175 ;
      RECT  21.86 44.7525 22.035 44.8175 ;
      RECT  21.86 45.3825 21.925 45.5175 ;
      RECT  21.285 44.2375 22.17 44.3025 ;
      RECT  22.0475 45.02 22.1125 45.155 ;
      RECT  21.34 44.9175 21.41 45.0525 ;
      RECT  21.61 44.5275 21.675 44.6625 ;
      RECT  21.86 44.9175 21.925 45.0525 ;
      RECT  21.7925 44.5275 21.8575 44.6625 ;
      RECT  21.345 44.9175 21.41 45.0525 ;
      RECT  21.53 45.3825 21.595 45.5175 ;
      RECT  21.86 44.7525 21.925 45.3825 ;
      RECT  21.3075 44.2375 21.4425 44.3025 ;
      RECT  21.425 44.5275 21.49 44.6625 ;
      RECT  22.235 44.9175 22.3 45.0525 ;
      RECT  22.75 44.9175 22.82 45.0525 ;
      RECT  22.13 44.7525 22.3 44.8175 ;
      RECT  21.99 44.3775 22.875 44.4425 ;
      RECT  22.045 45.3825 22.115 45.5825 ;
      RECT  22.75 45.3825 22.815 45.5175 ;
      RECT  22.3025 44.5275 22.3675 44.6625 ;
      RECT  22.485 44.5275 22.55 44.6625 ;
      RECT  22.75 44.9175 22.815 45.0525 ;
      RECT  22.7175 44.2375 22.8525 44.3025 ;
      RECT  22.4775 45.1175 22.6125 45.1825 ;
      RECT  22.7 44.38 22.7525 44.4425 ;
      RECT  22.2525 45.2675 22.3875 45.3325 ;
      RECT  22.13 44.5275 22.2 44.8175 ;
      RECT  22.235 44.7525 22.3 45.4925 ;
      RECT  22.75 45.3825 22.82 45.5825 ;
      RECT  22.67 44.5275 22.735 44.6625 ;
      RECT  21.995 44.38 22.0475 44.4425 ;
      RECT  21.99 45.5825 22.875 45.6475 ;
      RECT  22.0475 45.02 22.1125 45.155 ;
      RECT  22.365 44.2375 22.5 44.3025 ;
      RECT  22.67 44.5275 22.74 44.8175 ;
      RECT  22.3475 44.3775 22.4825 44.4425 ;
      RECT  22.05 45.3825 22.115 45.5175 ;
      RECT  22.565 44.7525 22.74 44.8175 ;
      RECT  22.565 45.3825 22.63 45.5175 ;
      RECT  21.99 44.2375 22.875 44.3025 ;
      RECT  22.7525 45.02 22.8175 45.155 ;
      RECT  22.045 44.9175 22.115 45.0525 ;
      RECT  22.315 44.5275 22.38 44.6625 ;
      RECT  22.565 44.9175 22.63 45.0525 ;
      RECT  22.4975 44.5275 22.5625 44.6625 ;
      RECT  22.05 44.9175 22.115 45.0525 ;
      RECT  22.235 45.3825 22.3 45.5175 ;
      RECT  22.565 44.7525 22.63 45.3825 ;
      RECT  22.0125 44.2375 22.1475 44.3025 ;
      RECT  22.13 44.5275 22.195 44.6625 ;
      RECT  21.375 44.3775 22.785 44.4425 ;
      RECT  20.12 20.7075 20.185 20.8425 ;
      RECT  20.635 20.7075 20.705 20.8425 ;
      RECT  20.015 20.5425 20.185 20.6075 ;
      RECT  19.875 20.1675 20.76 20.2325 ;
      RECT  19.93 21.1725 20.0 21.3725 ;
      RECT  20.635 21.1725 20.7 21.3075 ;
      RECT  20.1875 20.3175 20.2525 20.4525 ;
      RECT  20.37 20.3175 20.435 20.4525 ;
      RECT  20.635 20.7075 20.7 20.8425 ;
      RECT  20.6025 20.0275 20.7375 20.0925 ;
      RECT  20.3625 20.9075 20.4975 20.9725 ;
      RECT  20.585 20.17 20.6375 20.2325 ;
      RECT  20.1375 21.0575 20.2725 21.1225 ;
      RECT  20.015 20.3175 20.085 20.6075 ;
      RECT  20.12 20.5425 20.185 21.2825 ;
      RECT  20.635 21.1725 20.705 21.3725 ;
      RECT  20.555 20.3175 20.62 20.4525 ;
      RECT  19.88 20.17 19.9325 20.2325 ;
      RECT  19.875 21.3725 20.76 21.4375 ;
      RECT  19.9325 20.81 19.9975 20.945 ;
      RECT  20.25 20.0275 20.385 20.0925 ;
      RECT  20.555 20.3175 20.625 20.6075 ;
      RECT  20.2325 20.1675 20.3675 20.2325 ;
      RECT  19.935 21.1725 20.0 21.3075 ;
      RECT  20.45 20.5425 20.625 20.6075 ;
      RECT  20.45 21.1725 20.515 21.3075 ;
      RECT  19.875 20.0275 20.76 20.0925 ;
      RECT  20.6375 20.81 20.7025 20.945 ;
      RECT  19.93 20.7075 20.0 20.8425 ;
      RECT  20.2 20.3175 20.265 20.4525 ;
      RECT  20.45 20.7075 20.515 20.8425 ;
      RECT  20.3825 20.3175 20.4475 20.4525 ;
      RECT  19.935 20.7075 20.0 20.8425 ;
      RECT  20.12 21.1725 20.185 21.3075 ;
      RECT  20.45 20.5425 20.515 21.1725 ;
      RECT  19.8975 20.0275 20.0325 20.0925 ;
      RECT  20.015 20.3175 20.08 20.4525 ;
      RECT  20.12 22.1025 20.185 21.9675 ;
      RECT  20.635 22.1025 20.705 21.9675 ;
      RECT  20.015 22.2675 20.185 22.2025 ;
      RECT  19.875 22.6425 20.76 22.5775 ;
      RECT  19.93 21.6375 20.0 21.4375 ;
      RECT  20.635 21.6375 20.7 21.5025 ;
      RECT  20.1875 22.4925 20.2525 22.3575 ;
      RECT  20.37 22.4925 20.435 22.3575 ;
      RECT  20.635 22.1025 20.7 21.9675 ;
      RECT  20.6025 22.7825 20.7375 22.7175 ;
      RECT  20.3625 21.9025 20.4975 21.8375 ;
      RECT  20.585 22.64 20.6375 22.5775 ;
      RECT  20.1375 21.7525 20.2725 21.6875 ;
      RECT  20.015 22.4925 20.085 22.2025 ;
      RECT  20.12 22.2675 20.185 21.5275 ;
      RECT  20.635 21.6375 20.705 21.4375 ;
      RECT  20.555 22.4925 20.62 22.3575 ;
      RECT  19.88 22.64 19.9325 22.5775 ;
      RECT  19.875 21.4375 20.76 21.3725 ;
      RECT  19.9325 22.0 19.9975 21.865 ;
      RECT  20.25 22.7825 20.385 22.7175 ;
      RECT  20.555 22.4925 20.625 22.2025 ;
      RECT  20.2325 22.6425 20.3675 22.5775 ;
      RECT  19.935 21.6375 20.0 21.5025 ;
      RECT  20.45 22.2675 20.625 22.2025 ;
      RECT  20.45 21.6375 20.515 21.5025 ;
      RECT  19.875 22.7825 20.76 22.7175 ;
      RECT  20.6375 22.0 20.7025 21.865 ;
      RECT  19.93 22.1025 20.0 21.9675 ;
      RECT  20.2 22.4925 20.265 22.3575 ;
      RECT  20.45 22.1025 20.515 21.9675 ;
      RECT  20.3825 22.4925 20.4475 22.3575 ;
      RECT  19.935 22.1025 20.0 21.9675 ;
      RECT  20.12 21.6375 20.185 21.5025 ;
      RECT  20.45 22.2675 20.515 21.6375 ;
      RECT  19.8975 22.7825 20.0325 22.7175 ;
      RECT  20.015 22.4925 20.08 22.3575 ;
      RECT  20.12 23.3975 20.185 23.5325 ;
      RECT  20.635 23.3975 20.705 23.5325 ;
      RECT  20.015 23.2325 20.185 23.2975 ;
      RECT  19.875 22.8575 20.76 22.9225 ;
      RECT  19.93 23.8625 20.0 24.0625 ;
      RECT  20.635 23.8625 20.7 23.9975 ;
      RECT  20.1875 23.0075 20.2525 23.1425 ;
      RECT  20.37 23.0075 20.435 23.1425 ;
      RECT  20.635 23.3975 20.7 23.5325 ;
      RECT  20.6025 22.7175 20.7375 22.7825 ;
      RECT  20.3625 23.5975 20.4975 23.6625 ;
      RECT  20.585 22.86 20.6375 22.9225 ;
      RECT  20.1375 23.7475 20.2725 23.8125 ;
      RECT  20.015 23.0075 20.085 23.2975 ;
      RECT  20.12 23.2325 20.185 23.9725 ;
      RECT  20.635 23.8625 20.705 24.0625 ;
      RECT  20.555 23.0075 20.62 23.1425 ;
      RECT  19.88 22.86 19.9325 22.9225 ;
      RECT  19.875 24.0625 20.76 24.1275 ;
      RECT  19.9325 23.5 19.9975 23.635 ;
      RECT  20.25 22.7175 20.385 22.7825 ;
      RECT  20.555 23.0075 20.625 23.2975 ;
      RECT  20.2325 22.8575 20.3675 22.9225 ;
      RECT  19.935 23.8625 20.0 23.9975 ;
      RECT  20.45 23.2325 20.625 23.2975 ;
      RECT  20.45 23.8625 20.515 23.9975 ;
      RECT  19.875 22.7175 20.76 22.7825 ;
      RECT  20.6375 23.5 20.7025 23.635 ;
      RECT  19.93 23.3975 20.0 23.5325 ;
      RECT  20.2 23.0075 20.265 23.1425 ;
      RECT  20.45 23.3975 20.515 23.5325 ;
      RECT  20.3825 23.0075 20.4475 23.1425 ;
      RECT  19.935 23.3975 20.0 23.5325 ;
      RECT  20.12 23.8625 20.185 23.9975 ;
      RECT  20.45 23.2325 20.515 23.8625 ;
      RECT  19.8975 22.7175 20.0325 22.7825 ;
      RECT  20.015 23.0075 20.08 23.1425 ;
      RECT  20.12 24.7925 20.185 24.6575 ;
      RECT  20.635 24.7925 20.705 24.6575 ;
      RECT  20.015 24.9575 20.185 24.8925 ;
      RECT  19.875 25.3325 20.76 25.2675 ;
      RECT  19.93 24.3275 20.0 24.1275 ;
      RECT  20.635 24.3275 20.7 24.1925 ;
      RECT  20.1875 25.1825 20.2525 25.0475 ;
      RECT  20.37 25.1825 20.435 25.0475 ;
      RECT  20.635 24.7925 20.7 24.6575 ;
      RECT  20.6025 25.4725 20.7375 25.4075 ;
      RECT  20.3625 24.5925 20.4975 24.5275 ;
      RECT  20.585 25.33 20.6375 25.2675 ;
      RECT  20.1375 24.4425 20.2725 24.3775 ;
      RECT  20.015 25.1825 20.085 24.8925 ;
      RECT  20.12 24.9575 20.185 24.2175 ;
      RECT  20.635 24.3275 20.705 24.1275 ;
      RECT  20.555 25.1825 20.62 25.0475 ;
      RECT  19.88 25.33 19.9325 25.2675 ;
      RECT  19.875 24.1275 20.76 24.0625 ;
      RECT  19.9325 24.69 19.9975 24.555 ;
      RECT  20.25 25.4725 20.385 25.4075 ;
      RECT  20.555 25.1825 20.625 24.8925 ;
      RECT  20.2325 25.3325 20.3675 25.2675 ;
      RECT  19.935 24.3275 20.0 24.1925 ;
      RECT  20.45 24.9575 20.625 24.8925 ;
      RECT  20.45 24.3275 20.515 24.1925 ;
      RECT  19.875 25.4725 20.76 25.4075 ;
      RECT  20.6375 24.69 20.7025 24.555 ;
      RECT  19.93 24.7925 20.0 24.6575 ;
      RECT  20.2 25.1825 20.265 25.0475 ;
      RECT  20.45 24.7925 20.515 24.6575 ;
      RECT  20.3825 25.1825 20.4475 25.0475 ;
      RECT  19.935 24.7925 20.0 24.6575 ;
      RECT  20.12 24.3275 20.185 24.1925 ;
      RECT  20.45 24.9575 20.515 24.3275 ;
      RECT  19.8975 25.4725 20.0325 25.4075 ;
      RECT  20.015 25.1825 20.08 25.0475 ;
      RECT  20.12 26.0875 20.185 26.2225 ;
      RECT  20.635 26.0875 20.705 26.2225 ;
      RECT  20.015 25.9225 20.185 25.9875 ;
      RECT  19.875 25.5475 20.76 25.6125 ;
      RECT  19.93 26.5525 20.0 26.7525 ;
      RECT  20.635 26.5525 20.7 26.6875 ;
      RECT  20.1875 25.6975 20.2525 25.8325 ;
      RECT  20.37 25.6975 20.435 25.8325 ;
      RECT  20.635 26.0875 20.7 26.2225 ;
      RECT  20.6025 25.4075 20.7375 25.4725 ;
      RECT  20.3625 26.2875 20.4975 26.3525 ;
      RECT  20.585 25.55 20.6375 25.6125 ;
      RECT  20.1375 26.4375 20.2725 26.5025 ;
      RECT  20.015 25.6975 20.085 25.9875 ;
      RECT  20.12 25.9225 20.185 26.6625 ;
      RECT  20.635 26.5525 20.705 26.7525 ;
      RECT  20.555 25.6975 20.62 25.8325 ;
      RECT  19.88 25.55 19.9325 25.6125 ;
      RECT  19.875 26.7525 20.76 26.8175 ;
      RECT  19.9325 26.19 19.9975 26.325 ;
      RECT  20.25 25.4075 20.385 25.4725 ;
      RECT  20.555 25.6975 20.625 25.9875 ;
      RECT  20.2325 25.5475 20.3675 25.6125 ;
      RECT  19.935 26.5525 20.0 26.6875 ;
      RECT  20.45 25.9225 20.625 25.9875 ;
      RECT  20.45 26.5525 20.515 26.6875 ;
      RECT  19.875 25.4075 20.76 25.4725 ;
      RECT  20.6375 26.19 20.7025 26.325 ;
      RECT  19.93 26.0875 20.0 26.2225 ;
      RECT  20.2 25.6975 20.265 25.8325 ;
      RECT  20.45 26.0875 20.515 26.2225 ;
      RECT  20.3825 25.6975 20.4475 25.8325 ;
      RECT  19.935 26.0875 20.0 26.2225 ;
      RECT  20.12 26.5525 20.185 26.6875 ;
      RECT  20.45 25.9225 20.515 26.5525 ;
      RECT  19.8975 25.4075 20.0325 25.4725 ;
      RECT  20.015 25.6975 20.08 25.8325 ;
      RECT  20.12 27.4825 20.185 27.3475 ;
      RECT  20.635 27.4825 20.705 27.3475 ;
      RECT  20.015 27.6475 20.185 27.5825 ;
      RECT  19.875 28.0225 20.76 27.9575 ;
      RECT  19.93 27.0175 20.0 26.8175 ;
      RECT  20.635 27.0175 20.7 26.8825 ;
      RECT  20.1875 27.8725 20.2525 27.7375 ;
      RECT  20.37 27.8725 20.435 27.7375 ;
      RECT  20.635 27.4825 20.7 27.3475 ;
      RECT  20.6025 28.1625 20.7375 28.0975 ;
      RECT  20.3625 27.2825 20.4975 27.2175 ;
      RECT  20.585 28.02 20.6375 27.9575 ;
      RECT  20.1375 27.1325 20.2725 27.0675 ;
      RECT  20.015 27.8725 20.085 27.5825 ;
      RECT  20.12 27.6475 20.185 26.9075 ;
      RECT  20.635 27.0175 20.705 26.8175 ;
      RECT  20.555 27.8725 20.62 27.7375 ;
      RECT  19.88 28.02 19.9325 27.9575 ;
      RECT  19.875 26.8175 20.76 26.7525 ;
      RECT  19.9325 27.38 19.9975 27.245 ;
      RECT  20.25 28.1625 20.385 28.0975 ;
      RECT  20.555 27.8725 20.625 27.5825 ;
      RECT  20.2325 28.0225 20.3675 27.9575 ;
      RECT  19.935 27.0175 20.0 26.8825 ;
      RECT  20.45 27.6475 20.625 27.5825 ;
      RECT  20.45 27.0175 20.515 26.8825 ;
      RECT  19.875 28.1625 20.76 28.0975 ;
      RECT  20.6375 27.38 20.7025 27.245 ;
      RECT  19.93 27.4825 20.0 27.3475 ;
      RECT  20.2 27.8725 20.265 27.7375 ;
      RECT  20.45 27.4825 20.515 27.3475 ;
      RECT  20.3825 27.8725 20.4475 27.7375 ;
      RECT  19.935 27.4825 20.0 27.3475 ;
      RECT  20.12 27.0175 20.185 26.8825 ;
      RECT  20.45 27.6475 20.515 27.0175 ;
      RECT  19.8975 28.1625 20.0325 28.0975 ;
      RECT  20.015 27.8725 20.08 27.7375 ;
      RECT  20.12 28.7775 20.185 28.9125 ;
      RECT  20.635 28.7775 20.705 28.9125 ;
      RECT  20.015 28.6125 20.185 28.6775 ;
      RECT  19.875 28.2375 20.76 28.3025 ;
      RECT  19.93 29.2425 20.0 29.4425 ;
      RECT  20.635 29.2425 20.7 29.3775 ;
      RECT  20.1875 28.3875 20.2525 28.5225 ;
      RECT  20.37 28.3875 20.435 28.5225 ;
      RECT  20.635 28.7775 20.7 28.9125 ;
      RECT  20.6025 28.0975 20.7375 28.1625 ;
      RECT  20.3625 28.9775 20.4975 29.0425 ;
      RECT  20.585 28.24 20.6375 28.3025 ;
      RECT  20.1375 29.1275 20.2725 29.1925 ;
      RECT  20.015 28.3875 20.085 28.6775 ;
      RECT  20.12 28.6125 20.185 29.3525 ;
      RECT  20.635 29.2425 20.705 29.4425 ;
      RECT  20.555 28.3875 20.62 28.5225 ;
      RECT  19.88 28.24 19.9325 28.3025 ;
      RECT  19.875 29.4425 20.76 29.5075 ;
      RECT  19.9325 28.88 19.9975 29.015 ;
      RECT  20.25 28.0975 20.385 28.1625 ;
      RECT  20.555 28.3875 20.625 28.6775 ;
      RECT  20.2325 28.2375 20.3675 28.3025 ;
      RECT  19.935 29.2425 20.0 29.3775 ;
      RECT  20.45 28.6125 20.625 28.6775 ;
      RECT  20.45 29.2425 20.515 29.3775 ;
      RECT  19.875 28.0975 20.76 28.1625 ;
      RECT  20.6375 28.88 20.7025 29.015 ;
      RECT  19.93 28.7775 20.0 28.9125 ;
      RECT  20.2 28.3875 20.265 28.5225 ;
      RECT  20.45 28.7775 20.515 28.9125 ;
      RECT  20.3825 28.3875 20.4475 28.5225 ;
      RECT  19.935 28.7775 20.0 28.9125 ;
      RECT  20.12 29.2425 20.185 29.3775 ;
      RECT  20.45 28.6125 20.515 29.2425 ;
      RECT  19.8975 28.0975 20.0325 28.1625 ;
      RECT  20.015 28.3875 20.08 28.5225 ;
      RECT  20.12 30.1725 20.185 30.0375 ;
      RECT  20.635 30.1725 20.705 30.0375 ;
      RECT  20.015 30.3375 20.185 30.2725 ;
      RECT  19.875 30.7125 20.76 30.6475 ;
      RECT  19.93 29.7075 20.0 29.5075 ;
      RECT  20.635 29.7075 20.7 29.5725 ;
      RECT  20.1875 30.5625 20.2525 30.4275 ;
      RECT  20.37 30.5625 20.435 30.4275 ;
      RECT  20.635 30.1725 20.7 30.0375 ;
      RECT  20.6025 30.8525 20.7375 30.7875 ;
      RECT  20.3625 29.9725 20.4975 29.9075 ;
      RECT  20.585 30.71 20.6375 30.6475 ;
      RECT  20.1375 29.8225 20.2725 29.7575 ;
      RECT  20.015 30.5625 20.085 30.2725 ;
      RECT  20.12 30.3375 20.185 29.5975 ;
      RECT  20.635 29.7075 20.705 29.5075 ;
      RECT  20.555 30.5625 20.62 30.4275 ;
      RECT  19.88 30.71 19.9325 30.6475 ;
      RECT  19.875 29.5075 20.76 29.4425 ;
      RECT  19.9325 30.07 19.9975 29.935 ;
      RECT  20.25 30.8525 20.385 30.7875 ;
      RECT  20.555 30.5625 20.625 30.2725 ;
      RECT  20.2325 30.7125 20.3675 30.6475 ;
      RECT  19.935 29.7075 20.0 29.5725 ;
      RECT  20.45 30.3375 20.625 30.2725 ;
      RECT  20.45 29.7075 20.515 29.5725 ;
      RECT  19.875 30.8525 20.76 30.7875 ;
      RECT  20.6375 30.07 20.7025 29.935 ;
      RECT  19.93 30.1725 20.0 30.0375 ;
      RECT  20.2 30.5625 20.265 30.4275 ;
      RECT  20.45 30.1725 20.515 30.0375 ;
      RECT  20.3825 30.5625 20.4475 30.4275 ;
      RECT  19.935 30.1725 20.0 30.0375 ;
      RECT  20.12 29.7075 20.185 29.5725 ;
      RECT  20.45 30.3375 20.515 29.7075 ;
      RECT  19.8975 30.8525 20.0325 30.7875 ;
      RECT  20.015 30.5625 20.08 30.4275 ;
      RECT  20.12 31.4675 20.185 31.6025 ;
      RECT  20.635 31.4675 20.705 31.6025 ;
      RECT  20.015 31.3025 20.185 31.3675 ;
      RECT  19.875 30.9275 20.76 30.9925 ;
      RECT  19.93 31.9325 20.0 32.1325 ;
      RECT  20.635 31.9325 20.7 32.0675 ;
      RECT  20.1875 31.0775 20.2525 31.2125 ;
      RECT  20.37 31.0775 20.435 31.2125 ;
      RECT  20.635 31.4675 20.7 31.6025 ;
      RECT  20.6025 30.7875 20.7375 30.8525 ;
      RECT  20.3625 31.6675 20.4975 31.7325 ;
      RECT  20.585 30.93 20.6375 30.9925 ;
      RECT  20.1375 31.8175 20.2725 31.8825 ;
      RECT  20.015 31.0775 20.085 31.3675 ;
      RECT  20.12 31.3025 20.185 32.0425 ;
      RECT  20.635 31.9325 20.705 32.1325 ;
      RECT  20.555 31.0775 20.62 31.2125 ;
      RECT  19.88 30.93 19.9325 30.9925 ;
      RECT  19.875 32.1325 20.76 32.1975 ;
      RECT  19.9325 31.57 19.9975 31.705 ;
      RECT  20.25 30.7875 20.385 30.8525 ;
      RECT  20.555 31.0775 20.625 31.3675 ;
      RECT  20.2325 30.9275 20.3675 30.9925 ;
      RECT  19.935 31.9325 20.0 32.0675 ;
      RECT  20.45 31.3025 20.625 31.3675 ;
      RECT  20.45 31.9325 20.515 32.0675 ;
      RECT  19.875 30.7875 20.76 30.8525 ;
      RECT  20.6375 31.57 20.7025 31.705 ;
      RECT  19.93 31.4675 20.0 31.6025 ;
      RECT  20.2 31.0775 20.265 31.2125 ;
      RECT  20.45 31.4675 20.515 31.6025 ;
      RECT  20.3825 31.0775 20.4475 31.2125 ;
      RECT  19.935 31.4675 20.0 31.6025 ;
      RECT  20.12 31.9325 20.185 32.0675 ;
      RECT  20.45 31.3025 20.515 31.9325 ;
      RECT  19.8975 30.7875 20.0325 30.8525 ;
      RECT  20.015 31.0775 20.08 31.2125 ;
      RECT  20.12 32.8625 20.185 32.7275 ;
      RECT  20.635 32.8625 20.705 32.7275 ;
      RECT  20.015 33.0275 20.185 32.9625 ;
      RECT  19.875 33.4025 20.76 33.3375 ;
      RECT  19.93 32.3975 20.0 32.1975 ;
      RECT  20.635 32.3975 20.7 32.2625 ;
      RECT  20.1875 33.2525 20.2525 33.1175 ;
      RECT  20.37 33.2525 20.435 33.1175 ;
      RECT  20.635 32.8625 20.7 32.7275 ;
      RECT  20.6025 33.5425 20.7375 33.4775 ;
      RECT  20.3625 32.6625 20.4975 32.5975 ;
      RECT  20.585 33.4 20.6375 33.3375 ;
      RECT  20.1375 32.5125 20.2725 32.4475 ;
      RECT  20.015 33.2525 20.085 32.9625 ;
      RECT  20.12 33.0275 20.185 32.2875 ;
      RECT  20.635 32.3975 20.705 32.1975 ;
      RECT  20.555 33.2525 20.62 33.1175 ;
      RECT  19.88 33.4 19.9325 33.3375 ;
      RECT  19.875 32.1975 20.76 32.1325 ;
      RECT  19.9325 32.76 19.9975 32.625 ;
      RECT  20.25 33.5425 20.385 33.4775 ;
      RECT  20.555 33.2525 20.625 32.9625 ;
      RECT  20.2325 33.4025 20.3675 33.3375 ;
      RECT  19.935 32.3975 20.0 32.2625 ;
      RECT  20.45 33.0275 20.625 32.9625 ;
      RECT  20.45 32.3975 20.515 32.2625 ;
      RECT  19.875 33.5425 20.76 33.4775 ;
      RECT  20.6375 32.76 20.7025 32.625 ;
      RECT  19.93 32.8625 20.0 32.7275 ;
      RECT  20.2 33.2525 20.265 33.1175 ;
      RECT  20.45 32.8625 20.515 32.7275 ;
      RECT  20.3825 33.2525 20.4475 33.1175 ;
      RECT  19.935 32.8625 20.0 32.7275 ;
      RECT  20.12 32.3975 20.185 32.2625 ;
      RECT  20.45 33.0275 20.515 32.3975 ;
      RECT  19.8975 33.5425 20.0325 33.4775 ;
      RECT  20.015 33.2525 20.08 33.1175 ;
      RECT  20.12 34.1575 20.185 34.2925 ;
      RECT  20.635 34.1575 20.705 34.2925 ;
      RECT  20.015 33.9925 20.185 34.0575 ;
      RECT  19.875 33.6175 20.76 33.6825 ;
      RECT  19.93 34.6225 20.0 34.8225 ;
      RECT  20.635 34.6225 20.7 34.7575 ;
      RECT  20.1875 33.7675 20.2525 33.9025 ;
      RECT  20.37 33.7675 20.435 33.9025 ;
      RECT  20.635 34.1575 20.7 34.2925 ;
      RECT  20.6025 33.4775 20.7375 33.5425 ;
      RECT  20.3625 34.3575 20.4975 34.4225 ;
      RECT  20.585 33.62 20.6375 33.6825 ;
      RECT  20.1375 34.5075 20.2725 34.5725 ;
      RECT  20.015 33.7675 20.085 34.0575 ;
      RECT  20.12 33.9925 20.185 34.7325 ;
      RECT  20.635 34.6225 20.705 34.8225 ;
      RECT  20.555 33.7675 20.62 33.9025 ;
      RECT  19.88 33.62 19.9325 33.6825 ;
      RECT  19.875 34.8225 20.76 34.8875 ;
      RECT  19.9325 34.26 19.9975 34.395 ;
      RECT  20.25 33.4775 20.385 33.5425 ;
      RECT  20.555 33.7675 20.625 34.0575 ;
      RECT  20.2325 33.6175 20.3675 33.6825 ;
      RECT  19.935 34.6225 20.0 34.7575 ;
      RECT  20.45 33.9925 20.625 34.0575 ;
      RECT  20.45 34.6225 20.515 34.7575 ;
      RECT  19.875 33.4775 20.76 33.5425 ;
      RECT  20.6375 34.26 20.7025 34.395 ;
      RECT  19.93 34.1575 20.0 34.2925 ;
      RECT  20.2 33.7675 20.265 33.9025 ;
      RECT  20.45 34.1575 20.515 34.2925 ;
      RECT  20.3825 33.7675 20.4475 33.9025 ;
      RECT  19.935 34.1575 20.0 34.2925 ;
      RECT  20.12 34.6225 20.185 34.7575 ;
      RECT  20.45 33.9925 20.515 34.6225 ;
      RECT  19.8975 33.4775 20.0325 33.5425 ;
      RECT  20.015 33.7675 20.08 33.9025 ;
      RECT  20.12 35.5525 20.185 35.4175 ;
      RECT  20.635 35.5525 20.705 35.4175 ;
      RECT  20.015 35.7175 20.185 35.6525 ;
      RECT  19.875 36.0925 20.76 36.0275 ;
      RECT  19.93 35.0875 20.0 34.8875 ;
      RECT  20.635 35.0875 20.7 34.9525 ;
      RECT  20.1875 35.9425 20.2525 35.8075 ;
      RECT  20.37 35.9425 20.435 35.8075 ;
      RECT  20.635 35.5525 20.7 35.4175 ;
      RECT  20.6025 36.2325 20.7375 36.1675 ;
      RECT  20.3625 35.3525 20.4975 35.2875 ;
      RECT  20.585 36.09 20.6375 36.0275 ;
      RECT  20.1375 35.2025 20.2725 35.1375 ;
      RECT  20.015 35.9425 20.085 35.6525 ;
      RECT  20.12 35.7175 20.185 34.9775 ;
      RECT  20.635 35.0875 20.705 34.8875 ;
      RECT  20.555 35.9425 20.62 35.8075 ;
      RECT  19.88 36.09 19.9325 36.0275 ;
      RECT  19.875 34.8875 20.76 34.8225 ;
      RECT  19.9325 35.45 19.9975 35.315 ;
      RECT  20.25 36.2325 20.385 36.1675 ;
      RECT  20.555 35.9425 20.625 35.6525 ;
      RECT  20.2325 36.0925 20.3675 36.0275 ;
      RECT  19.935 35.0875 20.0 34.9525 ;
      RECT  20.45 35.7175 20.625 35.6525 ;
      RECT  20.45 35.0875 20.515 34.9525 ;
      RECT  19.875 36.2325 20.76 36.1675 ;
      RECT  20.6375 35.45 20.7025 35.315 ;
      RECT  19.93 35.5525 20.0 35.4175 ;
      RECT  20.2 35.9425 20.265 35.8075 ;
      RECT  20.45 35.5525 20.515 35.4175 ;
      RECT  20.3825 35.9425 20.4475 35.8075 ;
      RECT  19.935 35.5525 20.0 35.4175 ;
      RECT  20.12 35.0875 20.185 34.9525 ;
      RECT  20.45 35.7175 20.515 35.0875 ;
      RECT  19.8975 36.2325 20.0325 36.1675 ;
      RECT  20.015 35.9425 20.08 35.8075 ;
      RECT  20.12 36.8475 20.185 36.9825 ;
      RECT  20.635 36.8475 20.705 36.9825 ;
      RECT  20.015 36.6825 20.185 36.7475 ;
      RECT  19.875 36.3075 20.76 36.3725 ;
      RECT  19.93 37.3125 20.0 37.5125 ;
      RECT  20.635 37.3125 20.7 37.4475 ;
      RECT  20.1875 36.4575 20.2525 36.5925 ;
      RECT  20.37 36.4575 20.435 36.5925 ;
      RECT  20.635 36.8475 20.7 36.9825 ;
      RECT  20.6025 36.1675 20.7375 36.2325 ;
      RECT  20.3625 37.0475 20.4975 37.1125 ;
      RECT  20.585 36.31 20.6375 36.3725 ;
      RECT  20.1375 37.1975 20.2725 37.2625 ;
      RECT  20.015 36.4575 20.085 36.7475 ;
      RECT  20.12 36.6825 20.185 37.4225 ;
      RECT  20.635 37.3125 20.705 37.5125 ;
      RECT  20.555 36.4575 20.62 36.5925 ;
      RECT  19.88 36.31 19.9325 36.3725 ;
      RECT  19.875 37.5125 20.76 37.5775 ;
      RECT  19.9325 36.95 19.9975 37.085 ;
      RECT  20.25 36.1675 20.385 36.2325 ;
      RECT  20.555 36.4575 20.625 36.7475 ;
      RECT  20.2325 36.3075 20.3675 36.3725 ;
      RECT  19.935 37.3125 20.0 37.4475 ;
      RECT  20.45 36.6825 20.625 36.7475 ;
      RECT  20.45 37.3125 20.515 37.4475 ;
      RECT  19.875 36.1675 20.76 36.2325 ;
      RECT  20.6375 36.95 20.7025 37.085 ;
      RECT  19.93 36.8475 20.0 36.9825 ;
      RECT  20.2 36.4575 20.265 36.5925 ;
      RECT  20.45 36.8475 20.515 36.9825 ;
      RECT  20.3825 36.4575 20.4475 36.5925 ;
      RECT  19.935 36.8475 20.0 36.9825 ;
      RECT  20.12 37.3125 20.185 37.4475 ;
      RECT  20.45 36.6825 20.515 37.3125 ;
      RECT  19.8975 36.1675 20.0325 36.2325 ;
      RECT  20.015 36.4575 20.08 36.5925 ;
      RECT  20.12 38.2425 20.185 38.1075 ;
      RECT  20.635 38.2425 20.705 38.1075 ;
      RECT  20.015 38.4075 20.185 38.3425 ;
      RECT  19.875 38.7825 20.76 38.7175 ;
      RECT  19.93 37.7775 20.0 37.5775 ;
      RECT  20.635 37.7775 20.7 37.6425 ;
      RECT  20.1875 38.6325 20.2525 38.4975 ;
      RECT  20.37 38.6325 20.435 38.4975 ;
      RECT  20.635 38.2425 20.7 38.1075 ;
      RECT  20.6025 38.9225 20.7375 38.8575 ;
      RECT  20.3625 38.0425 20.4975 37.9775 ;
      RECT  20.585 38.78 20.6375 38.7175 ;
      RECT  20.1375 37.8925 20.2725 37.8275 ;
      RECT  20.015 38.6325 20.085 38.3425 ;
      RECT  20.12 38.4075 20.185 37.6675 ;
      RECT  20.635 37.7775 20.705 37.5775 ;
      RECT  20.555 38.6325 20.62 38.4975 ;
      RECT  19.88 38.78 19.9325 38.7175 ;
      RECT  19.875 37.5775 20.76 37.5125 ;
      RECT  19.9325 38.14 19.9975 38.005 ;
      RECT  20.25 38.9225 20.385 38.8575 ;
      RECT  20.555 38.6325 20.625 38.3425 ;
      RECT  20.2325 38.7825 20.3675 38.7175 ;
      RECT  19.935 37.7775 20.0 37.6425 ;
      RECT  20.45 38.4075 20.625 38.3425 ;
      RECT  20.45 37.7775 20.515 37.6425 ;
      RECT  19.875 38.9225 20.76 38.8575 ;
      RECT  20.6375 38.14 20.7025 38.005 ;
      RECT  19.93 38.2425 20.0 38.1075 ;
      RECT  20.2 38.6325 20.265 38.4975 ;
      RECT  20.45 38.2425 20.515 38.1075 ;
      RECT  20.3825 38.6325 20.4475 38.4975 ;
      RECT  19.935 38.2425 20.0 38.1075 ;
      RECT  20.12 37.7775 20.185 37.6425 ;
      RECT  20.45 38.4075 20.515 37.7775 ;
      RECT  19.8975 38.9225 20.0325 38.8575 ;
      RECT  20.015 38.6325 20.08 38.4975 ;
      RECT  20.12 39.5375 20.185 39.6725 ;
      RECT  20.635 39.5375 20.705 39.6725 ;
      RECT  20.015 39.3725 20.185 39.4375 ;
      RECT  19.875 38.9975 20.76 39.0625 ;
      RECT  19.93 40.0025 20.0 40.2025 ;
      RECT  20.635 40.0025 20.7 40.1375 ;
      RECT  20.1875 39.1475 20.2525 39.2825 ;
      RECT  20.37 39.1475 20.435 39.2825 ;
      RECT  20.635 39.5375 20.7 39.6725 ;
      RECT  20.6025 38.8575 20.7375 38.9225 ;
      RECT  20.3625 39.7375 20.4975 39.8025 ;
      RECT  20.585 39.0 20.6375 39.0625 ;
      RECT  20.1375 39.8875 20.2725 39.9525 ;
      RECT  20.015 39.1475 20.085 39.4375 ;
      RECT  20.12 39.3725 20.185 40.1125 ;
      RECT  20.635 40.0025 20.705 40.2025 ;
      RECT  20.555 39.1475 20.62 39.2825 ;
      RECT  19.88 39.0 19.9325 39.0625 ;
      RECT  19.875 40.2025 20.76 40.2675 ;
      RECT  19.9325 39.64 19.9975 39.775 ;
      RECT  20.25 38.8575 20.385 38.9225 ;
      RECT  20.555 39.1475 20.625 39.4375 ;
      RECT  20.2325 38.9975 20.3675 39.0625 ;
      RECT  19.935 40.0025 20.0 40.1375 ;
      RECT  20.45 39.3725 20.625 39.4375 ;
      RECT  20.45 40.0025 20.515 40.1375 ;
      RECT  19.875 38.8575 20.76 38.9225 ;
      RECT  20.6375 39.64 20.7025 39.775 ;
      RECT  19.93 39.5375 20.0 39.6725 ;
      RECT  20.2 39.1475 20.265 39.2825 ;
      RECT  20.45 39.5375 20.515 39.6725 ;
      RECT  20.3825 39.1475 20.4475 39.2825 ;
      RECT  19.935 39.5375 20.0 39.6725 ;
      RECT  20.12 40.0025 20.185 40.1375 ;
      RECT  20.45 39.3725 20.515 40.0025 ;
      RECT  19.8975 38.8575 20.0325 38.9225 ;
      RECT  20.015 39.1475 20.08 39.2825 ;
      RECT  20.12 40.9325 20.185 40.7975 ;
      RECT  20.635 40.9325 20.705 40.7975 ;
      RECT  20.015 41.0975 20.185 41.0325 ;
      RECT  19.875 41.4725 20.76 41.4075 ;
      RECT  19.93 40.4675 20.0 40.2675 ;
      RECT  20.635 40.4675 20.7 40.3325 ;
      RECT  20.1875 41.3225 20.2525 41.1875 ;
      RECT  20.37 41.3225 20.435 41.1875 ;
      RECT  20.635 40.9325 20.7 40.7975 ;
      RECT  20.6025 41.6125 20.7375 41.5475 ;
      RECT  20.3625 40.7325 20.4975 40.6675 ;
      RECT  20.585 41.47 20.6375 41.4075 ;
      RECT  20.1375 40.5825 20.2725 40.5175 ;
      RECT  20.015 41.3225 20.085 41.0325 ;
      RECT  20.12 41.0975 20.185 40.3575 ;
      RECT  20.635 40.4675 20.705 40.2675 ;
      RECT  20.555 41.3225 20.62 41.1875 ;
      RECT  19.88 41.47 19.9325 41.4075 ;
      RECT  19.875 40.2675 20.76 40.2025 ;
      RECT  19.9325 40.83 19.9975 40.695 ;
      RECT  20.25 41.6125 20.385 41.5475 ;
      RECT  20.555 41.3225 20.625 41.0325 ;
      RECT  20.2325 41.4725 20.3675 41.4075 ;
      RECT  19.935 40.4675 20.0 40.3325 ;
      RECT  20.45 41.0975 20.625 41.0325 ;
      RECT  20.45 40.4675 20.515 40.3325 ;
      RECT  19.875 41.6125 20.76 41.5475 ;
      RECT  20.6375 40.83 20.7025 40.695 ;
      RECT  19.93 40.9325 20.0 40.7975 ;
      RECT  20.2 41.3225 20.265 41.1875 ;
      RECT  20.45 40.9325 20.515 40.7975 ;
      RECT  20.3825 41.3225 20.4475 41.1875 ;
      RECT  19.935 40.9325 20.0 40.7975 ;
      RECT  20.12 40.4675 20.185 40.3325 ;
      RECT  20.45 41.0975 20.515 40.4675 ;
      RECT  19.8975 41.6125 20.0325 41.5475 ;
      RECT  20.015 41.3225 20.08 41.1875 ;
      RECT  20.12 42.2275 20.185 42.3625 ;
      RECT  20.635 42.2275 20.705 42.3625 ;
      RECT  20.015 42.0625 20.185 42.1275 ;
      RECT  19.875 41.6875 20.76 41.7525 ;
      RECT  19.93 42.6925 20.0 42.8925 ;
      RECT  20.635 42.6925 20.7 42.8275 ;
      RECT  20.1875 41.8375 20.2525 41.9725 ;
      RECT  20.37 41.8375 20.435 41.9725 ;
      RECT  20.635 42.2275 20.7 42.3625 ;
      RECT  20.6025 41.5475 20.7375 41.6125 ;
      RECT  20.3625 42.4275 20.4975 42.4925 ;
      RECT  20.585 41.69 20.6375 41.7525 ;
      RECT  20.1375 42.5775 20.2725 42.6425 ;
      RECT  20.015 41.8375 20.085 42.1275 ;
      RECT  20.12 42.0625 20.185 42.8025 ;
      RECT  20.635 42.6925 20.705 42.8925 ;
      RECT  20.555 41.8375 20.62 41.9725 ;
      RECT  19.88 41.69 19.9325 41.7525 ;
      RECT  19.875 42.8925 20.76 42.9575 ;
      RECT  19.9325 42.33 19.9975 42.465 ;
      RECT  20.25 41.5475 20.385 41.6125 ;
      RECT  20.555 41.8375 20.625 42.1275 ;
      RECT  20.2325 41.6875 20.3675 41.7525 ;
      RECT  19.935 42.6925 20.0 42.8275 ;
      RECT  20.45 42.0625 20.625 42.1275 ;
      RECT  20.45 42.6925 20.515 42.8275 ;
      RECT  19.875 41.5475 20.76 41.6125 ;
      RECT  20.6375 42.33 20.7025 42.465 ;
      RECT  19.93 42.2275 20.0 42.3625 ;
      RECT  20.2 41.8375 20.265 41.9725 ;
      RECT  20.45 42.2275 20.515 42.3625 ;
      RECT  20.3825 41.8375 20.4475 41.9725 ;
      RECT  19.935 42.2275 20.0 42.3625 ;
      RECT  20.12 42.6925 20.185 42.8275 ;
      RECT  20.45 42.0625 20.515 42.6925 ;
      RECT  19.8975 41.5475 20.0325 41.6125 ;
      RECT  20.015 41.8375 20.08 41.9725 ;
      RECT  20.12 43.6225 20.185 43.4875 ;
      RECT  20.635 43.6225 20.705 43.4875 ;
      RECT  20.015 43.7875 20.185 43.7225 ;
      RECT  19.875 44.1625 20.76 44.0975 ;
      RECT  19.93 43.1575 20.0 42.9575 ;
      RECT  20.635 43.1575 20.7 43.0225 ;
      RECT  20.1875 44.0125 20.2525 43.8775 ;
      RECT  20.37 44.0125 20.435 43.8775 ;
      RECT  20.635 43.6225 20.7 43.4875 ;
      RECT  20.6025 44.3025 20.7375 44.2375 ;
      RECT  20.3625 43.4225 20.4975 43.3575 ;
      RECT  20.585 44.16 20.6375 44.0975 ;
      RECT  20.1375 43.2725 20.2725 43.2075 ;
      RECT  20.015 44.0125 20.085 43.7225 ;
      RECT  20.12 43.7875 20.185 43.0475 ;
      RECT  20.635 43.1575 20.705 42.9575 ;
      RECT  20.555 44.0125 20.62 43.8775 ;
      RECT  19.88 44.16 19.9325 44.0975 ;
      RECT  19.875 42.9575 20.76 42.8925 ;
      RECT  19.9325 43.52 19.9975 43.385 ;
      RECT  20.25 44.3025 20.385 44.2375 ;
      RECT  20.555 44.0125 20.625 43.7225 ;
      RECT  20.2325 44.1625 20.3675 44.0975 ;
      RECT  19.935 43.1575 20.0 43.0225 ;
      RECT  20.45 43.7875 20.625 43.7225 ;
      RECT  20.45 43.1575 20.515 43.0225 ;
      RECT  19.875 44.3025 20.76 44.2375 ;
      RECT  20.6375 43.52 20.7025 43.385 ;
      RECT  19.93 43.6225 20.0 43.4875 ;
      RECT  20.2 44.0125 20.265 43.8775 ;
      RECT  20.45 43.6225 20.515 43.4875 ;
      RECT  20.3825 44.0125 20.4475 43.8775 ;
      RECT  19.935 43.6225 20.0 43.4875 ;
      RECT  20.12 43.1575 20.185 43.0225 ;
      RECT  20.45 43.7875 20.515 43.1575 ;
      RECT  19.8975 44.3025 20.0325 44.2375 ;
      RECT  20.015 44.0125 20.08 43.8775 ;
      RECT  20.12 44.9175 20.185 45.0525 ;
      RECT  20.635 44.9175 20.705 45.0525 ;
      RECT  20.015 44.7525 20.185 44.8175 ;
      RECT  19.875 44.3775 20.76 44.4425 ;
      RECT  19.93 45.3825 20.0 45.5825 ;
      RECT  20.635 45.3825 20.7 45.5175 ;
      RECT  20.1875 44.5275 20.2525 44.6625 ;
      RECT  20.37 44.5275 20.435 44.6625 ;
      RECT  20.635 44.9175 20.7 45.0525 ;
      RECT  20.6025 44.2375 20.7375 44.3025 ;
      RECT  20.3625 45.1175 20.4975 45.1825 ;
      RECT  20.585 44.38 20.6375 44.4425 ;
      RECT  20.1375 45.2675 20.2725 45.3325 ;
      RECT  20.015 44.5275 20.085 44.8175 ;
      RECT  20.12 44.7525 20.185 45.4925 ;
      RECT  20.635 45.3825 20.705 45.5825 ;
      RECT  20.555 44.5275 20.62 44.6625 ;
      RECT  19.88 44.38 19.9325 44.4425 ;
      RECT  19.875 45.5825 20.76 45.6475 ;
      RECT  19.9325 45.02 19.9975 45.155 ;
      RECT  20.25 44.2375 20.385 44.3025 ;
      RECT  20.555 44.5275 20.625 44.8175 ;
      RECT  20.2325 44.3775 20.3675 44.4425 ;
      RECT  19.935 45.3825 20.0 45.5175 ;
      RECT  20.45 44.7525 20.625 44.8175 ;
      RECT  20.45 45.3825 20.515 45.5175 ;
      RECT  19.875 44.2375 20.76 44.3025 ;
      RECT  20.6375 45.02 20.7025 45.155 ;
      RECT  19.93 44.9175 20.0 45.0525 ;
      RECT  20.2 44.5275 20.265 44.6625 ;
      RECT  20.45 44.9175 20.515 45.0525 ;
      RECT  20.3825 44.5275 20.4475 44.6625 ;
      RECT  19.935 44.9175 20.0 45.0525 ;
      RECT  20.12 45.3825 20.185 45.5175 ;
      RECT  20.45 44.7525 20.515 45.3825 ;
      RECT  19.8975 44.2375 20.0325 44.3025 ;
      RECT  20.015 44.5275 20.08 44.6625 ;
      RECT  19.965 20.1675 20.67 20.2325 ;
      RECT  19.965 22.5775 20.67 22.6425 ;
      RECT  19.965 22.8575 20.67 22.9225 ;
      RECT  19.965 25.2675 20.67 25.3325 ;
      RECT  19.965 25.5475 20.67 25.6125 ;
      RECT  19.965 27.9575 20.67 28.0225 ;
      RECT  19.965 28.2375 20.67 28.3025 ;
      RECT  19.965 30.6475 20.67 30.7125 ;
      RECT  19.965 30.9275 20.67 30.9925 ;
      RECT  19.965 33.3375 20.67 33.4025 ;
      RECT  19.965 33.6175 20.67 33.6825 ;
      RECT  19.965 36.0275 20.67 36.0925 ;
      RECT  19.965 36.3075 20.67 36.3725 ;
      RECT  19.965 38.7175 20.67 38.7825 ;
      RECT  19.965 38.9975 20.67 39.0625 ;
      RECT  19.965 41.4075 20.67 41.4725 ;
      RECT  19.965 41.6875 20.67 41.7525 ;
      RECT  19.965 44.0975 20.67 44.1625 ;
      RECT  19.965 44.3775 20.67 44.4425 ;
      RECT  22.94 20.7075 23.005 20.8425 ;
      RECT  23.455 20.7075 23.525 20.8425 ;
      RECT  22.835 20.5425 23.005 20.6075 ;
      RECT  22.695 20.1675 23.58 20.2325 ;
      RECT  22.75 21.1725 22.82 21.3725 ;
      RECT  23.455 21.1725 23.52 21.3075 ;
      RECT  23.0075 20.3175 23.0725 20.4525 ;
      RECT  23.19 20.3175 23.255 20.4525 ;
      RECT  23.455 20.7075 23.52 20.8425 ;
      RECT  23.4225 20.0275 23.5575 20.0925 ;
      RECT  23.1825 20.9075 23.3175 20.9725 ;
      RECT  23.405 20.17 23.4575 20.2325 ;
      RECT  22.9575 21.0575 23.0925 21.1225 ;
      RECT  22.835 20.3175 22.905 20.6075 ;
      RECT  22.94 20.5425 23.005 21.2825 ;
      RECT  23.455 21.1725 23.525 21.3725 ;
      RECT  23.375 20.3175 23.44 20.4525 ;
      RECT  22.7 20.17 22.7525 20.2325 ;
      RECT  22.695 21.3725 23.58 21.4375 ;
      RECT  22.7525 20.81 22.8175 20.945 ;
      RECT  23.07 20.0275 23.205 20.0925 ;
      RECT  23.375 20.3175 23.445 20.6075 ;
      RECT  23.0525 20.1675 23.1875 20.2325 ;
      RECT  22.755 21.1725 22.82 21.3075 ;
      RECT  23.27 20.5425 23.445 20.6075 ;
      RECT  23.27 21.1725 23.335 21.3075 ;
      RECT  22.695 20.0275 23.58 20.0925 ;
      RECT  23.4575 20.81 23.5225 20.945 ;
      RECT  22.75 20.7075 22.82 20.8425 ;
      RECT  23.02 20.3175 23.085 20.4525 ;
      RECT  23.27 20.7075 23.335 20.8425 ;
      RECT  23.2025 20.3175 23.2675 20.4525 ;
      RECT  22.755 20.7075 22.82 20.8425 ;
      RECT  22.94 21.1725 23.005 21.3075 ;
      RECT  23.27 20.5425 23.335 21.1725 ;
      RECT  22.7175 20.0275 22.8525 20.0925 ;
      RECT  22.835 20.3175 22.9 20.4525 ;
      RECT  22.94 22.1025 23.005 21.9675 ;
      RECT  23.455 22.1025 23.525 21.9675 ;
      RECT  22.835 22.2675 23.005 22.2025 ;
      RECT  22.695 22.6425 23.58 22.5775 ;
      RECT  22.75 21.6375 22.82 21.4375 ;
      RECT  23.455 21.6375 23.52 21.5025 ;
      RECT  23.0075 22.4925 23.0725 22.3575 ;
      RECT  23.19 22.4925 23.255 22.3575 ;
      RECT  23.455 22.1025 23.52 21.9675 ;
      RECT  23.4225 22.7825 23.5575 22.7175 ;
      RECT  23.1825 21.9025 23.3175 21.8375 ;
      RECT  23.405 22.64 23.4575 22.5775 ;
      RECT  22.9575 21.7525 23.0925 21.6875 ;
      RECT  22.835 22.4925 22.905 22.2025 ;
      RECT  22.94 22.2675 23.005 21.5275 ;
      RECT  23.455 21.6375 23.525 21.4375 ;
      RECT  23.375 22.4925 23.44 22.3575 ;
      RECT  22.7 22.64 22.7525 22.5775 ;
      RECT  22.695 21.4375 23.58 21.3725 ;
      RECT  22.7525 22.0 22.8175 21.865 ;
      RECT  23.07 22.7825 23.205 22.7175 ;
      RECT  23.375 22.4925 23.445 22.2025 ;
      RECT  23.0525 22.6425 23.1875 22.5775 ;
      RECT  22.755 21.6375 22.82 21.5025 ;
      RECT  23.27 22.2675 23.445 22.2025 ;
      RECT  23.27 21.6375 23.335 21.5025 ;
      RECT  22.695 22.7825 23.58 22.7175 ;
      RECT  23.4575 22.0 23.5225 21.865 ;
      RECT  22.75 22.1025 22.82 21.9675 ;
      RECT  23.02 22.4925 23.085 22.3575 ;
      RECT  23.27 22.1025 23.335 21.9675 ;
      RECT  23.2025 22.4925 23.2675 22.3575 ;
      RECT  22.755 22.1025 22.82 21.9675 ;
      RECT  22.94 21.6375 23.005 21.5025 ;
      RECT  23.27 22.2675 23.335 21.6375 ;
      RECT  22.7175 22.7825 22.8525 22.7175 ;
      RECT  22.835 22.4925 22.9 22.3575 ;
      RECT  22.94 23.3975 23.005 23.5325 ;
      RECT  23.455 23.3975 23.525 23.5325 ;
      RECT  22.835 23.2325 23.005 23.2975 ;
      RECT  22.695 22.8575 23.58 22.9225 ;
      RECT  22.75 23.8625 22.82 24.0625 ;
      RECT  23.455 23.8625 23.52 23.9975 ;
      RECT  23.0075 23.0075 23.0725 23.1425 ;
      RECT  23.19 23.0075 23.255 23.1425 ;
      RECT  23.455 23.3975 23.52 23.5325 ;
      RECT  23.4225 22.7175 23.5575 22.7825 ;
      RECT  23.1825 23.5975 23.3175 23.6625 ;
      RECT  23.405 22.86 23.4575 22.9225 ;
      RECT  22.9575 23.7475 23.0925 23.8125 ;
      RECT  22.835 23.0075 22.905 23.2975 ;
      RECT  22.94 23.2325 23.005 23.9725 ;
      RECT  23.455 23.8625 23.525 24.0625 ;
      RECT  23.375 23.0075 23.44 23.1425 ;
      RECT  22.7 22.86 22.7525 22.9225 ;
      RECT  22.695 24.0625 23.58 24.1275 ;
      RECT  22.7525 23.5 22.8175 23.635 ;
      RECT  23.07 22.7175 23.205 22.7825 ;
      RECT  23.375 23.0075 23.445 23.2975 ;
      RECT  23.0525 22.8575 23.1875 22.9225 ;
      RECT  22.755 23.8625 22.82 23.9975 ;
      RECT  23.27 23.2325 23.445 23.2975 ;
      RECT  23.27 23.8625 23.335 23.9975 ;
      RECT  22.695 22.7175 23.58 22.7825 ;
      RECT  23.4575 23.5 23.5225 23.635 ;
      RECT  22.75 23.3975 22.82 23.5325 ;
      RECT  23.02 23.0075 23.085 23.1425 ;
      RECT  23.27 23.3975 23.335 23.5325 ;
      RECT  23.2025 23.0075 23.2675 23.1425 ;
      RECT  22.755 23.3975 22.82 23.5325 ;
      RECT  22.94 23.8625 23.005 23.9975 ;
      RECT  23.27 23.2325 23.335 23.8625 ;
      RECT  22.7175 22.7175 22.8525 22.7825 ;
      RECT  22.835 23.0075 22.9 23.1425 ;
      RECT  22.94 24.7925 23.005 24.6575 ;
      RECT  23.455 24.7925 23.525 24.6575 ;
      RECT  22.835 24.9575 23.005 24.8925 ;
      RECT  22.695 25.3325 23.58 25.2675 ;
      RECT  22.75 24.3275 22.82 24.1275 ;
      RECT  23.455 24.3275 23.52 24.1925 ;
      RECT  23.0075 25.1825 23.0725 25.0475 ;
      RECT  23.19 25.1825 23.255 25.0475 ;
      RECT  23.455 24.7925 23.52 24.6575 ;
      RECT  23.4225 25.4725 23.5575 25.4075 ;
      RECT  23.1825 24.5925 23.3175 24.5275 ;
      RECT  23.405 25.33 23.4575 25.2675 ;
      RECT  22.9575 24.4425 23.0925 24.3775 ;
      RECT  22.835 25.1825 22.905 24.8925 ;
      RECT  22.94 24.9575 23.005 24.2175 ;
      RECT  23.455 24.3275 23.525 24.1275 ;
      RECT  23.375 25.1825 23.44 25.0475 ;
      RECT  22.7 25.33 22.7525 25.2675 ;
      RECT  22.695 24.1275 23.58 24.0625 ;
      RECT  22.7525 24.69 22.8175 24.555 ;
      RECT  23.07 25.4725 23.205 25.4075 ;
      RECT  23.375 25.1825 23.445 24.8925 ;
      RECT  23.0525 25.3325 23.1875 25.2675 ;
      RECT  22.755 24.3275 22.82 24.1925 ;
      RECT  23.27 24.9575 23.445 24.8925 ;
      RECT  23.27 24.3275 23.335 24.1925 ;
      RECT  22.695 25.4725 23.58 25.4075 ;
      RECT  23.4575 24.69 23.5225 24.555 ;
      RECT  22.75 24.7925 22.82 24.6575 ;
      RECT  23.02 25.1825 23.085 25.0475 ;
      RECT  23.27 24.7925 23.335 24.6575 ;
      RECT  23.2025 25.1825 23.2675 25.0475 ;
      RECT  22.755 24.7925 22.82 24.6575 ;
      RECT  22.94 24.3275 23.005 24.1925 ;
      RECT  23.27 24.9575 23.335 24.3275 ;
      RECT  22.7175 25.4725 22.8525 25.4075 ;
      RECT  22.835 25.1825 22.9 25.0475 ;
      RECT  22.94 26.0875 23.005 26.2225 ;
      RECT  23.455 26.0875 23.525 26.2225 ;
      RECT  22.835 25.9225 23.005 25.9875 ;
      RECT  22.695 25.5475 23.58 25.6125 ;
      RECT  22.75 26.5525 22.82 26.7525 ;
      RECT  23.455 26.5525 23.52 26.6875 ;
      RECT  23.0075 25.6975 23.0725 25.8325 ;
      RECT  23.19 25.6975 23.255 25.8325 ;
      RECT  23.455 26.0875 23.52 26.2225 ;
      RECT  23.4225 25.4075 23.5575 25.4725 ;
      RECT  23.1825 26.2875 23.3175 26.3525 ;
      RECT  23.405 25.55 23.4575 25.6125 ;
      RECT  22.9575 26.4375 23.0925 26.5025 ;
      RECT  22.835 25.6975 22.905 25.9875 ;
      RECT  22.94 25.9225 23.005 26.6625 ;
      RECT  23.455 26.5525 23.525 26.7525 ;
      RECT  23.375 25.6975 23.44 25.8325 ;
      RECT  22.7 25.55 22.7525 25.6125 ;
      RECT  22.695 26.7525 23.58 26.8175 ;
      RECT  22.7525 26.19 22.8175 26.325 ;
      RECT  23.07 25.4075 23.205 25.4725 ;
      RECT  23.375 25.6975 23.445 25.9875 ;
      RECT  23.0525 25.5475 23.1875 25.6125 ;
      RECT  22.755 26.5525 22.82 26.6875 ;
      RECT  23.27 25.9225 23.445 25.9875 ;
      RECT  23.27 26.5525 23.335 26.6875 ;
      RECT  22.695 25.4075 23.58 25.4725 ;
      RECT  23.4575 26.19 23.5225 26.325 ;
      RECT  22.75 26.0875 22.82 26.2225 ;
      RECT  23.02 25.6975 23.085 25.8325 ;
      RECT  23.27 26.0875 23.335 26.2225 ;
      RECT  23.2025 25.6975 23.2675 25.8325 ;
      RECT  22.755 26.0875 22.82 26.2225 ;
      RECT  22.94 26.5525 23.005 26.6875 ;
      RECT  23.27 25.9225 23.335 26.5525 ;
      RECT  22.7175 25.4075 22.8525 25.4725 ;
      RECT  22.835 25.6975 22.9 25.8325 ;
      RECT  22.94 27.4825 23.005 27.3475 ;
      RECT  23.455 27.4825 23.525 27.3475 ;
      RECT  22.835 27.6475 23.005 27.5825 ;
      RECT  22.695 28.0225 23.58 27.9575 ;
      RECT  22.75 27.0175 22.82 26.8175 ;
      RECT  23.455 27.0175 23.52 26.8825 ;
      RECT  23.0075 27.8725 23.0725 27.7375 ;
      RECT  23.19 27.8725 23.255 27.7375 ;
      RECT  23.455 27.4825 23.52 27.3475 ;
      RECT  23.4225 28.1625 23.5575 28.0975 ;
      RECT  23.1825 27.2825 23.3175 27.2175 ;
      RECT  23.405 28.02 23.4575 27.9575 ;
      RECT  22.9575 27.1325 23.0925 27.0675 ;
      RECT  22.835 27.8725 22.905 27.5825 ;
      RECT  22.94 27.6475 23.005 26.9075 ;
      RECT  23.455 27.0175 23.525 26.8175 ;
      RECT  23.375 27.8725 23.44 27.7375 ;
      RECT  22.7 28.02 22.7525 27.9575 ;
      RECT  22.695 26.8175 23.58 26.7525 ;
      RECT  22.7525 27.38 22.8175 27.245 ;
      RECT  23.07 28.1625 23.205 28.0975 ;
      RECT  23.375 27.8725 23.445 27.5825 ;
      RECT  23.0525 28.0225 23.1875 27.9575 ;
      RECT  22.755 27.0175 22.82 26.8825 ;
      RECT  23.27 27.6475 23.445 27.5825 ;
      RECT  23.27 27.0175 23.335 26.8825 ;
      RECT  22.695 28.1625 23.58 28.0975 ;
      RECT  23.4575 27.38 23.5225 27.245 ;
      RECT  22.75 27.4825 22.82 27.3475 ;
      RECT  23.02 27.8725 23.085 27.7375 ;
      RECT  23.27 27.4825 23.335 27.3475 ;
      RECT  23.2025 27.8725 23.2675 27.7375 ;
      RECT  22.755 27.4825 22.82 27.3475 ;
      RECT  22.94 27.0175 23.005 26.8825 ;
      RECT  23.27 27.6475 23.335 27.0175 ;
      RECT  22.7175 28.1625 22.8525 28.0975 ;
      RECT  22.835 27.8725 22.9 27.7375 ;
      RECT  22.94 28.7775 23.005 28.9125 ;
      RECT  23.455 28.7775 23.525 28.9125 ;
      RECT  22.835 28.6125 23.005 28.6775 ;
      RECT  22.695 28.2375 23.58 28.3025 ;
      RECT  22.75 29.2425 22.82 29.4425 ;
      RECT  23.455 29.2425 23.52 29.3775 ;
      RECT  23.0075 28.3875 23.0725 28.5225 ;
      RECT  23.19 28.3875 23.255 28.5225 ;
      RECT  23.455 28.7775 23.52 28.9125 ;
      RECT  23.4225 28.0975 23.5575 28.1625 ;
      RECT  23.1825 28.9775 23.3175 29.0425 ;
      RECT  23.405 28.24 23.4575 28.3025 ;
      RECT  22.9575 29.1275 23.0925 29.1925 ;
      RECT  22.835 28.3875 22.905 28.6775 ;
      RECT  22.94 28.6125 23.005 29.3525 ;
      RECT  23.455 29.2425 23.525 29.4425 ;
      RECT  23.375 28.3875 23.44 28.5225 ;
      RECT  22.7 28.24 22.7525 28.3025 ;
      RECT  22.695 29.4425 23.58 29.5075 ;
      RECT  22.7525 28.88 22.8175 29.015 ;
      RECT  23.07 28.0975 23.205 28.1625 ;
      RECT  23.375 28.3875 23.445 28.6775 ;
      RECT  23.0525 28.2375 23.1875 28.3025 ;
      RECT  22.755 29.2425 22.82 29.3775 ;
      RECT  23.27 28.6125 23.445 28.6775 ;
      RECT  23.27 29.2425 23.335 29.3775 ;
      RECT  22.695 28.0975 23.58 28.1625 ;
      RECT  23.4575 28.88 23.5225 29.015 ;
      RECT  22.75 28.7775 22.82 28.9125 ;
      RECT  23.02 28.3875 23.085 28.5225 ;
      RECT  23.27 28.7775 23.335 28.9125 ;
      RECT  23.2025 28.3875 23.2675 28.5225 ;
      RECT  22.755 28.7775 22.82 28.9125 ;
      RECT  22.94 29.2425 23.005 29.3775 ;
      RECT  23.27 28.6125 23.335 29.2425 ;
      RECT  22.7175 28.0975 22.8525 28.1625 ;
      RECT  22.835 28.3875 22.9 28.5225 ;
      RECT  22.94 30.1725 23.005 30.0375 ;
      RECT  23.455 30.1725 23.525 30.0375 ;
      RECT  22.835 30.3375 23.005 30.2725 ;
      RECT  22.695 30.7125 23.58 30.6475 ;
      RECT  22.75 29.7075 22.82 29.5075 ;
      RECT  23.455 29.7075 23.52 29.5725 ;
      RECT  23.0075 30.5625 23.0725 30.4275 ;
      RECT  23.19 30.5625 23.255 30.4275 ;
      RECT  23.455 30.1725 23.52 30.0375 ;
      RECT  23.4225 30.8525 23.5575 30.7875 ;
      RECT  23.1825 29.9725 23.3175 29.9075 ;
      RECT  23.405 30.71 23.4575 30.6475 ;
      RECT  22.9575 29.8225 23.0925 29.7575 ;
      RECT  22.835 30.5625 22.905 30.2725 ;
      RECT  22.94 30.3375 23.005 29.5975 ;
      RECT  23.455 29.7075 23.525 29.5075 ;
      RECT  23.375 30.5625 23.44 30.4275 ;
      RECT  22.7 30.71 22.7525 30.6475 ;
      RECT  22.695 29.5075 23.58 29.4425 ;
      RECT  22.7525 30.07 22.8175 29.935 ;
      RECT  23.07 30.8525 23.205 30.7875 ;
      RECT  23.375 30.5625 23.445 30.2725 ;
      RECT  23.0525 30.7125 23.1875 30.6475 ;
      RECT  22.755 29.7075 22.82 29.5725 ;
      RECT  23.27 30.3375 23.445 30.2725 ;
      RECT  23.27 29.7075 23.335 29.5725 ;
      RECT  22.695 30.8525 23.58 30.7875 ;
      RECT  23.4575 30.07 23.5225 29.935 ;
      RECT  22.75 30.1725 22.82 30.0375 ;
      RECT  23.02 30.5625 23.085 30.4275 ;
      RECT  23.27 30.1725 23.335 30.0375 ;
      RECT  23.2025 30.5625 23.2675 30.4275 ;
      RECT  22.755 30.1725 22.82 30.0375 ;
      RECT  22.94 29.7075 23.005 29.5725 ;
      RECT  23.27 30.3375 23.335 29.7075 ;
      RECT  22.7175 30.8525 22.8525 30.7875 ;
      RECT  22.835 30.5625 22.9 30.4275 ;
      RECT  22.94 31.4675 23.005 31.6025 ;
      RECT  23.455 31.4675 23.525 31.6025 ;
      RECT  22.835 31.3025 23.005 31.3675 ;
      RECT  22.695 30.9275 23.58 30.9925 ;
      RECT  22.75 31.9325 22.82 32.1325 ;
      RECT  23.455 31.9325 23.52 32.0675 ;
      RECT  23.0075 31.0775 23.0725 31.2125 ;
      RECT  23.19 31.0775 23.255 31.2125 ;
      RECT  23.455 31.4675 23.52 31.6025 ;
      RECT  23.4225 30.7875 23.5575 30.8525 ;
      RECT  23.1825 31.6675 23.3175 31.7325 ;
      RECT  23.405 30.93 23.4575 30.9925 ;
      RECT  22.9575 31.8175 23.0925 31.8825 ;
      RECT  22.835 31.0775 22.905 31.3675 ;
      RECT  22.94 31.3025 23.005 32.0425 ;
      RECT  23.455 31.9325 23.525 32.1325 ;
      RECT  23.375 31.0775 23.44 31.2125 ;
      RECT  22.7 30.93 22.7525 30.9925 ;
      RECT  22.695 32.1325 23.58 32.1975 ;
      RECT  22.7525 31.57 22.8175 31.705 ;
      RECT  23.07 30.7875 23.205 30.8525 ;
      RECT  23.375 31.0775 23.445 31.3675 ;
      RECT  23.0525 30.9275 23.1875 30.9925 ;
      RECT  22.755 31.9325 22.82 32.0675 ;
      RECT  23.27 31.3025 23.445 31.3675 ;
      RECT  23.27 31.9325 23.335 32.0675 ;
      RECT  22.695 30.7875 23.58 30.8525 ;
      RECT  23.4575 31.57 23.5225 31.705 ;
      RECT  22.75 31.4675 22.82 31.6025 ;
      RECT  23.02 31.0775 23.085 31.2125 ;
      RECT  23.27 31.4675 23.335 31.6025 ;
      RECT  23.2025 31.0775 23.2675 31.2125 ;
      RECT  22.755 31.4675 22.82 31.6025 ;
      RECT  22.94 31.9325 23.005 32.0675 ;
      RECT  23.27 31.3025 23.335 31.9325 ;
      RECT  22.7175 30.7875 22.8525 30.8525 ;
      RECT  22.835 31.0775 22.9 31.2125 ;
      RECT  22.94 32.8625 23.005 32.7275 ;
      RECT  23.455 32.8625 23.525 32.7275 ;
      RECT  22.835 33.0275 23.005 32.9625 ;
      RECT  22.695 33.4025 23.58 33.3375 ;
      RECT  22.75 32.3975 22.82 32.1975 ;
      RECT  23.455 32.3975 23.52 32.2625 ;
      RECT  23.0075 33.2525 23.0725 33.1175 ;
      RECT  23.19 33.2525 23.255 33.1175 ;
      RECT  23.455 32.8625 23.52 32.7275 ;
      RECT  23.4225 33.5425 23.5575 33.4775 ;
      RECT  23.1825 32.6625 23.3175 32.5975 ;
      RECT  23.405 33.4 23.4575 33.3375 ;
      RECT  22.9575 32.5125 23.0925 32.4475 ;
      RECT  22.835 33.2525 22.905 32.9625 ;
      RECT  22.94 33.0275 23.005 32.2875 ;
      RECT  23.455 32.3975 23.525 32.1975 ;
      RECT  23.375 33.2525 23.44 33.1175 ;
      RECT  22.7 33.4 22.7525 33.3375 ;
      RECT  22.695 32.1975 23.58 32.1325 ;
      RECT  22.7525 32.76 22.8175 32.625 ;
      RECT  23.07 33.5425 23.205 33.4775 ;
      RECT  23.375 33.2525 23.445 32.9625 ;
      RECT  23.0525 33.4025 23.1875 33.3375 ;
      RECT  22.755 32.3975 22.82 32.2625 ;
      RECT  23.27 33.0275 23.445 32.9625 ;
      RECT  23.27 32.3975 23.335 32.2625 ;
      RECT  22.695 33.5425 23.58 33.4775 ;
      RECT  23.4575 32.76 23.5225 32.625 ;
      RECT  22.75 32.8625 22.82 32.7275 ;
      RECT  23.02 33.2525 23.085 33.1175 ;
      RECT  23.27 32.8625 23.335 32.7275 ;
      RECT  23.2025 33.2525 23.2675 33.1175 ;
      RECT  22.755 32.8625 22.82 32.7275 ;
      RECT  22.94 32.3975 23.005 32.2625 ;
      RECT  23.27 33.0275 23.335 32.3975 ;
      RECT  22.7175 33.5425 22.8525 33.4775 ;
      RECT  22.835 33.2525 22.9 33.1175 ;
      RECT  22.94 34.1575 23.005 34.2925 ;
      RECT  23.455 34.1575 23.525 34.2925 ;
      RECT  22.835 33.9925 23.005 34.0575 ;
      RECT  22.695 33.6175 23.58 33.6825 ;
      RECT  22.75 34.6225 22.82 34.8225 ;
      RECT  23.455 34.6225 23.52 34.7575 ;
      RECT  23.0075 33.7675 23.0725 33.9025 ;
      RECT  23.19 33.7675 23.255 33.9025 ;
      RECT  23.455 34.1575 23.52 34.2925 ;
      RECT  23.4225 33.4775 23.5575 33.5425 ;
      RECT  23.1825 34.3575 23.3175 34.4225 ;
      RECT  23.405 33.62 23.4575 33.6825 ;
      RECT  22.9575 34.5075 23.0925 34.5725 ;
      RECT  22.835 33.7675 22.905 34.0575 ;
      RECT  22.94 33.9925 23.005 34.7325 ;
      RECT  23.455 34.6225 23.525 34.8225 ;
      RECT  23.375 33.7675 23.44 33.9025 ;
      RECT  22.7 33.62 22.7525 33.6825 ;
      RECT  22.695 34.8225 23.58 34.8875 ;
      RECT  22.7525 34.26 22.8175 34.395 ;
      RECT  23.07 33.4775 23.205 33.5425 ;
      RECT  23.375 33.7675 23.445 34.0575 ;
      RECT  23.0525 33.6175 23.1875 33.6825 ;
      RECT  22.755 34.6225 22.82 34.7575 ;
      RECT  23.27 33.9925 23.445 34.0575 ;
      RECT  23.27 34.6225 23.335 34.7575 ;
      RECT  22.695 33.4775 23.58 33.5425 ;
      RECT  23.4575 34.26 23.5225 34.395 ;
      RECT  22.75 34.1575 22.82 34.2925 ;
      RECT  23.02 33.7675 23.085 33.9025 ;
      RECT  23.27 34.1575 23.335 34.2925 ;
      RECT  23.2025 33.7675 23.2675 33.9025 ;
      RECT  22.755 34.1575 22.82 34.2925 ;
      RECT  22.94 34.6225 23.005 34.7575 ;
      RECT  23.27 33.9925 23.335 34.6225 ;
      RECT  22.7175 33.4775 22.8525 33.5425 ;
      RECT  22.835 33.7675 22.9 33.9025 ;
      RECT  22.94 35.5525 23.005 35.4175 ;
      RECT  23.455 35.5525 23.525 35.4175 ;
      RECT  22.835 35.7175 23.005 35.6525 ;
      RECT  22.695 36.0925 23.58 36.0275 ;
      RECT  22.75 35.0875 22.82 34.8875 ;
      RECT  23.455 35.0875 23.52 34.9525 ;
      RECT  23.0075 35.9425 23.0725 35.8075 ;
      RECT  23.19 35.9425 23.255 35.8075 ;
      RECT  23.455 35.5525 23.52 35.4175 ;
      RECT  23.4225 36.2325 23.5575 36.1675 ;
      RECT  23.1825 35.3525 23.3175 35.2875 ;
      RECT  23.405 36.09 23.4575 36.0275 ;
      RECT  22.9575 35.2025 23.0925 35.1375 ;
      RECT  22.835 35.9425 22.905 35.6525 ;
      RECT  22.94 35.7175 23.005 34.9775 ;
      RECT  23.455 35.0875 23.525 34.8875 ;
      RECT  23.375 35.9425 23.44 35.8075 ;
      RECT  22.7 36.09 22.7525 36.0275 ;
      RECT  22.695 34.8875 23.58 34.8225 ;
      RECT  22.7525 35.45 22.8175 35.315 ;
      RECT  23.07 36.2325 23.205 36.1675 ;
      RECT  23.375 35.9425 23.445 35.6525 ;
      RECT  23.0525 36.0925 23.1875 36.0275 ;
      RECT  22.755 35.0875 22.82 34.9525 ;
      RECT  23.27 35.7175 23.445 35.6525 ;
      RECT  23.27 35.0875 23.335 34.9525 ;
      RECT  22.695 36.2325 23.58 36.1675 ;
      RECT  23.4575 35.45 23.5225 35.315 ;
      RECT  22.75 35.5525 22.82 35.4175 ;
      RECT  23.02 35.9425 23.085 35.8075 ;
      RECT  23.27 35.5525 23.335 35.4175 ;
      RECT  23.2025 35.9425 23.2675 35.8075 ;
      RECT  22.755 35.5525 22.82 35.4175 ;
      RECT  22.94 35.0875 23.005 34.9525 ;
      RECT  23.27 35.7175 23.335 35.0875 ;
      RECT  22.7175 36.2325 22.8525 36.1675 ;
      RECT  22.835 35.9425 22.9 35.8075 ;
      RECT  22.94 36.8475 23.005 36.9825 ;
      RECT  23.455 36.8475 23.525 36.9825 ;
      RECT  22.835 36.6825 23.005 36.7475 ;
      RECT  22.695 36.3075 23.58 36.3725 ;
      RECT  22.75 37.3125 22.82 37.5125 ;
      RECT  23.455 37.3125 23.52 37.4475 ;
      RECT  23.0075 36.4575 23.0725 36.5925 ;
      RECT  23.19 36.4575 23.255 36.5925 ;
      RECT  23.455 36.8475 23.52 36.9825 ;
      RECT  23.4225 36.1675 23.5575 36.2325 ;
      RECT  23.1825 37.0475 23.3175 37.1125 ;
      RECT  23.405 36.31 23.4575 36.3725 ;
      RECT  22.9575 37.1975 23.0925 37.2625 ;
      RECT  22.835 36.4575 22.905 36.7475 ;
      RECT  22.94 36.6825 23.005 37.4225 ;
      RECT  23.455 37.3125 23.525 37.5125 ;
      RECT  23.375 36.4575 23.44 36.5925 ;
      RECT  22.7 36.31 22.7525 36.3725 ;
      RECT  22.695 37.5125 23.58 37.5775 ;
      RECT  22.7525 36.95 22.8175 37.085 ;
      RECT  23.07 36.1675 23.205 36.2325 ;
      RECT  23.375 36.4575 23.445 36.7475 ;
      RECT  23.0525 36.3075 23.1875 36.3725 ;
      RECT  22.755 37.3125 22.82 37.4475 ;
      RECT  23.27 36.6825 23.445 36.7475 ;
      RECT  23.27 37.3125 23.335 37.4475 ;
      RECT  22.695 36.1675 23.58 36.2325 ;
      RECT  23.4575 36.95 23.5225 37.085 ;
      RECT  22.75 36.8475 22.82 36.9825 ;
      RECT  23.02 36.4575 23.085 36.5925 ;
      RECT  23.27 36.8475 23.335 36.9825 ;
      RECT  23.2025 36.4575 23.2675 36.5925 ;
      RECT  22.755 36.8475 22.82 36.9825 ;
      RECT  22.94 37.3125 23.005 37.4475 ;
      RECT  23.27 36.6825 23.335 37.3125 ;
      RECT  22.7175 36.1675 22.8525 36.2325 ;
      RECT  22.835 36.4575 22.9 36.5925 ;
      RECT  22.94 38.2425 23.005 38.1075 ;
      RECT  23.455 38.2425 23.525 38.1075 ;
      RECT  22.835 38.4075 23.005 38.3425 ;
      RECT  22.695 38.7825 23.58 38.7175 ;
      RECT  22.75 37.7775 22.82 37.5775 ;
      RECT  23.455 37.7775 23.52 37.6425 ;
      RECT  23.0075 38.6325 23.0725 38.4975 ;
      RECT  23.19 38.6325 23.255 38.4975 ;
      RECT  23.455 38.2425 23.52 38.1075 ;
      RECT  23.4225 38.9225 23.5575 38.8575 ;
      RECT  23.1825 38.0425 23.3175 37.9775 ;
      RECT  23.405 38.78 23.4575 38.7175 ;
      RECT  22.9575 37.8925 23.0925 37.8275 ;
      RECT  22.835 38.6325 22.905 38.3425 ;
      RECT  22.94 38.4075 23.005 37.6675 ;
      RECT  23.455 37.7775 23.525 37.5775 ;
      RECT  23.375 38.6325 23.44 38.4975 ;
      RECT  22.7 38.78 22.7525 38.7175 ;
      RECT  22.695 37.5775 23.58 37.5125 ;
      RECT  22.7525 38.14 22.8175 38.005 ;
      RECT  23.07 38.9225 23.205 38.8575 ;
      RECT  23.375 38.6325 23.445 38.3425 ;
      RECT  23.0525 38.7825 23.1875 38.7175 ;
      RECT  22.755 37.7775 22.82 37.6425 ;
      RECT  23.27 38.4075 23.445 38.3425 ;
      RECT  23.27 37.7775 23.335 37.6425 ;
      RECT  22.695 38.9225 23.58 38.8575 ;
      RECT  23.4575 38.14 23.5225 38.005 ;
      RECT  22.75 38.2425 22.82 38.1075 ;
      RECT  23.02 38.6325 23.085 38.4975 ;
      RECT  23.27 38.2425 23.335 38.1075 ;
      RECT  23.2025 38.6325 23.2675 38.4975 ;
      RECT  22.755 38.2425 22.82 38.1075 ;
      RECT  22.94 37.7775 23.005 37.6425 ;
      RECT  23.27 38.4075 23.335 37.7775 ;
      RECT  22.7175 38.9225 22.8525 38.8575 ;
      RECT  22.835 38.6325 22.9 38.4975 ;
      RECT  22.94 39.5375 23.005 39.6725 ;
      RECT  23.455 39.5375 23.525 39.6725 ;
      RECT  22.835 39.3725 23.005 39.4375 ;
      RECT  22.695 38.9975 23.58 39.0625 ;
      RECT  22.75 40.0025 22.82 40.2025 ;
      RECT  23.455 40.0025 23.52 40.1375 ;
      RECT  23.0075 39.1475 23.0725 39.2825 ;
      RECT  23.19 39.1475 23.255 39.2825 ;
      RECT  23.455 39.5375 23.52 39.6725 ;
      RECT  23.4225 38.8575 23.5575 38.9225 ;
      RECT  23.1825 39.7375 23.3175 39.8025 ;
      RECT  23.405 39.0 23.4575 39.0625 ;
      RECT  22.9575 39.8875 23.0925 39.9525 ;
      RECT  22.835 39.1475 22.905 39.4375 ;
      RECT  22.94 39.3725 23.005 40.1125 ;
      RECT  23.455 40.0025 23.525 40.2025 ;
      RECT  23.375 39.1475 23.44 39.2825 ;
      RECT  22.7 39.0 22.7525 39.0625 ;
      RECT  22.695 40.2025 23.58 40.2675 ;
      RECT  22.7525 39.64 22.8175 39.775 ;
      RECT  23.07 38.8575 23.205 38.9225 ;
      RECT  23.375 39.1475 23.445 39.4375 ;
      RECT  23.0525 38.9975 23.1875 39.0625 ;
      RECT  22.755 40.0025 22.82 40.1375 ;
      RECT  23.27 39.3725 23.445 39.4375 ;
      RECT  23.27 40.0025 23.335 40.1375 ;
      RECT  22.695 38.8575 23.58 38.9225 ;
      RECT  23.4575 39.64 23.5225 39.775 ;
      RECT  22.75 39.5375 22.82 39.6725 ;
      RECT  23.02 39.1475 23.085 39.2825 ;
      RECT  23.27 39.5375 23.335 39.6725 ;
      RECT  23.2025 39.1475 23.2675 39.2825 ;
      RECT  22.755 39.5375 22.82 39.6725 ;
      RECT  22.94 40.0025 23.005 40.1375 ;
      RECT  23.27 39.3725 23.335 40.0025 ;
      RECT  22.7175 38.8575 22.8525 38.9225 ;
      RECT  22.835 39.1475 22.9 39.2825 ;
      RECT  22.94 40.9325 23.005 40.7975 ;
      RECT  23.455 40.9325 23.525 40.7975 ;
      RECT  22.835 41.0975 23.005 41.0325 ;
      RECT  22.695 41.4725 23.58 41.4075 ;
      RECT  22.75 40.4675 22.82 40.2675 ;
      RECT  23.455 40.4675 23.52 40.3325 ;
      RECT  23.0075 41.3225 23.0725 41.1875 ;
      RECT  23.19 41.3225 23.255 41.1875 ;
      RECT  23.455 40.9325 23.52 40.7975 ;
      RECT  23.4225 41.6125 23.5575 41.5475 ;
      RECT  23.1825 40.7325 23.3175 40.6675 ;
      RECT  23.405 41.47 23.4575 41.4075 ;
      RECT  22.9575 40.5825 23.0925 40.5175 ;
      RECT  22.835 41.3225 22.905 41.0325 ;
      RECT  22.94 41.0975 23.005 40.3575 ;
      RECT  23.455 40.4675 23.525 40.2675 ;
      RECT  23.375 41.3225 23.44 41.1875 ;
      RECT  22.7 41.47 22.7525 41.4075 ;
      RECT  22.695 40.2675 23.58 40.2025 ;
      RECT  22.7525 40.83 22.8175 40.695 ;
      RECT  23.07 41.6125 23.205 41.5475 ;
      RECT  23.375 41.3225 23.445 41.0325 ;
      RECT  23.0525 41.4725 23.1875 41.4075 ;
      RECT  22.755 40.4675 22.82 40.3325 ;
      RECT  23.27 41.0975 23.445 41.0325 ;
      RECT  23.27 40.4675 23.335 40.3325 ;
      RECT  22.695 41.6125 23.58 41.5475 ;
      RECT  23.4575 40.83 23.5225 40.695 ;
      RECT  22.75 40.9325 22.82 40.7975 ;
      RECT  23.02 41.3225 23.085 41.1875 ;
      RECT  23.27 40.9325 23.335 40.7975 ;
      RECT  23.2025 41.3225 23.2675 41.1875 ;
      RECT  22.755 40.9325 22.82 40.7975 ;
      RECT  22.94 40.4675 23.005 40.3325 ;
      RECT  23.27 41.0975 23.335 40.4675 ;
      RECT  22.7175 41.6125 22.8525 41.5475 ;
      RECT  22.835 41.3225 22.9 41.1875 ;
      RECT  22.94 42.2275 23.005 42.3625 ;
      RECT  23.455 42.2275 23.525 42.3625 ;
      RECT  22.835 42.0625 23.005 42.1275 ;
      RECT  22.695 41.6875 23.58 41.7525 ;
      RECT  22.75 42.6925 22.82 42.8925 ;
      RECT  23.455 42.6925 23.52 42.8275 ;
      RECT  23.0075 41.8375 23.0725 41.9725 ;
      RECT  23.19 41.8375 23.255 41.9725 ;
      RECT  23.455 42.2275 23.52 42.3625 ;
      RECT  23.4225 41.5475 23.5575 41.6125 ;
      RECT  23.1825 42.4275 23.3175 42.4925 ;
      RECT  23.405 41.69 23.4575 41.7525 ;
      RECT  22.9575 42.5775 23.0925 42.6425 ;
      RECT  22.835 41.8375 22.905 42.1275 ;
      RECT  22.94 42.0625 23.005 42.8025 ;
      RECT  23.455 42.6925 23.525 42.8925 ;
      RECT  23.375 41.8375 23.44 41.9725 ;
      RECT  22.7 41.69 22.7525 41.7525 ;
      RECT  22.695 42.8925 23.58 42.9575 ;
      RECT  22.7525 42.33 22.8175 42.465 ;
      RECT  23.07 41.5475 23.205 41.6125 ;
      RECT  23.375 41.8375 23.445 42.1275 ;
      RECT  23.0525 41.6875 23.1875 41.7525 ;
      RECT  22.755 42.6925 22.82 42.8275 ;
      RECT  23.27 42.0625 23.445 42.1275 ;
      RECT  23.27 42.6925 23.335 42.8275 ;
      RECT  22.695 41.5475 23.58 41.6125 ;
      RECT  23.4575 42.33 23.5225 42.465 ;
      RECT  22.75 42.2275 22.82 42.3625 ;
      RECT  23.02 41.8375 23.085 41.9725 ;
      RECT  23.27 42.2275 23.335 42.3625 ;
      RECT  23.2025 41.8375 23.2675 41.9725 ;
      RECT  22.755 42.2275 22.82 42.3625 ;
      RECT  22.94 42.6925 23.005 42.8275 ;
      RECT  23.27 42.0625 23.335 42.6925 ;
      RECT  22.7175 41.5475 22.8525 41.6125 ;
      RECT  22.835 41.8375 22.9 41.9725 ;
      RECT  22.94 43.6225 23.005 43.4875 ;
      RECT  23.455 43.6225 23.525 43.4875 ;
      RECT  22.835 43.7875 23.005 43.7225 ;
      RECT  22.695 44.1625 23.58 44.0975 ;
      RECT  22.75 43.1575 22.82 42.9575 ;
      RECT  23.455 43.1575 23.52 43.0225 ;
      RECT  23.0075 44.0125 23.0725 43.8775 ;
      RECT  23.19 44.0125 23.255 43.8775 ;
      RECT  23.455 43.6225 23.52 43.4875 ;
      RECT  23.4225 44.3025 23.5575 44.2375 ;
      RECT  23.1825 43.4225 23.3175 43.3575 ;
      RECT  23.405 44.16 23.4575 44.0975 ;
      RECT  22.9575 43.2725 23.0925 43.2075 ;
      RECT  22.835 44.0125 22.905 43.7225 ;
      RECT  22.94 43.7875 23.005 43.0475 ;
      RECT  23.455 43.1575 23.525 42.9575 ;
      RECT  23.375 44.0125 23.44 43.8775 ;
      RECT  22.7 44.16 22.7525 44.0975 ;
      RECT  22.695 42.9575 23.58 42.8925 ;
      RECT  22.7525 43.52 22.8175 43.385 ;
      RECT  23.07 44.3025 23.205 44.2375 ;
      RECT  23.375 44.0125 23.445 43.7225 ;
      RECT  23.0525 44.1625 23.1875 44.0975 ;
      RECT  22.755 43.1575 22.82 43.0225 ;
      RECT  23.27 43.7875 23.445 43.7225 ;
      RECT  23.27 43.1575 23.335 43.0225 ;
      RECT  22.695 44.3025 23.58 44.2375 ;
      RECT  23.4575 43.52 23.5225 43.385 ;
      RECT  22.75 43.6225 22.82 43.4875 ;
      RECT  23.02 44.0125 23.085 43.8775 ;
      RECT  23.27 43.6225 23.335 43.4875 ;
      RECT  23.2025 44.0125 23.2675 43.8775 ;
      RECT  22.755 43.6225 22.82 43.4875 ;
      RECT  22.94 43.1575 23.005 43.0225 ;
      RECT  23.27 43.7875 23.335 43.1575 ;
      RECT  22.7175 44.3025 22.8525 44.2375 ;
      RECT  22.835 44.0125 22.9 43.8775 ;
      RECT  22.94 44.9175 23.005 45.0525 ;
      RECT  23.455 44.9175 23.525 45.0525 ;
      RECT  22.835 44.7525 23.005 44.8175 ;
      RECT  22.695 44.3775 23.58 44.4425 ;
      RECT  22.75 45.3825 22.82 45.5825 ;
      RECT  23.455 45.3825 23.52 45.5175 ;
      RECT  23.0075 44.5275 23.0725 44.6625 ;
      RECT  23.19 44.5275 23.255 44.6625 ;
      RECT  23.455 44.9175 23.52 45.0525 ;
      RECT  23.4225 44.2375 23.5575 44.3025 ;
      RECT  23.1825 45.1175 23.3175 45.1825 ;
      RECT  23.405 44.38 23.4575 44.4425 ;
      RECT  22.9575 45.2675 23.0925 45.3325 ;
      RECT  22.835 44.5275 22.905 44.8175 ;
      RECT  22.94 44.7525 23.005 45.4925 ;
      RECT  23.455 45.3825 23.525 45.5825 ;
      RECT  23.375 44.5275 23.44 44.6625 ;
      RECT  22.7 44.38 22.7525 44.4425 ;
      RECT  22.695 45.5825 23.58 45.6475 ;
      RECT  22.7525 45.02 22.8175 45.155 ;
      RECT  23.07 44.2375 23.205 44.3025 ;
      RECT  23.375 44.5275 23.445 44.8175 ;
      RECT  23.0525 44.3775 23.1875 44.4425 ;
      RECT  22.755 45.3825 22.82 45.5175 ;
      RECT  23.27 44.7525 23.445 44.8175 ;
      RECT  23.27 45.3825 23.335 45.5175 ;
      RECT  22.695 44.2375 23.58 44.3025 ;
      RECT  23.4575 45.02 23.5225 45.155 ;
      RECT  22.75 44.9175 22.82 45.0525 ;
      RECT  23.02 44.5275 23.085 44.6625 ;
      RECT  23.27 44.9175 23.335 45.0525 ;
      RECT  23.2025 44.5275 23.2675 44.6625 ;
      RECT  22.755 44.9175 22.82 45.0525 ;
      RECT  22.94 45.3825 23.005 45.5175 ;
      RECT  23.27 44.7525 23.335 45.3825 ;
      RECT  22.7175 44.2375 22.8525 44.3025 ;
      RECT  22.835 44.5275 22.9 44.6625 ;
      RECT  22.785 20.1675 23.49 20.2325 ;
      RECT  22.785 22.5775 23.49 22.6425 ;
      RECT  22.785 22.8575 23.49 22.9225 ;
      RECT  22.785 25.2675 23.49 25.3325 ;
      RECT  22.785 25.5475 23.49 25.6125 ;
      RECT  22.785 27.9575 23.49 28.0225 ;
      RECT  22.785 28.2375 23.49 28.3025 ;
      RECT  22.785 30.6475 23.49 30.7125 ;
      RECT  22.785 30.9275 23.49 30.9925 ;
      RECT  22.785 33.3375 23.49 33.4025 ;
      RECT  22.785 33.6175 23.49 33.6825 ;
      RECT  22.785 36.0275 23.49 36.0925 ;
      RECT  22.785 36.3075 23.49 36.3725 ;
      RECT  22.785 38.7175 23.49 38.7825 ;
      RECT  22.785 38.9975 23.49 39.0625 ;
      RECT  22.785 41.4075 23.49 41.4725 ;
      RECT  22.785 41.6875 23.49 41.7525 ;
      RECT  22.785 44.0975 23.49 44.1625 ;
      RECT  22.785 44.3775 23.49 44.4425 ;
      RECT  19.77 22.5775 23.685 22.6425 ;
      RECT  19.77 22.8575 23.685 22.9225 ;
      RECT  19.77 25.2675 23.685 25.3325 ;
      RECT  19.77 25.5475 23.685 25.6125 ;
      RECT  19.77 27.9575 23.685 28.0225 ;
      RECT  19.77 28.2375 23.685 28.3025 ;
      RECT  19.77 30.6475 23.685 30.7125 ;
      RECT  19.77 30.9275 23.685 30.9925 ;
      RECT  19.77 33.3375 23.685 33.4025 ;
      RECT  19.77 33.6175 23.685 33.6825 ;
      RECT  19.77 36.0275 23.685 36.0925 ;
      RECT  19.77 36.3075 23.685 36.3725 ;
      RECT  19.77 38.7175 23.685 38.7825 ;
      RECT  19.77 38.9975 23.685 39.0625 ;
      RECT  19.77 41.4075 23.685 41.4725 ;
      RECT  19.77 41.6875 23.685 41.7525 ;
      RECT  19.77 44.0975 23.685 44.1625 ;
      RECT  21.01 18.5025 21.075 18.6375 ;
      RECT  20.795 18.5025 20.86 18.6375 ;
      RECT  21.01 19.0525 21.075 19.1875 ;
      RECT  20.795 19.0525 20.86 19.1875 ;
      RECT  21.225 19.0525 21.29 19.1875 ;
      RECT  21.01 19.0525 21.075 19.1875 ;
      RECT  20.67 18.17 21.375 18.235 ;
      RECT  21.715 18.5025 21.78 18.6375 ;
      RECT  21.5 18.5025 21.565 18.6375 ;
      RECT  21.715 19.0525 21.78 19.1875 ;
      RECT  21.5 19.0525 21.565 19.1875 ;
      RECT  21.93 19.0525 21.995 19.1875 ;
      RECT  21.715 19.0525 21.78 19.1875 ;
      RECT  21.375 18.17 22.08 18.235 ;
      RECT  22.42 18.5025 22.485 18.6375 ;
      RECT  22.205 18.5025 22.27 18.6375 ;
      RECT  22.42 19.0525 22.485 19.1875 ;
      RECT  22.205 19.0525 22.27 19.1875 ;
      RECT  22.635 19.0525 22.7 19.1875 ;
      RECT  22.42 19.0525 22.485 19.1875 ;
      RECT  22.08 18.17 22.785 18.235 ;
      RECT  19.77 18.17 22.785 18.235 ;
      RECT  21.8825 14.545 21.9475 15.24 ;
      RECT  21.3775 13.1525 22.005 13.2225 ;
      RECT  21.5075 16.5225 21.5725 16.7975 ;
      RECT  21.7925 16.98 21.8575 17.255 ;
      RECT  21.7925 17.3975 22.115 17.4625 ;
      RECT  21.5025 14.135 21.5675 14.27 ;
      RECT  21.5075 16.3575 21.7975 16.4225 ;
      RECT  22.0325 17.3275 22.0475 17.3975 ;
      RECT  21.66 13.2925 21.795 13.3575 ;
      RECT  21.6075 16.98 21.6725 17.255 ;
      RECT  21.695 14.2025 21.76 14.4 ;
      RECT  21.3775 13.0875 21.4425 13.2225 ;
      RECT  21.9675 17.0975 22.0325 17.2325 ;
      RECT  21.5075 14.4 21.5725 15.4975 ;
      RECT  21.8825 15.66 21.9475 16.5225 ;
      RECT  21.9675 17.2325 22.0325 17.4625 ;
      RECT  21.605 17.5275 21.67 17.5925 ;
      RECT  21.6375 16.1225 21.7025 16.2575 ;
      RECT  21.695 15.435 21.76 15.57 ;
      RECT  21.5075 15.66 21.5725 16.5275 ;
      RECT  21.6975 16.5225 21.7625 16.7975 ;
      RECT  21.6575 16.74 21.7275 17.0675 ;
      RECT  21.34 17.5275 22.115 17.5925 ;
      RECT  21.5075 15.4975 21.5725 16.0525 ;
      RECT  21.6925 13.575 21.7575 14.27 ;
      RECT  21.665 17.5275 21.8 17.5925 ;
      RECT  21.5075 14.335 22.005 14.4 ;
      RECT  21.6975 14.545 21.7625 15.24 ;
      RECT  21.6975 15.175 21.7625 15.37 ;
      RECT  21.695 13.2925 21.76 13.4275 ;
      RECT  21.8825 15.305 21.9475 15.5 ;
      RECT  21.6575 16.1575 21.9475 16.2225 ;
      RECT  21.6925 15.4975 21.7575 16.0525 ;
      RECT  21.885 14.545 21.95 14.68 ;
      RECT  21.8825 16.5225 21.9475 16.7975 ;
      RECT  21.7925 17.245 21.8575 17.3975 ;
      RECT  22.0475 17.3275 22.1125 17.4625 ;
      RECT  21.7525 16.3225 21.8175 16.4575 ;
      RECT  21.6975 15.305 21.9475 15.37 ;
      RECT  21.5075 13.575 21.5725 14.27 ;
      RECT  21.6975 15.4975 21.7625 16.0525 ;
      RECT  21.94 13.1525 22.005 14.4 ;
      RECT  21.8825 15.4975 21.9475 16.0525 ;
      RECT  21.6925 16.5225 21.7575 16.7975 ;
      RECT  22.5875 14.545 22.6525 15.24 ;
      RECT  22.0825 13.1525 22.71 13.2225 ;
      RECT  22.2125 16.5225 22.2775 16.7975 ;
      RECT  22.4975 16.98 22.5625 17.255 ;
      RECT  22.4975 17.3975 22.82 17.4625 ;
      RECT  22.2075 14.135 22.2725 14.27 ;
      RECT  22.2125 16.3575 22.5025 16.4225 ;
      RECT  22.7375 17.3275 22.7525 17.3975 ;
      RECT  22.365 13.2925 22.5 13.3575 ;
      RECT  22.3125 16.98 22.3775 17.255 ;
      RECT  22.4 14.2025 22.465 14.4 ;
      RECT  22.0825 13.0875 22.1475 13.2225 ;
      RECT  22.6725 17.0975 22.7375 17.2325 ;
      RECT  22.2125 14.4 22.2775 15.4975 ;
      RECT  22.5875 15.66 22.6525 16.5225 ;
      RECT  22.6725 17.2325 22.7375 17.4625 ;
      RECT  22.31 17.5275 22.375 17.5925 ;
      RECT  22.3425 16.1225 22.4075 16.2575 ;
      RECT  22.4 15.435 22.465 15.57 ;
      RECT  22.2125 15.66 22.2775 16.5275 ;
      RECT  22.4025 16.5225 22.4675 16.7975 ;
      RECT  22.3625 16.74 22.4325 17.0675 ;
      RECT  22.045 17.5275 22.82 17.5925 ;
      RECT  22.2125 15.4975 22.2775 16.0525 ;
      RECT  22.3975 13.575 22.4625 14.27 ;
      RECT  22.37 17.5275 22.505 17.5925 ;
      RECT  22.2125 14.335 22.71 14.4 ;
      RECT  22.4025 14.545 22.4675 15.24 ;
      RECT  22.4025 15.175 22.4675 15.37 ;
      RECT  22.4 13.2925 22.465 13.4275 ;
      RECT  22.5875 15.305 22.6525 15.5 ;
      RECT  22.3625 16.1575 22.6525 16.2225 ;
      RECT  22.3975 15.4975 22.4625 16.0525 ;
      RECT  22.59 14.545 22.655 14.68 ;
      RECT  22.5875 16.5225 22.6525 16.7975 ;
      RECT  22.4975 17.245 22.5625 17.3975 ;
      RECT  22.7525 17.3275 22.8175 17.4625 ;
      RECT  22.4575 16.3225 22.5225 16.4575 ;
      RECT  22.4025 15.305 22.6525 15.37 ;
      RECT  22.2125 13.575 22.2775 14.27 ;
      RECT  22.4025 15.4975 22.4675 16.0525 ;
      RECT  22.645 13.1525 22.71 14.4 ;
      RECT  22.5875 15.4975 22.6525 16.0525 ;
      RECT  22.3975 16.5225 22.4625 16.7975 ;
      RECT  19.77 17.5275 22.785 17.5925 ;
      RECT  21.6575 9.7225 21.82 9.7875 ;
      RECT  22.025 9.88 22.0475 10.015 ;
      RECT  21.41 9.515 21.42 9.65 ;
      RECT  21.42 9.515 21.485 9.65 ;
      RECT  21.42 8.6075 21.485 8.825 ;
      RECT  21.42 8.5425 22.01 8.6075 ;
      RECT  22.0475 9.31 22.1125 9.445 ;
      RECT  21.795 11.4275 21.86 11.8075 ;
      RECT  21.945 9.515 22.01 9.65 ;
      RECT  21.605 9.515 21.67 9.65 ;
      RECT  21.42 8.825 21.485 9.24 ;
      RECT  21.795 11.0125 21.86 11.4275 ;
      RECT  22.0275 11.8075 22.0475 11.9425 ;
      RECT  21.795 10.395 21.86 10.81 ;
      RECT  21.795 11.8075 21.86 11.9425 ;
      RECT  21.7925 9.88 21.8575 10.015 ;
      RECT  21.4775 8.2825 21.6125 8.3475 ;
      RECT  21.5275 12.0175 21.5925 12.1525 ;
      RECT  21.3425 10.8425 21.4075 10.9775 ;
      RECT  21.4025 9.88 21.415 10.015 ;
      RECT  21.4825 10.795 21.5475 10.93 ;
      RECT  21.47 10.795 21.485 10.93 ;
      RECT  22.0475 9.515 22.1125 9.65 ;
      RECT  21.6225 11.485 21.6875 11.62 ;
      RECT  21.96 9.88 22.025 10.015 ;
      RECT  21.755 9.5975 21.82 9.7225 ;
      RECT  21.42 11.8075 21.485 11.9425 ;
      RECT  21.3425 11.8075 21.4075 11.9425 ;
      RECT  21.5825 8.28 21.7175 8.345 ;
      RECT  21.41 9.88 21.42 10.015 ;
      RECT  21.525 12.0175 21.86 12.0825 ;
      RECT  21.42 9.88 21.485 10.015 ;
      RECT  21.34 9.345 22.115 9.41 ;
      RECT  21.645 8.6925 21.78 8.7575 ;
      RECT  21.7925 10.395 21.8575 10.53 ;
      RECT  21.6575 9.7225 21.7225 10.32 ;
      RECT  21.6775 8.6075 21.7425 8.7575 ;
      RECT  21.6225 9.515 21.6875 9.65 ;
      RECT  21.9625 11.8075 22.0275 11.9425 ;
      RECT  21.7625 9.515 21.8275 9.65 ;
      RECT  21.795 11.9425 21.86 12.0175 ;
      RECT  21.56 11.485 21.625 11.62 ;
      RECT  21.48 8.5425 21.615 8.6075 ;
      RECT  21.6575 10.235 21.7225 10.37 ;
      RECT  21.42 8.4125 22.01 8.4775 ;
      RECT  21.42 10.395 21.485 10.81 ;
      RECT  21.4025 9.515 21.415 9.65 ;
      RECT  21.945 8.6075 22.01 8.825 ;
      RECT  21.6225 9.105 21.6875 9.24 ;
      RECT  21.7625 9.105 21.8275 9.24 ;
      RECT  22.0475 11.8075 22.1125 11.9425 ;
      RECT  21.795 9.88 21.86 10.015 ;
      RECT  21.945 8.825 22.01 9.24 ;
      RECT  21.605 8.825 21.67 9.24 ;
      RECT  21.41 11.8075 21.42 11.9425 ;
      RECT  21.3425 9.515 21.4075 9.65 ;
      RECT  21.3425 9.31 21.4075 9.445 ;
      RECT  21.42 11.0125 21.485 11.4275 ;
      RECT  21.42 10.81 21.485 11.0125 ;
      RECT  21.4075 10.8425 21.55 10.9775 ;
      RECT  21.76 9.515 21.825 9.65 ;
      RECT  21.4025 11.8075 21.415 11.9425 ;
      RECT  22.0475 9.88 22.1125 10.015 ;
      RECT  22.005 9.515 22.0475 9.65 ;
      RECT  21.3425 9.88 21.4075 10.015 ;
      RECT  21.76 8.825 21.825 9.24 ;
      RECT  22.3625 9.7225 22.525 9.7875 ;
      RECT  22.73 9.88 22.7525 10.015 ;
      RECT  22.115 9.515 22.125 9.65 ;
      RECT  22.125 9.515 22.19 9.65 ;
      RECT  22.125 8.6075 22.19 8.825 ;
      RECT  22.125 8.5425 22.715 8.6075 ;
      RECT  22.7525 9.31 22.8175 9.445 ;
      RECT  22.5 11.4275 22.565 11.8075 ;
      RECT  22.65 9.515 22.715 9.65 ;
      RECT  22.31 9.515 22.375 9.65 ;
      RECT  22.125 8.825 22.19 9.24 ;
      RECT  22.5 11.0125 22.565 11.4275 ;
      RECT  22.7325 11.8075 22.7525 11.9425 ;
      RECT  22.5 10.395 22.565 10.81 ;
      RECT  22.5 11.8075 22.565 11.9425 ;
      RECT  22.4975 9.88 22.5625 10.015 ;
      RECT  22.1825 8.2825 22.3175 8.3475 ;
      RECT  22.2325 12.0175 22.2975 12.1525 ;
      RECT  22.0475 10.8425 22.1125 10.9775 ;
      RECT  22.1075 9.88 22.12 10.015 ;
      RECT  22.1875 10.795 22.2525 10.93 ;
      RECT  22.175 10.795 22.19 10.93 ;
      RECT  22.7525 9.515 22.8175 9.65 ;
      RECT  22.3275 11.485 22.3925 11.62 ;
      RECT  22.665 9.88 22.73 10.015 ;
      RECT  22.46 9.5975 22.525 9.7225 ;
      RECT  22.125 11.8075 22.19 11.9425 ;
      RECT  22.0475 11.8075 22.1125 11.9425 ;
      RECT  22.2875 8.28 22.4225 8.345 ;
      RECT  22.115 9.88 22.125 10.015 ;
      RECT  22.23 12.0175 22.565 12.0825 ;
      RECT  22.125 9.88 22.19 10.015 ;
      RECT  22.045 9.345 22.82 9.41 ;
      RECT  22.35 8.6925 22.485 8.7575 ;
      RECT  22.4975 10.395 22.5625 10.53 ;
      RECT  22.3625 9.7225 22.4275 10.32 ;
      RECT  22.3825 8.6075 22.4475 8.7575 ;
      RECT  22.3275 9.515 22.3925 9.65 ;
      RECT  22.6675 11.8075 22.7325 11.9425 ;
      RECT  22.4675 9.515 22.5325 9.65 ;
      RECT  22.5 11.9425 22.565 12.0175 ;
      RECT  22.265 11.485 22.33 11.62 ;
      RECT  22.185 8.5425 22.32 8.6075 ;
      RECT  22.3625 10.235 22.4275 10.37 ;
      RECT  22.125 8.4125 22.715 8.4775 ;
      RECT  22.125 10.395 22.19 10.81 ;
      RECT  22.1075 9.515 22.12 9.65 ;
      RECT  22.65 8.6075 22.715 8.825 ;
      RECT  22.3275 9.105 22.3925 9.24 ;
      RECT  22.4675 9.105 22.5325 9.24 ;
      RECT  22.7525 11.8075 22.8175 11.9425 ;
      RECT  22.5 9.88 22.565 10.015 ;
      RECT  22.65 8.825 22.715 9.24 ;
      RECT  22.31 8.825 22.375 9.24 ;
      RECT  22.115 11.8075 22.125 11.9425 ;
      RECT  22.0475 9.515 22.1125 9.65 ;
      RECT  22.0475 9.31 22.1125 9.445 ;
      RECT  22.125 11.0125 22.19 11.4275 ;
      RECT  22.125 10.81 22.19 11.0125 ;
      RECT  22.1125 10.8425 22.255 10.9775 ;
      RECT  22.465 9.515 22.53 9.65 ;
      RECT  22.1075 11.8075 22.12 11.9425 ;
      RECT  22.7525 9.88 22.8175 10.015 ;
      RECT  22.71 9.515 22.7525 9.65 ;
      RECT  22.0475 9.88 22.1125 10.015 ;
      RECT  22.465 8.825 22.53 9.24 ;
      RECT  19.77 8.4125 22.785 8.4775 ;
      RECT  19.77 17.5925 22.785 17.5275 ;
      RECT  19.77 18.235 22.785 18.17 ;
      RECT  19.77 8.4775 22.785 8.4125 ;
      RECT  11.4775 23.7675 11.5425 23.9025 ;
      RECT  11.2625 23.7675 11.3275 23.9025 ;
      RECT  11.4775 22.8525 11.5425 22.9875 ;
      RECT  11.2625 22.8525 11.3275 22.9875 ;
      RECT  11.2425 23.345 11.3775 23.41 ;
      RECT  11.51 23.345 11.575 23.41 ;
      RECT  11.17 24.0625 11.8575 24.1275 ;
      RECT  11.17 22.7175 11.8575 22.7825 ;
      RECT  11.4775 24.4225 11.5425 24.2875 ;
      RECT  11.2625 24.4225 11.3275 24.2875 ;
      RECT  11.4775 25.3375 11.5425 25.2025 ;
      RECT  11.2625 25.3375 11.3275 25.2025 ;
      RECT  11.2425 24.845 11.3775 24.78 ;
      RECT  11.51 24.845 11.575 24.78 ;
      RECT  11.17 24.1275 11.8575 24.0625 ;
      RECT  11.17 25.4725 11.8575 25.4075 ;
      RECT  13.005 23.7675 13.07 23.9025 ;
      RECT  12.79 23.7675 12.855 23.9025 ;
      RECT  13.22 23.7675 13.285 23.9025 ;
      RECT  13.005 23.7675 13.07 23.9025 ;
      RECT  12.79 22.8975 12.855 23.0325 ;
      RECT  13.22 22.8975 13.285 23.0325 ;
      RECT  12.8625 23.145 12.9975 23.21 ;
      RECT  13.0775 23.425 13.2125 23.49 ;
      RECT  13.35 23.6375 13.415 23.7025 ;
      RECT  12.6975 24.0625 13.6 24.1275 ;
      RECT  12.6975 22.7175 13.6 22.7825 ;
      RECT  13.9075 23.7675 13.9725 23.9025 ;
      RECT  13.6925 23.7675 13.7575 23.9025 ;
      RECT  13.9075 22.8525 13.9725 22.9875 ;
      RECT  13.6925 22.8525 13.7575 22.9875 ;
      RECT  13.6725 23.345 13.8075 23.41 ;
      RECT  13.94 23.345 14.005 23.41 ;
      RECT  13.6 24.0625 14.2875 24.1275 ;
      RECT  13.6 22.7175 14.2875 22.7825 ;
      RECT  12.8625 23.145 12.9975 23.21 ;
      RECT  13.0775 23.425 13.2125 23.49 ;
      RECT  13.94 23.345 14.005 23.41 ;
      RECT  12.6975 24.0625 14.2875 24.1275 ;
      RECT  12.6975 22.7175 14.2875 22.7825 ;
      RECT  13.005 24.4225 13.07 24.2875 ;
      RECT  12.79 24.4225 12.855 24.2875 ;
      RECT  13.22 24.4225 13.285 24.2875 ;
      RECT  13.005 24.4225 13.07 24.2875 ;
      RECT  12.79 25.2925 12.855 25.1575 ;
      RECT  13.22 25.2925 13.285 25.1575 ;
      RECT  12.8625 25.045 12.9975 24.98 ;
      RECT  13.0775 24.765 13.2125 24.7 ;
      RECT  13.35 24.5525 13.415 24.4875 ;
      RECT  12.6975 24.1275 13.6 24.0625 ;
      RECT  12.6975 25.4725 13.6 25.4075 ;
      RECT  13.9075 24.4225 13.9725 24.2875 ;
      RECT  13.6925 24.4225 13.7575 24.2875 ;
      RECT  13.9075 25.3375 13.9725 25.2025 ;
      RECT  13.6925 25.3375 13.7575 25.2025 ;
      RECT  13.6725 24.845 13.8075 24.78 ;
      RECT  13.94 24.845 14.005 24.78 ;
      RECT  13.6 24.1275 14.2875 24.0625 ;
      RECT  13.6 25.4725 14.2875 25.4075 ;
      RECT  12.8625 25.045 12.9975 24.98 ;
      RECT  13.0775 24.765 13.2125 24.7 ;
      RECT  13.94 24.845 14.005 24.78 ;
      RECT  12.6975 24.1275 14.2875 24.0625 ;
      RECT  12.6975 25.4725 14.2875 25.4075 ;
      RECT  13.005 26.4575 13.07 26.5925 ;
      RECT  12.79 26.4575 12.855 26.5925 ;
      RECT  13.22 26.4575 13.285 26.5925 ;
      RECT  13.005 26.4575 13.07 26.5925 ;
      RECT  12.79 25.5875 12.855 25.7225 ;
      RECT  13.22 25.5875 13.285 25.7225 ;
      RECT  12.8625 25.835 12.9975 25.9 ;
      RECT  13.0775 26.115 13.2125 26.18 ;
      RECT  13.35 26.3275 13.415 26.3925 ;
      RECT  12.6975 26.7525 13.6 26.8175 ;
      RECT  12.6975 25.4075 13.6 25.4725 ;
      RECT  13.9075 26.4575 13.9725 26.5925 ;
      RECT  13.6925 26.4575 13.7575 26.5925 ;
      RECT  13.9075 25.5425 13.9725 25.6775 ;
      RECT  13.6925 25.5425 13.7575 25.6775 ;
      RECT  13.6725 26.035 13.8075 26.1 ;
      RECT  13.94 26.035 14.005 26.1 ;
      RECT  13.6 26.7525 14.2875 26.8175 ;
      RECT  13.6 25.4075 14.2875 25.4725 ;
      RECT  12.8625 25.835 12.9975 25.9 ;
      RECT  13.0775 26.115 13.2125 26.18 ;
      RECT  13.94 26.035 14.005 26.1 ;
      RECT  12.6975 26.7525 14.2875 26.8175 ;
      RECT  12.6975 25.4075 14.2875 25.4725 ;
      RECT  13.005 27.1125 13.07 26.9775 ;
      RECT  12.79 27.1125 12.855 26.9775 ;
      RECT  13.22 27.1125 13.285 26.9775 ;
      RECT  13.005 27.1125 13.07 26.9775 ;
      RECT  12.79 27.9825 12.855 27.8475 ;
      RECT  13.22 27.9825 13.285 27.8475 ;
      RECT  12.8625 27.735 12.9975 27.67 ;
      RECT  13.0775 27.455 13.2125 27.39 ;
      RECT  13.35 27.2425 13.415 27.1775 ;
      RECT  12.6975 26.8175 13.6 26.7525 ;
      RECT  12.6975 28.1625 13.6 28.0975 ;
      RECT  13.9075 27.1125 13.9725 26.9775 ;
      RECT  13.6925 27.1125 13.7575 26.9775 ;
      RECT  13.9075 28.0275 13.9725 27.8925 ;
      RECT  13.6925 28.0275 13.7575 27.8925 ;
      RECT  13.6725 27.535 13.8075 27.47 ;
      RECT  13.94 27.535 14.005 27.47 ;
      RECT  13.6 26.8175 14.2875 26.7525 ;
      RECT  13.6 28.1625 14.2875 28.0975 ;
      RECT  12.8625 27.735 12.9975 27.67 ;
      RECT  13.0775 27.455 13.2125 27.39 ;
      RECT  13.94 27.535 14.005 27.47 ;
      RECT  12.6975 26.8175 14.2875 26.7525 ;
      RECT  12.6975 28.1625 14.2875 28.0975 ;
      RECT  13.94 23.345 14.005 23.41 ;
      RECT  13.94 24.78 14.005 24.845 ;
      RECT  13.94 26.035 14.005 26.1 ;
      RECT  13.94 27.47 14.005 27.535 ;
      RECT  11.4775 31.8375 11.5425 31.9725 ;
      RECT  11.2625 31.8375 11.3275 31.9725 ;
      RECT  11.4775 30.9225 11.5425 31.0575 ;
      RECT  11.2625 30.9225 11.3275 31.0575 ;
      RECT  11.2425 31.415 11.3775 31.48 ;
      RECT  11.51 31.415 11.575 31.48 ;
      RECT  11.17 32.1325 11.8575 32.1975 ;
      RECT  11.17 30.7875 11.8575 30.8525 ;
      RECT  11.4775 32.4925 11.5425 32.3575 ;
      RECT  11.2625 32.4925 11.3275 32.3575 ;
      RECT  11.4775 33.4075 11.5425 33.2725 ;
      RECT  11.2625 33.4075 11.3275 33.2725 ;
      RECT  11.2425 32.915 11.3775 32.85 ;
      RECT  11.51 32.915 11.575 32.85 ;
      RECT  11.17 32.1975 11.8575 32.1325 ;
      RECT  11.17 33.5425 11.8575 33.4775 ;
      RECT  13.005 31.8375 13.07 31.9725 ;
      RECT  12.79 31.8375 12.855 31.9725 ;
      RECT  13.22 31.8375 13.285 31.9725 ;
      RECT  13.005 31.8375 13.07 31.9725 ;
      RECT  12.79 30.9675 12.855 31.1025 ;
      RECT  13.22 30.9675 13.285 31.1025 ;
      RECT  12.8625 31.215 12.9975 31.28 ;
      RECT  13.0775 31.495 13.2125 31.56 ;
      RECT  13.35 31.7075 13.415 31.7725 ;
      RECT  12.6975 32.1325 13.6 32.1975 ;
      RECT  12.6975 30.7875 13.6 30.8525 ;
      RECT  13.9075 31.8375 13.9725 31.9725 ;
      RECT  13.6925 31.8375 13.7575 31.9725 ;
      RECT  13.9075 30.9225 13.9725 31.0575 ;
      RECT  13.6925 30.9225 13.7575 31.0575 ;
      RECT  13.6725 31.415 13.8075 31.48 ;
      RECT  13.94 31.415 14.005 31.48 ;
      RECT  13.6 32.1325 14.2875 32.1975 ;
      RECT  13.6 30.7875 14.2875 30.8525 ;
      RECT  12.8625 31.215 12.9975 31.28 ;
      RECT  13.0775 31.495 13.2125 31.56 ;
      RECT  13.94 31.415 14.005 31.48 ;
      RECT  12.6975 32.1325 14.2875 32.1975 ;
      RECT  12.6975 30.7875 14.2875 30.8525 ;
      RECT  13.005 32.4925 13.07 32.3575 ;
      RECT  12.79 32.4925 12.855 32.3575 ;
      RECT  13.22 32.4925 13.285 32.3575 ;
      RECT  13.005 32.4925 13.07 32.3575 ;
      RECT  12.79 33.3625 12.855 33.2275 ;
      RECT  13.22 33.3625 13.285 33.2275 ;
      RECT  12.8625 33.115 12.9975 33.05 ;
      RECT  13.0775 32.835 13.2125 32.77 ;
      RECT  13.35 32.6225 13.415 32.5575 ;
      RECT  12.6975 32.1975 13.6 32.1325 ;
      RECT  12.6975 33.5425 13.6 33.4775 ;
      RECT  13.9075 32.4925 13.9725 32.3575 ;
      RECT  13.6925 32.4925 13.7575 32.3575 ;
      RECT  13.9075 33.4075 13.9725 33.2725 ;
      RECT  13.6925 33.4075 13.7575 33.2725 ;
      RECT  13.6725 32.915 13.8075 32.85 ;
      RECT  13.94 32.915 14.005 32.85 ;
      RECT  13.6 32.1975 14.2875 32.1325 ;
      RECT  13.6 33.5425 14.2875 33.4775 ;
      RECT  12.8625 33.115 12.9975 33.05 ;
      RECT  13.0775 32.835 13.2125 32.77 ;
      RECT  13.94 32.915 14.005 32.85 ;
      RECT  12.6975 32.1975 14.2875 32.1325 ;
      RECT  12.6975 33.5425 14.2875 33.4775 ;
      RECT  13.005 34.5275 13.07 34.6625 ;
      RECT  12.79 34.5275 12.855 34.6625 ;
      RECT  13.22 34.5275 13.285 34.6625 ;
      RECT  13.005 34.5275 13.07 34.6625 ;
      RECT  12.79 33.6575 12.855 33.7925 ;
      RECT  13.22 33.6575 13.285 33.7925 ;
      RECT  12.8625 33.905 12.9975 33.97 ;
      RECT  13.0775 34.185 13.2125 34.25 ;
      RECT  13.35 34.3975 13.415 34.4625 ;
      RECT  12.6975 34.8225 13.6 34.8875 ;
      RECT  12.6975 33.4775 13.6 33.5425 ;
      RECT  13.9075 34.5275 13.9725 34.6625 ;
      RECT  13.6925 34.5275 13.7575 34.6625 ;
      RECT  13.9075 33.6125 13.9725 33.7475 ;
      RECT  13.6925 33.6125 13.7575 33.7475 ;
      RECT  13.6725 34.105 13.8075 34.17 ;
      RECT  13.94 34.105 14.005 34.17 ;
      RECT  13.6 34.8225 14.2875 34.8875 ;
      RECT  13.6 33.4775 14.2875 33.5425 ;
      RECT  12.8625 33.905 12.9975 33.97 ;
      RECT  13.0775 34.185 13.2125 34.25 ;
      RECT  13.94 34.105 14.005 34.17 ;
      RECT  12.6975 34.8225 14.2875 34.8875 ;
      RECT  12.6975 33.4775 14.2875 33.5425 ;
      RECT  13.005 35.1825 13.07 35.0475 ;
      RECT  12.79 35.1825 12.855 35.0475 ;
      RECT  13.22 35.1825 13.285 35.0475 ;
      RECT  13.005 35.1825 13.07 35.0475 ;
      RECT  12.79 36.0525 12.855 35.9175 ;
      RECT  13.22 36.0525 13.285 35.9175 ;
      RECT  12.8625 35.805 12.9975 35.74 ;
      RECT  13.0775 35.525 13.2125 35.46 ;
      RECT  13.35 35.3125 13.415 35.2475 ;
      RECT  12.6975 34.8875 13.6 34.8225 ;
      RECT  12.6975 36.2325 13.6 36.1675 ;
      RECT  13.9075 35.1825 13.9725 35.0475 ;
      RECT  13.6925 35.1825 13.7575 35.0475 ;
      RECT  13.9075 36.0975 13.9725 35.9625 ;
      RECT  13.6925 36.0975 13.7575 35.9625 ;
      RECT  13.6725 35.605 13.8075 35.54 ;
      RECT  13.94 35.605 14.005 35.54 ;
      RECT  13.6 34.8875 14.2875 34.8225 ;
      RECT  13.6 36.2325 14.2875 36.1675 ;
      RECT  12.8625 35.805 12.9975 35.74 ;
      RECT  13.0775 35.525 13.2125 35.46 ;
      RECT  13.94 35.605 14.005 35.54 ;
      RECT  12.6975 34.8875 14.2875 34.8225 ;
      RECT  12.6975 36.2325 14.2875 36.1675 ;
      RECT  13.94 31.415 14.005 31.48 ;
      RECT  13.94 32.85 14.005 32.915 ;
      RECT  13.94 34.105 14.005 34.17 ;
      RECT  13.94 35.54 14.005 35.605 ;
      RECT  15.855 23.7675 15.92 23.9025 ;
      RECT  15.64 23.7675 15.705 23.9025 ;
      RECT  16.07 23.7675 16.135 23.9025 ;
      RECT  15.855 23.7675 15.92 23.9025 ;
      RECT  15.64 22.8975 15.705 23.0325 ;
      RECT  16.07 22.8975 16.135 23.0325 ;
      RECT  15.7125 23.145 15.8475 23.21 ;
      RECT  15.9275 23.425 16.0625 23.49 ;
      RECT  16.2 23.6375 16.265 23.7025 ;
      RECT  15.5475 24.0625 16.45 24.1275 ;
      RECT  15.5475 22.7175 16.45 22.7825 ;
      RECT  16.7575 23.7675 16.8225 23.9025 ;
      RECT  16.5425 23.7675 16.6075 23.9025 ;
      RECT  16.7575 22.8525 16.8225 22.9875 ;
      RECT  16.5425 22.8525 16.6075 22.9875 ;
      RECT  16.5225 23.345 16.6575 23.41 ;
      RECT  16.79 23.345 16.855 23.41 ;
      RECT  16.45 24.0625 17.1375 24.1275 ;
      RECT  16.45 22.7175 17.1375 22.7825 ;
      RECT  15.7125 23.145 15.8475 23.21 ;
      RECT  15.9275 23.425 16.0625 23.49 ;
      RECT  16.79 23.345 16.855 23.41 ;
      RECT  15.5475 24.0625 17.1375 24.1275 ;
      RECT  15.5475 22.7175 17.1375 22.7825 ;
      RECT  15.855 24.4225 15.92 24.2875 ;
      RECT  15.64 24.4225 15.705 24.2875 ;
      RECT  16.07 24.4225 16.135 24.2875 ;
      RECT  15.855 24.4225 15.92 24.2875 ;
      RECT  15.64 25.2925 15.705 25.1575 ;
      RECT  16.07 25.2925 16.135 25.1575 ;
      RECT  15.7125 25.045 15.8475 24.98 ;
      RECT  15.9275 24.765 16.0625 24.7 ;
      RECT  16.2 24.5525 16.265 24.4875 ;
      RECT  15.5475 24.1275 16.45 24.0625 ;
      RECT  15.5475 25.4725 16.45 25.4075 ;
      RECT  16.7575 24.4225 16.8225 24.2875 ;
      RECT  16.5425 24.4225 16.6075 24.2875 ;
      RECT  16.7575 25.3375 16.8225 25.2025 ;
      RECT  16.5425 25.3375 16.6075 25.2025 ;
      RECT  16.5225 24.845 16.6575 24.78 ;
      RECT  16.79 24.845 16.855 24.78 ;
      RECT  16.45 24.1275 17.1375 24.0625 ;
      RECT  16.45 25.4725 17.1375 25.4075 ;
      RECT  15.7125 25.045 15.8475 24.98 ;
      RECT  15.9275 24.765 16.0625 24.7 ;
      RECT  16.79 24.845 16.855 24.78 ;
      RECT  15.5475 24.1275 17.1375 24.0625 ;
      RECT  15.5475 25.4725 17.1375 25.4075 ;
      RECT  15.855 26.4575 15.92 26.5925 ;
      RECT  15.64 26.4575 15.705 26.5925 ;
      RECT  16.07 26.4575 16.135 26.5925 ;
      RECT  15.855 26.4575 15.92 26.5925 ;
      RECT  15.64 25.5875 15.705 25.7225 ;
      RECT  16.07 25.5875 16.135 25.7225 ;
      RECT  15.7125 25.835 15.8475 25.9 ;
      RECT  15.9275 26.115 16.0625 26.18 ;
      RECT  16.2 26.3275 16.265 26.3925 ;
      RECT  15.5475 26.7525 16.45 26.8175 ;
      RECT  15.5475 25.4075 16.45 25.4725 ;
      RECT  16.7575 26.4575 16.8225 26.5925 ;
      RECT  16.5425 26.4575 16.6075 26.5925 ;
      RECT  16.7575 25.5425 16.8225 25.6775 ;
      RECT  16.5425 25.5425 16.6075 25.6775 ;
      RECT  16.5225 26.035 16.6575 26.1 ;
      RECT  16.79 26.035 16.855 26.1 ;
      RECT  16.45 26.7525 17.1375 26.8175 ;
      RECT  16.45 25.4075 17.1375 25.4725 ;
      RECT  15.7125 25.835 15.8475 25.9 ;
      RECT  15.9275 26.115 16.0625 26.18 ;
      RECT  16.79 26.035 16.855 26.1 ;
      RECT  15.5475 26.7525 17.1375 26.8175 ;
      RECT  15.5475 25.4075 17.1375 25.4725 ;
      RECT  15.855 27.1125 15.92 26.9775 ;
      RECT  15.64 27.1125 15.705 26.9775 ;
      RECT  16.07 27.1125 16.135 26.9775 ;
      RECT  15.855 27.1125 15.92 26.9775 ;
      RECT  15.64 27.9825 15.705 27.8475 ;
      RECT  16.07 27.9825 16.135 27.8475 ;
      RECT  15.7125 27.735 15.8475 27.67 ;
      RECT  15.9275 27.455 16.0625 27.39 ;
      RECT  16.2 27.2425 16.265 27.1775 ;
      RECT  15.5475 26.8175 16.45 26.7525 ;
      RECT  15.5475 28.1625 16.45 28.0975 ;
      RECT  16.7575 27.1125 16.8225 26.9775 ;
      RECT  16.5425 27.1125 16.6075 26.9775 ;
      RECT  16.7575 28.0275 16.8225 27.8925 ;
      RECT  16.5425 28.0275 16.6075 27.8925 ;
      RECT  16.5225 27.535 16.6575 27.47 ;
      RECT  16.79 27.535 16.855 27.47 ;
      RECT  16.45 26.8175 17.1375 26.7525 ;
      RECT  16.45 28.1625 17.1375 28.0975 ;
      RECT  15.7125 27.735 15.8475 27.67 ;
      RECT  15.9275 27.455 16.0625 27.39 ;
      RECT  16.79 27.535 16.855 27.47 ;
      RECT  15.5475 26.8175 17.1375 26.7525 ;
      RECT  15.5475 28.1625 17.1375 28.0975 ;
      RECT  15.855 29.1475 15.92 29.2825 ;
      RECT  15.64 29.1475 15.705 29.2825 ;
      RECT  16.07 29.1475 16.135 29.2825 ;
      RECT  15.855 29.1475 15.92 29.2825 ;
      RECT  15.64 28.2775 15.705 28.4125 ;
      RECT  16.07 28.2775 16.135 28.4125 ;
      RECT  15.7125 28.525 15.8475 28.59 ;
      RECT  15.9275 28.805 16.0625 28.87 ;
      RECT  16.2 29.0175 16.265 29.0825 ;
      RECT  15.5475 29.4425 16.45 29.5075 ;
      RECT  15.5475 28.0975 16.45 28.1625 ;
      RECT  16.7575 29.1475 16.8225 29.2825 ;
      RECT  16.5425 29.1475 16.6075 29.2825 ;
      RECT  16.7575 28.2325 16.8225 28.3675 ;
      RECT  16.5425 28.2325 16.6075 28.3675 ;
      RECT  16.5225 28.725 16.6575 28.79 ;
      RECT  16.79 28.725 16.855 28.79 ;
      RECT  16.45 29.4425 17.1375 29.5075 ;
      RECT  16.45 28.0975 17.1375 28.1625 ;
      RECT  15.7125 28.525 15.8475 28.59 ;
      RECT  15.9275 28.805 16.0625 28.87 ;
      RECT  16.79 28.725 16.855 28.79 ;
      RECT  15.5475 29.4425 17.1375 29.5075 ;
      RECT  15.5475 28.0975 17.1375 28.1625 ;
      RECT  15.855 29.8025 15.92 29.6675 ;
      RECT  15.64 29.8025 15.705 29.6675 ;
      RECT  16.07 29.8025 16.135 29.6675 ;
      RECT  15.855 29.8025 15.92 29.6675 ;
      RECT  15.64 30.6725 15.705 30.5375 ;
      RECT  16.07 30.6725 16.135 30.5375 ;
      RECT  15.7125 30.425 15.8475 30.36 ;
      RECT  15.9275 30.145 16.0625 30.08 ;
      RECT  16.2 29.9325 16.265 29.8675 ;
      RECT  15.5475 29.5075 16.45 29.4425 ;
      RECT  15.5475 30.8525 16.45 30.7875 ;
      RECT  16.7575 29.8025 16.8225 29.6675 ;
      RECT  16.5425 29.8025 16.6075 29.6675 ;
      RECT  16.7575 30.7175 16.8225 30.5825 ;
      RECT  16.5425 30.7175 16.6075 30.5825 ;
      RECT  16.5225 30.225 16.6575 30.16 ;
      RECT  16.79 30.225 16.855 30.16 ;
      RECT  16.45 29.5075 17.1375 29.4425 ;
      RECT  16.45 30.8525 17.1375 30.7875 ;
      RECT  15.7125 30.425 15.8475 30.36 ;
      RECT  15.9275 30.145 16.0625 30.08 ;
      RECT  16.79 30.225 16.855 30.16 ;
      RECT  15.5475 29.5075 17.1375 29.4425 ;
      RECT  15.5475 30.8525 17.1375 30.7875 ;
      RECT  15.855 31.8375 15.92 31.9725 ;
      RECT  15.64 31.8375 15.705 31.9725 ;
      RECT  16.07 31.8375 16.135 31.9725 ;
      RECT  15.855 31.8375 15.92 31.9725 ;
      RECT  15.64 30.9675 15.705 31.1025 ;
      RECT  16.07 30.9675 16.135 31.1025 ;
      RECT  15.7125 31.215 15.8475 31.28 ;
      RECT  15.9275 31.495 16.0625 31.56 ;
      RECT  16.2 31.7075 16.265 31.7725 ;
      RECT  15.5475 32.1325 16.45 32.1975 ;
      RECT  15.5475 30.7875 16.45 30.8525 ;
      RECT  16.7575 31.8375 16.8225 31.9725 ;
      RECT  16.5425 31.8375 16.6075 31.9725 ;
      RECT  16.7575 30.9225 16.8225 31.0575 ;
      RECT  16.5425 30.9225 16.6075 31.0575 ;
      RECT  16.5225 31.415 16.6575 31.48 ;
      RECT  16.79 31.415 16.855 31.48 ;
      RECT  16.45 32.1325 17.1375 32.1975 ;
      RECT  16.45 30.7875 17.1375 30.8525 ;
      RECT  15.7125 31.215 15.8475 31.28 ;
      RECT  15.9275 31.495 16.0625 31.56 ;
      RECT  16.79 31.415 16.855 31.48 ;
      RECT  15.5475 32.1325 17.1375 32.1975 ;
      RECT  15.5475 30.7875 17.1375 30.8525 ;
      RECT  15.855 32.4925 15.92 32.3575 ;
      RECT  15.64 32.4925 15.705 32.3575 ;
      RECT  16.07 32.4925 16.135 32.3575 ;
      RECT  15.855 32.4925 15.92 32.3575 ;
      RECT  15.64 33.3625 15.705 33.2275 ;
      RECT  16.07 33.3625 16.135 33.2275 ;
      RECT  15.7125 33.115 15.8475 33.05 ;
      RECT  15.9275 32.835 16.0625 32.77 ;
      RECT  16.2 32.6225 16.265 32.5575 ;
      RECT  15.5475 32.1975 16.45 32.1325 ;
      RECT  15.5475 33.5425 16.45 33.4775 ;
      RECT  16.7575 32.4925 16.8225 32.3575 ;
      RECT  16.5425 32.4925 16.6075 32.3575 ;
      RECT  16.7575 33.4075 16.8225 33.2725 ;
      RECT  16.5425 33.4075 16.6075 33.2725 ;
      RECT  16.5225 32.915 16.6575 32.85 ;
      RECT  16.79 32.915 16.855 32.85 ;
      RECT  16.45 32.1975 17.1375 32.1325 ;
      RECT  16.45 33.5425 17.1375 33.4775 ;
      RECT  15.7125 33.115 15.8475 33.05 ;
      RECT  15.9275 32.835 16.0625 32.77 ;
      RECT  16.79 32.915 16.855 32.85 ;
      RECT  15.5475 32.1975 17.1375 32.1325 ;
      RECT  15.5475 33.5425 17.1375 33.4775 ;
      RECT  15.855 34.5275 15.92 34.6625 ;
      RECT  15.64 34.5275 15.705 34.6625 ;
      RECT  16.07 34.5275 16.135 34.6625 ;
      RECT  15.855 34.5275 15.92 34.6625 ;
      RECT  15.64 33.6575 15.705 33.7925 ;
      RECT  16.07 33.6575 16.135 33.7925 ;
      RECT  15.7125 33.905 15.8475 33.97 ;
      RECT  15.9275 34.185 16.0625 34.25 ;
      RECT  16.2 34.3975 16.265 34.4625 ;
      RECT  15.5475 34.8225 16.45 34.8875 ;
      RECT  15.5475 33.4775 16.45 33.5425 ;
      RECT  16.7575 34.5275 16.8225 34.6625 ;
      RECT  16.5425 34.5275 16.6075 34.6625 ;
      RECT  16.7575 33.6125 16.8225 33.7475 ;
      RECT  16.5425 33.6125 16.6075 33.7475 ;
      RECT  16.5225 34.105 16.6575 34.17 ;
      RECT  16.79 34.105 16.855 34.17 ;
      RECT  16.45 34.8225 17.1375 34.8875 ;
      RECT  16.45 33.4775 17.1375 33.5425 ;
      RECT  15.7125 33.905 15.8475 33.97 ;
      RECT  15.9275 34.185 16.0625 34.25 ;
      RECT  16.79 34.105 16.855 34.17 ;
      RECT  15.5475 34.8225 17.1375 34.8875 ;
      RECT  15.5475 33.4775 17.1375 33.5425 ;
      RECT  15.855 35.1825 15.92 35.0475 ;
      RECT  15.64 35.1825 15.705 35.0475 ;
      RECT  16.07 35.1825 16.135 35.0475 ;
      RECT  15.855 35.1825 15.92 35.0475 ;
      RECT  15.64 36.0525 15.705 35.9175 ;
      RECT  16.07 36.0525 16.135 35.9175 ;
      RECT  15.7125 35.805 15.8475 35.74 ;
      RECT  15.9275 35.525 16.0625 35.46 ;
      RECT  16.2 35.3125 16.265 35.2475 ;
      RECT  15.5475 34.8875 16.45 34.8225 ;
      RECT  15.5475 36.2325 16.45 36.1675 ;
      RECT  16.7575 35.1825 16.8225 35.0475 ;
      RECT  16.5425 35.1825 16.6075 35.0475 ;
      RECT  16.7575 36.0975 16.8225 35.9625 ;
      RECT  16.5425 36.0975 16.6075 35.9625 ;
      RECT  16.5225 35.605 16.6575 35.54 ;
      RECT  16.79 35.605 16.855 35.54 ;
      RECT  16.45 34.8875 17.1375 34.8225 ;
      RECT  16.45 36.2325 17.1375 36.1675 ;
      RECT  15.7125 35.805 15.8475 35.74 ;
      RECT  15.9275 35.525 16.0625 35.46 ;
      RECT  16.79 35.605 16.855 35.54 ;
      RECT  15.5475 34.8875 17.1375 34.8225 ;
      RECT  15.5475 36.2325 17.1375 36.1675 ;
      RECT  15.855 37.2175 15.92 37.3525 ;
      RECT  15.64 37.2175 15.705 37.3525 ;
      RECT  16.07 37.2175 16.135 37.3525 ;
      RECT  15.855 37.2175 15.92 37.3525 ;
      RECT  15.64 36.3475 15.705 36.4825 ;
      RECT  16.07 36.3475 16.135 36.4825 ;
      RECT  15.7125 36.595 15.8475 36.66 ;
      RECT  15.9275 36.875 16.0625 36.94 ;
      RECT  16.2 37.0875 16.265 37.1525 ;
      RECT  15.5475 37.5125 16.45 37.5775 ;
      RECT  15.5475 36.1675 16.45 36.2325 ;
      RECT  16.7575 37.2175 16.8225 37.3525 ;
      RECT  16.5425 37.2175 16.6075 37.3525 ;
      RECT  16.7575 36.3025 16.8225 36.4375 ;
      RECT  16.5425 36.3025 16.6075 36.4375 ;
      RECT  16.5225 36.795 16.6575 36.86 ;
      RECT  16.79 36.795 16.855 36.86 ;
      RECT  16.45 37.5125 17.1375 37.5775 ;
      RECT  16.45 36.1675 17.1375 36.2325 ;
      RECT  15.7125 36.595 15.8475 36.66 ;
      RECT  15.9275 36.875 16.0625 36.94 ;
      RECT  16.79 36.795 16.855 36.86 ;
      RECT  15.5475 37.5125 17.1375 37.5775 ;
      RECT  15.5475 36.1675 17.1375 36.2325 ;
      RECT  15.855 37.8725 15.92 37.7375 ;
      RECT  15.64 37.8725 15.705 37.7375 ;
      RECT  16.07 37.8725 16.135 37.7375 ;
      RECT  15.855 37.8725 15.92 37.7375 ;
      RECT  15.64 38.7425 15.705 38.6075 ;
      RECT  16.07 38.7425 16.135 38.6075 ;
      RECT  15.7125 38.495 15.8475 38.43 ;
      RECT  15.9275 38.215 16.0625 38.15 ;
      RECT  16.2 38.0025 16.265 37.9375 ;
      RECT  15.5475 37.5775 16.45 37.5125 ;
      RECT  15.5475 38.9225 16.45 38.8575 ;
      RECT  16.7575 37.8725 16.8225 37.7375 ;
      RECT  16.5425 37.8725 16.6075 37.7375 ;
      RECT  16.7575 38.7875 16.8225 38.6525 ;
      RECT  16.5425 38.7875 16.6075 38.6525 ;
      RECT  16.5225 38.295 16.6575 38.23 ;
      RECT  16.79 38.295 16.855 38.23 ;
      RECT  16.45 37.5775 17.1375 37.5125 ;
      RECT  16.45 38.9225 17.1375 38.8575 ;
      RECT  15.7125 38.495 15.8475 38.43 ;
      RECT  15.9275 38.215 16.0625 38.15 ;
      RECT  16.79 38.295 16.855 38.23 ;
      RECT  15.5475 37.5775 17.1375 37.5125 ;
      RECT  15.5475 38.9225 17.1375 38.8575 ;
      RECT  15.855 39.9075 15.92 40.0425 ;
      RECT  15.64 39.9075 15.705 40.0425 ;
      RECT  16.07 39.9075 16.135 40.0425 ;
      RECT  15.855 39.9075 15.92 40.0425 ;
      RECT  15.64 39.0375 15.705 39.1725 ;
      RECT  16.07 39.0375 16.135 39.1725 ;
      RECT  15.7125 39.285 15.8475 39.35 ;
      RECT  15.9275 39.565 16.0625 39.63 ;
      RECT  16.2 39.7775 16.265 39.8425 ;
      RECT  15.5475 40.2025 16.45 40.2675 ;
      RECT  15.5475 38.8575 16.45 38.9225 ;
      RECT  16.7575 39.9075 16.8225 40.0425 ;
      RECT  16.5425 39.9075 16.6075 40.0425 ;
      RECT  16.7575 38.9925 16.8225 39.1275 ;
      RECT  16.5425 38.9925 16.6075 39.1275 ;
      RECT  16.5225 39.485 16.6575 39.55 ;
      RECT  16.79 39.485 16.855 39.55 ;
      RECT  16.45 40.2025 17.1375 40.2675 ;
      RECT  16.45 38.8575 17.1375 38.9225 ;
      RECT  15.7125 39.285 15.8475 39.35 ;
      RECT  15.9275 39.565 16.0625 39.63 ;
      RECT  16.79 39.485 16.855 39.55 ;
      RECT  15.5475 40.2025 17.1375 40.2675 ;
      RECT  15.5475 38.8575 17.1375 38.9225 ;
      RECT  15.855 40.5625 15.92 40.4275 ;
      RECT  15.64 40.5625 15.705 40.4275 ;
      RECT  16.07 40.5625 16.135 40.4275 ;
      RECT  15.855 40.5625 15.92 40.4275 ;
      RECT  15.64 41.4325 15.705 41.2975 ;
      RECT  16.07 41.4325 16.135 41.2975 ;
      RECT  15.7125 41.185 15.8475 41.12 ;
      RECT  15.9275 40.905 16.0625 40.84 ;
      RECT  16.2 40.6925 16.265 40.6275 ;
      RECT  15.5475 40.2675 16.45 40.2025 ;
      RECT  15.5475 41.6125 16.45 41.5475 ;
      RECT  16.7575 40.5625 16.8225 40.4275 ;
      RECT  16.5425 40.5625 16.6075 40.4275 ;
      RECT  16.7575 41.4775 16.8225 41.3425 ;
      RECT  16.5425 41.4775 16.6075 41.3425 ;
      RECT  16.5225 40.985 16.6575 40.92 ;
      RECT  16.79 40.985 16.855 40.92 ;
      RECT  16.45 40.2675 17.1375 40.2025 ;
      RECT  16.45 41.6125 17.1375 41.5475 ;
      RECT  15.7125 41.185 15.8475 41.12 ;
      RECT  15.9275 40.905 16.0625 40.84 ;
      RECT  16.79 40.985 16.855 40.92 ;
      RECT  15.5475 40.2675 17.1375 40.2025 ;
      RECT  15.5475 41.6125 17.1375 41.5475 ;
      RECT  15.855 42.5975 15.92 42.7325 ;
      RECT  15.64 42.5975 15.705 42.7325 ;
      RECT  16.07 42.5975 16.135 42.7325 ;
      RECT  15.855 42.5975 15.92 42.7325 ;
      RECT  15.64 41.7275 15.705 41.8625 ;
      RECT  16.07 41.7275 16.135 41.8625 ;
      RECT  15.7125 41.975 15.8475 42.04 ;
      RECT  15.9275 42.255 16.0625 42.32 ;
      RECT  16.2 42.4675 16.265 42.5325 ;
      RECT  15.5475 42.8925 16.45 42.9575 ;
      RECT  15.5475 41.5475 16.45 41.6125 ;
      RECT  16.7575 42.5975 16.8225 42.7325 ;
      RECT  16.5425 42.5975 16.6075 42.7325 ;
      RECT  16.7575 41.6825 16.8225 41.8175 ;
      RECT  16.5425 41.6825 16.6075 41.8175 ;
      RECT  16.5225 42.175 16.6575 42.24 ;
      RECT  16.79 42.175 16.855 42.24 ;
      RECT  16.45 42.8925 17.1375 42.9575 ;
      RECT  16.45 41.5475 17.1375 41.6125 ;
      RECT  15.7125 41.975 15.8475 42.04 ;
      RECT  15.9275 42.255 16.0625 42.32 ;
      RECT  16.79 42.175 16.855 42.24 ;
      RECT  15.5475 42.8925 17.1375 42.9575 ;
      RECT  15.5475 41.5475 17.1375 41.6125 ;
      RECT  15.855 43.2525 15.92 43.1175 ;
      RECT  15.64 43.2525 15.705 43.1175 ;
      RECT  16.07 43.2525 16.135 43.1175 ;
      RECT  15.855 43.2525 15.92 43.1175 ;
      RECT  15.64 44.1225 15.705 43.9875 ;
      RECT  16.07 44.1225 16.135 43.9875 ;
      RECT  15.7125 43.875 15.8475 43.81 ;
      RECT  15.9275 43.595 16.0625 43.53 ;
      RECT  16.2 43.3825 16.265 43.3175 ;
      RECT  15.5475 42.9575 16.45 42.8925 ;
      RECT  15.5475 44.3025 16.45 44.2375 ;
      RECT  16.7575 43.2525 16.8225 43.1175 ;
      RECT  16.5425 43.2525 16.6075 43.1175 ;
      RECT  16.7575 44.1675 16.8225 44.0325 ;
      RECT  16.5425 44.1675 16.6075 44.0325 ;
      RECT  16.5225 43.675 16.6575 43.61 ;
      RECT  16.79 43.675 16.855 43.61 ;
      RECT  16.45 42.9575 17.1375 42.8925 ;
      RECT  16.45 44.3025 17.1375 44.2375 ;
      RECT  15.7125 43.875 15.8475 43.81 ;
      RECT  15.9275 43.595 16.0625 43.53 ;
      RECT  16.79 43.675 16.855 43.61 ;
      RECT  15.5475 42.9575 17.1375 42.8925 ;
      RECT  15.5475 44.3025 17.1375 44.2375 ;
      RECT  16.79 23.345 16.855 23.41 ;
      RECT  16.79 24.78 16.855 24.845 ;
      RECT  16.79 26.035 16.855 26.1 ;
      RECT  16.79 27.47 16.855 27.535 ;
      RECT  16.79 28.725 16.855 28.79 ;
      RECT  16.79 30.16 16.855 30.225 ;
      RECT  16.79 31.415 16.855 31.48 ;
      RECT  16.79 32.85 16.855 32.915 ;
      RECT  16.79 34.105 16.855 34.17 ;
      RECT  16.79 35.54 16.855 35.605 ;
      RECT  16.79 36.795 16.855 36.86 ;
      RECT  16.79 38.23 16.855 38.295 ;
      RECT  16.79 39.485 16.855 39.55 ;
      RECT  16.79 40.92 16.855 40.985 ;
      RECT  16.79 42.175 16.855 42.24 ;
      RECT  16.79 43.61 16.855 43.675 ;
      RECT  17.4775 23.7675 17.5425 23.9025 ;
      RECT  17.2625 23.7675 17.3275 23.9025 ;
      RECT  17.6925 23.7675 17.7575 23.9025 ;
      RECT  17.4775 23.7675 17.5425 23.9025 ;
      RECT  17.2625 22.8975 17.3275 23.0325 ;
      RECT  17.6925 22.8975 17.7575 23.0325 ;
      RECT  17.335 23.145 17.47 23.21 ;
      RECT  17.55 23.425 17.685 23.49 ;
      RECT  17.8225 23.6375 17.8875 23.7025 ;
      RECT  17.17 24.0625 18.0725 24.1275 ;
      RECT  17.17 22.7175 18.0725 22.7825 ;
      RECT  18.38 23.7675 18.445 23.9025 ;
      RECT  18.165 23.7675 18.23 23.9025 ;
      RECT  18.38 22.8525 18.445 22.9875 ;
      RECT  18.165 22.8525 18.23 22.9875 ;
      RECT  18.145 23.345 18.28 23.41 ;
      RECT  18.4125 23.345 18.4775 23.41 ;
      RECT  18.0725 24.0625 18.76 24.1275 ;
      RECT  18.0725 22.7175 18.76 22.7825 ;
      RECT  17.335 23.145 17.47 23.21 ;
      RECT  17.55 23.425 17.685 23.49 ;
      RECT  18.4125 23.345 18.4775 23.41 ;
      RECT  17.17 24.0625 18.76 24.1275 ;
      RECT  17.17 22.7175 18.76 22.7825 ;
      RECT  17.4775 24.4225 17.5425 24.2875 ;
      RECT  17.2625 24.4225 17.3275 24.2875 ;
      RECT  17.6925 24.4225 17.7575 24.2875 ;
      RECT  17.4775 24.4225 17.5425 24.2875 ;
      RECT  17.2625 25.2925 17.3275 25.1575 ;
      RECT  17.6925 25.2925 17.7575 25.1575 ;
      RECT  17.335 25.045 17.47 24.98 ;
      RECT  17.55 24.765 17.685 24.7 ;
      RECT  17.8225 24.5525 17.8875 24.4875 ;
      RECT  17.17 24.1275 18.0725 24.0625 ;
      RECT  17.17 25.4725 18.0725 25.4075 ;
      RECT  18.38 24.4225 18.445 24.2875 ;
      RECT  18.165 24.4225 18.23 24.2875 ;
      RECT  18.38 25.3375 18.445 25.2025 ;
      RECT  18.165 25.3375 18.23 25.2025 ;
      RECT  18.145 24.845 18.28 24.78 ;
      RECT  18.4125 24.845 18.4775 24.78 ;
      RECT  18.0725 24.1275 18.76 24.0625 ;
      RECT  18.0725 25.4725 18.76 25.4075 ;
      RECT  17.335 25.045 17.47 24.98 ;
      RECT  17.55 24.765 17.685 24.7 ;
      RECT  18.4125 24.845 18.4775 24.78 ;
      RECT  17.17 24.1275 18.76 24.0625 ;
      RECT  17.17 25.4725 18.76 25.4075 ;
      RECT  17.4775 26.4575 17.5425 26.5925 ;
      RECT  17.2625 26.4575 17.3275 26.5925 ;
      RECT  17.6925 26.4575 17.7575 26.5925 ;
      RECT  17.4775 26.4575 17.5425 26.5925 ;
      RECT  17.2625 25.5875 17.3275 25.7225 ;
      RECT  17.6925 25.5875 17.7575 25.7225 ;
      RECT  17.335 25.835 17.47 25.9 ;
      RECT  17.55 26.115 17.685 26.18 ;
      RECT  17.8225 26.3275 17.8875 26.3925 ;
      RECT  17.17 26.7525 18.0725 26.8175 ;
      RECT  17.17 25.4075 18.0725 25.4725 ;
      RECT  18.38 26.4575 18.445 26.5925 ;
      RECT  18.165 26.4575 18.23 26.5925 ;
      RECT  18.38 25.5425 18.445 25.6775 ;
      RECT  18.165 25.5425 18.23 25.6775 ;
      RECT  18.145 26.035 18.28 26.1 ;
      RECT  18.4125 26.035 18.4775 26.1 ;
      RECT  18.0725 26.7525 18.76 26.8175 ;
      RECT  18.0725 25.4075 18.76 25.4725 ;
      RECT  17.335 25.835 17.47 25.9 ;
      RECT  17.55 26.115 17.685 26.18 ;
      RECT  18.4125 26.035 18.4775 26.1 ;
      RECT  17.17 26.7525 18.76 26.8175 ;
      RECT  17.17 25.4075 18.76 25.4725 ;
      RECT  17.4775 27.1125 17.5425 26.9775 ;
      RECT  17.2625 27.1125 17.3275 26.9775 ;
      RECT  17.6925 27.1125 17.7575 26.9775 ;
      RECT  17.4775 27.1125 17.5425 26.9775 ;
      RECT  17.2625 27.9825 17.3275 27.8475 ;
      RECT  17.6925 27.9825 17.7575 27.8475 ;
      RECT  17.335 27.735 17.47 27.67 ;
      RECT  17.55 27.455 17.685 27.39 ;
      RECT  17.8225 27.2425 17.8875 27.1775 ;
      RECT  17.17 26.8175 18.0725 26.7525 ;
      RECT  17.17 28.1625 18.0725 28.0975 ;
      RECT  18.38 27.1125 18.445 26.9775 ;
      RECT  18.165 27.1125 18.23 26.9775 ;
      RECT  18.38 28.0275 18.445 27.8925 ;
      RECT  18.165 28.0275 18.23 27.8925 ;
      RECT  18.145 27.535 18.28 27.47 ;
      RECT  18.4125 27.535 18.4775 27.47 ;
      RECT  18.0725 26.8175 18.76 26.7525 ;
      RECT  18.0725 28.1625 18.76 28.0975 ;
      RECT  17.335 27.735 17.47 27.67 ;
      RECT  17.55 27.455 17.685 27.39 ;
      RECT  18.4125 27.535 18.4775 27.47 ;
      RECT  17.17 26.8175 18.76 26.7525 ;
      RECT  17.17 28.1625 18.76 28.0975 ;
      RECT  17.4775 29.1475 17.5425 29.2825 ;
      RECT  17.2625 29.1475 17.3275 29.2825 ;
      RECT  17.6925 29.1475 17.7575 29.2825 ;
      RECT  17.4775 29.1475 17.5425 29.2825 ;
      RECT  17.2625 28.2775 17.3275 28.4125 ;
      RECT  17.6925 28.2775 17.7575 28.4125 ;
      RECT  17.335 28.525 17.47 28.59 ;
      RECT  17.55 28.805 17.685 28.87 ;
      RECT  17.8225 29.0175 17.8875 29.0825 ;
      RECT  17.17 29.4425 18.0725 29.5075 ;
      RECT  17.17 28.0975 18.0725 28.1625 ;
      RECT  18.38 29.1475 18.445 29.2825 ;
      RECT  18.165 29.1475 18.23 29.2825 ;
      RECT  18.38 28.2325 18.445 28.3675 ;
      RECT  18.165 28.2325 18.23 28.3675 ;
      RECT  18.145 28.725 18.28 28.79 ;
      RECT  18.4125 28.725 18.4775 28.79 ;
      RECT  18.0725 29.4425 18.76 29.5075 ;
      RECT  18.0725 28.0975 18.76 28.1625 ;
      RECT  17.335 28.525 17.47 28.59 ;
      RECT  17.55 28.805 17.685 28.87 ;
      RECT  18.4125 28.725 18.4775 28.79 ;
      RECT  17.17 29.4425 18.76 29.5075 ;
      RECT  17.17 28.0975 18.76 28.1625 ;
      RECT  17.4775 29.8025 17.5425 29.6675 ;
      RECT  17.2625 29.8025 17.3275 29.6675 ;
      RECT  17.6925 29.8025 17.7575 29.6675 ;
      RECT  17.4775 29.8025 17.5425 29.6675 ;
      RECT  17.2625 30.6725 17.3275 30.5375 ;
      RECT  17.6925 30.6725 17.7575 30.5375 ;
      RECT  17.335 30.425 17.47 30.36 ;
      RECT  17.55 30.145 17.685 30.08 ;
      RECT  17.8225 29.9325 17.8875 29.8675 ;
      RECT  17.17 29.5075 18.0725 29.4425 ;
      RECT  17.17 30.8525 18.0725 30.7875 ;
      RECT  18.38 29.8025 18.445 29.6675 ;
      RECT  18.165 29.8025 18.23 29.6675 ;
      RECT  18.38 30.7175 18.445 30.5825 ;
      RECT  18.165 30.7175 18.23 30.5825 ;
      RECT  18.145 30.225 18.28 30.16 ;
      RECT  18.4125 30.225 18.4775 30.16 ;
      RECT  18.0725 29.5075 18.76 29.4425 ;
      RECT  18.0725 30.8525 18.76 30.7875 ;
      RECT  17.335 30.425 17.47 30.36 ;
      RECT  17.55 30.145 17.685 30.08 ;
      RECT  18.4125 30.225 18.4775 30.16 ;
      RECT  17.17 29.5075 18.76 29.4425 ;
      RECT  17.17 30.8525 18.76 30.7875 ;
      RECT  17.4775 31.8375 17.5425 31.9725 ;
      RECT  17.2625 31.8375 17.3275 31.9725 ;
      RECT  17.6925 31.8375 17.7575 31.9725 ;
      RECT  17.4775 31.8375 17.5425 31.9725 ;
      RECT  17.2625 30.9675 17.3275 31.1025 ;
      RECT  17.6925 30.9675 17.7575 31.1025 ;
      RECT  17.335 31.215 17.47 31.28 ;
      RECT  17.55 31.495 17.685 31.56 ;
      RECT  17.8225 31.7075 17.8875 31.7725 ;
      RECT  17.17 32.1325 18.0725 32.1975 ;
      RECT  17.17 30.7875 18.0725 30.8525 ;
      RECT  18.38 31.8375 18.445 31.9725 ;
      RECT  18.165 31.8375 18.23 31.9725 ;
      RECT  18.38 30.9225 18.445 31.0575 ;
      RECT  18.165 30.9225 18.23 31.0575 ;
      RECT  18.145 31.415 18.28 31.48 ;
      RECT  18.4125 31.415 18.4775 31.48 ;
      RECT  18.0725 32.1325 18.76 32.1975 ;
      RECT  18.0725 30.7875 18.76 30.8525 ;
      RECT  17.335 31.215 17.47 31.28 ;
      RECT  17.55 31.495 17.685 31.56 ;
      RECT  18.4125 31.415 18.4775 31.48 ;
      RECT  17.17 32.1325 18.76 32.1975 ;
      RECT  17.17 30.7875 18.76 30.8525 ;
      RECT  17.4775 32.4925 17.5425 32.3575 ;
      RECT  17.2625 32.4925 17.3275 32.3575 ;
      RECT  17.6925 32.4925 17.7575 32.3575 ;
      RECT  17.4775 32.4925 17.5425 32.3575 ;
      RECT  17.2625 33.3625 17.3275 33.2275 ;
      RECT  17.6925 33.3625 17.7575 33.2275 ;
      RECT  17.335 33.115 17.47 33.05 ;
      RECT  17.55 32.835 17.685 32.77 ;
      RECT  17.8225 32.6225 17.8875 32.5575 ;
      RECT  17.17 32.1975 18.0725 32.1325 ;
      RECT  17.17 33.5425 18.0725 33.4775 ;
      RECT  18.38 32.4925 18.445 32.3575 ;
      RECT  18.165 32.4925 18.23 32.3575 ;
      RECT  18.38 33.4075 18.445 33.2725 ;
      RECT  18.165 33.4075 18.23 33.2725 ;
      RECT  18.145 32.915 18.28 32.85 ;
      RECT  18.4125 32.915 18.4775 32.85 ;
      RECT  18.0725 32.1975 18.76 32.1325 ;
      RECT  18.0725 33.5425 18.76 33.4775 ;
      RECT  17.335 33.115 17.47 33.05 ;
      RECT  17.55 32.835 17.685 32.77 ;
      RECT  18.4125 32.915 18.4775 32.85 ;
      RECT  17.17 32.1975 18.76 32.1325 ;
      RECT  17.17 33.5425 18.76 33.4775 ;
      RECT  17.4775 34.5275 17.5425 34.6625 ;
      RECT  17.2625 34.5275 17.3275 34.6625 ;
      RECT  17.6925 34.5275 17.7575 34.6625 ;
      RECT  17.4775 34.5275 17.5425 34.6625 ;
      RECT  17.2625 33.6575 17.3275 33.7925 ;
      RECT  17.6925 33.6575 17.7575 33.7925 ;
      RECT  17.335 33.905 17.47 33.97 ;
      RECT  17.55 34.185 17.685 34.25 ;
      RECT  17.8225 34.3975 17.8875 34.4625 ;
      RECT  17.17 34.8225 18.0725 34.8875 ;
      RECT  17.17 33.4775 18.0725 33.5425 ;
      RECT  18.38 34.5275 18.445 34.6625 ;
      RECT  18.165 34.5275 18.23 34.6625 ;
      RECT  18.38 33.6125 18.445 33.7475 ;
      RECT  18.165 33.6125 18.23 33.7475 ;
      RECT  18.145 34.105 18.28 34.17 ;
      RECT  18.4125 34.105 18.4775 34.17 ;
      RECT  18.0725 34.8225 18.76 34.8875 ;
      RECT  18.0725 33.4775 18.76 33.5425 ;
      RECT  17.335 33.905 17.47 33.97 ;
      RECT  17.55 34.185 17.685 34.25 ;
      RECT  18.4125 34.105 18.4775 34.17 ;
      RECT  17.17 34.8225 18.76 34.8875 ;
      RECT  17.17 33.4775 18.76 33.5425 ;
      RECT  17.4775 35.1825 17.5425 35.0475 ;
      RECT  17.2625 35.1825 17.3275 35.0475 ;
      RECT  17.6925 35.1825 17.7575 35.0475 ;
      RECT  17.4775 35.1825 17.5425 35.0475 ;
      RECT  17.2625 36.0525 17.3275 35.9175 ;
      RECT  17.6925 36.0525 17.7575 35.9175 ;
      RECT  17.335 35.805 17.47 35.74 ;
      RECT  17.55 35.525 17.685 35.46 ;
      RECT  17.8225 35.3125 17.8875 35.2475 ;
      RECT  17.17 34.8875 18.0725 34.8225 ;
      RECT  17.17 36.2325 18.0725 36.1675 ;
      RECT  18.38 35.1825 18.445 35.0475 ;
      RECT  18.165 35.1825 18.23 35.0475 ;
      RECT  18.38 36.0975 18.445 35.9625 ;
      RECT  18.165 36.0975 18.23 35.9625 ;
      RECT  18.145 35.605 18.28 35.54 ;
      RECT  18.4125 35.605 18.4775 35.54 ;
      RECT  18.0725 34.8875 18.76 34.8225 ;
      RECT  18.0725 36.2325 18.76 36.1675 ;
      RECT  17.335 35.805 17.47 35.74 ;
      RECT  17.55 35.525 17.685 35.46 ;
      RECT  18.4125 35.605 18.4775 35.54 ;
      RECT  17.17 34.8875 18.76 34.8225 ;
      RECT  17.17 36.2325 18.76 36.1675 ;
      RECT  17.4775 37.2175 17.5425 37.3525 ;
      RECT  17.2625 37.2175 17.3275 37.3525 ;
      RECT  17.6925 37.2175 17.7575 37.3525 ;
      RECT  17.4775 37.2175 17.5425 37.3525 ;
      RECT  17.2625 36.3475 17.3275 36.4825 ;
      RECT  17.6925 36.3475 17.7575 36.4825 ;
      RECT  17.335 36.595 17.47 36.66 ;
      RECT  17.55 36.875 17.685 36.94 ;
      RECT  17.8225 37.0875 17.8875 37.1525 ;
      RECT  17.17 37.5125 18.0725 37.5775 ;
      RECT  17.17 36.1675 18.0725 36.2325 ;
      RECT  18.38 37.2175 18.445 37.3525 ;
      RECT  18.165 37.2175 18.23 37.3525 ;
      RECT  18.38 36.3025 18.445 36.4375 ;
      RECT  18.165 36.3025 18.23 36.4375 ;
      RECT  18.145 36.795 18.28 36.86 ;
      RECT  18.4125 36.795 18.4775 36.86 ;
      RECT  18.0725 37.5125 18.76 37.5775 ;
      RECT  18.0725 36.1675 18.76 36.2325 ;
      RECT  17.335 36.595 17.47 36.66 ;
      RECT  17.55 36.875 17.685 36.94 ;
      RECT  18.4125 36.795 18.4775 36.86 ;
      RECT  17.17 37.5125 18.76 37.5775 ;
      RECT  17.17 36.1675 18.76 36.2325 ;
      RECT  17.4775 37.8725 17.5425 37.7375 ;
      RECT  17.2625 37.8725 17.3275 37.7375 ;
      RECT  17.6925 37.8725 17.7575 37.7375 ;
      RECT  17.4775 37.8725 17.5425 37.7375 ;
      RECT  17.2625 38.7425 17.3275 38.6075 ;
      RECT  17.6925 38.7425 17.7575 38.6075 ;
      RECT  17.335 38.495 17.47 38.43 ;
      RECT  17.55 38.215 17.685 38.15 ;
      RECT  17.8225 38.0025 17.8875 37.9375 ;
      RECT  17.17 37.5775 18.0725 37.5125 ;
      RECT  17.17 38.9225 18.0725 38.8575 ;
      RECT  18.38 37.8725 18.445 37.7375 ;
      RECT  18.165 37.8725 18.23 37.7375 ;
      RECT  18.38 38.7875 18.445 38.6525 ;
      RECT  18.165 38.7875 18.23 38.6525 ;
      RECT  18.145 38.295 18.28 38.23 ;
      RECT  18.4125 38.295 18.4775 38.23 ;
      RECT  18.0725 37.5775 18.76 37.5125 ;
      RECT  18.0725 38.9225 18.76 38.8575 ;
      RECT  17.335 38.495 17.47 38.43 ;
      RECT  17.55 38.215 17.685 38.15 ;
      RECT  18.4125 38.295 18.4775 38.23 ;
      RECT  17.17 37.5775 18.76 37.5125 ;
      RECT  17.17 38.9225 18.76 38.8575 ;
      RECT  17.4775 39.9075 17.5425 40.0425 ;
      RECT  17.2625 39.9075 17.3275 40.0425 ;
      RECT  17.6925 39.9075 17.7575 40.0425 ;
      RECT  17.4775 39.9075 17.5425 40.0425 ;
      RECT  17.2625 39.0375 17.3275 39.1725 ;
      RECT  17.6925 39.0375 17.7575 39.1725 ;
      RECT  17.335 39.285 17.47 39.35 ;
      RECT  17.55 39.565 17.685 39.63 ;
      RECT  17.8225 39.7775 17.8875 39.8425 ;
      RECT  17.17 40.2025 18.0725 40.2675 ;
      RECT  17.17 38.8575 18.0725 38.9225 ;
      RECT  18.38 39.9075 18.445 40.0425 ;
      RECT  18.165 39.9075 18.23 40.0425 ;
      RECT  18.38 38.9925 18.445 39.1275 ;
      RECT  18.165 38.9925 18.23 39.1275 ;
      RECT  18.145 39.485 18.28 39.55 ;
      RECT  18.4125 39.485 18.4775 39.55 ;
      RECT  18.0725 40.2025 18.76 40.2675 ;
      RECT  18.0725 38.8575 18.76 38.9225 ;
      RECT  17.335 39.285 17.47 39.35 ;
      RECT  17.55 39.565 17.685 39.63 ;
      RECT  18.4125 39.485 18.4775 39.55 ;
      RECT  17.17 40.2025 18.76 40.2675 ;
      RECT  17.17 38.8575 18.76 38.9225 ;
      RECT  17.4775 40.5625 17.5425 40.4275 ;
      RECT  17.2625 40.5625 17.3275 40.4275 ;
      RECT  17.6925 40.5625 17.7575 40.4275 ;
      RECT  17.4775 40.5625 17.5425 40.4275 ;
      RECT  17.2625 41.4325 17.3275 41.2975 ;
      RECT  17.6925 41.4325 17.7575 41.2975 ;
      RECT  17.335 41.185 17.47 41.12 ;
      RECT  17.55 40.905 17.685 40.84 ;
      RECT  17.8225 40.6925 17.8875 40.6275 ;
      RECT  17.17 40.2675 18.0725 40.2025 ;
      RECT  17.17 41.6125 18.0725 41.5475 ;
      RECT  18.38 40.5625 18.445 40.4275 ;
      RECT  18.165 40.5625 18.23 40.4275 ;
      RECT  18.38 41.4775 18.445 41.3425 ;
      RECT  18.165 41.4775 18.23 41.3425 ;
      RECT  18.145 40.985 18.28 40.92 ;
      RECT  18.4125 40.985 18.4775 40.92 ;
      RECT  18.0725 40.2675 18.76 40.2025 ;
      RECT  18.0725 41.6125 18.76 41.5475 ;
      RECT  17.335 41.185 17.47 41.12 ;
      RECT  17.55 40.905 17.685 40.84 ;
      RECT  18.4125 40.985 18.4775 40.92 ;
      RECT  17.17 40.2675 18.76 40.2025 ;
      RECT  17.17 41.6125 18.76 41.5475 ;
      RECT  17.4775 42.5975 17.5425 42.7325 ;
      RECT  17.2625 42.5975 17.3275 42.7325 ;
      RECT  17.6925 42.5975 17.7575 42.7325 ;
      RECT  17.4775 42.5975 17.5425 42.7325 ;
      RECT  17.2625 41.7275 17.3275 41.8625 ;
      RECT  17.6925 41.7275 17.7575 41.8625 ;
      RECT  17.335 41.975 17.47 42.04 ;
      RECT  17.55 42.255 17.685 42.32 ;
      RECT  17.8225 42.4675 17.8875 42.5325 ;
      RECT  17.17 42.8925 18.0725 42.9575 ;
      RECT  17.17 41.5475 18.0725 41.6125 ;
      RECT  18.38 42.5975 18.445 42.7325 ;
      RECT  18.165 42.5975 18.23 42.7325 ;
      RECT  18.38 41.6825 18.445 41.8175 ;
      RECT  18.165 41.6825 18.23 41.8175 ;
      RECT  18.145 42.175 18.28 42.24 ;
      RECT  18.4125 42.175 18.4775 42.24 ;
      RECT  18.0725 42.8925 18.76 42.9575 ;
      RECT  18.0725 41.5475 18.76 41.6125 ;
      RECT  17.335 41.975 17.47 42.04 ;
      RECT  17.55 42.255 17.685 42.32 ;
      RECT  18.4125 42.175 18.4775 42.24 ;
      RECT  17.17 42.8925 18.76 42.9575 ;
      RECT  17.17 41.5475 18.76 41.6125 ;
      RECT  17.4775 43.2525 17.5425 43.1175 ;
      RECT  17.2625 43.2525 17.3275 43.1175 ;
      RECT  17.6925 43.2525 17.7575 43.1175 ;
      RECT  17.4775 43.2525 17.5425 43.1175 ;
      RECT  17.2625 44.1225 17.3275 43.9875 ;
      RECT  17.6925 44.1225 17.7575 43.9875 ;
      RECT  17.335 43.875 17.47 43.81 ;
      RECT  17.55 43.595 17.685 43.53 ;
      RECT  17.8225 43.3825 17.8875 43.3175 ;
      RECT  17.17 42.9575 18.0725 42.8925 ;
      RECT  17.17 44.3025 18.0725 44.2375 ;
      RECT  18.38 43.2525 18.445 43.1175 ;
      RECT  18.165 43.2525 18.23 43.1175 ;
      RECT  18.38 44.1675 18.445 44.0325 ;
      RECT  18.165 44.1675 18.23 44.0325 ;
      RECT  18.145 43.675 18.28 43.61 ;
      RECT  18.4125 43.675 18.4775 43.61 ;
      RECT  18.0725 42.9575 18.76 42.8925 ;
      RECT  18.0725 44.3025 18.76 44.2375 ;
      RECT  17.335 43.875 17.47 43.81 ;
      RECT  17.55 43.595 17.685 43.53 ;
      RECT  18.4125 43.675 18.4775 43.61 ;
      RECT  17.17 42.9575 18.76 42.8925 ;
      RECT  17.17 44.3025 18.76 44.2375 ;
      RECT  17.335 23.145 17.47 23.21 ;
      RECT  17.335 24.98 17.47 25.045 ;
      RECT  17.335 25.835 17.47 25.9 ;
      RECT  17.335 27.67 17.47 27.735 ;
      RECT  17.335 28.525 17.47 28.59 ;
      RECT  17.335 30.36 17.47 30.425 ;
      RECT  17.335 31.215 17.47 31.28 ;
      RECT  17.335 33.05 17.47 33.115 ;
      RECT  17.335 33.905 17.47 33.97 ;
      RECT  17.335 35.74 17.47 35.805 ;
      RECT  17.335 36.595 17.47 36.66 ;
      RECT  17.335 38.43 17.47 38.495 ;
      RECT  17.335 39.285 17.47 39.35 ;
      RECT  17.335 41.12 17.47 41.185 ;
      RECT  17.335 41.975 17.47 42.04 ;
      RECT  17.335 43.81 17.47 43.875 ;
      RECT  18.4125 23.345 18.4775 23.41 ;
      RECT  18.4125 24.78 18.4775 24.845 ;
      RECT  18.4125 26.035 18.4775 26.1 ;
      RECT  18.4125 27.47 18.4775 27.535 ;
      RECT  18.4125 28.725 18.4775 28.79 ;
      RECT  18.4125 30.16 18.4775 30.225 ;
      RECT  18.4125 31.415 18.4775 31.48 ;
      RECT  18.4125 32.85 18.4775 32.915 ;
      RECT  18.4125 34.105 18.4775 34.17 ;
      RECT  18.4125 35.54 18.4775 35.605 ;
      RECT  18.4125 36.795 18.4775 36.86 ;
      RECT  18.4125 38.23 18.4775 38.295 ;
      RECT  18.4125 39.485 18.4775 39.55 ;
      RECT  18.4125 40.92 18.4775 40.985 ;
      RECT  18.4125 42.175 18.4775 42.24 ;
      RECT  18.4125 43.61 18.4775 43.675 ;
      RECT  18.29 21.7325 18.355 21.5975 ;
      RECT  18.075 21.7325 18.14 21.5975 ;
      RECT  18.29 22.6475 18.355 22.5125 ;
      RECT  18.075 22.6475 18.14 22.5125 ;
      RECT  18.055 22.155 18.19 22.09 ;
      RECT  18.3225 22.155 18.3875 22.09 ;
      RECT  17.9825 21.4375 18.67 21.3725 ;
      RECT  17.9825 22.7825 18.67 22.7175 ;
      RECT  18.9775 21.7325 19.0425 21.5975 ;
      RECT  18.7625 21.7325 18.8275 21.5975 ;
      RECT  18.9775 22.6475 19.0425 22.5125 ;
      RECT  18.7625 22.6475 18.8275 22.5125 ;
      RECT  18.7425 22.155 18.8775 22.09 ;
      RECT  19.01 22.155 19.075 22.09 ;
      RECT  18.67 21.4375 19.135 21.3725 ;
      RECT  18.67 22.7825 19.135 22.7175 ;
      RECT  18.055 22.155 18.19 22.09 ;
      RECT  19.01 22.155 19.075 22.09 ;
      RECT  17.9825 21.4375 19.135 21.3725 ;
      RECT  17.9825 22.7825 19.135 22.7175 ;
      RECT  18.4125 23.345 18.4775 23.41 ;
      RECT  18.4125 24.78 18.4775 24.845 ;
      RECT  18.4125 26.035 18.4775 26.1 ;
      RECT  18.4125 27.47 18.4775 27.535 ;
      RECT  18.4125 28.725 18.4775 28.79 ;
      RECT  18.4125 30.16 18.4775 30.225 ;
      RECT  18.4125 31.415 18.4775 31.48 ;
      RECT  18.4125 32.85 18.4775 32.915 ;
      RECT  18.4125 34.105 18.4775 34.17 ;
      RECT  18.4125 35.54 18.4775 35.605 ;
      RECT  18.4125 36.795 18.4775 36.86 ;
      RECT  18.4125 38.23 18.4775 38.295 ;
      RECT  18.4125 39.485 18.4775 39.55 ;
      RECT  18.4125 40.92 18.4775 40.985 ;
      RECT  18.4125 42.175 18.4775 42.24 ;
      RECT  18.4125 43.61 18.4775 43.675 ;
      RECT  19.01 22.09 19.075 22.155 ;
      RECT  0.0 -0.065 2.86 0.065 ;
      POLYGON  1.8475 1.4425 1.8475 2.2675 2.3925 2.2675 2.3925 2.2025 1.9125 2.2025 1.9125 1.8575 2.1075 1.8575 2.1075 1.4425 1.8475 1.4425 ;
      RECT  2.6325 1.0475 2.71 1.1825 ;
      POLYGON  0.4175 0.335 0.4175 0.975 0.7175 0.975 0.7175 1.8625 0.6475 1.8625 0.6475 1.9275 0.7825 1.9275 0.7825 1.7975 1.3725 1.7975 1.3725 2.1475 1.4375 2.1475 1.4375 1.6575 1.7175 1.6575 1.7175 2.0725 1.7825 2.0725 1.7825 1.5925 1.3725 1.5925 1.3725 1.7325 0.7825 1.7325 0.7825 0.91 0.4825 0.91 0.4825 0.4 1.3725 0.4 1.3725 0.7925 1.4375 0.7925 1.4375 0.335 0.4175 0.335 ;
      RECT  2.0475 0.5875 2.1125 0.8625 ;
      POLYGON  0.5175 1.3825 0.5175 2.0575 1.1625 2.0575 1.1625 1.9225 1.0975 1.9225 1.0975 1.9925 0.5825 1.9925 0.5825 1.7975 0.6075 1.7975 0.6075 1.3825 0.5175 1.3825 ;
      POLYGON  2.6425 0.2175 2.6425 0.9175 2.5375 0.9175 2.5375 0.9825 2.6425 0.9825 2.6425 1.6475 2.3125 1.6475 2.3125 1.7125 2.6425 1.7125 2.6425 2.2375 2.7075 2.2375 2.7075 0.2175 2.6425 0.2175 ;
      POLYGON  1.7775 0.9275 1.7775 1.1425 1.5475 1.1425 1.5475 1.015 1.4125 1.015 1.4125 1.4625 1.1725 1.4625 1.1725 1.6675 1.3075 1.6675 1.3075 1.5275 1.4775 1.5275 1.4775 1.2075 1.9725 1.2075 1.9725 0.9925 2.1875 0.9925 2.1875 1.1925 2.3225 1.1925 2.3225 1.1275 2.2525 1.1275 2.2525 0.9275 1.7775 0.9275 ;
      POLYGON  0.1675 1.2675 0.1675 2.405 0.1 2.405 0.1 2.535 2.86 2.535 2.86 2.405 2.5225 2.405 2.5225 1.9075 2.4575 1.9075 2.4575 2.405 1.6225 2.405 1.6225 1.7225 1.5575 1.7225 1.5575 2.405 1.0575 2.405 1.0575 2.2525 0.9225 2.2525 0.9225 2.405 0.2325 2.405 0.2325 1.2675 0.1675 1.2675 ;
      RECT  2.6425 0.915 2.7075 1.1275 ;
      POLYGON  2.1075 0.2275 2.1075 0.5025 2.2375 0.5025 2.2375 0.7625 2.3025 0.7625 2.3025 0.4375 2.1725 0.4375 2.1725 0.2275 2.1075 0.2275 ;
      RECT  0.245 1.0375 0.3225 1.1725 ;
      RECT  1.7775 0.9275 1.9725 1.2075 ;
      POLYGON  0.3875 1.1175 0.3875 2.1875 1.2925 2.1875 1.2925 1.8625 1.2275 1.8625 1.2275 2.1225 0.4525 2.1225 0.4525 1.1825 0.5375 1.1825 0.5375 1.1175 0.3875 1.1175 ;
      POLYGON  0.1 -0.065 0.1 0.065 0.1675 0.065 0.1675 0.845 0.2325 0.845 0.2325 0.065 0.9175 0.065 0.9175 0.235 1.0525 0.235 1.0525 0.065 1.5575 0.065 1.5575 0.7925 1.6225 0.7925 1.6225 0.065 1.9225 0.065 1.9225 0.4675 1.9875 0.4675 1.9875 0.065 2.4075 0.065 2.4075 0.9875 2.4725 0.9875 2.4725 0.065 2.76 0.065 2.76 -0.065 0.1 -0.065 ;
      POLYGON  1.2175 0.685 1.2175 0.95 0.9425 0.95 0.9425 1.015 1.2175 1.015 1.2175 1.3975 1.2825 1.3975 1.2825 0.95 1.6125 0.95 1.6125 1.0775 1.6775 1.0775 1.6775 0.885 1.2825 0.885 1.2825 0.685 1.2175 0.685 ;
      POLYGON  2.0525 1.0575 2.0525 1.3225 2.5025 1.3225 2.5025 1.5175 2.3025 1.5175 2.3025 1.5825 2.5675 1.5825 2.5675 1.0575 2.4025 1.0575 2.4025 1.1925 2.5025 1.1925 2.5025 1.2575 2.1175 1.2575 2.1175 1.0575 2.0525 1.0575 ;
      RECT  2.3275 1.7775 2.3925 2.1275 ;
      RECT  0.0 2.405 2.76 2.535 ;
      POLYGON  0.5475 0.465 0.5475 0.845 0.6125 0.845 0.6125 0.53 1.2125 0.53 1.2125 0.465 0.5475 0.465 ;
      POLYGON  2.1725 1.3875 2.1725 2.1375 2.2625 2.1375 2.2625 1.8625 2.2375 1.8625 2.2375 1.4525 2.4375 1.4525 2.4375 1.3875 2.1725 1.3875 ;
      RECT  3.4475 2.0125 3.5125 2.1475 ;
      RECT  3.2325 2.0125 3.2975 2.1475 ;
      RECT  3.4475 0.1475 3.5125 0.2825 ;
      RECT  3.2325 0.1475 3.2975 0.2825 ;
      RECT  3.2125 1.115 3.3475 1.18 ;
      RECT  3.48 1.115 3.545 1.18 ;
      RECT  3.14 2.4425 3.8275 2.5075 ;
      RECT  3.14 -0.0325 3.8275 0.0325 ;
      RECT  4.165 2.0125 4.23 2.1475 ;
      RECT  3.92 2.0125 3.985 2.1475 ;
      RECT  4.41 2.0125 4.475 2.1475 ;
      RECT  4.165 0.1475 4.23 0.2825 ;
      RECT  3.92 0.1475 3.985 0.2825 ;
      RECT  4.41 0.1475 4.475 0.2825 ;
      RECT  3.9 1.115 4.035 1.18 ;
      RECT  4.1975 1.115 4.2625 1.18 ;
      RECT  3.8275 2.4425 4.79 2.5075 ;
      RECT  3.8275 -0.0325 4.79 0.0325 ;
      RECT  0.0 2.405 4.79 2.535 ;
      RECT  0.0 -0.065 4.79 0.065 ;
      RECT  0.0 5.015 2.86 4.885 ;
      POLYGON  1.8475 3.5075 1.8475 2.6825 2.3925 2.6825 2.3925 2.7475 1.9125 2.7475 1.9125 3.0925 2.1075 3.0925 2.1075 3.5075 1.8475 3.5075 ;
      RECT  2.6325 3.9025 2.71 3.7675 ;
      POLYGON  0.4175 4.615 0.4175 3.975 0.7175 3.975 0.7175 3.0875 0.6475 3.0875 0.6475 3.0225 0.7825 3.0225 0.7825 3.1525 1.3725 3.1525 1.3725 2.8025 1.4375 2.8025 1.4375 3.2925 1.7175 3.2925 1.7175 2.8775 1.7825 2.8775 1.7825 3.3575 1.3725 3.3575 1.3725 3.2175 0.7825 3.2175 0.7825 4.04 0.4825 4.04 0.4825 4.55 1.3725 4.55 1.3725 4.1575 1.4375 4.1575 1.4375 4.615 0.4175 4.615 ;
      RECT  2.0475 4.3625 2.1125 4.0875 ;
      POLYGON  0.5175 3.5675 0.5175 2.8925 1.1625 2.8925 1.1625 3.0275 1.0975 3.0275 1.0975 2.9575 0.5825 2.9575 0.5825 3.1525 0.6075 3.1525 0.6075 3.5675 0.5175 3.5675 ;
      POLYGON  2.6425 4.7325 2.6425 4.0325 2.5375 4.0325 2.5375 3.9675 2.6425 3.9675 2.6425 3.3025 2.3125 3.3025 2.3125 3.2375 2.6425 3.2375 2.6425 2.7125 2.7075 2.7125 2.7075 4.7325 2.6425 4.7325 ;
      POLYGON  1.7775 4.0225 1.7775 3.8075 1.5475 3.8075 1.5475 3.935 1.4125 3.935 1.4125 3.4875 1.1725 3.4875 1.1725 3.2825 1.3075 3.2825 1.3075 3.4225 1.4775 3.4225 1.4775 3.7425 1.9725 3.7425 1.9725 3.9575 2.1875 3.9575 2.1875 3.7575 2.3225 3.7575 2.3225 3.8225 2.2525 3.8225 2.2525 4.0225 1.7775 4.0225 ;
      POLYGON  0.1675 3.6825 0.1675 2.545 0.1 2.545 0.1 2.415 2.86 2.415 2.86 2.545 2.5225 2.545 2.5225 3.0425 2.4575 3.0425 2.4575 2.545 1.6225 2.545 1.6225 3.2275 1.5575 3.2275 1.5575 2.545 1.0575 2.545 1.0575 2.6975 0.9225 2.6975 0.9225 2.545 0.2325 2.545 0.2325 3.6825 0.1675 3.6825 ;
      RECT  2.6425 4.035 2.7075 3.8225 ;
      POLYGON  2.1075 4.7225 2.1075 4.4475 2.2375 4.4475 2.2375 4.1875 2.3025 4.1875 2.3025 4.5125 2.1725 4.5125 2.1725 4.7225 2.1075 4.7225 ;
      RECT  0.245 3.9125 0.3225 3.7775 ;
      RECT  1.7775 4.0225 1.9725 3.7425 ;
      POLYGON  0.3875 3.8325 0.3875 2.7625 1.2925 2.7625 1.2925 3.0875 1.2275 3.0875 1.2275 2.8275 0.4525 2.8275 0.4525 3.7675 0.5375 3.7675 0.5375 3.8325 0.3875 3.8325 ;
      POLYGON  0.1 5.015 0.1 4.885 0.1675 4.885 0.1675 4.105 0.2325 4.105 0.2325 4.885 0.9175 4.885 0.9175 4.715 1.0525 4.715 1.0525 4.885 1.5575 4.885 1.5575 4.1575 1.6225 4.1575 1.6225 4.885 1.9225 4.885 1.9225 4.4825 1.9875 4.4825 1.9875 4.885 2.4075 4.885 2.4075 3.9625 2.4725 3.9625 2.4725 4.885 2.76 4.885 2.76 5.015 0.1 5.015 ;
      POLYGON  1.2175 4.265 1.2175 4.0 0.9425 4.0 0.9425 3.935 1.2175 3.935 1.2175 3.5525 1.2825 3.5525 1.2825 4.0 1.6125 4.0 1.6125 3.8725 1.6775 3.8725 1.6775 4.065 1.2825 4.065 1.2825 4.265 1.2175 4.265 ;
      POLYGON  2.0525 3.8925 2.0525 3.6275 2.5025 3.6275 2.5025 3.4325 2.3025 3.4325 2.3025 3.3675 2.5675 3.3675 2.5675 3.8925 2.4025 3.8925 2.4025 3.7575 2.5025 3.7575 2.5025 3.6925 2.1175 3.6925 2.1175 3.8925 2.0525 3.8925 ;
      RECT  2.3275 3.1725 2.3925 2.8225 ;
      RECT  0.0 2.545 2.76 2.415 ;
      POLYGON  0.5475 4.485 0.5475 4.105 0.6125 4.105 0.6125 4.42 1.2125 4.42 1.2125 4.485 0.5475 4.485 ;
      POLYGON  2.1725 3.5625 2.1725 2.8125 2.2625 2.8125 2.2625 3.0875 2.2375 3.0875 2.2375 3.4975 2.4375 3.4975 2.4375 3.5625 2.1725 3.5625 ;
      RECT  3.4475 2.9375 3.5125 2.8025 ;
      RECT  3.2325 2.9375 3.2975 2.8025 ;
      RECT  3.4475 4.8025 3.5125 4.6675 ;
      RECT  3.2325 4.8025 3.2975 4.6675 ;
      RECT  3.2125 3.835 3.3475 3.77 ;
      RECT  3.48 3.835 3.545 3.77 ;
      RECT  3.14 2.5075 3.8275 2.4425 ;
      RECT  3.14 4.9825 3.8275 4.9175 ;
      RECT  4.165 2.9375 4.23 2.8025 ;
      RECT  3.92 2.9375 3.985 2.8025 ;
      RECT  4.41 2.9375 4.475 2.8025 ;
      RECT  4.165 4.8025 4.23 4.6675 ;
      RECT  3.92 4.8025 3.985 4.6675 ;
      RECT  4.41 4.8025 4.475 4.6675 ;
      RECT  3.9 3.835 4.035 3.77 ;
      RECT  4.1975 3.835 4.2625 3.77 ;
      RECT  3.8275 2.5075 4.79 2.4425 ;
      RECT  3.8275 4.9825 4.79 4.9175 ;
      RECT  0.0 2.545 4.79 2.415 ;
      RECT  0.0 5.015 4.79 4.885 ;
      RECT  6.3575 2.1475 6.4225 2.2825 ;
      RECT  6.1425 2.1475 6.2075 2.2825 ;
      RECT  6.3575 0.1025 6.4225 0.2375 ;
      RECT  6.1425 0.1025 6.2075 0.2375 ;
      RECT  6.1225 1.16 6.2575 1.225 ;
      RECT  6.39 1.16 6.455 1.225 ;
      RECT  6.05 2.4425 6.7375 2.5075 ;
      RECT  6.05 -0.0325 6.7375 0.0325 ;
      RECT  7.045 2.0125 7.11 2.1475 ;
      RECT  6.83 2.0125 6.895 2.1475 ;
      RECT  7.045 0.1475 7.11 0.2825 ;
      RECT  6.83 0.1475 6.895 0.2825 ;
      RECT  6.81 1.115 6.945 1.18 ;
      RECT  7.0775 1.115 7.1425 1.18 ;
      RECT  6.7375 2.4425 7.2025 2.5075 ;
      RECT  6.7375 -0.0325 7.2025 0.0325 ;
      RECT  7.54 1.945 7.605 2.08 ;
      RECT  7.785 1.945 7.85 2.08 ;
      RECT  7.295 1.945 7.36 2.08 ;
      RECT  7.54 0.17 7.605 0.305 ;
      RECT  7.785 0.17 7.85 0.305 ;
      RECT  7.295 0.17 7.36 0.305 ;
      RECT  7.275 1.0925 7.41 1.1575 ;
      RECT  7.5725 1.0925 7.6375 1.1575 ;
      RECT  7.2025 2.4425 7.9425 2.5075 ;
      RECT  7.2025 -0.0325 7.9425 0.0325 ;
      RECT  8.28 1.7475 9.415 1.8125 ;
      RECT  8.555 1.8775 8.62 2.0125 ;
      RECT  8.035 1.8775 8.1 2.0125 ;
      RECT  9.105 1.8775 9.17 2.0125 ;
      RECT  8.28 0.3925 9.415 0.4575 ;
      RECT  8.035 0.1925 8.1 0.3275 ;
      RECT  9.105 0.1925 9.17 0.3275 ;
      RECT  8.555 0.1925 8.62 0.3275 ;
      RECT  8.015 1.07 8.15 1.135 ;
      RECT  8.8475 1.07 8.9125 1.135 ;
      RECT  7.9425 2.4425 9.5275 2.5075 ;
      RECT  7.9425 -0.0325 9.5275 0.0325 ;
      RECT  6.1225 1.16 6.2575 1.225 ;
      RECT  8.8475 1.07 8.9125 1.135 ;
      RECT  6.05 2.4425 9.5275 2.5075 ;
      RECT  6.05 -0.0325 9.5275 0.0325 ;
      RECT  6.3575 2.8025 6.4225 2.6675 ;
      RECT  6.1425 2.8025 6.2075 2.6675 ;
      RECT  6.3575 4.8475 6.4225 4.7125 ;
      RECT  6.1425 4.8475 6.2075 4.7125 ;
      RECT  6.1225 3.79 6.2575 3.725 ;
      RECT  6.39 3.79 6.455 3.725 ;
      RECT  6.05 2.5075 6.7375 2.4425 ;
      RECT  6.05 4.9825 6.7375 4.9175 ;
      RECT  7.045 2.8025 7.11 2.6675 ;
      RECT  6.83 2.8025 6.895 2.6675 ;
      RECT  7.26 2.8025 7.325 2.6675 ;
      RECT  7.045 2.8025 7.11 2.6675 ;
      RECT  6.83 4.8025 6.895 4.6675 ;
      RECT  7.26 4.8025 7.325 4.6675 ;
      RECT  6.9025 4.555 7.0375 4.49 ;
      RECT  7.1175 4.275 7.2525 4.21 ;
      RECT  7.39 2.9325 7.455 2.8675 ;
      RECT  6.7375 2.5075 7.4875 2.4425 ;
      RECT  6.7375 4.9825 7.4875 4.9175 ;
      RECT  7.825 3.2025 8.44 3.1375 ;
      RECT  8.1 3.0725 8.165 2.9375 ;
      RECT  7.58 3.0725 7.645 2.9375 ;
      RECT  8.62 3.0725 8.685 2.9375 ;
      RECT  7.825 4.5575 8.44 4.4925 ;
      RECT  7.58 4.7575 7.645 4.6225 ;
      RECT  8.62 4.7575 8.685 4.6225 ;
      RECT  8.1 4.7575 8.165 4.6225 ;
      RECT  7.56 3.88 7.695 3.815 ;
      RECT  8.1325 3.88 8.1975 3.815 ;
      RECT  7.4875 2.5075 9.0 2.4425 ;
      RECT  7.4875 4.9825 9.0 4.9175 ;
      RECT  7.56 3.88 7.695 3.815 ;
      RECT  8.1325 3.88 8.1975 3.815 ;
      RECT  7.4875 2.5075 9.0 2.4425 ;
      RECT  7.4875 4.9825 9.0 4.9175 ;
      RECT  6.9025 4.555 7.0375 4.49 ;
      RECT  7.1175 4.275 7.2525 4.21 ;
      RECT  8.1325 3.88 8.1975 3.815 ;
      RECT  6.7375 2.5075 9.0 2.4425 ;
      RECT  6.7375 4.9825 9.0 4.9175 ;
      RECT  6.3575 7.0975 6.4225 7.2325 ;
      RECT  6.1425 7.0975 6.2075 7.2325 ;
      RECT  6.5725 7.0975 6.6375 7.2325 ;
      RECT  6.3575 7.0975 6.4225 7.2325 ;
      RECT  6.1425 5.0975 6.2075 5.2325 ;
      RECT  6.5725 5.0975 6.6375 5.2325 ;
      RECT  6.215 5.345 6.35 5.41 ;
      RECT  6.43 5.625 6.565 5.69 ;
      RECT  6.7025 6.9675 6.7675 7.0325 ;
      RECT  6.05 7.3925 6.8 7.4575 ;
      RECT  6.05 4.9175 6.8 4.9825 ;
      RECT  7.1375 6.6975 7.7525 6.7625 ;
      RECT  7.4125 6.8275 7.4775 6.9625 ;
      RECT  6.8925 6.8275 6.9575 6.9625 ;
      RECT  7.9325 6.8275 7.9975 6.9625 ;
      RECT  7.1375 5.3425 7.7525 5.4075 ;
      RECT  6.8925 5.1425 6.9575 5.2775 ;
      RECT  7.9325 5.1425 7.9975 5.2775 ;
      RECT  7.4125 5.1425 7.4775 5.2775 ;
      RECT  6.8725 6.02 7.0075 6.085 ;
      RECT  7.445 6.02 7.51 6.085 ;
      RECT  6.8 7.3925 8.3125 7.4575 ;
      RECT  6.8 4.9175 8.3125 4.9825 ;
      RECT  6.8725 6.02 7.0075 6.085 ;
      RECT  7.445 6.02 7.51 6.085 ;
      RECT  6.8 7.3925 8.3125 7.4575 ;
      RECT  6.8 4.9175 8.3125 4.9825 ;
      RECT  6.215 5.345 6.35 5.41 ;
      RECT  6.43 5.625 6.565 5.69 ;
      RECT  7.445 6.02 7.51 6.085 ;
      RECT  6.05 7.3925 8.3125 7.4575 ;
      RECT  6.05 4.9175 8.3125 4.9825 ;
      RECT  6.3575 7.7525 6.4225 7.6175 ;
      RECT  6.1425 7.7525 6.2075 7.6175 ;
      RECT  6.3575 9.7975 6.4225 9.6625 ;
      RECT  6.1425 9.7975 6.2075 9.6625 ;
      RECT  6.1225 8.74 6.2575 8.675 ;
      RECT  6.39 8.74 6.455 8.675 ;
      RECT  6.05 7.4575 6.7375 7.3925 ;
      RECT  6.05 9.9325 6.7375 9.8675 ;
      RECT  7.045 7.7525 7.11 7.6175 ;
      RECT  6.83 7.7525 6.895 7.6175 ;
      RECT  7.045 9.7975 7.11 9.6625 ;
      RECT  6.83 9.7975 6.895 9.6625 ;
      RECT  6.81 8.74 6.945 8.675 ;
      RECT  7.0775 8.74 7.1425 8.675 ;
      RECT  6.7375 7.4575 7.2025 7.3925 ;
      RECT  6.7375 9.9325 7.2025 9.8675 ;
      RECT  7.51 7.8875 7.575 7.7525 ;
      RECT  7.295 7.8875 7.36 7.7525 ;
      RECT  7.51 9.7525 7.575 9.6175 ;
      RECT  7.295 9.7525 7.36 9.6175 ;
      RECT  7.275 8.785 7.41 8.72 ;
      RECT  7.5425 8.785 7.6075 8.72 ;
      RECT  7.2025 7.4575 7.6675 7.3925 ;
      RECT  7.2025 9.9325 7.6675 9.8675 ;
      RECT  8.005 7.955 8.07 7.82 ;
      RECT  8.25 7.955 8.315 7.82 ;
      RECT  7.76 7.955 7.825 7.82 ;
      RECT  8.005 9.73 8.07 9.595 ;
      RECT  8.25 9.73 8.315 9.595 ;
      RECT  7.76 9.73 7.825 9.595 ;
      RECT  7.74 8.8075 7.875 8.7425 ;
      RECT  8.0375 8.8075 8.1025 8.7425 ;
      RECT  7.6675 7.4575 8.4075 7.3925 ;
      RECT  7.6675 9.9325 8.4075 9.8675 ;
      RECT  6.1225 8.74 6.2575 8.675 ;
      RECT  8.0375 8.8075 8.1025 8.7425 ;
      RECT  6.05 7.4575 8.4075 7.3925 ;
      RECT  6.05 9.9325 8.4075 9.8675 ;
      RECT  6.3575 16.9975 6.4225 17.1325 ;
      RECT  6.1425 16.9975 6.2075 17.1325 ;
      RECT  6.3575 14.9525 6.4225 15.0875 ;
      RECT  6.1425 14.9525 6.2075 15.0875 ;
      RECT  6.1225 16.01 6.2575 16.075 ;
      RECT  6.39 16.01 6.455 16.075 ;
      RECT  6.05 17.2925 6.7375 17.3575 ;
      RECT  6.05 14.8175 6.7375 14.8825 ;
      RECT  6.3575 12.0475 6.4225 12.1825 ;
      RECT  6.1425 12.0475 6.2075 12.1825 ;
      RECT  6.5725 12.0475 6.6375 12.1825 ;
      RECT  6.3575 12.0475 6.4225 12.1825 ;
      RECT  6.7875 12.0475 6.8525 12.1825 ;
      RECT  6.5725 12.0475 6.6375 12.1825 ;
      RECT  6.1425 10.0475 6.2075 10.1825 ;
      RECT  6.7875 10.0475 6.8525 10.1825 ;
      RECT  6.1475 10.295 6.2825 10.36 ;
      RECT  6.43 10.435 6.565 10.5 ;
      RECT  6.7125 10.575 6.8475 10.64 ;
      RECT  6.9175 11.9175 6.9825 11.9825 ;
      RECT  6.05 12.3425 7.015 12.4075 ;
      RECT  6.05 9.8675 7.015 9.9325 ;
      RECT  7.3525 11.6025 7.9375 11.6675 ;
      RECT  7.6275 11.7325 7.6925 11.8675 ;
      RECT  7.1075 11.7325 7.1725 11.8675 ;
      RECT  7.3525 10.3075 7.9375 10.3725 ;
      RECT  7.6275 10.1075 7.6925 10.2425 ;
      RECT  7.1075 10.1075 7.1725 10.2425 ;
      RECT  7.0875 10.955 7.2225 11.02 ;
      RECT  7.645 10.955 7.71 11.02 ;
      RECT  7.015 12.3425 8.2525 12.4075 ;
      RECT  7.015 9.8675 8.2525 9.9325 ;
      RECT  7.0875 10.955 7.2225 11.02 ;
      RECT  7.645 10.955 7.71 11.02 ;
      RECT  7.015 12.3425 8.2525 12.4075 ;
      RECT  7.015 9.8675 8.2525 9.9325 ;
      RECT  6.1475 10.295 6.2825 10.36 ;
      RECT  6.43 10.435 6.565 10.5 ;
      RECT  6.7125 10.575 6.8475 10.64 ;
      RECT  7.645 10.955 7.71 11.02 ;
      RECT  6.05 12.3425 8.2525 12.4075 ;
      RECT  6.05 9.8675 8.2525 9.9325 ;
      RECT  6.3575 17.6525 6.4225 17.5175 ;
      RECT  6.1425 17.6525 6.2075 17.5175 ;
      RECT  6.5725 17.6525 6.6375 17.5175 ;
      RECT  6.3575 17.6525 6.4225 17.5175 ;
      RECT  6.7875 17.6525 6.8525 17.5175 ;
      RECT  6.5725 17.6525 6.6375 17.5175 ;
      RECT  6.1425 19.6525 6.2075 19.5175 ;
      RECT  6.7875 19.6525 6.8525 19.5175 ;
      RECT  6.1475 19.405 6.2825 19.34 ;
      RECT  6.43 19.265 6.565 19.2 ;
      RECT  6.7125 19.125 6.8475 19.06 ;
      RECT  6.9175 17.7825 6.9825 17.7175 ;
      RECT  6.05 17.3575 7.015 17.2925 ;
      RECT  6.05 19.8325 7.015 19.7675 ;
      RECT  7.3225 17.7875 7.3875 17.6525 ;
      RECT  7.1075 17.7875 7.1725 17.6525 ;
      RECT  7.3225 19.6525 7.3875 19.5175 ;
      RECT  7.1075 19.6525 7.1725 19.5175 ;
      RECT  7.0875 18.685 7.2225 18.62 ;
      RECT  7.355 18.685 7.42 18.62 ;
      RECT  7.015 17.3575 7.7025 17.2925 ;
      RECT  7.015 19.8325 7.7025 19.7675 ;
      RECT  7.0875 18.685 7.2225 18.62 ;
      RECT  7.355 18.685 7.42 18.62 ;
      RECT  7.015 17.3575 7.7025 17.2925 ;
      RECT  7.015 19.8325 7.7025 19.7675 ;
      RECT  6.1475 19.405 6.2825 19.34 ;
      RECT  6.43 19.265 6.565 19.2 ;
      RECT  6.7125 19.125 6.8475 19.06 ;
      RECT  7.355 18.685 7.42 18.62 ;
      RECT  6.05 17.3575 7.7025 17.2925 ;
      RECT  6.05 19.8325 7.7025 19.7675 ;
      RECT  3.13 21.5525 3.065 21.6875 ;
      RECT  3.345 21.5525 3.28 21.6875 ;
      RECT  3.13 20.1625 3.065 20.2975 ;
      RECT  3.345 20.1625 3.28 20.2975 ;
      RECT  3.365 20.8925 3.23 20.9575 ;
      RECT  3.0975 20.8925 3.0325 20.9575 ;
      RECT  3.4375 21.8475 2.75 21.9125 ;
      RECT  3.4375 20.0275 2.75 20.0925 ;
      RECT  2.4425 21.5525 2.3775 21.6875 ;
      RECT  2.6575 21.5525 2.5925 21.6875 ;
      RECT  2.4425 20.1625 2.3775 20.2975 ;
      RECT  2.6575 20.1625 2.5925 20.2975 ;
      RECT  2.6775 20.8925 2.5425 20.9575 ;
      RECT  2.41 20.8925 2.345 20.9575 ;
      RECT  2.75 21.8475 2.0625 21.9125 ;
      RECT  2.75 20.0275 2.0625 20.0925 ;
      RECT  1.755 21.5525 1.69 21.6875 ;
      RECT  1.97 21.5525 1.905 21.6875 ;
      RECT  1.755 20.1625 1.69 20.2975 ;
      RECT  1.97 20.1625 1.905 20.2975 ;
      RECT  1.99 20.8925 1.855 20.9575 ;
      RECT  1.7225 20.8925 1.6575 20.9575 ;
      RECT  2.0625 21.8475 1.375 21.9125 ;
      RECT  2.0625 20.0275 1.375 20.0925 ;
      RECT  1.0675 21.5525 1.0025 21.6875 ;
      RECT  1.2825 21.5525 1.2175 21.6875 ;
      RECT  1.0675 20.1625 1.0025 20.2975 ;
      RECT  1.2825 20.1625 1.2175 20.2975 ;
      RECT  1.3025 20.8925 1.1675 20.9575 ;
      RECT  1.035 20.8925 0.97 20.9575 ;
      RECT  1.375 21.8475 0.6875 21.9125 ;
      RECT  1.375 20.0275 0.6875 20.0925 ;
      RECT  0.38 21.5525 0.315 21.6875 ;
      RECT  0.595 21.5525 0.53 21.6875 ;
      RECT  0.38 20.1625 0.315 20.2975 ;
      RECT  0.595 20.1625 0.53 20.2975 ;
      RECT  0.615 20.8925 0.48 20.9575 ;
      RECT  0.3475 20.8925 0.2825 20.9575 ;
      RECT  0.6875 21.8475 0.0 21.9125 ;
      RECT  0.6875 20.0275 0.0 20.0925 ;
      RECT  3.13 22.2075 3.065 22.0725 ;
      RECT  3.345 22.2075 3.28 22.0725 ;
      RECT  3.13 23.5975 3.065 23.4625 ;
      RECT  3.345 23.5975 3.28 23.4625 ;
      RECT  3.365 22.8675 3.23 22.8025 ;
      RECT  3.0975 22.8675 3.0325 22.8025 ;
      RECT  3.4375 21.9125 2.75 21.8475 ;
      RECT  3.4375 23.7325 2.75 23.6675 ;
      RECT  2.4425 22.2075 2.3775 22.0725 ;
      RECT  2.6575 22.2075 2.5925 22.0725 ;
      RECT  2.4425 23.5975 2.3775 23.4625 ;
      RECT  2.6575 23.5975 2.5925 23.4625 ;
      RECT  2.6775 22.8675 2.5425 22.8025 ;
      RECT  2.41 22.8675 2.345 22.8025 ;
      RECT  2.75 21.9125 2.0625 21.8475 ;
      RECT  2.75 23.7325 2.0625 23.6675 ;
      RECT  1.755 22.2075 1.69 22.0725 ;
      RECT  1.97 22.2075 1.905 22.0725 ;
      RECT  1.755 23.5975 1.69 23.4625 ;
      RECT  1.97 23.5975 1.905 23.4625 ;
      RECT  1.99 22.8675 1.855 22.8025 ;
      RECT  1.7225 22.8675 1.6575 22.8025 ;
      RECT  2.0625 21.9125 1.375 21.8475 ;
      RECT  2.0625 23.7325 1.375 23.6675 ;
      RECT  1.0675 22.2075 1.0025 22.0725 ;
      RECT  1.2825 22.2075 1.2175 22.0725 ;
      RECT  1.0675 23.5975 1.0025 23.4625 ;
      RECT  1.2825 23.5975 1.2175 23.4625 ;
      RECT  1.3025 22.8675 1.1675 22.8025 ;
      RECT  1.035 22.8675 0.97 22.8025 ;
      RECT  1.375 21.9125 0.6875 21.8475 ;
      RECT  1.375 23.7325 0.6875 23.6675 ;
      RECT  0.38 22.2075 0.315 22.0725 ;
      RECT  0.595 22.2075 0.53 22.0725 ;
      RECT  0.38 23.5975 0.315 23.4625 ;
      RECT  0.595 23.5975 0.53 23.4625 ;
      RECT  0.615 22.8675 0.48 22.8025 ;
      RECT  0.3475 22.8675 0.2825 22.8025 ;
      RECT  0.6875 21.9125 0.0 21.8475 ;
      RECT  0.6875 23.7325 0.0 23.6675 ;
      RECT  3.13 25.1925 3.065 25.3275 ;
      RECT  3.345 25.1925 3.28 25.3275 ;
      RECT  3.13 23.8025 3.065 23.9375 ;
      RECT  3.345 23.8025 3.28 23.9375 ;
      RECT  3.365 24.5325 3.23 24.5975 ;
      RECT  3.0975 24.5325 3.0325 24.5975 ;
      RECT  3.4375 25.4875 2.75 25.5525 ;
      RECT  3.4375 23.6675 2.75 23.7325 ;
      RECT  2.4425 25.1925 2.3775 25.3275 ;
      RECT  2.6575 25.1925 2.5925 25.3275 ;
      RECT  2.4425 23.8025 2.3775 23.9375 ;
      RECT  2.6575 23.8025 2.5925 23.9375 ;
      RECT  2.6775 24.5325 2.5425 24.5975 ;
      RECT  2.41 24.5325 2.345 24.5975 ;
      RECT  2.75 25.4875 2.0625 25.5525 ;
      RECT  2.75 23.6675 2.0625 23.7325 ;
      RECT  1.755 25.1925 1.69 25.3275 ;
      RECT  1.97 25.1925 1.905 25.3275 ;
      RECT  1.755 23.8025 1.69 23.9375 ;
      RECT  1.97 23.8025 1.905 23.9375 ;
      RECT  1.99 24.5325 1.855 24.5975 ;
      RECT  1.7225 24.5325 1.6575 24.5975 ;
      RECT  2.0625 25.4875 1.375 25.5525 ;
      RECT  2.0625 23.6675 1.375 23.7325 ;
      RECT  1.0675 25.1925 1.0025 25.3275 ;
      RECT  1.2825 25.1925 1.2175 25.3275 ;
      RECT  1.0675 23.8025 1.0025 23.9375 ;
      RECT  1.2825 23.8025 1.2175 23.9375 ;
      RECT  1.3025 24.5325 1.1675 24.5975 ;
      RECT  1.035 24.5325 0.97 24.5975 ;
      RECT  1.375 25.4875 0.6875 25.5525 ;
      RECT  1.375 23.6675 0.6875 23.7325 ;
      RECT  0.38 25.1925 0.315 25.3275 ;
      RECT  0.595 25.1925 0.53 25.3275 ;
      RECT  0.38 23.8025 0.315 23.9375 ;
      RECT  0.595 23.8025 0.53 23.9375 ;
      RECT  0.615 24.5325 0.48 24.5975 ;
      RECT  0.3475 24.5325 0.2825 24.5975 ;
      RECT  0.6875 25.4875 0.0 25.5525 ;
      RECT  0.6875 23.6675 0.0 23.7325 ;
      RECT  3.13 25.8475 3.065 25.7125 ;
      RECT  3.345 25.8475 3.28 25.7125 ;
      RECT  3.13 27.2375 3.065 27.1025 ;
      RECT  3.345 27.2375 3.28 27.1025 ;
      RECT  3.365 26.5075 3.23 26.4425 ;
      RECT  3.0975 26.5075 3.0325 26.4425 ;
      RECT  3.4375 25.5525 2.75 25.4875 ;
      RECT  3.4375 27.3725 2.75 27.3075 ;
      RECT  2.4425 25.8475 2.3775 25.7125 ;
      RECT  2.6575 25.8475 2.5925 25.7125 ;
      RECT  2.4425 27.2375 2.3775 27.1025 ;
      RECT  2.6575 27.2375 2.5925 27.1025 ;
      RECT  2.6775 26.5075 2.5425 26.4425 ;
      RECT  2.41 26.5075 2.345 26.4425 ;
      RECT  2.75 25.5525 2.0625 25.4875 ;
      RECT  2.75 27.3725 2.0625 27.3075 ;
      RECT  1.755 25.8475 1.69 25.7125 ;
      RECT  1.97 25.8475 1.905 25.7125 ;
      RECT  1.755 27.2375 1.69 27.1025 ;
      RECT  1.97 27.2375 1.905 27.1025 ;
      RECT  1.99 26.5075 1.855 26.4425 ;
      RECT  1.7225 26.5075 1.6575 26.4425 ;
      RECT  2.0625 25.5525 1.375 25.4875 ;
      RECT  2.0625 27.3725 1.375 27.3075 ;
      RECT  1.0675 25.8475 1.0025 25.7125 ;
      RECT  1.2825 25.8475 1.2175 25.7125 ;
      RECT  1.0675 27.2375 1.0025 27.1025 ;
      RECT  1.2825 27.2375 1.2175 27.1025 ;
      RECT  1.3025 26.5075 1.1675 26.4425 ;
      RECT  1.035 26.5075 0.97 26.4425 ;
      RECT  1.375 25.5525 0.6875 25.4875 ;
      RECT  1.375 27.3725 0.6875 27.3075 ;
      RECT  0.38 25.8475 0.315 25.7125 ;
      RECT  0.595 25.8475 0.53 25.7125 ;
      RECT  0.38 27.2375 0.315 27.1025 ;
      RECT  0.595 27.2375 0.53 27.1025 ;
      RECT  0.615 26.5075 0.48 26.4425 ;
      RECT  0.3475 26.5075 0.2825 26.4425 ;
      RECT  0.6875 25.5525 0.0 25.4875 ;
      RECT  0.6875 27.3725 0.0 27.3075 ;
      RECT  3.13 28.8325 3.065 28.9675 ;
      RECT  3.345 28.8325 3.28 28.9675 ;
      RECT  3.13 27.4425 3.065 27.5775 ;
      RECT  3.345 27.4425 3.28 27.5775 ;
      RECT  3.365 28.1725 3.23 28.2375 ;
      RECT  3.0975 28.1725 3.0325 28.2375 ;
      RECT  3.4375 29.1275 2.75 29.1925 ;
      RECT  3.4375 27.3075 2.75 27.3725 ;
      RECT  2.4425 28.8325 2.3775 28.9675 ;
      RECT  2.6575 28.8325 2.5925 28.9675 ;
      RECT  2.4425 27.4425 2.3775 27.5775 ;
      RECT  2.6575 27.4425 2.5925 27.5775 ;
      RECT  2.6775 28.1725 2.5425 28.2375 ;
      RECT  2.41 28.1725 2.345 28.2375 ;
      RECT  2.75 29.1275 2.0625 29.1925 ;
      RECT  2.75 27.3075 2.0625 27.3725 ;
      RECT  1.755 28.8325 1.69 28.9675 ;
      RECT  1.97 28.8325 1.905 28.9675 ;
      RECT  1.755 27.4425 1.69 27.5775 ;
      RECT  1.97 27.4425 1.905 27.5775 ;
      RECT  1.99 28.1725 1.855 28.2375 ;
      RECT  1.7225 28.1725 1.6575 28.2375 ;
      RECT  2.0625 29.1275 1.375 29.1925 ;
      RECT  2.0625 27.3075 1.375 27.3725 ;
      RECT  1.0675 28.8325 1.0025 28.9675 ;
      RECT  1.2825 28.8325 1.2175 28.9675 ;
      RECT  1.0675 27.4425 1.0025 27.5775 ;
      RECT  1.2825 27.4425 1.2175 27.5775 ;
      RECT  1.3025 28.1725 1.1675 28.2375 ;
      RECT  1.035 28.1725 0.97 28.2375 ;
      RECT  1.375 29.1275 0.6875 29.1925 ;
      RECT  1.375 27.3075 0.6875 27.3725 ;
      RECT  0.38 28.8325 0.315 28.9675 ;
      RECT  0.595 28.8325 0.53 28.9675 ;
      RECT  0.38 27.4425 0.315 27.5775 ;
      RECT  0.595 27.4425 0.53 27.5775 ;
      RECT  0.615 28.1725 0.48 28.2375 ;
      RECT  0.3475 28.1725 0.2825 28.2375 ;
      RECT  0.6875 29.1275 0.0 29.1925 ;
      RECT  0.6875 27.3075 0.0 27.3725 ;
      RECT  3.13 29.4875 3.065 29.3525 ;
      RECT  3.345 29.4875 3.28 29.3525 ;
      RECT  3.13 30.8775 3.065 30.7425 ;
      RECT  3.345 30.8775 3.28 30.7425 ;
      RECT  3.365 30.1475 3.23 30.0825 ;
      RECT  3.0975 30.1475 3.0325 30.0825 ;
      RECT  3.4375 29.1925 2.75 29.1275 ;
      RECT  3.4375 31.0125 2.75 30.9475 ;
      RECT  2.4425 29.4875 2.3775 29.3525 ;
      RECT  2.6575 29.4875 2.5925 29.3525 ;
      RECT  2.4425 30.8775 2.3775 30.7425 ;
      RECT  2.6575 30.8775 2.5925 30.7425 ;
      RECT  2.6775 30.1475 2.5425 30.0825 ;
      RECT  2.41 30.1475 2.345 30.0825 ;
      RECT  2.75 29.1925 2.0625 29.1275 ;
      RECT  2.75 31.0125 2.0625 30.9475 ;
      RECT  1.755 29.4875 1.69 29.3525 ;
      RECT  1.97 29.4875 1.905 29.3525 ;
      RECT  1.755 30.8775 1.69 30.7425 ;
      RECT  1.97 30.8775 1.905 30.7425 ;
      RECT  1.99 30.1475 1.855 30.0825 ;
      RECT  1.7225 30.1475 1.6575 30.0825 ;
      RECT  2.0625 29.1925 1.375 29.1275 ;
      RECT  2.0625 31.0125 1.375 30.9475 ;
      RECT  1.0675 29.4875 1.0025 29.3525 ;
      RECT  1.2825 29.4875 1.2175 29.3525 ;
      RECT  1.0675 30.8775 1.0025 30.7425 ;
      RECT  1.2825 30.8775 1.2175 30.7425 ;
      RECT  1.3025 30.1475 1.1675 30.0825 ;
      RECT  1.035 30.1475 0.97 30.0825 ;
      RECT  1.375 29.1925 0.6875 29.1275 ;
      RECT  1.375 31.0125 0.6875 30.9475 ;
      RECT  0.38 29.4875 0.315 29.3525 ;
      RECT  0.595 29.4875 0.53 29.3525 ;
      RECT  0.38 30.8775 0.315 30.7425 ;
      RECT  0.595 30.8775 0.53 30.7425 ;
      RECT  0.615 30.1475 0.48 30.0825 ;
      RECT  0.3475 30.1475 0.2825 30.0825 ;
      RECT  0.6875 29.1925 0.0 29.1275 ;
      RECT  0.6875 31.0125 0.0 30.9475 ;
      RECT  3.13 32.4725 3.065 32.6075 ;
      RECT  3.345 32.4725 3.28 32.6075 ;
      RECT  3.13 31.0825 3.065 31.2175 ;
      RECT  3.345 31.0825 3.28 31.2175 ;
      RECT  3.365 31.8125 3.23 31.8775 ;
      RECT  3.0975 31.8125 3.0325 31.8775 ;
      RECT  3.4375 32.7675 2.75 32.8325 ;
      RECT  3.4375 30.9475 2.75 31.0125 ;
      RECT  2.4425 32.4725 2.3775 32.6075 ;
      RECT  2.6575 32.4725 2.5925 32.6075 ;
      RECT  2.4425 31.0825 2.3775 31.2175 ;
      RECT  2.6575 31.0825 2.5925 31.2175 ;
      RECT  2.6775 31.8125 2.5425 31.8775 ;
      RECT  2.41 31.8125 2.345 31.8775 ;
      RECT  2.75 32.7675 2.0625 32.8325 ;
      RECT  2.75 30.9475 2.0625 31.0125 ;
      RECT  1.755 32.4725 1.69 32.6075 ;
      RECT  1.97 32.4725 1.905 32.6075 ;
      RECT  1.755 31.0825 1.69 31.2175 ;
      RECT  1.97 31.0825 1.905 31.2175 ;
      RECT  1.99 31.8125 1.855 31.8775 ;
      RECT  1.7225 31.8125 1.6575 31.8775 ;
      RECT  2.0625 32.7675 1.375 32.8325 ;
      RECT  2.0625 30.9475 1.375 31.0125 ;
      RECT  1.0675 32.4725 1.0025 32.6075 ;
      RECT  1.2825 32.4725 1.2175 32.6075 ;
      RECT  1.0675 31.0825 1.0025 31.2175 ;
      RECT  1.2825 31.0825 1.2175 31.2175 ;
      RECT  1.3025 31.8125 1.1675 31.8775 ;
      RECT  1.035 31.8125 0.97 31.8775 ;
      RECT  1.375 32.7675 0.6875 32.8325 ;
      RECT  1.375 30.9475 0.6875 31.0125 ;
      RECT  0.38 32.4725 0.315 32.6075 ;
      RECT  0.595 32.4725 0.53 32.6075 ;
      RECT  0.38 31.0825 0.315 31.2175 ;
      RECT  0.595 31.0825 0.53 31.2175 ;
      RECT  0.615 31.8125 0.48 31.8775 ;
      RECT  0.3475 31.8125 0.2825 31.8775 ;
      RECT  0.6875 32.7675 0.0 32.8325 ;
      RECT  0.6875 30.9475 0.0 31.0125 ;
      RECT  3.13 33.1275 3.065 32.9925 ;
      RECT  3.345 33.1275 3.28 32.9925 ;
      RECT  3.13 34.5175 3.065 34.3825 ;
      RECT  3.345 34.5175 3.28 34.3825 ;
      RECT  3.365 33.7875 3.23 33.7225 ;
      RECT  3.0975 33.7875 3.0325 33.7225 ;
      RECT  3.4375 32.8325 2.75 32.7675 ;
      RECT  3.4375 34.6525 2.75 34.5875 ;
      RECT  2.4425 33.1275 2.3775 32.9925 ;
      RECT  2.6575 33.1275 2.5925 32.9925 ;
      RECT  2.4425 34.5175 2.3775 34.3825 ;
      RECT  2.6575 34.5175 2.5925 34.3825 ;
      RECT  2.6775 33.7875 2.5425 33.7225 ;
      RECT  2.41 33.7875 2.345 33.7225 ;
      RECT  2.75 32.8325 2.0625 32.7675 ;
      RECT  2.75 34.6525 2.0625 34.5875 ;
      RECT  1.755 33.1275 1.69 32.9925 ;
      RECT  1.97 33.1275 1.905 32.9925 ;
      RECT  1.755 34.5175 1.69 34.3825 ;
      RECT  1.97 34.5175 1.905 34.3825 ;
      RECT  1.99 33.7875 1.855 33.7225 ;
      RECT  1.7225 33.7875 1.6575 33.7225 ;
      RECT  2.0625 32.8325 1.375 32.7675 ;
      RECT  2.0625 34.6525 1.375 34.5875 ;
      RECT  1.0675 33.1275 1.0025 32.9925 ;
      RECT  1.2825 33.1275 1.2175 32.9925 ;
      RECT  1.0675 34.5175 1.0025 34.3825 ;
      RECT  1.2825 34.5175 1.2175 34.3825 ;
      RECT  1.3025 33.7875 1.1675 33.7225 ;
      RECT  1.035 33.7875 0.97 33.7225 ;
      RECT  1.375 32.8325 0.6875 32.7675 ;
      RECT  1.375 34.6525 0.6875 34.5875 ;
      RECT  0.38 33.1275 0.315 32.9925 ;
      RECT  0.595 33.1275 0.53 32.9925 ;
      RECT  0.38 34.5175 0.315 34.3825 ;
      RECT  0.595 34.5175 0.53 34.3825 ;
      RECT  0.615 33.7875 0.48 33.7225 ;
      RECT  0.3475 33.7875 0.2825 33.7225 ;
      RECT  0.6875 32.8325 0.0 32.7675 ;
      RECT  0.6875 34.6525 0.0 34.5875 ;
      RECT  3.13 36.1125 3.065 36.2475 ;
      RECT  3.345 36.1125 3.28 36.2475 ;
      RECT  3.13 34.7225 3.065 34.8575 ;
      RECT  3.345 34.7225 3.28 34.8575 ;
      RECT  3.365 35.4525 3.23 35.5175 ;
      RECT  3.0975 35.4525 3.0325 35.5175 ;
      RECT  3.4375 36.4075 2.75 36.4725 ;
      RECT  3.4375 34.5875 2.75 34.6525 ;
      RECT  2.4425 36.1125 2.3775 36.2475 ;
      RECT  2.6575 36.1125 2.5925 36.2475 ;
      RECT  2.4425 34.7225 2.3775 34.8575 ;
      RECT  2.6575 34.7225 2.5925 34.8575 ;
      RECT  2.6775 35.4525 2.5425 35.5175 ;
      RECT  2.41 35.4525 2.345 35.5175 ;
      RECT  2.75 36.4075 2.0625 36.4725 ;
      RECT  2.75 34.5875 2.0625 34.6525 ;
      RECT  1.755 36.1125 1.69 36.2475 ;
      RECT  1.97 36.1125 1.905 36.2475 ;
      RECT  1.755 34.7225 1.69 34.8575 ;
      RECT  1.97 34.7225 1.905 34.8575 ;
      RECT  1.99 35.4525 1.855 35.5175 ;
      RECT  1.7225 35.4525 1.6575 35.5175 ;
      RECT  2.0625 36.4075 1.375 36.4725 ;
      RECT  2.0625 34.5875 1.375 34.6525 ;
      RECT  1.0675 36.1125 1.0025 36.2475 ;
      RECT  1.2825 36.1125 1.2175 36.2475 ;
      RECT  1.0675 34.7225 1.0025 34.8575 ;
      RECT  1.2825 34.7225 1.2175 34.8575 ;
      RECT  1.3025 35.4525 1.1675 35.5175 ;
      RECT  1.035 35.4525 0.97 35.5175 ;
      RECT  1.375 36.4075 0.6875 36.4725 ;
      RECT  1.375 34.5875 0.6875 34.6525 ;
      RECT  0.38 36.1125 0.315 36.2475 ;
      RECT  0.595 36.1125 0.53 36.2475 ;
      RECT  0.38 34.7225 0.315 34.8575 ;
      RECT  0.595 34.7225 0.53 34.8575 ;
      RECT  0.615 35.4525 0.48 35.5175 ;
      RECT  0.3475 35.4525 0.2825 35.5175 ;
      RECT  0.6875 36.4075 0.0 36.4725 ;
      RECT  0.6875 34.5875 0.0 34.6525 ;
      RECT  6.3575 12.7025 6.4225 12.5675 ;
      RECT  6.1425 12.7025 6.2075 12.5675 ;
      RECT  6.5725 12.7025 6.6375 12.5675 ;
      RECT  6.3575 12.7025 6.4225 12.5675 ;
      RECT  6.1425 14.7025 6.2075 14.5675 ;
      RECT  6.5725 14.7025 6.6375 14.5675 ;
      RECT  6.215 14.455 6.35 14.39 ;
      RECT  6.43 14.175 6.565 14.11 ;
      RECT  6.7025 12.8325 6.7675 12.7675 ;
      RECT  6.05 12.4075 6.9525 12.3425 ;
      RECT  6.05 14.8825 6.9525 14.8175 ;
      RECT  7.26 12.7025 7.325 12.5675 ;
      RECT  7.045 12.7025 7.11 12.5675 ;
      RECT  7.26 14.7475 7.325 14.6125 ;
      RECT  7.045 14.7475 7.11 14.6125 ;
      RECT  7.025 13.69 7.16 13.625 ;
      RECT  7.2925 13.69 7.3575 13.625 ;
      RECT  6.9525 12.4075 7.64 12.3425 ;
      RECT  6.9525 14.8825 7.64 14.8175 ;
      RECT  7.9475 12.7025 8.0125 12.5675 ;
      RECT  7.7325 12.7025 7.7975 12.5675 ;
      RECT  7.9475 14.7475 8.0125 14.6125 ;
      RECT  7.7325 14.7475 7.7975 14.6125 ;
      RECT  7.7125 13.69 7.8475 13.625 ;
      RECT  7.98 13.69 8.045 13.625 ;
      RECT  7.64 12.4075 8.105 12.3425 ;
      RECT  7.64 14.8825 8.105 14.8175 ;
      RECT  7.025 13.69 7.16 13.625 ;
      RECT  7.98 13.69 8.045 13.625 ;
      RECT  6.9525 12.4075 8.105 12.3425 ;
      RECT  6.9525 14.8825 8.105 14.8175 ;
      RECT  6.8075 36.635 9.6675 36.765 ;
      POLYGON  8.655 38.1425 8.655 38.9675 9.2 38.9675 9.2 38.9025 8.72 38.9025 8.72 38.5575 8.915 38.5575 8.915 38.1425 8.655 38.1425 ;
      RECT  9.44 37.7475 9.5175 37.8825 ;
      POLYGON  7.225 37.035 7.225 37.675 7.525 37.675 7.525 38.5625 7.455 38.5625 7.455 38.6275 7.59 38.6275 7.59 38.4975 8.18 38.4975 8.18 38.8475 8.245 38.8475 8.245 38.3575 8.525 38.3575 8.525 38.7725 8.59 38.7725 8.59 38.2925 8.18 38.2925 8.18 38.4325 7.59 38.4325 7.59 37.61 7.29 37.61 7.29 37.1 8.18 37.1 8.18 37.4925 8.245 37.4925 8.245 37.035 7.225 37.035 ;
      RECT  8.855 37.2875 8.92 37.5625 ;
      POLYGON  7.325 38.0825 7.325 38.7575 7.97 38.7575 7.97 38.6225 7.905 38.6225 7.905 38.6925 7.39 38.6925 7.39 38.4975 7.415 38.4975 7.415 38.0825 7.325 38.0825 ;
      POLYGON  9.45 36.9175 9.45 37.6175 9.345 37.6175 9.345 37.6825 9.45 37.6825 9.45 38.3475 9.12 38.3475 9.12 38.4125 9.45 38.4125 9.45 38.9375 9.515 38.9375 9.515 36.9175 9.45 36.9175 ;
      POLYGON  8.585 37.6275 8.585 37.8425 8.355 37.8425 8.355 37.715 8.22 37.715 8.22 38.1625 7.98 38.1625 7.98 38.3675 8.115 38.3675 8.115 38.2275 8.285 38.2275 8.285 37.9075 8.78 37.9075 8.78 37.6925 8.995 37.6925 8.995 37.8925 9.13 37.8925 9.13 37.8275 9.06 37.8275 9.06 37.6275 8.585 37.6275 ;
      POLYGON  6.975 37.9675 6.975 39.105 6.9075 39.105 6.9075 39.235 9.6675 39.235 9.6675 39.105 9.33 39.105 9.33 38.6075 9.265 38.6075 9.265 39.105 8.43 39.105 8.43 38.4225 8.365 38.4225 8.365 39.105 7.865 39.105 7.865 38.9525 7.73 38.9525 7.73 39.105 7.04 39.105 7.04 37.9675 6.975 37.9675 ;
      RECT  9.45 37.615 9.515 37.8275 ;
      POLYGON  8.915 36.9275 8.915 37.2025 9.045 37.2025 9.045 37.4625 9.11 37.4625 9.11 37.1375 8.98 37.1375 8.98 36.9275 8.915 36.9275 ;
      RECT  7.0525 37.7375 7.13 37.8725 ;
      RECT  8.585 37.6275 8.78 37.9075 ;
      POLYGON  7.195 37.8175 7.195 38.8875 8.1 38.8875 8.1 38.5625 8.035 38.5625 8.035 38.8225 7.26 38.8225 7.26 37.8825 7.345 37.8825 7.345 37.8175 7.195 37.8175 ;
      POLYGON  6.9075 36.635 6.9075 36.765 6.975 36.765 6.975 37.545 7.04 37.545 7.04 36.765 7.725 36.765 7.725 36.935 7.86 36.935 7.86 36.765 8.365 36.765 8.365 37.4925 8.43 37.4925 8.43 36.765 8.73 36.765 8.73 37.1675 8.795 37.1675 8.795 36.765 9.215 36.765 9.215 37.6875 9.28 37.6875 9.28 36.765 9.5675 36.765 9.5675 36.635 6.9075 36.635 ;
      POLYGON  8.025 37.385 8.025 37.65 7.75 37.65 7.75 37.715 8.025 37.715 8.025 38.0975 8.09 38.0975 8.09 37.65 8.42 37.65 8.42 37.7775 8.485 37.7775 8.485 37.585 8.09 37.585 8.09 37.385 8.025 37.385 ;
      POLYGON  8.86 37.7575 8.86 38.0225 9.31 38.0225 9.31 38.2175 9.11 38.2175 9.11 38.2825 9.375 38.2825 9.375 37.7575 9.21 37.7575 9.21 37.8925 9.31 37.8925 9.31 37.9575 8.925 37.9575 8.925 37.7575 8.86 37.7575 ;
      RECT  9.135 38.4775 9.2 38.8275 ;
      RECT  6.8075 39.105 9.5675 39.235 ;
      POLYGON  7.355 37.165 7.355 37.545 7.42 37.545 7.42 37.23 8.02 37.23 8.02 37.165 7.355 37.165 ;
      POLYGON  8.98 38.0875 8.98 38.8375 9.07 38.8375 9.07 38.5625 9.045 38.5625 9.045 38.1525 9.245 38.1525 9.245 38.0875 8.98 38.0875 ;
      RECT  6.8075 41.715 9.6675 41.585 ;
      POLYGON  8.655 40.2075 8.655 39.3825 9.2 39.3825 9.2 39.4475 8.72 39.4475 8.72 39.7925 8.915 39.7925 8.915 40.2075 8.655 40.2075 ;
      RECT  9.44 40.6025 9.5175 40.4675 ;
      POLYGON  7.225 41.315 7.225 40.675 7.525 40.675 7.525 39.7875 7.455 39.7875 7.455 39.7225 7.59 39.7225 7.59 39.8525 8.18 39.8525 8.18 39.5025 8.245 39.5025 8.245 39.9925 8.525 39.9925 8.525 39.5775 8.59 39.5775 8.59 40.0575 8.18 40.0575 8.18 39.9175 7.59 39.9175 7.59 40.74 7.29 40.74 7.29 41.25 8.18 41.25 8.18 40.8575 8.245 40.8575 8.245 41.315 7.225 41.315 ;
      RECT  8.855 41.0625 8.92 40.7875 ;
      POLYGON  7.325 40.2675 7.325 39.5925 7.97 39.5925 7.97 39.7275 7.905 39.7275 7.905 39.6575 7.39 39.6575 7.39 39.8525 7.415 39.8525 7.415 40.2675 7.325 40.2675 ;
      POLYGON  9.45 41.4325 9.45 40.7325 9.345 40.7325 9.345 40.6675 9.45 40.6675 9.45 40.0025 9.12 40.0025 9.12 39.9375 9.45 39.9375 9.45 39.4125 9.515 39.4125 9.515 41.4325 9.45 41.4325 ;
      POLYGON  8.585 40.7225 8.585 40.5075 8.355 40.5075 8.355 40.635 8.22 40.635 8.22 40.1875 7.98 40.1875 7.98 39.9825 8.115 39.9825 8.115 40.1225 8.285 40.1225 8.285 40.4425 8.78 40.4425 8.78 40.6575 8.995 40.6575 8.995 40.4575 9.13 40.4575 9.13 40.5225 9.06 40.5225 9.06 40.7225 8.585 40.7225 ;
      POLYGON  6.975 40.3825 6.975 39.245 6.9075 39.245 6.9075 39.115 9.6675 39.115 9.6675 39.245 9.33 39.245 9.33 39.7425 9.265 39.7425 9.265 39.245 8.43 39.245 8.43 39.9275 8.365 39.9275 8.365 39.245 7.865 39.245 7.865 39.3975 7.73 39.3975 7.73 39.245 7.04 39.245 7.04 40.3825 6.975 40.3825 ;
      RECT  9.45 40.735 9.515 40.5225 ;
      POLYGON  8.915 41.4225 8.915 41.1475 9.045 41.1475 9.045 40.8875 9.11 40.8875 9.11 41.2125 8.98 41.2125 8.98 41.4225 8.915 41.4225 ;
      RECT  7.0525 40.6125 7.13 40.4775 ;
      RECT  8.585 40.7225 8.78 40.4425 ;
      POLYGON  7.195 40.5325 7.195 39.4625 8.1 39.4625 8.1 39.7875 8.035 39.7875 8.035 39.5275 7.26 39.5275 7.26 40.4675 7.345 40.4675 7.345 40.5325 7.195 40.5325 ;
      POLYGON  6.9075 41.715 6.9075 41.585 6.975 41.585 6.975 40.805 7.04 40.805 7.04 41.585 7.725 41.585 7.725 41.415 7.86 41.415 7.86 41.585 8.365 41.585 8.365 40.8575 8.43 40.8575 8.43 41.585 8.73 41.585 8.73 41.1825 8.795 41.1825 8.795 41.585 9.215 41.585 9.215 40.6625 9.28 40.6625 9.28 41.585 9.5675 41.585 9.5675 41.715 6.9075 41.715 ;
      POLYGON  8.025 40.965 8.025 40.7 7.75 40.7 7.75 40.635 8.025 40.635 8.025 40.2525 8.09 40.2525 8.09 40.7 8.42 40.7 8.42 40.5725 8.485 40.5725 8.485 40.765 8.09 40.765 8.09 40.965 8.025 40.965 ;
      POLYGON  8.86 40.5925 8.86 40.3275 9.31 40.3275 9.31 40.1325 9.11 40.1325 9.11 40.0675 9.375 40.0675 9.375 40.5925 9.21 40.5925 9.21 40.4575 9.31 40.4575 9.31 40.3925 8.925 40.3925 8.925 40.5925 8.86 40.5925 ;
      RECT  9.135 39.8725 9.2 39.5225 ;
      RECT  6.8075 39.245 9.5675 39.115 ;
      POLYGON  7.355 41.185 7.355 40.805 7.42 40.805 7.42 41.12 8.02 41.12 8.02 41.185 7.355 41.185 ;
      POLYGON  8.98 40.2625 8.98 39.5125 9.07 39.5125 9.07 39.7875 9.045 39.7875 9.045 40.1975 9.245 40.1975 9.245 40.2625 8.98 40.2625 ;
      RECT  6.8075 41.585 9.6675 41.715 ;
      POLYGON  8.655 43.0925 8.655 43.9175 9.2 43.9175 9.2 43.8525 8.72 43.8525 8.72 43.5075 8.915 43.5075 8.915 43.0925 8.655 43.0925 ;
      RECT  9.44 42.6975 9.5175 42.8325 ;
      POLYGON  7.225 41.985 7.225 42.625 7.525 42.625 7.525 43.5125 7.455 43.5125 7.455 43.5775 7.59 43.5775 7.59 43.4475 8.18 43.4475 8.18 43.7975 8.245 43.7975 8.245 43.3075 8.525 43.3075 8.525 43.7225 8.59 43.7225 8.59 43.2425 8.18 43.2425 8.18 43.3825 7.59 43.3825 7.59 42.56 7.29 42.56 7.29 42.05 8.18 42.05 8.18 42.4425 8.245 42.4425 8.245 41.985 7.225 41.985 ;
      RECT  8.855 42.2375 8.92 42.5125 ;
      POLYGON  7.325 43.0325 7.325 43.7075 7.97 43.7075 7.97 43.5725 7.905 43.5725 7.905 43.6425 7.39 43.6425 7.39 43.4475 7.415 43.4475 7.415 43.0325 7.325 43.0325 ;
      POLYGON  9.45 41.8675 9.45 42.5675 9.345 42.5675 9.345 42.6325 9.45 42.6325 9.45 43.2975 9.12 43.2975 9.12 43.3625 9.45 43.3625 9.45 43.8875 9.515 43.8875 9.515 41.8675 9.45 41.8675 ;
      POLYGON  8.585 42.5775 8.585 42.7925 8.355 42.7925 8.355 42.665 8.22 42.665 8.22 43.1125 7.98 43.1125 7.98 43.3175 8.115 43.3175 8.115 43.1775 8.285 43.1775 8.285 42.8575 8.78 42.8575 8.78 42.6425 8.995 42.6425 8.995 42.8425 9.13 42.8425 9.13 42.7775 9.06 42.7775 9.06 42.5775 8.585 42.5775 ;
      POLYGON  6.975 42.9175 6.975 44.055 6.9075 44.055 6.9075 44.185 9.6675 44.185 9.6675 44.055 9.33 44.055 9.33 43.5575 9.265 43.5575 9.265 44.055 8.43 44.055 8.43 43.3725 8.365 43.3725 8.365 44.055 7.865 44.055 7.865 43.9025 7.73 43.9025 7.73 44.055 7.04 44.055 7.04 42.9175 6.975 42.9175 ;
      RECT  9.45 42.565 9.515 42.7775 ;
      POLYGON  8.915 41.8775 8.915 42.1525 9.045 42.1525 9.045 42.4125 9.11 42.4125 9.11 42.0875 8.98 42.0875 8.98 41.8775 8.915 41.8775 ;
      RECT  7.0525 42.6875 7.13 42.8225 ;
      RECT  8.585 42.5775 8.78 42.8575 ;
      POLYGON  7.195 42.7675 7.195 43.8375 8.1 43.8375 8.1 43.5125 8.035 43.5125 8.035 43.7725 7.26 43.7725 7.26 42.8325 7.345 42.8325 7.345 42.7675 7.195 42.7675 ;
      POLYGON  6.9075 41.585 6.9075 41.715 6.975 41.715 6.975 42.495 7.04 42.495 7.04 41.715 7.725 41.715 7.725 41.885 7.86 41.885 7.86 41.715 8.365 41.715 8.365 42.4425 8.43 42.4425 8.43 41.715 8.73 41.715 8.73 42.1175 8.795 42.1175 8.795 41.715 9.215 41.715 9.215 42.6375 9.28 42.6375 9.28 41.715 9.5675 41.715 9.5675 41.585 6.9075 41.585 ;
      POLYGON  8.025 42.335 8.025 42.6 7.75 42.6 7.75 42.665 8.025 42.665 8.025 43.0475 8.09 43.0475 8.09 42.6 8.42 42.6 8.42 42.7275 8.485 42.7275 8.485 42.535 8.09 42.535 8.09 42.335 8.025 42.335 ;
      POLYGON  8.86 42.7075 8.86 42.9725 9.31 42.9725 9.31 43.1675 9.11 43.1675 9.11 43.2325 9.375 43.2325 9.375 42.7075 9.21 42.7075 9.21 42.8425 9.31 42.8425 9.31 42.9075 8.925 42.9075 8.925 42.7075 8.86 42.7075 ;
      RECT  9.135 43.4275 9.2 43.7775 ;
      RECT  6.8075 44.055 9.5675 44.185 ;
      POLYGON  7.355 42.115 7.355 42.495 7.42 42.495 7.42 42.18 8.02 42.18 8.02 42.115 7.355 42.115 ;
      POLYGON  8.98 43.0375 8.98 43.7875 9.07 43.7875 9.07 43.5125 9.045 43.5125 9.045 43.1025 9.245 43.1025 9.245 43.0375 8.98 43.0375 ;
      RECT  6.8075 46.665 9.6675 46.535 ;
      POLYGON  8.655 45.1575 8.655 44.3325 9.2 44.3325 9.2 44.3975 8.72 44.3975 8.72 44.7425 8.915 44.7425 8.915 45.1575 8.655 45.1575 ;
      RECT  9.44 45.5525 9.5175 45.4175 ;
      POLYGON  7.225 46.265 7.225 45.625 7.525 45.625 7.525 44.7375 7.455 44.7375 7.455 44.6725 7.59 44.6725 7.59 44.8025 8.18 44.8025 8.18 44.4525 8.245 44.4525 8.245 44.9425 8.525 44.9425 8.525 44.5275 8.59 44.5275 8.59 45.0075 8.18 45.0075 8.18 44.8675 7.59 44.8675 7.59 45.69 7.29 45.69 7.29 46.2 8.18 46.2 8.18 45.8075 8.245 45.8075 8.245 46.265 7.225 46.265 ;
      RECT  8.855 46.0125 8.92 45.7375 ;
      POLYGON  7.325 45.2175 7.325 44.5425 7.97 44.5425 7.97 44.6775 7.905 44.6775 7.905 44.6075 7.39 44.6075 7.39 44.8025 7.415 44.8025 7.415 45.2175 7.325 45.2175 ;
      POLYGON  9.45 46.3825 9.45 45.6825 9.345 45.6825 9.345 45.6175 9.45 45.6175 9.45 44.9525 9.12 44.9525 9.12 44.8875 9.45 44.8875 9.45 44.3625 9.515 44.3625 9.515 46.3825 9.45 46.3825 ;
      POLYGON  8.585 45.6725 8.585 45.4575 8.355 45.4575 8.355 45.585 8.22 45.585 8.22 45.1375 7.98 45.1375 7.98 44.9325 8.115 44.9325 8.115 45.0725 8.285 45.0725 8.285 45.3925 8.78 45.3925 8.78 45.6075 8.995 45.6075 8.995 45.4075 9.13 45.4075 9.13 45.4725 9.06 45.4725 9.06 45.6725 8.585 45.6725 ;
      POLYGON  6.975 45.3325 6.975 44.195 6.9075 44.195 6.9075 44.065 9.6675 44.065 9.6675 44.195 9.33 44.195 9.33 44.6925 9.265 44.6925 9.265 44.195 8.43 44.195 8.43 44.8775 8.365 44.8775 8.365 44.195 7.865 44.195 7.865 44.3475 7.73 44.3475 7.73 44.195 7.04 44.195 7.04 45.3325 6.975 45.3325 ;
      RECT  9.45 45.685 9.515 45.4725 ;
      POLYGON  8.915 46.3725 8.915 46.0975 9.045 46.0975 9.045 45.8375 9.11 45.8375 9.11 46.1625 8.98 46.1625 8.98 46.3725 8.915 46.3725 ;
      RECT  7.0525 45.5625 7.13 45.4275 ;
      RECT  8.585 45.6725 8.78 45.3925 ;
      POLYGON  7.195 45.4825 7.195 44.4125 8.1 44.4125 8.1 44.7375 8.035 44.7375 8.035 44.4775 7.26 44.4775 7.26 45.4175 7.345 45.4175 7.345 45.4825 7.195 45.4825 ;
      POLYGON  6.9075 46.665 6.9075 46.535 6.975 46.535 6.975 45.755 7.04 45.755 7.04 46.535 7.725 46.535 7.725 46.365 7.86 46.365 7.86 46.535 8.365 46.535 8.365 45.8075 8.43 45.8075 8.43 46.535 8.73 46.535 8.73 46.1325 8.795 46.1325 8.795 46.535 9.215 46.535 9.215 45.6125 9.28 45.6125 9.28 46.535 9.5675 46.535 9.5675 46.665 6.9075 46.665 ;
      POLYGON  8.025 45.915 8.025 45.65 7.75 45.65 7.75 45.585 8.025 45.585 8.025 45.2025 8.09 45.2025 8.09 45.65 8.42 45.65 8.42 45.5225 8.485 45.5225 8.485 45.715 8.09 45.715 8.09 45.915 8.025 45.915 ;
      POLYGON  8.86 45.5425 8.86 45.2775 9.31 45.2775 9.31 45.0825 9.11 45.0825 9.11 45.0175 9.375 45.0175 9.375 45.5425 9.21 45.5425 9.21 45.4075 9.31 45.4075 9.31 45.3425 8.925 45.3425 8.925 45.5425 8.86 45.5425 ;
      RECT  9.135 44.8225 9.2 44.4725 ;
      RECT  6.8075 44.195 9.5675 44.065 ;
      POLYGON  7.355 46.135 7.355 45.755 7.42 45.755 7.42 46.07 8.02 46.07 8.02 46.135 7.355 46.135 ;
      POLYGON  8.98 45.2125 8.98 44.4625 9.07 44.4625 9.07 44.7375 9.045 44.7375 9.045 45.1475 9.245 45.1475 9.245 45.2125 8.98 45.2125 ;
      RECT  12.5275 -0.065 15.3875 0.065 ;
      POLYGON  14.375 1.4425 14.375 2.2675 14.92 2.2675 14.92 2.2025 14.44 2.2025 14.44 1.8575 14.635 1.8575 14.635 1.4425 14.375 1.4425 ;
      RECT  15.16 1.0475 15.2375 1.1825 ;
      POLYGON  12.945 0.335 12.945 0.975 13.245 0.975 13.245 1.8625 13.175 1.8625 13.175 1.9275 13.31 1.9275 13.31 1.7975 13.9 1.7975 13.9 2.1475 13.965 2.1475 13.965 1.6575 14.245 1.6575 14.245 2.0725 14.31 2.0725 14.31 1.5925 13.9 1.5925 13.9 1.7325 13.31 1.7325 13.31 0.91 13.01 0.91 13.01 0.4 13.9 0.4 13.9 0.7925 13.965 0.7925 13.965 0.335 12.945 0.335 ;
      RECT  14.575 0.5875 14.64 0.8625 ;
      POLYGON  13.045 1.3825 13.045 2.0575 13.69 2.0575 13.69 1.9225 13.625 1.9225 13.625 1.9925 13.11 1.9925 13.11 1.7975 13.135 1.7975 13.135 1.3825 13.045 1.3825 ;
      POLYGON  15.17 0.2175 15.17 0.9175 15.065 0.9175 15.065 0.9825 15.17 0.9825 15.17 1.6475 14.84 1.6475 14.84 1.7125 15.17 1.7125 15.17 2.2375 15.235 2.2375 15.235 0.2175 15.17 0.2175 ;
      POLYGON  14.305 0.9275 14.305 1.1425 14.075 1.1425 14.075 1.015 13.94 1.015 13.94 1.4625 13.7 1.4625 13.7 1.6675 13.835 1.6675 13.835 1.5275 14.005 1.5275 14.005 1.2075 14.5 1.2075 14.5 0.9925 14.715 0.9925 14.715 1.1925 14.85 1.1925 14.85 1.1275 14.78 1.1275 14.78 0.9275 14.305 0.9275 ;
      POLYGON  12.695 1.2675 12.695 2.405 12.6275 2.405 12.6275 2.535 15.3875 2.535 15.3875 2.405 15.05 2.405 15.05 1.9075 14.985 1.9075 14.985 2.405 14.15 2.405 14.15 1.7225 14.085 1.7225 14.085 2.405 13.585 2.405 13.585 2.2525 13.45 2.2525 13.45 2.405 12.76 2.405 12.76 1.2675 12.695 1.2675 ;
      RECT  15.17 0.915 15.235 1.1275 ;
      POLYGON  14.635 0.2275 14.635 0.5025 14.765 0.5025 14.765 0.7625 14.83 0.7625 14.83 0.4375 14.7 0.4375 14.7 0.2275 14.635 0.2275 ;
      RECT  12.7725 1.0375 12.85 1.1725 ;
      RECT  14.305 0.9275 14.5 1.2075 ;
      POLYGON  12.915 1.1175 12.915 2.1875 13.82 2.1875 13.82 1.8625 13.755 1.8625 13.755 2.1225 12.98 2.1225 12.98 1.1825 13.065 1.1825 13.065 1.1175 12.915 1.1175 ;
      POLYGON  12.6275 -0.065 12.6275 0.065 12.695 0.065 12.695 0.845 12.76 0.845 12.76 0.065 13.445 0.065 13.445 0.235 13.58 0.235 13.58 0.065 14.085 0.065 14.085 0.7925 14.15 0.7925 14.15 0.065 14.45 0.065 14.45 0.4675 14.515 0.4675 14.515 0.065 14.935 0.065 14.935 0.9875 15.0 0.9875 15.0 0.065 15.2875 0.065 15.2875 -0.065 12.6275 -0.065 ;
      POLYGON  13.745 0.685 13.745 0.95 13.47 0.95 13.47 1.015 13.745 1.015 13.745 1.3975 13.81 1.3975 13.81 0.95 14.14 0.95 14.14 1.0775 14.205 1.0775 14.205 0.885 13.81 0.885 13.81 0.685 13.745 0.685 ;
      POLYGON  14.58 1.0575 14.58 1.3225 15.03 1.3225 15.03 1.5175 14.83 1.5175 14.83 1.5825 15.095 1.5825 15.095 1.0575 14.93 1.0575 14.93 1.1925 15.03 1.1925 15.03 1.2575 14.645 1.2575 14.645 1.0575 14.58 1.0575 ;
      RECT  14.855 1.7775 14.92 2.1275 ;
      RECT  12.5275 2.405 15.2875 2.535 ;
      POLYGON  13.075 0.465 13.075 0.845 13.14 0.845 13.14 0.53 13.74 0.53 13.74 0.465 13.075 0.465 ;
      POLYGON  14.7 1.3875 14.7 2.1375 14.79 2.1375 14.79 1.8625 14.765 1.8625 14.765 1.4525 14.965 1.4525 14.965 1.3875 14.7 1.3875 ;
      RECT  15.3875 -0.065 18.2475 0.065 ;
      POLYGON  17.235 1.4425 17.235 2.2675 17.78 2.2675 17.78 2.2025 17.3 2.2025 17.3 1.8575 17.495 1.8575 17.495 1.4425 17.235 1.4425 ;
      RECT  18.02 1.0475 18.0975 1.1825 ;
      POLYGON  15.805 0.335 15.805 0.975 16.105 0.975 16.105 1.8625 16.035 1.8625 16.035 1.9275 16.17 1.9275 16.17 1.7975 16.76 1.7975 16.76 2.1475 16.825 2.1475 16.825 1.6575 17.105 1.6575 17.105 2.0725 17.17 2.0725 17.17 1.5925 16.76 1.5925 16.76 1.7325 16.17 1.7325 16.17 0.91 15.87 0.91 15.87 0.4 16.76 0.4 16.76 0.7925 16.825 0.7925 16.825 0.335 15.805 0.335 ;
      RECT  17.435 0.5875 17.5 0.8625 ;
      POLYGON  15.905 1.3825 15.905 2.0575 16.55 2.0575 16.55 1.9225 16.485 1.9225 16.485 1.9925 15.97 1.9925 15.97 1.7975 15.995 1.7975 15.995 1.3825 15.905 1.3825 ;
      POLYGON  18.03 0.2175 18.03 0.9175 17.925 0.9175 17.925 0.9825 18.03 0.9825 18.03 1.6475 17.7 1.6475 17.7 1.7125 18.03 1.7125 18.03 2.2375 18.095 2.2375 18.095 0.2175 18.03 0.2175 ;
      POLYGON  17.165 0.9275 17.165 1.1425 16.935 1.1425 16.935 1.015 16.8 1.015 16.8 1.4625 16.56 1.4625 16.56 1.6675 16.695 1.6675 16.695 1.5275 16.865 1.5275 16.865 1.2075 17.36 1.2075 17.36 0.9925 17.575 0.9925 17.575 1.1925 17.71 1.1925 17.71 1.1275 17.64 1.1275 17.64 0.9275 17.165 0.9275 ;
      POLYGON  15.555 1.2675 15.555 2.405 15.4875 2.405 15.4875 2.535 18.2475 2.535 18.2475 2.405 17.91 2.405 17.91 1.9075 17.845 1.9075 17.845 2.405 17.01 2.405 17.01 1.7225 16.945 1.7225 16.945 2.405 16.445 2.405 16.445 2.2525 16.31 2.2525 16.31 2.405 15.62 2.405 15.62 1.2675 15.555 1.2675 ;
      RECT  18.03 0.915 18.095 1.1275 ;
      POLYGON  17.495 0.2275 17.495 0.5025 17.625 0.5025 17.625 0.7625 17.69 0.7625 17.69 0.4375 17.56 0.4375 17.56 0.2275 17.495 0.2275 ;
      RECT  15.6325 1.0375 15.71 1.1725 ;
      RECT  17.165 0.9275 17.36 1.2075 ;
      POLYGON  15.775 1.1175 15.775 2.1875 16.68 2.1875 16.68 1.8625 16.615 1.8625 16.615 2.1225 15.84 2.1225 15.84 1.1825 15.925 1.1825 15.925 1.1175 15.775 1.1175 ;
      POLYGON  15.4875 -0.065 15.4875 0.065 15.555 0.065 15.555 0.845 15.62 0.845 15.62 0.065 16.305 0.065 16.305 0.235 16.44 0.235 16.44 0.065 16.945 0.065 16.945 0.7925 17.01 0.7925 17.01 0.065 17.31 0.065 17.31 0.4675 17.375 0.4675 17.375 0.065 17.795 0.065 17.795 0.9875 17.86 0.9875 17.86 0.065 18.1475 0.065 18.1475 -0.065 15.4875 -0.065 ;
      POLYGON  16.605 0.685 16.605 0.95 16.33 0.95 16.33 1.015 16.605 1.015 16.605 1.3975 16.67 1.3975 16.67 0.95 17.0 0.95 17.0 1.0775 17.065 1.0775 17.065 0.885 16.67 0.885 16.67 0.685 16.605 0.685 ;
      POLYGON  17.44 1.0575 17.44 1.3225 17.89 1.3225 17.89 1.5175 17.69 1.5175 17.69 1.5825 17.955 1.5825 17.955 1.0575 17.79 1.0575 17.79 1.1925 17.89 1.1925 17.89 1.2575 17.505 1.2575 17.505 1.0575 17.44 1.0575 ;
      RECT  17.715 1.7775 17.78 2.1275 ;
      RECT  15.3875 2.405 18.1475 2.535 ;
      POLYGON  15.935 0.465 15.935 0.845 16.0 0.845 16.0 0.53 16.6 0.53 16.6 0.465 15.935 0.465 ;
      POLYGON  17.56 1.3875 17.56 2.1375 17.65 2.1375 17.65 1.8625 17.625 1.8625 17.625 1.4525 17.825 1.4525 17.825 1.3875 17.56 1.3875 ;
   LAYER  metal2 ;
      RECT  22.05 22.725 22.11 22.7825 ;
      RECT  21.34 23.5 21.41 23.635 ;
      RECT  21.525 22.65 21.595 24.195 ;
      RECT  22.0125 22.715 22.1475 22.785 ;
      RECT  22.045 22.65 22.115 24.195 ;
      RECT  21.34 22.65 21.41 24.195 ;
      RECT  21.79 23.0075 21.86 23.1425 ;
      RECT  22.045 22.7175 22.115 24.1275 ;
      RECT  21.595 23.0075 21.665 23.1425 ;
      RECT  21.5325 22.725 21.5875 22.7775 ;
      RECT  21.6875 24.0275 21.7575 24.1625 ;
      RECT  21.345 22.72 21.405 22.7775 ;
      RECT  22.045 23.5 22.115 23.635 ;
      RECT  21.3075 22.715 21.4425 22.785 ;
      RECT  21.8675 22.7175 21.925 22.7775 ;
      RECT  21.86 22.65 21.93 24.195 ;
      RECT  22.05 25.465 22.11 25.4075 ;
      RECT  21.34 24.69 21.41 24.555 ;
      RECT  21.525 25.54 21.595 23.995 ;
      RECT  22.0125 25.475 22.1475 25.405 ;
      RECT  22.045 25.54 22.115 23.995 ;
      RECT  21.34 25.54 21.41 23.995 ;
      RECT  21.79 25.1825 21.86 25.0475 ;
      RECT  22.045 25.4725 22.115 24.0625 ;
      RECT  21.595 25.1825 21.665 25.0475 ;
      RECT  21.5325 25.465 21.5875 25.4125 ;
      RECT  21.6875 24.1625 21.7575 24.0275 ;
      RECT  21.345 25.47 21.405 25.4125 ;
      RECT  22.045 24.69 22.115 24.555 ;
      RECT  21.3075 25.475 21.4425 25.405 ;
      RECT  21.8675 25.4725 21.925 25.4125 ;
      RECT  21.86 25.54 21.93 23.995 ;
      RECT  22.05 25.415 22.11 25.4725 ;
      RECT  21.34 26.19 21.41 26.325 ;
      RECT  21.525 25.34 21.595 26.885 ;
      RECT  22.0125 25.405 22.1475 25.475 ;
      RECT  22.045 25.34 22.115 26.885 ;
      RECT  21.34 25.34 21.41 26.885 ;
      RECT  21.79 25.6975 21.86 25.8325 ;
      RECT  22.045 25.4075 22.115 26.8175 ;
      RECT  21.595 25.6975 21.665 25.8325 ;
      RECT  21.5325 25.415 21.5875 25.4675 ;
      RECT  21.6875 26.7175 21.7575 26.8525 ;
      RECT  21.345 25.41 21.405 25.4675 ;
      RECT  22.045 26.19 22.115 26.325 ;
      RECT  21.3075 25.405 21.4425 25.475 ;
      RECT  21.8675 25.4075 21.925 25.4675 ;
      RECT  21.86 25.34 21.93 26.885 ;
      RECT  22.05 28.155 22.11 28.0975 ;
      RECT  21.34 27.38 21.41 27.245 ;
      RECT  21.525 28.23 21.595 26.685 ;
      RECT  22.0125 28.165 22.1475 28.095 ;
      RECT  22.045 28.23 22.115 26.685 ;
      RECT  21.34 28.23 21.41 26.685 ;
      RECT  21.79 27.8725 21.86 27.7375 ;
      RECT  22.045 28.1625 22.115 26.7525 ;
      RECT  21.595 27.8725 21.665 27.7375 ;
      RECT  21.5325 28.155 21.5875 28.1025 ;
      RECT  21.6875 26.8525 21.7575 26.7175 ;
      RECT  21.345 28.16 21.405 28.1025 ;
      RECT  22.045 27.38 22.115 27.245 ;
      RECT  21.3075 28.165 21.4425 28.095 ;
      RECT  21.8675 28.1625 21.925 28.1025 ;
      RECT  21.86 28.23 21.93 26.685 ;
      RECT  22.05 28.105 22.11 28.1625 ;
      RECT  21.34 28.88 21.41 29.015 ;
      RECT  21.525 28.03 21.595 29.575 ;
      RECT  22.0125 28.095 22.1475 28.165 ;
      RECT  22.045 28.03 22.115 29.575 ;
      RECT  21.34 28.03 21.41 29.575 ;
      RECT  21.79 28.3875 21.86 28.5225 ;
      RECT  22.045 28.0975 22.115 29.5075 ;
      RECT  21.595 28.3875 21.665 28.5225 ;
      RECT  21.5325 28.105 21.5875 28.1575 ;
      RECT  21.6875 29.4075 21.7575 29.5425 ;
      RECT  21.345 28.1 21.405 28.1575 ;
      RECT  22.045 28.88 22.115 29.015 ;
      RECT  21.3075 28.095 21.4425 28.165 ;
      RECT  21.8675 28.0975 21.925 28.1575 ;
      RECT  21.86 28.03 21.93 29.575 ;
      RECT  22.05 30.845 22.11 30.7875 ;
      RECT  21.34 30.07 21.41 29.935 ;
      RECT  21.525 30.92 21.595 29.375 ;
      RECT  22.0125 30.855 22.1475 30.785 ;
      RECT  22.045 30.92 22.115 29.375 ;
      RECT  21.34 30.92 21.41 29.375 ;
      RECT  21.79 30.5625 21.86 30.4275 ;
      RECT  22.045 30.8525 22.115 29.4425 ;
      RECT  21.595 30.5625 21.665 30.4275 ;
      RECT  21.5325 30.845 21.5875 30.7925 ;
      RECT  21.6875 29.5425 21.7575 29.4075 ;
      RECT  21.345 30.85 21.405 30.7925 ;
      RECT  22.045 30.07 22.115 29.935 ;
      RECT  21.3075 30.855 21.4425 30.785 ;
      RECT  21.8675 30.8525 21.925 30.7925 ;
      RECT  21.86 30.92 21.93 29.375 ;
      RECT  22.05 30.795 22.11 30.8525 ;
      RECT  21.34 31.57 21.41 31.705 ;
      RECT  21.525 30.72 21.595 32.265 ;
      RECT  22.0125 30.785 22.1475 30.855 ;
      RECT  22.045 30.72 22.115 32.265 ;
      RECT  21.34 30.72 21.41 32.265 ;
      RECT  21.79 31.0775 21.86 31.2125 ;
      RECT  22.045 30.7875 22.115 32.1975 ;
      RECT  21.595 31.0775 21.665 31.2125 ;
      RECT  21.5325 30.795 21.5875 30.8475 ;
      RECT  21.6875 32.0975 21.7575 32.2325 ;
      RECT  21.345 30.79 21.405 30.8475 ;
      RECT  22.045 31.57 22.115 31.705 ;
      RECT  21.3075 30.785 21.4425 30.855 ;
      RECT  21.8675 30.7875 21.925 30.8475 ;
      RECT  21.86 30.72 21.93 32.265 ;
      RECT  22.05 33.535 22.11 33.4775 ;
      RECT  21.34 32.76 21.41 32.625 ;
      RECT  21.525 33.61 21.595 32.065 ;
      RECT  22.0125 33.545 22.1475 33.475 ;
      RECT  22.045 33.61 22.115 32.065 ;
      RECT  21.34 33.61 21.41 32.065 ;
      RECT  21.79 33.2525 21.86 33.1175 ;
      RECT  22.045 33.5425 22.115 32.1325 ;
      RECT  21.595 33.2525 21.665 33.1175 ;
      RECT  21.5325 33.535 21.5875 33.4825 ;
      RECT  21.6875 32.2325 21.7575 32.0975 ;
      RECT  21.345 33.54 21.405 33.4825 ;
      RECT  22.045 32.76 22.115 32.625 ;
      RECT  21.3075 33.545 21.4425 33.475 ;
      RECT  21.8675 33.5425 21.925 33.4825 ;
      RECT  21.86 33.61 21.93 32.065 ;
      RECT  22.05 33.485 22.11 33.5425 ;
      RECT  21.34 34.26 21.41 34.395 ;
      RECT  21.525 33.41 21.595 34.955 ;
      RECT  22.0125 33.475 22.1475 33.545 ;
      RECT  22.045 33.41 22.115 34.955 ;
      RECT  21.34 33.41 21.41 34.955 ;
      RECT  21.79 33.7675 21.86 33.9025 ;
      RECT  22.045 33.4775 22.115 34.8875 ;
      RECT  21.595 33.7675 21.665 33.9025 ;
      RECT  21.5325 33.485 21.5875 33.5375 ;
      RECT  21.6875 34.7875 21.7575 34.9225 ;
      RECT  21.345 33.48 21.405 33.5375 ;
      RECT  22.045 34.26 22.115 34.395 ;
      RECT  21.3075 33.475 21.4425 33.545 ;
      RECT  21.8675 33.4775 21.925 33.5375 ;
      RECT  21.86 33.41 21.93 34.955 ;
      RECT  22.05 36.225 22.11 36.1675 ;
      RECT  21.34 35.45 21.41 35.315 ;
      RECT  21.525 36.3 21.595 34.755 ;
      RECT  22.0125 36.235 22.1475 36.165 ;
      RECT  22.045 36.3 22.115 34.755 ;
      RECT  21.34 36.3 21.41 34.755 ;
      RECT  21.79 35.9425 21.86 35.8075 ;
      RECT  22.045 36.2325 22.115 34.8225 ;
      RECT  21.595 35.9425 21.665 35.8075 ;
      RECT  21.5325 36.225 21.5875 36.1725 ;
      RECT  21.6875 34.9225 21.7575 34.7875 ;
      RECT  21.345 36.23 21.405 36.1725 ;
      RECT  22.045 35.45 22.115 35.315 ;
      RECT  21.3075 36.235 21.4425 36.165 ;
      RECT  21.8675 36.2325 21.925 36.1725 ;
      RECT  21.86 36.3 21.93 34.755 ;
      RECT  22.05 36.175 22.11 36.2325 ;
      RECT  21.34 36.95 21.41 37.085 ;
      RECT  21.525 36.1 21.595 37.645 ;
      RECT  22.0125 36.165 22.1475 36.235 ;
      RECT  22.045 36.1 22.115 37.645 ;
      RECT  21.34 36.1 21.41 37.645 ;
      RECT  21.79 36.4575 21.86 36.5925 ;
      RECT  22.045 36.1675 22.115 37.5775 ;
      RECT  21.595 36.4575 21.665 36.5925 ;
      RECT  21.5325 36.175 21.5875 36.2275 ;
      RECT  21.6875 37.4775 21.7575 37.6125 ;
      RECT  21.345 36.17 21.405 36.2275 ;
      RECT  22.045 36.95 22.115 37.085 ;
      RECT  21.3075 36.165 21.4425 36.235 ;
      RECT  21.8675 36.1675 21.925 36.2275 ;
      RECT  21.86 36.1 21.93 37.645 ;
      RECT  22.05 38.915 22.11 38.8575 ;
      RECT  21.34 38.14 21.41 38.005 ;
      RECT  21.525 38.99 21.595 37.445 ;
      RECT  22.0125 38.925 22.1475 38.855 ;
      RECT  22.045 38.99 22.115 37.445 ;
      RECT  21.34 38.99 21.41 37.445 ;
      RECT  21.79 38.6325 21.86 38.4975 ;
      RECT  22.045 38.9225 22.115 37.5125 ;
      RECT  21.595 38.6325 21.665 38.4975 ;
      RECT  21.5325 38.915 21.5875 38.8625 ;
      RECT  21.6875 37.6125 21.7575 37.4775 ;
      RECT  21.345 38.92 21.405 38.8625 ;
      RECT  22.045 38.14 22.115 38.005 ;
      RECT  21.3075 38.925 21.4425 38.855 ;
      RECT  21.8675 38.9225 21.925 38.8625 ;
      RECT  21.86 38.99 21.93 37.445 ;
      RECT  22.05 38.865 22.11 38.9225 ;
      RECT  21.34 39.64 21.41 39.775 ;
      RECT  21.525 38.79 21.595 40.335 ;
      RECT  22.0125 38.855 22.1475 38.925 ;
      RECT  22.045 38.79 22.115 40.335 ;
      RECT  21.34 38.79 21.41 40.335 ;
      RECT  21.79 39.1475 21.86 39.2825 ;
      RECT  22.045 38.8575 22.115 40.2675 ;
      RECT  21.595 39.1475 21.665 39.2825 ;
      RECT  21.5325 38.865 21.5875 38.9175 ;
      RECT  21.6875 40.1675 21.7575 40.3025 ;
      RECT  21.345 38.86 21.405 38.9175 ;
      RECT  22.045 39.64 22.115 39.775 ;
      RECT  21.3075 38.855 21.4425 38.925 ;
      RECT  21.8675 38.8575 21.925 38.9175 ;
      RECT  21.86 38.79 21.93 40.335 ;
      RECT  22.05 41.605 22.11 41.5475 ;
      RECT  21.34 40.83 21.41 40.695 ;
      RECT  21.525 41.68 21.595 40.135 ;
      RECT  22.0125 41.615 22.1475 41.545 ;
      RECT  22.045 41.68 22.115 40.135 ;
      RECT  21.34 41.68 21.41 40.135 ;
      RECT  21.79 41.3225 21.86 41.1875 ;
      RECT  22.045 41.6125 22.115 40.2025 ;
      RECT  21.595 41.3225 21.665 41.1875 ;
      RECT  21.5325 41.605 21.5875 41.5525 ;
      RECT  21.6875 40.3025 21.7575 40.1675 ;
      RECT  21.345 41.61 21.405 41.5525 ;
      RECT  22.045 40.83 22.115 40.695 ;
      RECT  21.3075 41.615 21.4425 41.545 ;
      RECT  21.8675 41.6125 21.925 41.5525 ;
      RECT  21.86 41.68 21.93 40.135 ;
      RECT  22.05 41.555 22.11 41.6125 ;
      RECT  21.34 42.33 21.41 42.465 ;
      RECT  21.525 41.48 21.595 43.025 ;
      RECT  22.0125 41.545 22.1475 41.615 ;
      RECT  22.045 41.48 22.115 43.025 ;
      RECT  21.34 41.48 21.41 43.025 ;
      RECT  21.79 41.8375 21.86 41.9725 ;
      RECT  22.045 41.5475 22.115 42.9575 ;
      RECT  21.595 41.8375 21.665 41.9725 ;
      RECT  21.5325 41.555 21.5875 41.6075 ;
      RECT  21.6875 42.8575 21.7575 42.9925 ;
      RECT  21.345 41.55 21.405 41.6075 ;
      RECT  22.045 42.33 22.115 42.465 ;
      RECT  21.3075 41.545 21.4425 41.615 ;
      RECT  21.8675 41.5475 21.925 41.6075 ;
      RECT  21.86 41.48 21.93 43.025 ;
      RECT  22.05 44.295 22.11 44.2375 ;
      RECT  21.34 43.52 21.41 43.385 ;
      RECT  21.525 44.37 21.595 42.825 ;
      RECT  22.0125 44.305 22.1475 44.235 ;
      RECT  22.045 44.37 22.115 42.825 ;
      RECT  21.34 44.37 21.41 42.825 ;
      RECT  21.79 44.0125 21.86 43.8775 ;
      RECT  22.045 44.3025 22.115 42.8925 ;
      RECT  21.595 44.0125 21.665 43.8775 ;
      RECT  21.5325 44.295 21.5875 44.2425 ;
      RECT  21.6875 42.9925 21.7575 42.8575 ;
      RECT  21.345 44.3 21.405 44.2425 ;
      RECT  22.045 43.52 22.115 43.385 ;
      RECT  21.3075 44.305 21.4425 44.235 ;
      RECT  21.8675 44.3025 21.925 44.2425 ;
      RECT  21.86 44.37 21.93 42.825 ;
      RECT  22.755 22.725 22.815 22.7825 ;
      RECT  22.045 23.5 22.115 23.635 ;
      RECT  22.23 22.65 22.3 24.195 ;
      RECT  22.7175 22.715 22.8525 22.785 ;
      RECT  22.75 22.65 22.82 24.195 ;
      RECT  22.045 22.65 22.115 24.195 ;
      RECT  22.495 23.0075 22.565 23.1425 ;
      RECT  22.75 22.7175 22.82 24.1275 ;
      RECT  22.3 23.0075 22.37 23.1425 ;
      RECT  22.2375 22.725 22.2925 22.7775 ;
      RECT  22.3925 24.0275 22.4625 24.1625 ;
      RECT  22.05 22.72 22.11 22.7775 ;
      RECT  22.75 23.5 22.82 23.635 ;
      RECT  22.0125 22.715 22.1475 22.785 ;
      RECT  22.5725 22.7175 22.63 22.7775 ;
      RECT  22.565 22.65 22.635 24.195 ;
      RECT  22.755 25.465 22.815 25.4075 ;
      RECT  22.045 24.69 22.115 24.555 ;
      RECT  22.23 25.54 22.3 23.995 ;
      RECT  22.7175 25.475 22.8525 25.405 ;
      RECT  22.75 25.54 22.82 23.995 ;
      RECT  22.045 25.54 22.115 23.995 ;
      RECT  22.495 25.1825 22.565 25.0475 ;
      RECT  22.75 25.4725 22.82 24.0625 ;
      RECT  22.3 25.1825 22.37 25.0475 ;
      RECT  22.2375 25.465 22.2925 25.4125 ;
      RECT  22.3925 24.1625 22.4625 24.0275 ;
      RECT  22.05 25.47 22.11 25.4125 ;
      RECT  22.75 24.69 22.82 24.555 ;
      RECT  22.0125 25.475 22.1475 25.405 ;
      RECT  22.5725 25.4725 22.63 25.4125 ;
      RECT  22.565 25.54 22.635 23.995 ;
      RECT  22.755 25.415 22.815 25.4725 ;
      RECT  22.045 26.19 22.115 26.325 ;
      RECT  22.23 25.34 22.3 26.885 ;
      RECT  22.7175 25.405 22.8525 25.475 ;
      RECT  22.75 25.34 22.82 26.885 ;
      RECT  22.045 25.34 22.115 26.885 ;
      RECT  22.495 25.6975 22.565 25.8325 ;
      RECT  22.75 25.4075 22.82 26.8175 ;
      RECT  22.3 25.6975 22.37 25.8325 ;
      RECT  22.2375 25.415 22.2925 25.4675 ;
      RECT  22.3925 26.7175 22.4625 26.8525 ;
      RECT  22.05 25.41 22.11 25.4675 ;
      RECT  22.75 26.19 22.82 26.325 ;
      RECT  22.0125 25.405 22.1475 25.475 ;
      RECT  22.5725 25.4075 22.63 25.4675 ;
      RECT  22.565 25.34 22.635 26.885 ;
      RECT  22.755 28.155 22.815 28.0975 ;
      RECT  22.045 27.38 22.115 27.245 ;
      RECT  22.23 28.23 22.3 26.685 ;
      RECT  22.7175 28.165 22.8525 28.095 ;
      RECT  22.75 28.23 22.82 26.685 ;
      RECT  22.045 28.23 22.115 26.685 ;
      RECT  22.495 27.8725 22.565 27.7375 ;
      RECT  22.75 28.1625 22.82 26.7525 ;
      RECT  22.3 27.8725 22.37 27.7375 ;
      RECT  22.2375 28.155 22.2925 28.1025 ;
      RECT  22.3925 26.8525 22.4625 26.7175 ;
      RECT  22.05 28.16 22.11 28.1025 ;
      RECT  22.75 27.38 22.82 27.245 ;
      RECT  22.0125 28.165 22.1475 28.095 ;
      RECT  22.5725 28.1625 22.63 28.1025 ;
      RECT  22.565 28.23 22.635 26.685 ;
      RECT  22.755 28.105 22.815 28.1625 ;
      RECT  22.045 28.88 22.115 29.015 ;
      RECT  22.23 28.03 22.3 29.575 ;
      RECT  22.7175 28.095 22.8525 28.165 ;
      RECT  22.75 28.03 22.82 29.575 ;
      RECT  22.045 28.03 22.115 29.575 ;
      RECT  22.495 28.3875 22.565 28.5225 ;
      RECT  22.75 28.0975 22.82 29.5075 ;
      RECT  22.3 28.3875 22.37 28.5225 ;
      RECT  22.2375 28.105 22.2925 28.1575 ;
      RECT  22.3925 29.4075 22.4625 29.5425 ;
      RECT  22.05 28.1 22.11 28.1575 ;
      RECT  22.75 28.88 22.82 29.015 ;
      RECT  22.0125 28.095 22.1475 28.165 ;
      RECT  22.5725 28.0975 22.63 28.1575 ;
      RECT  22.565 28.03 22.635 29.575 ;
      RECT  22.755 30.845 22.815 30.7875 ;
      RECT  22.045 30.07 22.115 29.935 ;
      RECT  22.23 30.92 22.3 29.375 ;
      RECT  22.7175 30.855 22.8525 30.785 ;
      RECT  22.75 30.92 22.82 29.375 ;
      RECT  22.045 30.92 22.115 29.375 ;
      RECT  22.495 30.5625 22.565 30.4275 ;
      RECT  22.75 30.8525 22.82 29.4425 ;
      RECT  22.3 30.5625 22.37 30.4275 ;
      RECT  22.2375 30.845 22.2925 30.7925 ;
      RECT  22.3925 29.5425 22.4625 29.4075 ;
      RECT  22.05 30.85 22.11 30.7925 ;
      RECT  22.75 30.07 22.82 29.935 ;
      RECT  22.0125 30.855 22.1475 30.785 ;
      RECT  22.5725 30.8525 22.63 30.7925 ;
      RECT  22.565 30.92 22.635 29.375 ;
      RECT  22.755 30.795 22.815 30.8525 ;
      RECT  22.045 31.57 22.115 31.705 ;
      RECT  22.23 30.72 22.3 32.265 ;
      RECT  22.7175 30.785 22.8525 30.855 ;
      RECT  22.75 30.72 22.82 32.265 ;
      RECT  22.045 30.72 22.115 32.265 ;
      RECT  22.495 31.0775 22.565 31.2125 ;
      RECT  22.75 30.7875 22.82 32.1975 ;
      RECT  22.3 31.0775 22.37 31.2125 ;
      RECT  22.2375 30.795 22.2925 30.8475 ;
      RECT  22.3925 32.0975 22.4625 32.2325 ;
      RECT  22.05 30.79 22.11 30.8475 ;
      RECT  22.75 31.57 22.82 31.705 ;
      RECT  22.0125 30.785 22.1475 30.855 ;
      RECT  22.5725 30.7875 22.63 30.8475 ;
      RECT  22.565 30.72 22.635 32.265 ;
      RECT  22.755 33.535 22.815 33.4775 ;
      RECT  22.045 32.76 22.115 32.625 ;
      RECT  22.23 33.61 22.3 32.065 ;
      RECT  22.7175 33.545 22.8525 33.475 ;
      RECT  22.75 33.61 22.82 32.065 ;
      RECT  22.045 33.61 22.115 32.065 ;
      RECT  22.495 33.2525 22.565 33.1175 ;
      RECT  22.75 33.5425 22.82 32.1325 ;
      RECT  22.3 33.2525 22.37 33.1175 ;
      RECT  22.2375 33.535 22.2925 33.4825 ;
      RECT  22.3925 32.2325 22.4625 32.0975 ;
      RECT  22.05 33.54 22.11 33.4825 ;
      RECT  22.75 32.76 22.82 32.625 ;
      RECT  22.0125 33.545 22.1475 33.475 ;
      RECT  22.5725 33.5425 22.63 33.4825 ;
      RECT  22.565 33.61 22.635 32.065 ;
      RECT  22.755 33.485 22.815 33.5425 ;
      RECT  22.045 34.26 22.115 34.395 ;
      RECT  22.23 33.41 22.3 34.955 ;
      RECT  22.7175 33.475 22.8525 33.545 ;
      RECT  22.75 33.41 22.82 34.955 ;
      RECT  22.045 33.41 22.115 34.955 ;
      RECT  22.495 33.7675 22.565 33.9025 ;
      RECT  22.75 33.4775 22.82 34.8875 ;
      RECT  22.3 33.7675 22.37 33.9025 ;
      RECT  22.2375 33.485 22.2925 33.5375 ;
      RECT  22.3925 34.7875 22.4625 34.9225 ;
      RECT  22.05 33.48 22.11 33.5375 ;
      RECT  22.75 34.26 22.82 34.395 ;
      RECT  22.0125 33.475 22.1475 33.545 ;
      RECT  22.5725 33.4775 22.63 33.5375 ;
      RECT  22.565 33.41 22.635 34.955 ;
      RECT  22.755 36.225 22.815 36.1675 ;
      RECT  22.045 35.45 22.115 35.315 ;
      RECT  22.23 36.3 22.3 34.755 ;
      RECT  22.7175 36.235 22.8525 36.165 ;
      RECT  22.75 36.3 22.82 34.755 ;
      RECT  22.045 36.3 22.115 34.755 ;
      RECT  22.495 35.9425 22.565 35.8075 ;
      RECT  22.75 36.2325 22.82 34.8225 ;
      RECT  22.3 35.9425 22.37 35.8075 ;
      RECT  22.2375 36.225 22.2925 36.1725 ;
      RECT  22.3925 34.9225 22.4625 34.7875 ;
      RECT  22.05 36.23 22.11 36.1725 ;
      RECT  22.75 35.45 22.82 35.315 ;
      RECT  22.0125 36.235 22.1475 36.165 ;
      RECT  22.5725 36.2325 22.63 36.1725 ;
      RECT  22.565 36.3 22.635 34.755 ;
      RECT  22.755 36.175 22.815 36.2325 ;
      RECT  22.045 36.95 22.115 37.085 ;
      RECT  22.23 36.1 22.3 37.645 ;
      RECT  22.7175 36.165 22.8525 36.235 ;
      RECT  22.75 36.1 22.82 37.645 ;
      RECT  22.045 36.1 22.115 37.645 ;
      RECT  22.495 36.4575 22.565 36.5925 ;
      RECT  22.75 36.1675 22.82 37.5775 ;
      RECT  22.3 36.4575 22.37 36.5925 ;
      RECT  22.2375 36.175 22.2925 36.2275 ;
      RECT  22.3925 37.4775 22.4625 37.6125 ;
      RECT  22.05 36.17 22.11 36.2275 ;
      RECT  22.75 36.95 22.82 37.085 ;
      RECT  22.0125 36.165 22.1475 36.235 ;
      RECT  22.5725 36.1675 22.63 36.2275 ;
      RECT  22.565 36.1 22.635 37.645 ;
      RECT  22.755 38.915 22.815 38.8575 ;
      RECT  22.045 38.14 22.115 38.005 ;
      RECT  22.23 38.99 22.3 37.445 ;
      RECT  22.7175 38.925 22.8525 38.855 ;
      RECT  22.75 38.99 22.82 37.445 ;
      RECT  22.045 38.99 22.115 37.445 ;
      RECT  22.495 38.6325 22.565 38.4975 ;
      RECT  22.75 38.9225 22.82 37.5125 ;
      RECT  22.3 38.6325 22.37 38.4975 ;
      RECT  22.2375 38.915 22.2925 38.8625 ;
      RECT  22.3925 37.6125 22.4625 37.4775 ;
      RECT  22.05 38.92 22.11 38.8625 ;
      RECT  22.75 38.14 22.82 38.005 ;
      RECT  22.0125 38.925 22.1475 38.855 ;
      RECT  22.5725 38.9225 22.63 38.8625 ;
      RECT  22.565 38.99 22.635 37.445 ;
      RECT  22.755 38.865 22.815 38.9225 ;
      RECT  22.045 39.64 22.115 39.775 ;
      RECT  22.23 38.79 22.3 40.335 ;
      RECT  22.7175 38.855 22.8525 38.925 ;
      RECT  22.75 38.79 22.82 40.335 ;
      RECT  22.045 38.79 22.115 40.335 ;
      RECT  22.495 39.1475 22.565 39.2825 ;
      RECT  22.75 38.8575 22.82 40.2675 ;
      RECT  22.3 39.1475 22.37 39.2825 ;
      RECT  22.2375 38.865 22.2925 38.9175 ;
      RECT  22.3925 40.1675 22.4625 40.3025 ;
      RECT  22.05 38.86 22.11 38.9175 ;
      RECT  22.75 39.64 22.82 39.775 ;
      RECT  22.0125 38.855 22.1475 38.925 ;
      RECT  22.5725 38.8575 22.63 38.9175 ;
      RECT  22.565 38.79 22.635 40.335 ;
      RECT  22.755 41.605 22.815 41.5475 ;
      RECT  22.045 40.83 22.115 40.695 ;
      RECT  22.23 41.68 22.3 40.135 ;
      RECT  22.7175 41.615 22.8525 41.545 ;
      RECT  22.75 41.68 22.82 40.135 ;
      RECT  22.045 41.68 22.115 40.135 ;
      RECT  22.495 41.3225 22.565 41.1875 ;
      RECT  22.75 41.6125 22.82 40.2025 ;
      RECT  22.3 41.3225 22.37 41.1875 ;
      RECT  22.2375 41.605 22.2925 41.5525 ;
      RECT  22.3925 40.3025 22.4625 40.1675 ;
      RECT  22.05 41.61 22.11 41.5525 ;
      RECT  22.75 40.83 22.82 40.695 ;
      RECT  22.0125 41.615 22.1475 41.545 ;
      RECT  22.5725 41.6125 22.63 41.5525 ;
      RECT  22.565 41.68 22.635 40.135 ;
      RECT  22.755 41.555 22.815 41.6125 ;
      RECT  22.045 42.33 22.115 42.465 ;
      RECT  22.23 41.48 22.3 43.025 ;
      RECT  22.7175 41.545 22.8525 41.615 ;
      RECT  22.75 41.48 22.82 43.025 ;
      RECT  22.045 41.48 22.115 43.025 ;
      RECT  22.495 41.8375 22.565 41.9725 ;
      RECT  22.75 41.5475 22.82 42.9575 ;
      RECT  22.3 41.8375 22.37 41.9725 ;
      RECT  22.2375 41.555 22.2925 41.6075 ;
      RECT  22.3925 42.8575 22.4625 42.9925 ;
      RECT  22.05 41.55 22.11 41.6075 ;
      RECT  22.75 42.33 22.82 42.465 ;
      RECT  22.0125 41.545 22.1475 41.615 ;
      RECT  22.5725 41.5475 22.63 41.6075 ;
      RECT  22.565 41.48 22.635 43.025 ;
      RECT  22.755 44.295 22.815 44.2375 ;
      RECT  22.045 43.52 22.115 43.385 ;
      RECT  22.23 44.37 22.3 42.825 ;
      RECT  22.7175 44.305 22.8525 44.235 ;
      RECT  22.75 44.37 22.82 42.825 ;
      RECT  22.045 44.37 22.115 42.825 ;
      RECT  22.495 44.0125 22.565 43.8775 ;
      RECT  22.75 44.3025 22.82 42.8925 ;
      RECT  22.3 44.0125 22.37 43.8775 ;
      RECT  22.2375 44.295 22.2925 44.2425 ;
      RECT  22.3925 42.9925 22.4625 42.8575 ;
      RECT  22.05 44.3 22.11 44.2425 ;
      RECT  22.75 43.52 22.82 43.385 ;
      RECT  22.0125 44.305 22.1475 44.235 ;
      RECT  22.5725 44.3025 22.63 44.2425 ;
      RECT  22.565 44.37 22.635 42.825 ;
      RECT  21.525 22.75 21.595 44.27 ;
      RECT  21.86 22.75 21.93 44.27 ;
      RECT  22.23 22.75 22.3 44.27 ;
      RECT  22.565 22.75 22.635 44.27 ;
      RECT  21.6875 32.0975 21.7575 32.2325 ;
      RECT  22.3925 34.7875 22.4625 34.9225 ;
      RECT  22.3925 34.7875 22.4625 34.9225 ;
      RECT  21.6875 24.0275 21.7575 24.1625 ;
      RECT  21.6875 24.0275 21.7575 24.1625 ;
      RECT  21.6875 40.1675 21.7575 40.3025 ;
      RECT  22.3925 42.8575 22.4625 42.9925 ;
      RECT  22.3925 42.8575 22.4625 42.9925 ;
      RECT  22.3925 26.7175 22.4625 26.8525 ;
      RECT  22.3925 26.7175 22.4625 26.8525 ;
      RECT  21.6875 37.4775 21.7575 37.6125 ;
      RECT  21.6875 34.7875 21.7575 34.9225 ;
      RECT  21.6875 34.7875 21.7575 34.9225 ;
      RECT  21.6875 42.8575 21.7575 42.9925 ;
      RECT  21.6875 42.8575 21.7575 42.9925 ;
      RECT  21.6875 26.7175 21.7575 26.8525 ;
      RECT  21.6875 26.7175 21.7575 26.8525 ;
      RECT  22.3925 37.4775 22.4625 37.6125 ;
      RECT  22.3925 29.4075 22.4625 29.5425 ;
      RECT  22.3925 29.4075 22.4625 29.5425 ;
      RECT  22.3925 40.1675 22.4625 40.3025 ;
      RECT  22.3925 24.0275 22.4625 24.1625 ;
      RECT  22.3925 24.0275 22.4625 24.1625 ;
      RECT  22.3925 32.0975 22.4625 32.2325 ;
      RECT  21.6875 29.4075 21.7575 29.5425 ;
      RECT  21.6875 29.4075 21.7575 29.5425 ;
      RECT  22.0125 22.715 22.1475 22.785 ;
      RECT  21.3075 44.235 21.4425 44.305 ;
      RECT  21.3075 33.475 21.4425 33.545 ;
      RECT  21.3075 38.855 21.4425 38.925 ;
      RECT  22.0125 38.855 22.1475 38.925 ;
      RECT  21.3075 41.545 21.4425 41.615 ;
      RECT  22.0125 36.165 22.1475 36.235 ;
      RECT  21.3075 22.715 21.4425 22.785 ;
      RECT  22.0125 25.405 22.1475 25.475 ;
      RECT  21.3075 30.785 21.4425 30.855 ;
      RECT  22.0125 41.545 22.1475 41.615 ;
      RECT  21.3075 25.405 21.4425 25.475 ;
      RECT  22.0125 28.095 22.1475 28.165 ;
      RECT  21.3075 36.165 21.4425 36.235 ;
      RECT  22.0125 33.475 22.1475 33.545 ;
      RECT  22.0125 30.785 22.1475 30.855 ;
      RECT  21.3075 28.095 21.4425 28.165 ;
      RECT  22.0125 44.235 22.1475 44.305 ;
      RECT  21.345 20.035 21.405 20.0925 ;
      RECT  20.635 20.81 20.705 20.945 ;
      RECT  20.82 19.96 20.89 21.505 ;
      RECT  21.3075 20.025 21.4425 20.095 ;
      RECT  21.34 19.96 21.41 21.505 ;
      RECT  20.635 19.96 20.705 21.505 ;
      RECT  21.085 20.3175 21.155 20.4525 ;
      RECT  21.34 20.0275 21.41 21.4375 ;
      RECT  20.89 20.3175 20.96 20.4525 ;
      RECT  20.8275 20.035 20.8825 20.0875 ;
      RECT  20.9825 21.3375 21.0525 21.4725 ;
      RECT  20.64 20.03 20.7 20.0875 ;
      RECT  21.34 20.81 21.41 20.945 ;
      RECT  20.6025 20.025 20.7375 20.095 ;
      RECT  21.1625 20.0275 21.22 20.0875 ;
      RECT  21.155 19.96 21.225 21.505 ;
      RECT  21.345 22.775 21.405 22.7175 ;
      RECT  20.82 22.85 20.89 21.305 ;
      RECT  21.34 22.85 21.41 21.305 ;
      RECT  21.3075 22.785 21.4425 22.715 ;
      RECT  20.635 22.0 20.705 21.865 ;
      RECT  21.34 22.0 21.41 21.865 ;
      RECT  21.085 22.4925 21.155 22.3575 ;
      RECT  21.34 22.7825 21.41 21.3725 ;
      RECT  20.89 22.4925 20.96 22.3575 ;
      RECT  20.8275 22.775 20.8825 22.7225 ;
      RECT  20.6025 22.785 20.7375 22.715 ;
      RECT  20.64 22.78 20.7 22.7225 ;
      RECT  20.635 22.85 20.705 21.305 ;
      RECT  20.9825 21.4725 21.0525 21.3375 ;
      RECT  21.1625 22.7825 21.22 22.7225 ;
      RECT  21.155 22.85 21.225 21.305 ;
      RECT  21.345 22.725 21.405 22.7825 ;
      RECT  20.82 22.65 20.89 24.195 ;
      RECT  21.34 22.65 21.41 24.195 ;
      RECT  21.3075 22.715 21.4425 22.785 ;
      RECT  20.635 23.5 20.705 23.635 ;
      RECT  21.34 23.5 21.41 23.635 ;
      RECT  21.085 23.0075 21.155 23.1425 ;
      RECT  21.34 22.7175 21.41 24.1275 ;
      RECT  20.89 23.0075 20.96 23.1425 ;
      RECT  20.8275 22.725 20.8825 22.7775 ;
      RECT  20.6025 22.715 20.7375 22.785 ;
      RECT  20.64 22.72 20.7 22.7775 ;
      RECT  20.635 22.65 20.705 24.195 ;
      RECT  20.9825 24.0275 21.0525 24.1625 ;
      RECT  21.1625 22.7175 21.22 22.7775 ;
      RECT  21.155 22.65 21.225 24.195 ;
      RECT  21.345 25.465 21.405 25.4075 ;
      RECT  20.82 25.54 20.89 23.995 ;
      RECT  21.34 25.54 21.41 23.995 ;
      RECT  21.3075 25.475 21.4425 25.405 ;
      RECT  20.635 24.69 20.705 24.555 ;
      RECT  21.34 24.69 21.41 24.555 ;
      RECT  21.085 25.1825 21.155 25.0475 ;
      RECT  21.34 25.4725 21.41 24.0625 ;
      RECT  20.89 25.1825 20.96 25.0475 ;
      RECT  20.8275 25.465 20.8825 25.4125 ;
      RECT  20.6025 25.475 20.7375 25.405 ;
      RECT  20.64 25.47 20.7 25.4125 ;
      RECT  20.635 25.54 20.705 23.995 ;
      RECT  20.9825 24.1625 21.0525 24.0275 ;
      RECT  21.1625 25.4725 21.22 25.4125 ;
      RECT  21.155 25.54 21.225 23.995 ;
      RECT  21.345 25.415 21.405 25.4725 ;
      RECT  20.82 25.34 20.89 26.885 ;
      RECT  21.34 25.34 21.41 26.885 ;
      RECT  21.3075 25.405 21.4425 25.475 ;
      RECT  20.635 26.19 20.705 26.325 ;
      RECT  21.34 26.19 21.41 26.325 ;
      RECT  21.085 25.6975 21.155 25.8325 ;
      RECT  21.34 25.4075 21.41 26.8175 ;
      RECT  20.89 25.6975 20.96 25.8325 ;
      RECT  20.8275 25.415 20.8825 25.4675 ;
      RECT  20.6025 25.405 20.7375 25.475 ;
      RECT  20.64 25.41 20.7 25.4675 ;
      RECT  20.635 25.34 20.705 26.885 ;
      RECT  20.9825 26.7175 21.0525 26.8525 ;
      RECT  21.1625 25.4075 21.22 25.4675 ;
      RECT  21.155 25.34 21.225 26.885 ;
      RECT  21.345 28.155 21.405 28.0975 ;
      RECT  20.82 28.23 20.89 26.685 ;
      RECT  21.34 28.23 21.41 26.685 ;
      RECT  21.3075 28.165 21.4425 28.095 ;
      RECT  20.635 27.38 20.705 27.245 ;
      RECT  21.34 27.38 21.41 27.245 ;
      RECT  21.085 27.8725 21.155 27.7375 ;
      RECT  21.34 28.1625 21.41 26.7525 ;
      RECT  20.89 27.8725 20.96 27.7375 ;
      RECT  20.8275 28.155 20.8825 28.1025 ;
      RECT  20.6025 28.165 20.7375 28.095 ;
      RECT  20.64 28.16 20.7 28.1025 ;
      RECT  20.635 28.23 20.705 26.685 ;
      RECT  20.9825 26.8525 21.0525 26.7175 ;
      RECT  21.1625 28.1625 21.22 28.1025 ;
      RECT  21.155 28.23 21.225 26.685 ;
      RECT  21.345 28.105 21.405 28.1625 ;
      RECT  20.82 28.03 20.89 29.575 ;
      RECT  21.34 28.03 21.41 29.575 ;
      RECT  21.3075 28.095 21.4425 28.165 ;
      RECT  20.635 28.88 20.705 29.015 ;
      RECT  21.34 28.88 21.41 29.015 ;
      RECT  21.085 28.3875 21.155 28.5225 ;
      RECT  21.34 28.0975 21.41 29.5075 ;
      RECT  20.89 28.3875 20.96 28.5225 ;
      RECT  20.8275 28.105 20.8825 28.1575 ;
      RECT  20.6025 28.095 20.7375 28.165 ;
      RECT  20.64 28.1 20.7 28.1575 ;
      RECT  20.635 28.03 20.705 29.575 ;
      RECT  20.9825 29.4075 21.0525 29.5425 ;
      RECT  21.1625 28.0975 21.22 28.1575 ;
      RECT  21.155 28.03 21.225 29.575 ;
      RECT  21.345 30.845 21.405 30.7875 ;
      RECT  20.82 30.92 20.89 29.375 ;
      RECT  21.34 30.92 21.41 29.375 ;
      RECT  21.3075 30.855 21.4425 30.785 ;
      RECT  20.635 30.07 20.705 29.935 ;
      RECT  21.34 30.07 21.41 29.935 ;
      RECT  21.085 30.5625 21.155 30.4275 ;
      RECT  21.34 30.8525 21.41 29.4425 ;
      RECT  20.89 30.5625 20.96 30.4275 ;
      RECT  20.8275 30.845 20.8825 30.7925 ;
      RECT  20.6025 30.855 20.7375 30.785 ;
      RECT  20.64 30.85 20.7 30.7925 ;
      RECT  20.635 30.92 20.705 29.375 ;
      RECT  20.9825 29.5425 21.0525 29.4075 ;
      RECT  21.1625 30.8525 21.22 30.7925 ;
      RECT  21.155 30.92 21.225 29.375 ;
      RECT  21.345 30.795 21.405 30.8525 ;
      RECT  20.82 30.72 20.89 32.265 ;
      RECT  21.34 30.72 21.41 32.265 ;
      RECT  21.3075 30.785 21.4425 30.855 ;
      RECT  20.635 31.57 20.705 31.705 ;
      RECT  21.34 31.57 21.41 31.705 ;
      RECT  21.085 31.0775 21.155 31.2125 ;
      RECT  21.34 30.7875 21.41 32.1975 ;
      RECT  20.89 31.0775 20.96 31.2125 ;
      RECT  20.8275 30.795 20.8825 30.8475 ;
      RECT  20.6025 30.785 20.7375 30.855 ;
      RECT  20.64 30.79 20.7 30.8475 ;
      RECT  20.635 30.72 20.705 32.265 ;
      RECT  20.9825 32.0975 21.0525 32.2325 ;
      RECT  21.1625 30.7875 21.22 30.8475 ;
      RECT  21.155 30.72 21.225 32.265 ;
      RECT  21.345 33.535 21.405 33.4775 ;
      RECT  20.82 33.61 20.89 32.065 ;
      RECT  21.34 33.61 21.41 32.065 ;
      RECT  21.3075 33.545 21.4425 33.475 ;
      RECT  20.635 32.76 20.705 32.625 ;
      RECT  21.34 32.76 21.41 32.625 ;
      RECT  21.085 33.2525 21.155 33.1175 ;
      RECT  21.34 33.5425 21.41 32.1325 ;
      RECT  20.89 33.2525 20.96 33.1175 ;
      RECT  20.8275 33.535 20.8825 33.4825 ;
      RECT  20.6025 33.545 20.7375 33.475 ;
      RECT  20.64 33.54 20.7 33.4825 ;
      RECT  20.635 33.61 20.705 32.065 ;
      RECT  20.9825 32.2325 21.0525 32.0975 ;
      RECT  21.1625 33.5425 21.22 33.4825 ;
      RECT  21.155 33.61 21.225 32.065 ;
      RECT  21.345 33.485 21.405 33.5425 ;
      RECT  20.82 33.41 20.89 34.955 ;
      RECT  21.34 33.41 21.41 34.955 ;
      RECT  21.3075 33.475 21.4425 33.545 ;
      RECT  20.635 34.26 20.705 34.395 ;
      RECT  21.34 34.26 21.41 34.395 ;
      RECT  21.085 33.7675 21.155 33.9025 ;
      RECT  21.34 33.4775 21.41 34.8875 ;
      RECT  20.89 33.7675 20.96 33.9025 ;
      RECT  20.8275 33.485 20.8825 33.5375 ;
      RECT  20.6025 33.475 20.7375 33.545 ;
      RECT  20.64 33.48 20.7 33.5375 ;
      RECT  20.635 33.41 20.705 34.955 ;
      RECT  20.9825 34.7875 21.0525 34.9225 ;
      RECT  21.1625 33.4775 21.22 33.5375 ;
      RECT  21.155 33.41 21.225 34.955 ;
      RECT  21.345 36.225 21.405 36.1675 ;
      RECT  20.82 36.3 20.89 34.755 ;
      RECT  21.34 36.3 21.41 34.755 ;
      RECT  21.3075 36.235 21.4425 36.165 ;
      RECT  20.635 35.45 20.705 35.315 ;
      RECT  21.34 35.45 21.41 35.315 ;
      RECT  21.085 35.9425 21.155 35.8075 ;
      RECT  21.34 36.2325 21.41 34.8225 ;
      RECT  20.89 35.9425 20.96 35.8075 ;
      RECT  20.8275 36.225 20.8825 36.1725 ;
      RECT  20.6025 36.235 20.7375 36.165 ;
      RECT  20.64 36.23 20.7 36.1725 ;
      RECT  20.635 36.3 20.705 34.755 ;
      RECT  20.9825 34.9225 21.0525 34.7875 ;
      RECT  21.1625 36.2325 21.22 36.1725 ;
      RECT  21.155 36.3 21.225 34.755 ;
      RECT  21.345 36.175 21.405 36.2325 ;
      RECT  20.82 36.1 20.89 37.645 ;
      RECT  21.34 36.1 21.41 37.645 ;
      RECT  21.3075 36.165 21.4425 36.235 ;
      RECT  20.635 36.95 20.705 37.085 ;
      RECT  21.34 36.95 21.41 37.085 ;
      RECT  21.085 36.4575 21.155 36.5925 ;
      RECT  21.34 36.1675 21.41 37.5775 ;
      RECT  20.89 36.4575 20.96 36.5925 ;
      RECT  20.8275 36.175 20.8825 36.2275 ;
      RECT  20.6025 36.165 20.7375 36.235 ;
      RECT  20.64 36.17 20.7 36.2275 ;
      RECT  20.635 36.1 20.705 37.645 ;
      RECT  20.9825 37.4775 21.0525 37.6125 ;
      RECT  21.1625 36.1675 21.22 36.2275 ;
      RECT  21.155 36.1 21.225 37.645 ;
      RECT  21.345 38.915 21.405 38.8575 ;
      RECT  20.82 38.99 20.89 37.445 ;
      RECT  21.34 38.99 21.41 37.445 ;
      RECT  21.3075 38.925 21.4425 38.855 ;
      RECT  20.635 38.14 20.705 38.005 ;
      RECT  21.34 38.14 21.41 38.005 ;
      RECT  21.085 38.6325 21.155 38.4975 ;
      RECT  21.34 38.9225 21.41 37.5125 ;
      RECT  20.89 38.6325 20.96 38.4975 ;
      RECT  20.8275 38.915 20.8825 38.8625 ;
      RECT  20.6025 38.925 20.7375 38.855 ;
      RECT  20.64 38.92 20.7 38.8625 ;
      RECT  20.635 38.99 20.705 37.445 ;
      RECT  20.9825 37.6125 21.0525 37.4775 ;
      RECT  21.1625 38.9225 21.22 38.8625 ;
      RECT  21.155 38.99 21.225 37.445 ;
      RECT  21.345 38.865 21.405 38.9225 ;
      RECT  20.82 38.79 20.89 40.335 ;
      RECT  21.34 38.79 21.41 40.335 ;
      RECT  21.3075 38.855 21.4425 38.925 ;
      RECT  20.635 39.64 20.705 39.775 ;
      RECT  21.34 39.64 21.41 39.775 ;
      RECT  21.085 39.1475 21.155 39.2825 ;
      RECT  21.34 38.8575 21.41 40.2675 ;
      RECT  20.89 39.1475 20.96 39.2825 ;
      RECT  20.8275 38.865 20.8825 38.9175 ;
      RECT  20.6025 38.855 20.7375 38.925 ;
      RECT  20.64 38.86 20.7 38.9175 ;
      RECT  20.635 38.79 20.705 40.335 ;
      RECT  20.9825 40.1675 21.0525 40.3025 ;
      RECT  21.1625 38.8575 21.22 38.9175 ;
      RECT  21.155 38.79 21.225 40.335 ;
      RECT  21.345 41.605 21.405 41.5475 ;
      RECT  20.82 41.68 20.89 40.135 ;
      RECT  21.34 41.68 21.41 40.135 ;
      RECT  21.3075 41.615 21.4425 41.545 ;
      RECT  20.635 40.83 20.705 40.695 ;
      RECT  21.34 40.83 21.41 40.695 ;
      RECT  21.085 41.3225 21.155 41.1875 ;
      RECT  21.34 41.6125 21.41 40.2025 ;
      RECT  20.89 41.3225 20.96 41.1875 ;
      RECT  20.8275 41.605 20.8825 41.5525 ;
      RECT  20.6025 41.615 20.7375 41.545 ;
      RECT  20.64 41.61 20.7 41.5525 ;
      RECT  20.635 41.68 20.705 40.135 ;
      RECT  20.9825 40.3025 21.0525 40.1675 ;
      RECT  21.1625 41.6125 21.22 41.5525 ;
      RECT  21.155 41.68 21.225 40.135 ;
      RECT  21.345 41.555 21.405 41.6125 ;
      RECT  20.82 41.48 20.89 43.025 ;
      RECT  21.34 41.48 21.41 43.025 ;
      RECT  21.3075 41.545 21.4425 41.615 ;
      RECT  20.635 42.33 20.705 42.465 ;
      RECT  21.34 42.33 21.41 42.465 ;
      RECT  21.085 41.8375 21.155 41.9725 ;
      RECT  21.34 41.5475 21.41 42.9575 ;
      RECT  20.89 41.8375 20.96 41.9725 ;
      RECT  20.8275 41.555 20.8825 41.6075 ;
      RECT  20.6025 41.545 20.7375 41.615 ;
      RECT  20.64 41.55 20.7 41.6075 ;
      RECT  20.635 41.48 20.705 43.025 ;
      RECT  20.9825 42.8575 21.0525 42.9925 ;
      RECT  21.1625 41.5475 21.22 41.6075 ;
      RECT  21.155 41.48 21.225 43.025 ;
      RECT  21.345 44.295 21.405 44.2375 ;
      RECT  20.82 44.37 20.89 42.825 ;
      RECT  21.34 44.37 21.41 42.825 ;
      RECT  21.3075 44.305 21.4425 44.235 ;
      RECT  20.635 43.52 20.705 43.385 ;
      RECT  21.34 43.52 21.41 43.385 ;
      RECT  21.085 44.0125 21.155 43.8775 ;
      RECT  21.34 44.3025 21.41 42.8925 ;
      RECT  20.89 44.0125 20.96 43.8775 ;
      RECT  20.8275 44.295 20.8825 44.2425 ;
      RECT  20.6025 44.305 20.7375 44.235 ;
      RECT  20.64 44.3 20.7 44.2425 ;
      RECT  20.635 44.37 20.705 42.825 ;
      RECT  20.9825 42.9925 21.0525 42.8575 ;
      RECT  21.1625 44.3025 21.22 44.2425 ;
      RECT  21.155 44.37 21.225 42.825 ;
      RECT  21.345 44.245 21.405 44.3025 ;
      RECT  20.635 45.02 20.705 45.155 ;
      RECT  20.82 44.17 20.89 45.715 ;
      RECT  21.3075 44.235 21.4425 44.305 ;
      RECT  21.34 44.17 21.41 45.715 ;
      RECT  20.635 44.17 20.705 45.715 ;
      RECT  21.085 44.5275 21.155 44.6625 ;
      RECT  21.34 44.2375 21.41 45.6475 ;
      RECT  20.89 44.5275 20.96 44.6625 ;
      RECT  20.8275 44.245 20.8825 44.2975 ;
      RECT  20.9825 45.5475 21.0525 45.6825 ;
      RECT  20.64 44.24 20.7 44.2975 ;
      RECT  21.34 45.02 21.41 45.155 ;
      RECT  20.6025 44.235 20.7375 44.305 ;
      RECT  21.1625 44.2375 21.22 44.2975 ;
      RECT  21.155 44.17 21.225 45.715 ;
      RECT  20.82 20.06 20.89 45.615 ;
      RECT  21.155 20.06 21.225 45.615 ;
      RECT  20.9825 29.4075 21.0525 29.5425 ;
      RECT  20.9825 32.0975 21.0525 32.2325 ;
      RECT  20.9825 32.0975 21.0525 32.2325 ;
      RECT  20.9825 26.7175 21.0525 26.8525 ;
      RECT  20.9825 21.3375 21.0525 21.4725 ;
      RECT  20.9825 24.0275 21.0525 24.1625 ;
      RECT  20.9825 24.0275 21.0525 24.1625 ;
      RECT  20.9825 26.7175 21.0525 26.8525 ;
      RECT  20.9825 42.8575 21.0525 42.9925 ;
      RECT  20.9825 37.4775 21.0525 37.6125 ;
      RECT  20.9825 40.1675 21.0525 40.3025 ;
      RECT  20.9825 40.1675 21.0525 40.3025 ;
      RECT  20.9825 34.7875 21.0525 34.9225 ;
      RECT  20.6025 41.545 20.7375 41.615 ;
      RECT  20.6025 30.785 20.7375 30.855 ;
      RECT  20.6025 36.165 20.7375 36.235 ;
      RECT  20.6025 38.855 20.7375 38.925 ;
      RECT  20.6025 44.235 20.7375 44.305 ;
      RECT  20.6025 28.095 20.7375 28.165 ;
      RECT  20.6025 22.715 20.7375 22.785 ;
      RECT  20.6025 33.475 20.7375 33.545 ;
      RECT  20.6025 25.405 20.7375 25.475 ;
      RECT  22.05 22.775 22.11 22.7175 ;
      RECT  21.34 22.0 21.41 21.865 ;
      RECT  21.525 22.85 21.595 21.305 ;
      RECT  22.0125 22.785 22.1475 22.715 ;
      RECT  22.045 22.85 22.115 21.305 ;
      RECT  21.34 22.85 21.41 21.305 ;
      RECT  21.79 22.4925 21.86 22.3575 ;
      RECT  22.045 22.7825 22.115 21.3725 ;
      RECT  21.595 22.4925 21.665 22.3575 ;
      RECT  21.5325 22.775 21.5875 22.7225 ;
      RECT  21.6875 21.4725 21.7575 21.3375 ;
      RECT  21.345 22.78 21.405 22.7225 ;
      RECT  22.045 22.0 22.115 21.865 ;
      RECT  21.3075 22.785 21.4425 22.715 ;
      RECT  21.8675 22.7825 21.925 22.7225 ;
      RECT  21.86 22.85 21.93 21.305 ;
      RECT  22.755 22.775 22.815 22.7175 ;
      RECT  22.045 22.0 22.115 21.865 ;
      RECT  22.23 22.85 22.3 21.305 ;
      RECT  22.7175 22.785 22.8525 22.715 ;
      RECT  22.75 22.85 22.82 21.305 ;
      RECT  22.045 22.85 22.115 21.305 ;
      RECT  22.495 22.4925 22.565 22.3575 ;
      RECT  22.75 22.7825 22.82 21.3725 ;
      RECT  22.3 22.4925 22.37 22.3575 ;
      RECT  22.2375 22.775 22.2925 22.7225 ;
      RECT  22.3925 21.4725 22.4625 21.3375 ;
      RECT  22.05 22.78 22.11 22.7225 ;
      RECT  22.75 22.0 22.82 21.865 ;
      RECT  22.0125 22.785 22.1475 22.715 ;
      RECT  22.5725 22.7825 22.63 22.7225 ;
      RECT  22.565 22.85 22.635 21.305 ;
      RECT  22.3925 21.4725 22.4625 21.3375 ;
      RECT  21.6875 21.4725 21.7575 21.3375 ;
      RECT  22.0125 22.785 22.1475 22.715 ;
      RECT  21.3075 22.785 21.4425 22.715 ;
      RECT  22.05 20.035 22.11 20.0925 ;
      RECT  21.34 20.81 21.41 20.945 ;
      RECT  21.525 19.96 21.595 21.505 ;
      RECT  22.0125 20.025 22.1475 20.095 ;
      RECT  22.045 19.96 22.115 21.505 ;
      RECT  21.34 19.96 21.41 21.505 ;
      RECT  21.79 20.3175 21.86 20.4525 ;
      RECT  22.045 20.0275 22.115 21.4375 ;
      RECT  21.595 20.3175 21.665 20.4525 ;
      RECT  21.5325 20.035 21.5875 20.0875 ;
      RECT  21.6875 21.3375 21.7575 21.4725 ;
      RECT  21.345 20.03 21.405 20.0875 ;
      RECT  22.045 20.81 22.115 20.945 ;
      RECT  21.3075 20.025 21.4425 20.095 ;
      RECT  21.8675 20.0275 21.925 20.0875 ;
      RECT  21.86 19.96 21.93 21.505 ;
      RECT  22.755 20.035 22.815 20.0925 ;
      RECT  22.045 20.81 22.115 20.945 ;
      RECT  22.23 19.96 22.3 21.505 ;
      RECT  22.7175 20.025 22.8525 20.095 ;
      RECT  22.75 19.96 22.82 21.505 ;
      RECT  22.045 19.96 22.115 21.505 ;
      RECT  22.495 20.3175 22.565 20.4525 ;
      RECT  22.75 20.0275 22.82 21.4375 ;
      RECT  22.3 20.3175 22.37 20.4525 ;
      RECT  22.2375 20.035 22.2925 20.0875 ;
      RECT  22.3925 21.3375 22.4625 21.4725 ;
      RECT  22.05 20.03 22.11 20.0875 ;
      RECT  22.75 20.81 22.82 20.945 ;
      RECT  22.0125 20.025 22.1475 20.095 ;
      RECT  22.5725 20.0275 22.63 20.0875 ;
      RECT  22.565 19.96 22.635 21.505 ;
      RECT  22.3925 21.3375 22.4625 21.4725 ;
      RECT  21.6875 21.3375 21.7575 21.4725 ;
      RECT  22.0125 20.025 22.1475 20.095 ;
      RECT  21.3075 20.025 21.4425 20.095 ;
      RECT  22.05 44.245 22.11 44.3025 ;
      RECT  21.34 45.02 21.41 45.155 ;
      RECT  21.525 44.17 21.595 45.715 ;
      RECT  22.0125 44.235 22.1475 44.305 ;
      RECT  22.045 44.17 22.115 45.715 ;
      RECT  21.34 44.17 21.41 45.715 ;
      RECT  21.79 44.5275 21.86 44.6625 ;
      RECT  22.045 44.2375 22.115 45.6475 ;
      RECT  21.595 44.5275 21.665 44.6625 ;
      RECT  21.5325 44.245 21.5875 44.2975 ;
      RECT  21.6875 45.5475 21.7575 45.6825 ;
      RECT  21.345 44.24 21.405 44.2975 ;
      RECT  22.045 45.02 22.115 45.155 ;
      RECT  21.3075 44.235 21.4425 44.305 ;
      RECT  21.8675 44.2375 21.925 44.2975 ;
      RECT  21.86 44.17 21.93 45.715 ;
      RECT  22.755 44.245 22.815 44.3025 ;
      RECT  22.045 45.02 22.115 45.155 ;
      RECT  22.23 44.17 22.3 45.715 ;
      RECT  22.7175 44.235 22.8525 44.305 ;
      RECT  22.75 44.17 22.82 45.715 ;
      RECT  22.045 44.17 22.115 45.715 ;
      RECT  22.495 44.5275 22.565 44.6625 ;
      RECT  22.75 44.2375 22.82 45.6475 ;
      RECT  22.3 44.5275 22.37 44.6625 ;
      RECT  22.2375 44.245 22.2925 44.2975 ;
      RECT  22.3925 45.5475 22.4625 45.6825 ;
      RECT  22.05 44.24 22.11 44.2975 ;
      RECT  22.75 45.02 22.82 45.155 ;
      RECT  22.0125 44.235 22.1475 44.305 ;
      RECT  22.5725 44.2375 22.63 44.2975 ;
      RECT  22.565 44.17 22.635 45.715 ;
      RECT  22.3925 45.5475 22.4625 45.6825 ;
      RECT  21.6875 45.5475 21.7575 45.6825 ;
      RECT  22.0125 44.235 22.1475 44.305 ;
      RECT  21.3075 44.235 21.4425 44.305 ;
      RECT  20.64 20.035 20.7 20.0925 ;
      RECT  19.93 20.81 20.0 20.945 ;
      RECT  20.115 19.96 20.185 21.505 ;
      RECT  20.6025 20.025 20.7375 20.095 ;
      RECT  20.635 19.96 20.705 21.505 ;
      RECT  19.93 19.96 20.0 21.505 ;
      RECT  20.38 20.3175 20.45 20.4525 ;
      RECT  20.635 20.0275 20.705 21.4375 ;
      RECT  20.185 20.3175 20.255 20.4525 ;
      RECT  20.1225 20.035 20.1775 20.0875 ;
      RECT  20.2775 21.3375 20.3475 21.4725 ;
      RECT  19.935 20.03 19.995 20.0875 ;
      RECT  20.635 20.81 20.705 20.945 ;
      RECT  19.8975 20.025 20.0325 20.095 ;
      RECT  20.4575 20.0275 20.515 20.0875 ;
      RECT  20.45 19.96 20.52 21.505 ;
      RECT  20.64 22.775 20.7 22.7175 ;
      RECT  19.93 22.0 20.0 21.865 ;
      RECT  20.115 22.85 20.185 21.305 ;
      RECT  20.6025 22.785 20.7375 22.715 ;
      RECT  20.635 22.85 20.705 21.305 ;
      RECT  19.93 22.85 20.0 21.305 ;
      RECT  20.38 22.4925 20.45 22.3575 ;
      RECT  20.635 22.7825 20.705 21.3725 ;
      RECT  20.185 22.4925 20.255 22.3575 ;
      RECT  20.1225 22.775 20.1775 22.7225 ;
      RECT  20.2775 21.4725 20.3475 21.3375 ;
      RECT  19.935 22.78 19.995 22.7225 ;
      RECT  20.635 22.0 20.705 21.865 ;
      RECT  19.8975 22.785 20.0325 22.715 ;
      RECT  20.4575 22.7825 20.515 22.7225 ;
      RECT  20.45 22.85 20.52 21.305 ;
      RECT  20.64 22.725 20.7 22.7825 ;
      RECT  19.93 23.5 20.0 23.635 ;
      RECT  20.115 22.65 20.185 24.195 ;
      RECT  20.6025 22.715 20.7375 22.785 ;
      RECT  20.635 22.65 20.705 24.195 ;
      RECT  19.93 22.65 20.0 24.195 ;
      RECT  20.38 23.0075 20.45 23.1425 ;
      RECT  20.635 22.7175 20.705 24.1275 ;
      RECT  20.185 23.0075 20.255 23.1425 ;
      RECT  20.1225 22.725 20.1775 22.7775 ;
      RECT  20.2775 24.0275 20.3475 24.1625 ;
      RECT  19.935 22.72 19.995 22.7775 ;
      RECT  20.635 23.5 20.705 23.635 ;
      RECT  19.8975 22.715 20.0325 22.785 ;
      RECT  20.4575 22.7175 20.515 22.7775 ;
      RECT  20.45 22.65 20.52 24.195 ;
      RECT  20.64 25.465 20.7 25.4075 ;
      RECT  19.93 24.69 20.0 24.555 ;
      RECT  20.115 25.54 20.185 23.995 ;
      RECT  20.6025 25.475 20.7375 25.405 ;
      RECT  20.635 25.54 20.705 23.995 ;
      RECT  19.93 25.54 20.0 23.995 ;
      RECT  20.38 25.1825 20.45 25.0475 ;
      RECT  20.635 25.4725 20.705 24.0625 ;
      RECT  20.185 25.1825 20.255 25.0475 ;
      RECT  20.1225 25.465 20.1775 25.4125 ;
      RECT  20.2775 24.1625 20.3475 24.0275 ;
      RECT  19.935 25.47 19.995 25.4125 ;
      RECT  20.635 24.69 20.705 24.555 ;
      RECT  19.8975 25.475 20.0325 25.405 ;
      RECT  20.4575 25.4725 20.515 25.4125 ;
      RECT  20.45 25.54 20.52 23.995 ;
      RECT  20.64 25.415 20.7 25.4725 ;
      RECT  19.93 26.19 20.0 26.325 ;
      RECT  20.115 25.34 20.185 26.885 ;
      RECT  20.6025 25.405 20.7375 25.475 ;
      RECT  20.635 25.34 20.705 26.885 ;
      RECT  19.93 25.34 20.0 26.885 ;
      RECT  20.38 25.6975 20.45 25.8325 ;
      RECT  20.635 25.4075 20.705 26.8175 ;
      RECT  20.185 25.6975 20.255 25.8325 ;
      RECT  20.1225 25.415 20.1775 25.4675 ;
      RECT  20.2775 26.7175 20.3475 26.8525 ;
      RECT  19.935 25.41 19.995 25.4675 ;
      RECT  20.635 26.19 20.705 26.325 ;
      RECT  19.8975 25.405 20.0325 25.475 ;
      RECT  20.4575 25.4075 20.515 25.4675 ;
      RECT  20.45 25.34 20.52 26.885 ;
      RECT  20.64 28.155 20.7 28.0975 ;
      RECT  19.93 27.38 20.0 27.245 ;
      RECT  20.115 28.23 20.185 26.685 ;
      RECT  20.6025 28.165 20.7375 28.095 ;
      RECT  20.635 28.23 20.705 26.685 ;
      RECT  19.93 28.23 20.0 26.685 ;
      RECT  20.38 27.8725 20.45 27.7375 ;
      RECT  20.635 28.1625 20.705 26.7525 ;
      RECT  20.185 27.8725 20.255 27.7375 ;
      RECT  20.1225 28.155 20.1775 28.1025 ;
      RECT  20.2775 26.8525 20.3475 26.7175 ;
      RECT  19.935 28.16 19.995 28.1025 ;
      RECT  20.635 27.38 20.705 27.245 ;
      RECT  19.8975 28.165 20.0325 28.095 ;
      RECT  20.4575 28.1625 20.515 28.1025 ;
      RECT  20.45 28.23 20.52 26.685 ;
      RECT  20.64 28.105 20.7 28.1625 ;
      RECT  19.93 28.88 20.0 29.015 ;
      RECT  20.115 28.03 20.185 29.575 ;
      RECT  20.6025 28.095 20.7375 28.165 ;
      RECT  20.635 28.03 20.705 29.575 ;
      RECT  19.93 28.03 20.0 29.575 ;
      RECT  20.38 28.3875 20.45 28.5225 ;
      RECT  20.635 28.0975 20.705 29.5075 ;
      RECT  20.185 28.3875 20.255 28.5225 ;
      RECT  20.1225 28.105 20.1775 28.1575 ;
      RECT  20.2775 29.4075 20.3475 29.5425 ;
      RECT  19.935 28.1 19.995 28.1575 ;
      RECT  20.635 28.88 20.705 29.015 ;
      RECT  19.8975 28.095 20.0325 28.165 ;
      RECT  20.4575 28.0975 20.515 28.1575 ;
      RECT  20.45 28.03 20.52 29.575 ;
      RECT  20.64 30.845 20.7 30.7875 ;
      RECT  19.93 30.07 20.0 29.935 ;
      RECT  20.115 30.92 20.185 29.375 ;
      RECT  20.6025 30.855 20.7375 30.785 ;
      RECT  20.635 30.92 20.705 29.375 ;
      RECT  19.93 30.92 20.0 29.375 ;
      RECT  20.38 30.5625 20.45 30.4275 ;
      RECT  20.635 30.8525 20.705 29.4425 ;
      RECT  20.185 30.5625 20.255 30.4275 ;
      RECT  20.1225 30.845 20.1775 30.7925 ;
      RECT  20.2775 29.5425 20.3475 29.4075 ;
      RECT  19.935 30.85 19.995 30.7925 ;
      RECT  20.635 30.07 20.705 29.935 ;
      RECT  19.8975 30.855 20.0325 30.785 ;
      RECT  20.4575 30.8525 20.515 30.7925 ;
      RECT  20.45 30.92 20.52 29.375 ;
      RECT  20.64 30.795 20.7 30.8525 ;
      RECT  19.93 31.57 20.0 31.705 ;
      RECT  20.115 30.72 20.185 32.265 ;
      RECT  20.6025 30.785 20.7375 30.855 ;
      RECT  20.635 30.72 20.705 32.265 ;
      RECT  19.93 30.72 20.0 32.265 ;
      RECT  20.38 31.0775 20.45 31.2125 ;
      RECT  20.635 30.7875 20.705 32.1975 ;
      RECT  20.185 31.0775 20.255 31.2125 ;
      RECT  20.1225 30.795 20.1775 30.8475 ;
      RECT  20.2775 32.0975 20.3475 32.2325 ;
      RECT  19.935 30.79 19.995 30.8475 ;
      RECT  20.635 31.57 20.705 31.705 ;
      RECT  19.8975 30.785 20.0325 30.855 ;
      RECT  20.4575 30.7875 20.515 30.8475 ;
      RECT  20.45 30.72 20.52 32.265 ;
      RECT  20.64 33.535 20.7 33.4775 ;
      RECT  19.93 32.76 20.0 32.625 ;
      RECT  20.115 33.61 20.185 32.065 ;
      RECT  20.6025 33.545 20.7375 33.475 ;
      RECT  20.635 33.61 20.705 32.065 ;
      RECT  19.93 33.61 20.0 32.065 ;
      RECT  20.38 33.2525 20.45 33.1175 ;
      RECT  20.635 33.5425 20.705 32.1325 ;
      RECT  20.185 33.2525 20.255 33.1175 ;
      RECT  20.1225 33.535 20.1775 33.4825 ;
      RECT  20.2775 32.2325 20.3475 32.0975 ;
      RECT  19.935 33.54 19.995 33.4825 ;
      RECT  20.635 32.76 20.705 32.625 ;
      RECT  19.8975 33.545 20.0325 33.475 ;
      RECT  20.4575 33.5425 20.515 33.4825 ;
      RECT  20.45 33.61 20.52 32.065 ;
      RECT  20.64 33.485 20.7 33.5425 ;
      RECT  19.93 34.26 20.0 34.395 ;
      RECT  20.115 33.41 20.185 34.955 ;
      RECT  20.6025 33.475 20.7375 33.545 ;
      RECT  20.635 33.41 20.705 34.955 ;
      RECT  19.93 33.41 20.0 34.955 ;
      RECT  20.38 33.7675 20.45 33.9025 ;
      RECT  20.635 33.4775 20.705 34.8875 ;
      RECT  20.185 33.7675 20.255 33.9025 ;
      RECT  20.1225 33.485 20.1775 33.5375 ;
      RECT  20.2775 34.7875 20.3475 34.9225 ;
      RECT  19.935 33.48 19.995 33.5375 ;
      RECT  20.635 34.26 20.705 34.395 ;
      RECT  19.8975 33.475 20.0325 33.545 ;
      RECT  20.4575 33.4775 20.515 33.5375 ;
      RECT  20.45 33.41 20.52 34.955 ;
      RECT  20.64 36.225 20.7 36.1675 ;
      RECT  19.93 35.45 20.0 35.315 ;
      RECT  20.115 36.3 20.185 34.755 ;
      RECT  20.6025 36.235 20.7375 36.165 ;
      RECT  20.635 36.3 20.705 34.755 ;
      RECT  19.93 36.3 20.0 34.755 ;
      RECT  20.38 35.9425 20.45 35.8075 ;
      RECT  20.635 36.2325 20.705 34.8225 ;
      RECT  20.185 35.9425 20.255 35.8075 ;
      RECT  20.1225 36.225 20.1775 36.1725 ;
      RECT  20.2775 34.9225 20.3475 34.7875 ;
      RECT  19.935 36.23 19.995 36.1725 ;
      RECT  20.635 35.45 20.705 35.315 ;
      RECT  19.8975 36.235 20.0325 36.165 ;
      RECT  20.4575 36.2325 20.515 36.1725 ;
      RECT  20.45 36.3 20.52 34.755 ;
      RECT  20.64 36.175 20.7 36.2325 ;
      RECT  19.93 36.95 20.0 37.085 ;
      RECT  20.115 36.1 20.185 37.645 ;
      RECT  20.6025 36.165 20.7375 36.235 ;
      RECT  20.635 36.1 20.705 37.645 ;
      RECT  19.93 36.1 20.0 37.645 ;
      RECT  20.38 36.4575 20.45 36.5925 ;
      RECT  20.635 36.1675 20.705 37.5775 ;
      RECT  20.185 36.4575 20.255 36.5925 ;
      RECT  20.1225 36.175 20.1775 36.2275 ;
      RECT  20.2775 37.4775 20.3475 37.6125 ;
      RECT  19.935 36.17 19.995 36.2275 ;
      RECT  20.635 36.95 20.705 37.085 ;
      RECT  19.8975 36.165 20.0325 36.235 ;
      RECT  20.4575 36.1675 20.515 36.2275 ;
      RECT  20.45 36.1 20.52 37.645 ;
      RECT  20.64 38.915 20.7 38.8575 ;
      RECT  19.93 38.14 20.0 38.005 ;
      RECT  20.115 38.99 20.185 37.445 ;
      RECT  20.6025 38.925 20.7375 38.855 ;
      RECT  20.635 38.99 20.705 37.445 ;
      RECT  19.93 38.99 20.0 37.445 ;
      RECT  20.38 38.6325 20.45 38.4975 ;
      RECT  20.635 38.9225 20.705 37.5125 ;
      RECT  20.185 38.6325 20.255 38.4975 ;
      RECT  20.1225 38.915 20.1775 38.8625 ;
      RECT  20.2775 37.6125 20.3475 37.4775 ;
      RECT  19.935 38.92 19.995 38.8625 ;
      RECT  20.635 38.14 20.705 38.005 ;
      RECT  19.8975 38.925 20.0325 38.855 ;
      RECT  20.4575 38.9225 20.515 38.8625 ;
      RECT  20.45 38.99 20.52 37.445 ;
      RECT  20.64 38.865 20.7 38.9225 ;
      RECT  19.93 39.64 20.0 39.775 ;
      RECT  20.115 38.79 20.185 40.335 ;
      RECT  20.6025 38.855 20.7375 38.925 ;
      RECT  20.635 38.79 20.705 40.335 ;
      RECT  19.93 38.79 20.0 40.335 ;
      RECT  20.38 39.1475 20.45 39.2825 ;
      RECT  20.635 38.8575 20.705 40.2675 ;
      RECT  20.185 39.1475 20.255 39.2825 ;
      RECT  20.1225 38.865 20.1775 38.9175 ;
      RECT  20.2775 40.1675 20.3475 40.3025 ;
      RECT  19.935 38.86 19.995 38.9175 ;
      RECT  20.635 39.64 20.705 39.775 ;
      RECT  19.8975 38.855 20.0325 38.925 ;
      RECT  20.4575 38.8575 20.515 38.9175 ;
      RECT  20.45 38.79 20.52 40.335 ;
      RECT  20.64 41.605 20.7 41.5475 ;
      RECT  19.93 40.83 20.0 40.695 ;
      RECT  20.115 41.68 20.185 40.135 ;
      RECT  20.6025 41.615 20.7375 41.545 ;
      RECT  20.635 41.68 20.705 40.135 ;
      RECT  19.93 41.68 20.0 40.135 ;
      RECT  20.38 41.3225 20.45 41.1875 ;
      RECT  20.635 41.6125 20.705 40.2025 ;
      RECT  20.185 41.3225 20.255 41.1875 ;
      RECT  20.1225 41.605 20.1775 41.5525 ;
      RECT  20.2775 40.3025 20.3475 40.1675 ;
      RECT  19.935 41.61 19.995 41.5525 ;
      RECT  20.635 40.83 20.705 40.695 ;
      RECT  19.8975 41.615 20.0325 41.545 ;
      RECT  20.4575 41.6125 20.515 41.5525 ;
      RECT  20.45 41.68 20.52 40.135 ;
      RECT  20.64 41.555 20.7 41.6125 ;
      RECT  19.93 42.33 20.0 42.465 ;
      RECT  20.115 41.48 20.185 43.025 ;
      RECT  20.6025 41.545 20.7375 41.615 ;
      RECT  20.635 41.48 20.705 43.025 ;
      RECT  19.93 41.48 20.0 43.025 ;
      RECT  20.38 41.8375 20.45 41.9725 ;
      RECT  20.635 41.5475 20.705 42.9575 ;
      RECT  20.185 41.8375 20.255 41.9725 ;
      RECT  20.1225 41.555 20.1775 41.6075 ;
      RECT  20.2775 42.8575 20.3475 42.9925 ;
      RECT  19.935 41.55 19.995 41.6075 ;
      RECT  20.635 42.33 20.705 42.465 ;
      RECT  19.8975 41.545 20.0325 41.615 ;
      RECT  20.4575 41.5475 20.515 41.6075 ;
      RECT  20.45 41.48 20.52 43.025 ;
      RECT  20.64 44.295 20.7 44.2375 ;
      RECT  19.93 43.52 20.0 43.385 ;
      RECT  20.115 44.37 20.185 42.825 ;
      RECT  20.6025 44.305 20.7375 44.235 ;
      RECT  20.635 44.37 20.705 42.825 ;
      RECT  19.93 44.37 20.0 42.825 ;
      RECT  20.38 44.0125 20.45 43.8775 ;
      RECT  20.635 44.3025 20.705 42.8925 ;
      RECT  20.185 44.0125 20.255 43.8775 ;
      RECT  20.1225 44.295 20.1775 44.2425 ;
      RECT  20.2775 42.9925 20.3475 42.8575 ;
      RECT  19.935 44.3 19.995 44.2425 ;
      RECT  20.635 43.52 20.705 43.385 ;
      RECT  19.8975 44.305 20.0325 44.235 ;
      RECT  20.4575 44.3025 20.515 44.2425 ;
      RECT  20.45 44.37 20.52 42.825 ;
      RECT  20.64 44.245 20.7 44.3025 ;
      RECT  19.93 45.02 20.0 45.155 ;
      RECT  20.115 44.17 20.185 45.715 ;
      RECT  20.6025 44.235 20.7375 44.305 ;
      RECT  20.635 44.17 20.705 45.715 ;
      RECT  19.93 44.17 20.0 45.715 ;
      RECT  20.38 44.5275 20.45 44.6625 ;
      RECT  20.635 44.2375 20.705 45.6475 ;
      RECT  20.185 44.5275 20.255 44.6625 ;
      RECT  20.1225 44.245 20.1775 44.2975 ;
      RECT  20.2775 45.5475 20.3475 45.6825 ;
      RECT  19.935 44.24 19.995 44.2975 ;
      RECT  20.635 45.02 20.705 45.155 ;
      RECT  19.8975 44.235 20.0325 44.305 ;
      RECT  20.4575 44.2375 20.515 44.2975 ;
      RECT  20.45 44.17 20.52 45.715 ;
      RECT  20.2775 29.4075 20.3475 29.5425 ;
      RECT  20.2775 32.0975 20.3475 32.2325 ;
      RECT  20.2775 32.0975 20.3475 32.2325 ;
      RECT  20.2775 45.5475 20.3475 45.6825 ;
      RECT  20.2775 26.7175 20.3475 26.8525 ;
      RECT  20.2775 21.3375 20.3475 21.4725 ;
      RECT  20.2775 24.0275 20.3475 24.1625 ;
      RECT  20.2775 24.0275 20.3475 24.1625 ;
      RECT  20.2775 21.3375 20.3475 21.4725 ;
      RECT  20.2775 26.7175 20.3475 26.8525 ;
      RECT  20.2775 42.8575 20.3475 42.9925 ;
      RECT  20.2775 37.4775 20.3475 37.6125 ;
      RECT  20.2775 40.1675 20.3475 40.3025 ;
      RECT  20.2775 40.1675 20.3475 40.3025 ;
      RECT  20.2775 34.7875 20.3475 34.9225 ;
      RECT  19.8975 41.545 20.0325 41.615 ;
      RECT  19.8975 30.785 20.0325 30.855 ;
      RECT  19.8975 36.165 20.0325 36.235 ;
      RECT  19.8975 38.855 20.0325 38.925 ;
      RECT  19.8975 44.235 20.0325 44.305 ;
      RECT  19.8975 20.025 20.0325 20.095 ;
      RECT  19.8975 28.095 20.0325 28.165 ;
      RECT  19.8975 22.715 20.0325 22.785 ;
      RECT  19.8975 33.475 20.0325 33.545 ;
      RECT  19.8975 25.405 20.0325 25.475 ;
      RECT  23.46 20.035 23.52 20.0925 ;
      RECT  22.75 20.81 22.82 20.945 ;
      RECT  22.935 19.96 23.005 21.505 ;
      RECT  23.4225 20.025 23.5575 20.095 ;
      RECT  23.455 19.96 23.525 21.505 ;
      RECT  22.75 19.96 22.82 21.505 ;
      RECT  23.2 20.3175 23.27 20.4525 ;
      RECT  23.455 20.0275 23.525 21.4375 ;
      RECT  23.005 20.3175 23.075 20.4525 ;
      RECT  22.9425 20.035 22.9975 20.0875 ;
      RECT  23.0975 21.3375 23.1675 21.4725 ;
      RECT  22.755 20.03 22.815 20.0875 ;
      RECT  23.455 20.81 23.525 20.945 ;
      RECT  22.7175 20.025 22.8525 20.095 ;
      RECT  23.2775 20.0275 23.335 20.0875 ;
      RECT  23.27 19.96 23.34 21.505 ;
      RECT  23.46 22.775 23.52 22.7175 ;
      RECT  22.75 22.0 22.82 21.865 ;
      RECT  22.935 22.85 23.005 21.305 ;
      RECT  23.4225 22.785 23.5575 22.715 ;
      RECT  23.455 22.85 23.525 21.305 ;
      RECT  22.75 22.85 22.82 21.305 ;
      RECT  23.2 22.4925 23.27 22.3575 ;
      RECT  23.455 22.7825 23.525 21.3725 ;
      RECT  23.005 22.4925 23.075 22.3575 ;
      RECT  22.9425 22.775 22.9975 22.7225 ;
      RECT  23.0975 21.4725 23.1675 21.3375 ;
      RECT  22.755 22.78 22.815 22.7225 ;
      RECT  23.455 22.0 23.525 21.865 ;
      RECT  22.7175 22.785 22.8525 22.715 ;
      RECT  23.2775 22.7825 23.335 22.7225 ;
      RECT  23.27 22.85 23.34 21.305 ;
      RECT  23.46 22.725 23.52 22.7825 ;
      RECT  22.75 23.5 22.82 23.635 ;
      RECT  22.935 22.65 23.005 24.195 ;
      RECT  23.4225 22.715 23.5575 22.785 ;
      RECT  23.455 22.65 23.525 24.195 ;
      RECT  22.75 22.65 22.82 24.195 ;
      RECT  23.2 23.0075 23.27 23.1425 ;
      RECT  23.455 22.7175 23.525 24.1275 ;
      RECT  23.005 23.0075 23.075 23.1425 ;
      RECT  22.9425 22.725 22.9975 22.7775 ;
      RECT  23.0975 24.0275 23.1675 24.1625 ;
      RECT  22.755 22.72 22.815 22.7775 ;
      RECT  23.455 23.5 23.525 23.635 ;
      RECT  22.7175 22.715 22.8525 22.785 ;
      RECT  23.2775 22.7175 23.335 22.7775 ;
      RECT  23.27 22.65 23.34 24.195 ;
      RECT  23.46 25.465 23.52 25.4075 ;
      RECT  22.75 24.69 22.82 24.555 ;
      RECT  22.935 25.54 23.005 23.995 ;
      RECT  23.4225 25.475 23.5575 25.405 ;
      RECT  23.455 25.54 23.525 23.995 ;
      RECT  22.75 25.54 22.82 23.995 ;
      RECT  23.2 25.1825 23.27 25.0475 ;
      RECT  23.455 25.4725 23.525 24.0625 ;
      RECT  23.005 25.1825 23.075 25.0475 ;
      RECT  22.9425 25.465 22.9975 25.4125 ;
      RECT  23.0975 24.1625 23.1675 24.0275 ;
      RECT  22.755 25.47 22.815 25.4125 ;
      RECT  23.455 24.69 23.525 24.555 ;
      RECT  22.7175 25.475 22.8525 25.405 ;
      RECT  23.2775 25.4725 23.335 25.4125 ;
      RECT  23.27 25.54 23.34 23.995 ;
      RECT  23.46 25.415 23.52 25.4725 ;
      RECT  22.75 26.19 22.82 26.325 ;
      RECT  22.935 25.34 23.005 26.885 ;
      RECT  23.4225 25.405 23.5575 25.475 ;
      RECT  23.455 25.34 23.525 26.885 ;
      RECT  22.75 25.34 22.82 26.885 ;
      RECT  23.2 25.6975 23.27 25.8325 ;
      RECT  23.455 25.4075 23.525 26.8175 ;
      RECT  23.005 25.6975 23.075 25.8325 ;
      RECT  22.9425 25.415 22.9975 25.4675 ;
      RECT  23.0975 26.7175 23.1675 26.8525 ;
      RECT  22.755 25.41 22.815 25.4675 ;
      RECT  23.455 26.19 23.525 26.325 ;
      RECT  22.7175 25.405 22.8525 25.475 ;
      RECT  23.2775 25.4075 23.335 25.4675 ;
      RECT  23.27 25.34 23.34 26.885 ;
      RECT  23.46 28.155 23.52 28.0975 ;
      RECT  22.75 27.38 22.82 27.245 ;
      RECT  22.935 28.23 23.005 26.685 ;
      RECT  23.4225 28.165 23.5575 28.095 ;
      RECT  23.455 28.23 23.525 26.685 ;
      RECT  22.75 28.23 22.82 26.685 ;
      RECT  23.2 27.8725 23.27 27.7375 ;
      RECT  23.455 28.1625 23.525 26.7525 ;
      RECT  23.005 27.8725 23.075 27.7375 ;
      RECT  22.9425 28.155 22.9975 28.1025 ;
      RECT  23.0975 26.8525 23.1675 26.7175 ;
      RECT  22.755 28.16 22.815 28.1025 ;
      RECT  23.455 27.38 23.525 27.245 ;
      RECT  22.7175 28.165 22.8525 28.095 ;
      RECT  23.2775 28.1625 23.335 28.1025 ;
      RECT  23.27 28.23 23.34 26.685 ;
      RECT  23.46 28.105 23.52 28.1625 ;
      RECT  22.75 28.88 22.82 29.015 ;
      RECT  22.935 28.03 23.005 29.575 ;
      RECT  23.4225 28.095 23.5575 28.165 ;
      RECT  23.455 28.03 23.525 29.575 ;
      RECT  22.75 28.03 22.82 29.575 ;
      RECT  23.2 28.3875 23.27 28.5225 ;
      RECT  23.455 28.0975 23.525 29.5075 ;
      RECT  23.005 28.3875 23.075 28.5225 ;
      RECT  22.9425 28.105 22.9975 28.1575 ;
      RECT  23.0975 29.4075 23.1675 29.5425 ;
      RECT  22.755 28.1 22.815 28.1575 ;
      RECT  23.455 28.88 23.525 29.015 ;
      RECT  22.7175 28.095 22.8525 28.165 ;
      RECT  23.2775 28.0975 23.335 28.1575 ;
      RECT  23.27 28.03 23.34 29.575 ;
      RECT  23.46 30.845 23.52 30.7875 ;
      RECT  22.75 30.07 22.82 29.935 ;
      RECT  22.935 30.92 23.005 29.375 ;
      RECT  23.4225 30.855 23.5575 30.785 ;
      RECT  23.455 30.92 23.525 29.375 ;
      RECT  22.75 30.92 22.82 29.375 ;
      RECT  23.2 30.5625 23.27 30.4275 ;
      RECT  23.455 30.8525 23.525 29.4425 ;
      RECT  23.005 30.5625 23.075 30.4275 ;
      RECT  22.9425 30.845 22.9975 30.7925 ;
      RECT  23.0975 29.5425 23.1675 29.4075 ;
      RECT  22.755 30.85 22.815 30.7925 ;
      RECT  23.455 30.07 23.525 29.935 ;
      RECT  22.7175 30.855 22.8525 30.785 ;
      RECT  23.2775 30.8525 23.335 30.7925 ;
      RECT  23.27 30.92 23.34 29.375 ;
      RECT  23.46 30.795 23.52 30.8525 ;
      RECT  22.75 31.57 22.82 31.705 ;
      RECT  22.935 30.72 23.005 32.265 ;
      RECT  23.4225 30.785 23.5575 30.855 ;
      RECT  23.455 30.72 23.525 32.265 ;
      RECT  22.75 30.72 22.82 32.265 ;
      RECT  23.2 31.0775 23.27 31.2125 ;
      RECT  23.455 30.7875 23.525 32.1975 ;
      RECT  23.005 31.0775 23.075 31.2125 ;
      RECT  22.9425 30.795 22.9975 30.8475 ;
      RECT  23.0975 32.0975 23.1675 32.2325 ;
      RECT  22.755 30.79 22.815 30.8475 ;
      RECT  23.455 31.57 23.525 31.705 ;
      RECT  22.7175 30.785 22.8525 30.855 ;
      RECT  23.2775 30.7875 23.335 30.8475 ;
      RECT  23.27 30.72 23.34 32.265 ;
      RECT  23.46 33.535 23.52 33.4775 ;
      RECT  22.75 32.76 22.82 32.625 ;
      RECT  22.935 33.61 23.005 32.065 ;
      RECT  23.4225 33.545 23.5575 33.475 ;
      RECT  23.455 33.61 23.525 32.065 ;
      RECT  22.75 33.61 22.82 32.065 ;
      RECT  23.2 33.2525 23.27 33.1175 ;
      RECT  23.455 33.5425 23.525 32.1325 ;
      RECT  23.005 33.2525 23.075 33.1175 ;
      RECT  22.9425 33.535 22.9975 33.4825 ;
      RECT  23.0975 32.2325 23.1675 32.0975 ;
      RECT  22.755 33.54 22.815 33.4825 ;
      RECT  23.455 32.76 23.525 32.625 ;
      RECT  22.7175 33.545 22.8525 33.475 ;
      RECT  23.2775 33.5425 23.335 33.4825 ;
      RECT  23.27 33.61 23.34 32.065 ;
      RECT  23.46 33.485 23.52 33.5425 ;
      RECT  22.75 34.26 22.82 34.395 ;
      RECT  22.935 33.41 23.005 34.955 ;
      RECT  23.4225 33.475 23.5575 33.545 ;
      RECT  23.455 33.41 23.525 34.955 ;
      RECT  22.75 33.41 22.82 34.955 ;
      RECT  23.2 33.7675 23.27 33.9025 ;
      RECT  23.455 33.4775 23.525 34.8875 ;
      RECT  23.005 33.7675 23.075 33.9025 ;
      RECT  22.9425 33.485 22.9975 33.5375 ;
      RECT  23.0975 34.7875 23.1675 34.9225 ;
      RECT  22.755 33.48 22.815 33.5375 ;
      RECT  23.455 34.26 23.525 34.395 ;
      RECT  22.7175 33.475 22.8525 33.545 ;
      RECT  23.2775 33.4775 23.335 33.5375 ;
      RECT  23.27 33.41 23.34 34.955 ;
      RECT  23.46 36.225 23.52 36.1675 ;
      RECT  22.75 35.45 22.82 35.315 ;
      RECT  22.935 36.3 23.005 34.755 ;
      RECT  23.4225 36.235 23.5575 36.165 ;
      RECT  23.455 36.3 23.525 34.755 ;
      RECT  22.75 36.3 22.82 34.755 ;
      RECT  23.2 35.9425 23.27 35.8075 ;
      RECT  23.455 36.2325 23.525 34.8225 ;
      RECT  23.005 35.9425 23.075 35.8075 ;
      RECT  22.9425 36.225 22.9975 36.1725 ;
      RECT  23.0975 34.9225 23.1675 34.7875 ;
      RECT  22.755 36.23 22.815 36.1725 ;
      RECT  23.455 35.45 23.525 35.315 ;
      RECT  22.7175 36.235 22.8525 36.165 ;
      RECT  23.2775 36.2325 23.335 36.1725 ;
      RECT  23.27 36.3 23.34 34.755 ;
      RECT  23.46 36.175 23.52 36.2325 ;
      RECT  22.75 36.95 22.82 37.085 ;
      RECT  22.935 36.1 23.005 37.645 ;
      RECT  23.4225 36.165 23.5575 36.235 ;
      RECT  23.455 36.1 23.525 37.645 ;
      RECT  22.75 36.1 22.82 37.645 ;
      RECT  23.2 36.4575 23.27 36.5925 ;
      RECT  23.455 36.1675 23.525 37.5775 ;
      RECT  23.005 36.4575 23.075 36.5925 ;
      RECT  22.9425 36.175 22.9975 36.2275 ;
      RECT  23.0975 37.4775 23.1675 37.6125 ;
      RECT  22.755 36.17 22.815 36.2275 ;
      RECT  23.455 36.95 23.525 37.085 ;
      RECT  22.7175 36.165 22.8525 36.235 ;
      RECT  23.2775 36.1675 23.335 36.2275 ;
      RECT  23.27 36.1 23.34 37.645 ;
      RECT  23.46 38.915 23.52 38.8575 ;
      RECT  22.75 38.14 22.82 38.005 ;
      RECT  22.935 38.99 23.005 37.445 ;
      RECT  23.4225 38.925 23.5575 38.855 ;
      RECT  23.455 38.99 23.525 37.445 ;
      RECT  22.75 38.99 22.82 37.445 ;
      RECT  23.2 38.6325 23.27 38.4975 ;
      RECT  23.455 38.9225 23.525 37.5125 ;
      RECT  23.005 38.6325 23.075 38.4975 ;
      RECT  22.9425 38.915 22.9975 38.8625 ;
      RECT  23.0975 37.6125 23.1675 37.4775 ;
      RECT  22.755 38.92 22.815 38.8625 ;
      RECT  23.455 38.14 23.525 38.005 ;
      RECT  22.7175 38.925 22.8525 38.855 ;
      RECT  23.2775 38.9225 23.335 38.8625 ;
      RECT  23.27 38.99 23.34 37.445 ;
      RECT  23.46 38.865 23.52 38.9225 ;
      RECT  22.75 39.64 22.82 39.775 ;
      RECT  22.935 38.79 23.005 40.335 ;
      RECT  23.4225 38.855 23.5575 38.925 ;
      RECT  23.455 38.79 23.525 40.335 ;
      RECT  22.75 38.79 22.82 40.335 ;
      RECT  23.2 39.1475 23.27 39.2825 ;
      RECT  23.455 38.8575 23.525 40.2675 ;
      RECT  23.005 39.1475 23.075 39.2825 ;
      RECT  22.9425 38.865 22.9975 38.9175 ;
      RECT  23.0975 40.1675 23.1675 40.3025 ;
      RECT  22.755 38.86 22.815 38.9175 ;
      RECT  23.455 39.64 23.525 39.775 ;
      RECT  22.7175 38.855 22.8525 38.925 ;
      RECT  23.2775 38.8575 23.335 38.9175 ;
      RECT  23.27 38.79 23.34 40.335 ;
      RECT  23.46 41.605 23.52 41.5475 ;
      RECT  22.75 40.83 22.82 40.695 ;
      RECT  22.935 41.68 23.005 40.135 ;
      RECT  23.4225 41.615 23.5575 41.545 ;
      RECT  23.455 41.68 23.525 40.135 ;
      RECT  22.75 41.68 22.82 40.135 ;
      RECT  23.2 41.3225 23.27 41.1875 ;
      RECT  23.455 41.6125 23.525 40.2025 ;
      RECT  23.005 41.3225 23.075 41.1875 ;
      RECT  22.9425 41.605 22.9975 41.5525 ;
      RECT  23.0975 40.3025 23.1675 40.1675 ;
      RECT  22.755 41.61 22.815 41.5525 ;
      RECT  23.455 40.83 23.525 40.695 ;
      RECT  22.7175 41.615 22.8525 41.545 ;
      RECT  23.2775 41.6125 23.335 41.5525 ;
      RECT  23.27 41.68 23.34 40.135 ;
      RECT  23.46 41.555 23.52 41.6125 ;
      RECT  22.75 42.33 22.82 42.465 ;
      RECT  22.935 41.48 23.005 43.025 ;
      RECT  23.4225 41.545 23.5575 41.615 ;
      RECT  23.455 41.48 23.525 43.025 ;
      RECT  22.75 41.48 22.82 43.025 ;
      RECT  23.2 41.8375 23.27 41.9725 ;
      RECT  23.455 41.5475 23.525 42.9575 ;
      RECT  23.005 41.8375 23.075 41.9725 ;
      RECT  22.9425 41.555 22.9975 41.6075 ;
      RECT  23.0975 42.8575 23.1675 42.9925 ;
      RECT  22.755 41.55 22.815 41.6075 ;
      RECT  23.455 42.33 23.525 42.465 ;
      RECT  22.7175 41.545 22.8525 41.615 ;
      RECT  23.2775 41.5475 23.335 41.6075 ;
      RECT  23.27 41.48 23.34 43.025 ;
      RECT  23.46 44.295 23.52 44.2375 ;
      RECT  22.75 43.52 22.82 43.385 ;
      RECT  22.935 44.37 23.005 42.825 ;
      RECT  23.4225 44.305 23.5575 44.235 ;
      RECT  23.455 44.37 23.525 42.825 ;
      RECT  22.75 44.37 22.82 42.825 ;
      RECT  23.2 44.0125 23.27 43.8775 ;
      RECT  23.455 44.3025 23.525 42.8925 ;
      RECT  23.005 44.0125 23.075 43.8775 ;
      RECT  22.9425 44.295 22.9975 44.2425 ;
      RECT  23.0975 42.9925 23.1675 42.8575 ;
      RECT  22.755 44.3 22.815 44.2425 ;
      RECT  23.455 43.52 23.525 43.385 ;
      RECT  22.7175 44.305 22.8525 44.235 ;
      RECT  23.2775 44.3025 23.335 44.2425 ;
      RECT  23.27 44.37 23.34 42.825 ;
      RECT  23.46 44.245 23.52 44.3025 ;
      RECT  22.75 45.02 22.82 45.155 ;
      RECT  22.935 44.17 23.005 45.715 ;
      RECT  23.4225 44.235 23.5575 44.305 ;
      RECT  23.455 44.17 23.525 45.715 ;
      RECT  22.75 44.17 22.82 45.715 ;
      RECT  23.2 44.5275 23.27 44.6625 ;
      RECT  23.455 44.2375 23.525 45.6475 ;
      RECT  23.005 44.5275 23.075 44.6625 ;
      RECT  22.9425 44.245 22.9975 44.2975 ;
      RECT  23.0975 45.5475 23.1675 45.6825 ;
      RECT  22.755 44.24 22.815 44.2975 ;
      RECT  23.455 45.02 23.525 45.155 ;
      RECT  22.7175 44.235 22.8525 44.305 ;
      RECT  23.2775 44.2375 23.335 44.2975 ;
      RECT  23.27 44.17 23.34 45.715 ;
      RECT  23.0975 29.4075 23.1675 29.5425 ;
      RECT  23.0975 32.0975 23.1675 32.2325 ;
      RECT  23.0975 32.0975 23.1675 32.2325 ;
      RECT  23.0975 45.5475 23.1675 45.6825 ;
      RECT  23.0975 26.7175 23.1675 26.8525 ;
      RECT  23.0975 21.3375 23.1675 21.4725 ;
      RECT  23.0975 24.0275 23.1675 24.1625 ;
      RECT  23.0975 24.0275 23.1675 24.1625 ;
      RECT  23.0975 21.3375 23.1675 21.4725 ;
      RECT  23.0975 26.7175 23.1675 26.8525 ;
      RECT  23.0975 42.8575 23.1675 42.9925 ;
      RECT  23.0975 37.4775 23.1675 37.6125 ;
      RECT  23.0975 40.1675 23.1675 40.3025 ;
      RECT  23.0975 40.1675 23.1675 40.3025 ;
      RECT  23.0975 34.7875 23.1675 34.9225 ;
      RECT  22.7175 41.545 22.8525 41.615 ;
      RECT  22.7175 30.785 22.8525 30.855 ;
      RECT  22.7175 36.165 22.8525 36.235 ;
      RECT  22.7175 38.855 22.8525 38.925 ;
      RECT  22.7175 44.235 22.8525 44.305 ;
      RECT  22.7175 20.025 22.8525 20.095 ;
      RECT  22.7175 28.095 22.8525 28.165 ;
      RECT  22.7175 22.715 22.8525 22.785 ;
      RECT  22.7175 33.475 22.8525 33.545 ;
      RECT  22.7175 25.405 22.8525 25.475 ;
      RECT  20.82 20.06 20.89 45.615 ;
      RECT  21.155 20.06 21.225 45.615 ;
      RECT  21.525 20.06 21.595 45.615 ;
      RECT  21.86 20.06 21.93 45.615 ;
      RECT  22.23 20.06 22.3 45.615 ;
      RECT  22.565 20.06 22.635 45.615 ;
      RECT  20.9825 40.1675 21.0525 40.3025 ;
      RECT  20.9825 37.4775 21.0525 37.6125 ;
      RECT  20.9825 42.8575 21.0525 42.9925 ;
      RECT  20.9825 29.4075 21.0525 29.5425 ;
      RECT  20.9825 24.0275 21.0525 24.1625 ;
      RECT  20.9825 34.7875 21.0525 34.9225 ;
      RECT  20.9825 26.7175 21.0525 26.8525 ;
      RECT  20.9825 32.0975 21.0525 32.2325 ;
      RECT  20.9825 21.3375 21.0525 21.4725 ;
      RECT  20.6025 33.475 20.7375 33.545 ;
      RECT  20.6025 36.165 20.7375 36.235 ;
      RECT  20.6025 28.095 20.7375 28.165 ;
      RECT  20.6025 44.235 20.7375 44.305 ;
      RECT  20.6025 25.405 20.7375 25.475 ;
      RECT  20.6025 30.785 20.7375 30.855 ;
      RECT  20.6025 22.715 20.7375 22.785 ;
      RECT  20.6025 38.855 20.7375 38.925 ;
      RECT  20.6025 41.545 20.7375 41.615 ;
      RECT  20.775 18.215 20.845 19.555 ;
      RECT  21.2 18.215 21.27 19.555 ;
      RECT  21.48 18.215 21.55 19.555 ;
      RECT  21.905 18.215 21.975 19.555 ;
      RECT  22.185 18.215 22.255 19.555 ;
      RECT  22.61 18.215 22.68 19.555 ;
      RECT  20.775 18.215 20.845 19.555 ;
      RECT  21.2 18.215 21.27 19.555 ;
      RECT  21.48 18.215 21.55 19.555 ;
      RECT  21.905 18.215 21.975 19.555 ;
      RECT  22.185 18.215 22.255 19.555 ;
      RECT  22.61 18.215 22.68 19.555 ;
      RECT  21.86 12.825 21.93 17.71 ;
      RECT  21.8825 14.545 21.9525 14.68 ;
      RECT  21.5 14.135 21.57 14.27 ;
      RECT  21.6925 13.425 21.7625 15.435 ;
      RECT  21.6925 15.435 21.7625 15.57 ;
      RECT  21.6925 13.2925 21.7625 13.4275 ;
      RECT  22.045 17.3275 22.115 17.4625 ;
      RECT  21.525 12.825 21.595 17.71 ;
      RECT  21.375 12.825 21.445 13.2225 ;
      RECT  22.565 12.825 22.635 17.71 ;
      RECT  22.5875 14.545 22.6575 14.68 ;
      RECT  22.205 14.135 22.275 14.27 ;
      RECT  22.3975 13.425 22.4675 15.435 ;
      RECT  22.3975 15.435 22.4675 15.57 ;
      RECT  22.3975 13.2925 22.4675 13.4275 ;
      RECT  22.75 17.3275 22.82 17.4625 ;
      RECT  22.23 12.825 22.3 17.71 ;
      RECT  22.08 12.825 22.15 13.2225 ;
      RECT  21.375 12.825 21.445 13.2225 ;
      RECT  21.525 12.825 21.595 17.71 ;
      RECT  21.86 12.825 21.93 17.71 ;
      RECT  22.08 12.825 22.15 13.2225 ;
      RECT  22.23 12.825 22.3 17.71 ;
      RECT  22.565 12.825 22.635 17.71 ;
      RECT  21.48 8.61 21.55 10.93 ;
      RECT  21.76 9.515 21.83 9.65 ;
      RECT  21.62 9.24 21.69 9.515 ;
      RECT  21.34 11.8075 21.41 11.9425 ;
      RECT  21.79 9.88 21.86 10.015 ;
      RECT  21.79 10.395 21.86 10.53 ;
      RECT  22.045 9.88 22.115 10.015 ;
      RECT  21.62 9.515 21.69 11.6125 ;
      RECT  21.76 9.105 21.83 9.24 ;
      RECT  21.34 9.88 21.41 10.015 ;
      RECT  21.48 8.54 21.615 8.61 ;
      RECT  21.5825 8.2775 21.7175 8.3475 ;
      RECT  21.34 9.515 21.41 9.65 ;
      RECT  22.045 9.31 22.115 11.9425 ;
      RECT  21.76 9.24 21.83 9.515 ;
      RECT  21.525 12.0175 21.595 12.1525 ;
      RECT  21.62 11.485 21.69 11.62 ;
      RECT  21.86 9.88 21.93 12.32 ;
      RECT  21.525 12.02 21.595 12.32 ;
      RECT  21.5325 8.2775 21.725 8.3475 ;
      RECT  21.62 9.105 21.69 9.24 ;
      RECT  21.48 10.795 21.55 10.93 ;
      RECT  22.045 11.8075 22.115 11.9425 ;
      RECT  21.655 8.145 21.725 8.285 ;
      RECT  21.34 9.31 21.41 9.445 ;
      RECT  21.34 9.3075 21.41 11.9425 ;
      RECT  21.62 9.515 21.69 9.65 ;
      RECT  22.045 9.515 22.115 9.65 ;
      RECT  22.045 9.31 22.115 9.445 ;
      RECT  22.185 8.61 22.255 10.93 ;
      RECT  22.465 9.515 22.535 9.65 ;
      RECT  22.325 9.24 22.395 9.515 ;
      RECT  22.045 11.8075 22.115 11.9425 ;
      RECT  22.495 9.88 22.565 10.015 ;
      RECT  22.495 10.395 22.565 10.53 ;
      RECT  22.75 9.88 22.82 10.015 ;
      RECT  22.325 9.515 22.395 11.6125 ;
      RECT  22.465 9.105 22.535 9.24 ;
      RECT  22.045 9.88 22.115 10.015 ;
      RECT  22.185 8.54 22.32 8.61 ;
      RECT  22.2875 8.2775 22.4225 8.3475 ;
      RECT  22.045 9.515 22.115 9.65 ;
      RECT  22.75 9.31 22.82 11.9425 ;
      RECT  22.465 9.24 22.535 9.515 ;
      RECT  22.23 12.0175 22.3 12.1525 ;
      RECT  22.325 11.485 22.395 11.62 ;
      RECT  22.565 9.88 22.635 12.32 ;
      RECT  22.23 12.02 22.3 12.32 ;
      RECT  22.2375 8.2775 22.43 8.3475 ;
      RECT  22.325 9.105 22.395 9.24 ;
      RECT  22.185 10.795 22.255 10.93 ;
      RECT  22.75 11.8075 22.82 11.9425 ;
      RECT  22.36 8.145 22.43 8.285 ;
      RECT  22.045 9.31 22.115 9.445 ;
      RECT  22.045 9.3075 22.115 11.9425 ;
      RECT  22.325 9.515 22.395 9.65 ;
      RECT  22.75 9.515 22.82 9.65 ;
      RECT  22.75 9.31 22.82 9.445 ;
      RECT  21.655 8.145 21.725 8.285 ;
      RECT  22.36 8.145 22.43 8.285 ;
      RECT  21.525 12.02 21.595 12.32 ;
      RECT  21.86 9.88 21.93 12.32 ;
      RECT  22.23 12.02 22.3 12.32 ;
      RECT  22.565 9.88 22.635 12.32 ;
      RECT  20.775 19.555 20.845 18.215 ;
      RECT  21.2 19.555 21.27 18.215 ;
      RECT  21.48 19.555 21.55 18.215 ;
      RECT  21.905 19.555 21.975 18.215 ;
      RECT  22.185 19.555 22.255 18.215 ;
      RECT  22.61 19.555 22.68 18.215 ;
      RECT  21.375 13.2225 21.445 12.825 ;
      RECT  22.08 13.2225 22.15 12.825 ;
      RECT  21.655 8.285 21.725 8.145 ;
      RECT  22.36 8.285 22.43 8.145 ;
      RECT  10.75 23.31 10.82 23.445 ;
      RECT  10.89 24.745 10.96 24.88 ;
      RECT  10.75 31.38 10.82 31.515 ;
      RECT  10.89 32.815 10.96 32.95 ;
      RECT  9.98 22.75 10.05 36.2 ;
      RECT  10.12 22.75 10.19 36.2 ;
      RECT  10.26 22.75 10.33 36.2 ;
      RECT  10.4 22.75 10.47 36.2 ;
      RECT  17.55 22.75 17.62 44.27 ;
      RECT  9.98 22.75 10.05 36.2 ;
      RECT  10.12 22.75 10.19 36.2 ;
      RECT  10.26 22.75 10.33 36.2 ;
      RECT  10.4 22.75 10.47 36.2 ;
      RECT  18.0875 22.0875 18.1575 22.1575 ;
      RECT  21.375 12.825 21.445 13.2225 ;
      RECT  22.08 12.825 22.15 13.2225 ;
      RECT  21.655 8.145 21.725 8.285 ;
      RECT  22.36 8.145 22.43 8.285 ;
      RECT  9.98 22.75 10.05 36.2 ;
      RECT  10.12 22.75 10.19 36.2 ;
      RECT  10.26 22.75 10.33 36.2 ;
      RECT  10.4 22.75 10.47 36.2 ;
      RECT  18.93 8.145 19.0 20.06 ;
      RECT  19.21 8.145 19.28 20.06 ;
      RECT  19.07 8.145 19.14 20.06 ;
      RECT  19.35 8.145 19.42 20.06 ;
      RECT  2.0475 0.5875 2.1175 1.1925 ;
      RECT  2.6325 1.0475 2.71 1.1825 ;
      RECT  0.245 1.0375 0.3225 1.1725 ;
      RECT  1.82 1.0375 1.8975 1.1725 ;
      POLYGON  2.3225 1.9925 2.3225 2.1975 1.9775 2.1975 1.9775 2.2675 2.3925 2.2675 2.3925 1.9925 2.3225 1.9925 ;
      POLYGON  1.2075 1.4275 1.2075 1.7025 1.2225 1.7025 1.2225 1.9975 1.2925 1.9975 1.2925 1.4275 1.2075 1.4275 ;
      POLYGON  2.3325 1.4825 2.3325 1.7775 2.3275 1.7775 2.3275 1.9125 2.4025 1.9125 2.4025 1.4825 2.3325 1.4825 ;
      RECT  0.245 1.0375 0.3225 1.1725 ;
      RECT  4.4 0.7025 4.47 0.7725 ;
      RECT  3.705 1.5225 3.775 1.5925 ;
      RECT  1.82 1.0375 1.8975 1.1725 ;
      RECT  2.0475 4.3625 2.1175 3.7575 ;
      RECT  2.6325 3.9025 2.71 3.7675 ;
      RECT  0.245 3.9125 0.3225 3.7775 ;
      RECT  1.82 3.9125 1.8975 3.7775 ;
      POLYGON  2.3225 2.9575 2.3225 2.7525 1.9775 2.7525 1.9775 2.6825 2.3925 2.6825 2.3925 2.9575 2.3225 2.9575 ;
      POLYGON  1.2075 3.5225 1.2075 3.2475 1.2225 3.2475 1.2225 2.9525 1.2925 2.9525 1.2925 3.5225 1.2075 3.5225 ;
      POLYGON  2.3325 3.4675 2.3325 3.1725 2.3275 3.1725 2.3275 3.0375 2.4025 3.0375 2.4025 3.4675 2.3325 3.4675 ;
      RECT  0.245 3.9125 0.3225 3.7775 ;
      RECT  4.4 4.2475 4.47 4.1775 ;
      RECT  3.705 3.4275 3.775 3.3575 ;
      RECT  1.82 3.9125 1.8975 3.7775 ;
      RECT  0.245 1.0375 0.3225 1.1725 ;
      RECT  0.245 3.7775 0.3225 3.9125 ;
      RECT  4.4 0.7025 4.47 0.7725 ;
      RECT  3.705 1.5225 3.775 1.5925 ;
      RECT  4.4 4.1775 4.47 4.2475 ;
      RECT  3.705 3.3575 3.775 3.4275 ;
      RECT  1.82 0.0 1.89 4.95 ;
      RECT  3.365 20.06 3.295 20.925 ;
      RECT  0.3725 20.06 0.3025 35.485 ;
      RECT  0.245 1.0375 0.3225 1.1725 ;
      RECT  0.245 3.7775 0.3225 3.9125 ;
      RECT  6.155 1.1575 6.225 1.2275 ;
      RECT  3.295 20.06 3.365 20.925 ;
      RECT  7.3875 18.6175 9.6675 18.6875 ;
      RECT  7.6775 10.9525 9.6675 11.0225 ;
      RECT  8.0125 13.6225 9.6675 13.6925 ;
      RECT  8.07 8.74 9.6675 8.81 ;
      RECT  8.88 1.0675 9.6675 1.1375 ;
      RECT  8.855 37.2875 8.925 37.8925 ;
      RECT  9.44 37.7475 9.5175 37.8825 ;
      RECT  7.0525 37.7375 7.13 37.8725 ;
      RECT  8.6275 37.7375 8.705 37.8725 ;
      POLYGON  9.13 38.6925 9.13 38.8975 8.785 38.8975 8.785 38.9675 9.2 38.9675 9.2 38.6925 9.13 38.6925 ;
      POLYGON  8.015 38.1275 8.015 38.4025 8.03 38.4025 8.03 38.6975 8.1 38.6975 8.1 38.1275 8.015 38.1275 ;
      POLYGON  9.14 38.1825 9.14 38.4775 9.135 38.4775 9.135 38.6125 9.21 38.6125 9.21 38.1825 9.14 38.1825 ;
      RECT  8.855 41.0625 8.925 40.4575 ;
      RECT  9.44 40.6025 9.5175 40.4675 ;
      RECT  7.0525 40.6125 7.13 40.4775 ;
      RECT  8.6275 40.6125 8.705 40.4775 ;
      POLYGON  9.13 39.6575 9.13 39.4525 8.785 39.4525 8.785 39.3825 9.2 39.3825 9.2 39.6575 9.13 39.6575 ;
      POLYGON  8.015 40.2225 8.015 39.9475 8.03 39.9475 8.03 39.6525 8.1 39.6525 8.1 40.2225 8.015 40.2225 ;
      POLYGON  9.14 40.1675 9.14 39.8725 9.135 39.8725 9.135 39.7375 9.21 39.7375 9.21 40.1675 9.14 40.1675 ;
      RECT  8.855 42.2375 8.925 42.8425 ;
      RECT  9.44 42.6975 9.5175 42.8325 ;
      RECT  7.0525 42.6875 7.13 42.8225 ;
      RECT  8.6275 42.6875 8.705 42.8225 ;
      POLYGON  9.13 43.6425 9.13 43.8475 8.785 43.8475 8.785 43.9175 9.2 43.9175 9.2 43.6425 9.13 43.6425 ;
      POLYGON  8.015 43.0775 8.015 43.3525 8.03 43.3525 8.03 43.6475 8.1 43.6475 8.1 43.0775 8.015 43.0775 ;
      POLYGON  9.14 43.1325 9.14 43.4275 9.135 43.4275 9.135 43.5625 9.21 43.5625 9.21 43.1325 9.14 43.1325 ;
      RECT  8.855 46.0125 8.925 45.4075 ;
      RECT  9.44 45.5525 9.5175 45.4175 ;
      RECT  7.0525 45.5625 7.13 45.4275 ;
      RECT  8.6275 45.5625 8.705 45.4275 ;
      POLYGON  9.13 44.6075 9.13 44.4025 8.785 44.4025 8.785 44.3325 9.2 44.3325 9.2 44.6075 9.13 44.6075 ;
      POLYGON  8.015 45.1725 8.015 44.8975 8.03 44.8975 8.03 44.6025 8.1 44.6025 8.1 45.1725 8.015 45.1725 ;
      POLYGON  9.14 45.1175 9.14 44.8225 9.135 44.8225 9.135 44.6875 9.21 44.6875 9.21 45.1175 9.14 45.1175 ;
      RECT  7.0525 37.7375 7.13 37.8725 ;
      RECT  7.0525 40.4775 7.13 40.6125 ;
      RECT  7.0525 42.6875 7.13 42.8225 ;
      RECT  7.0525 45.4275 7.13 45.5625 ;
      RECT  9.44 37.7475 9.5175 37.8825 ;
      RECT  9.44 40.4675 9.5175 40.6025 ;
      RECT  9.44 42.6975 9.5175 42.8325 ;
      RECT  9.44 45.4175 9.5175 45.5525 ;
      RECT  14.575 0.5875 14.645 1.1925 ;
      RECT  15.16 1.0475 15.2375 1.1825 ;
      RECT  12.7725 1.0375 12.85 1.1725 ;
      RECT  14.3475 1.0375 14.425 1.1725 ;
      POLYGON  14.85 1.9925 14.85 2.1975 14.505 2.1975 14.505 2.2675 14.92 2.2675 14.92 1.9925 14.85 1.9925 ;
      POLYGON  13.735 1.4275 13.735 1.7025 13.75 1.7025 13.75 1.9975 13.82 1.9975 13.82 1.4275 13.735 1.4275 ;
      POLYGON  14.86 1.4825 14.86 1.7775 14.855 1.7775 14.855 1.9125 14.93 1.9125 14.93 1.4825 14.86 1.4825 ;
      RECT  17.435 0.5875 17.505 1.1925 ;
      RECT  18.02 1.0475 18.0975 1.1825 ;
      RECT  15.6325 1.0375 15.71 1.1725 ;
      RECT  17.2075 1.0375 17.285 1.1725 ;
      POLYGON  17.71 1.9925 17.71 2.1975 17.365 2.1975 17.365 2.2675 17.78 2.2675 17.78 1.9925 17.71 1.9925 ;
      POLYGON  16.595 1.4275 16.595 1.7025 16.61 1.7025 16.61 1.9975 16.68 1.9975 16.68 1.4275 16.595 1.4275 ;
      POLYGON  17.72 1.4825 17.72 1.7775 17.715 1.7775 17.715 1.9125 17.79 1.9125 17.79 1.4825 17.72 1.4825 ;
      RECT  12.7725 1.0375 12.85 1.1725 ;
      RECT  15.6325 1.0375 15.71 1.1725 ;
      RECT  15.16 1.0475 15.2375 1.1825 ;
      RECT  18.02 1.0475 18.0975 1.1825 ;
   LAYER  metal3 ;
      RECT  20.95 21.3375 21.085 21.4725 ;
      RECT  20.95 45.5475 21.085 45.6825 ;
      RECT  20.6025 19.9925 20.7375 20.1275 ;
      RECT  20.6025 44.2025 20.7375 44.3375 ;
      RECT  20.245 26.7175 20.38 26.8525 ;
      RECT  20.245 45.5475 20.38 45.6825 ;
      RECT  23.065 37.4775 23.2 37.6125 ;
      RECT  21.655 21.3375 21.79 21.4725 ;
      RECT  20.245 40.1675 20.38 40.3025 ;
      RECT  23.065 42.8575 23.2 42.9925 ;
      RECT  22.36 21.3375 22.495 21.4725 ;
      RECT  23.065 40.1675 23.2 40.3025 ;
      RECT  20.245 24.0275 20.38 24.1625 ;
      RECT  20.245 34.7875 20.38 34.9225 ;
      RECT  21.655 45.5475 21.79 45.6825 ;
      RECT  23.065 45.5475 23.2 45.6825 ;
      RECT  23.065 34.7875 23.2 34.9225 ;
      RECT  20.245 29.4075 20.38 29.5425 ;
      RECT  20.245 42.8575 20.38 42.9925 ;
      RECT  20.95 45.5475 21.085 45.6825 ;
      RECT  23.065 21.3375 23.2 21.4725 ;
      RECT  20.245 37.4775 20.38 37.6125 ;
      RECT  23.065 32.0975 23.2 32.2325 ;
      RECT  20.95 21.3375 21.085 21.4725 ;
      RECT  23.065 26.7175 23.2 26.8525 ;
      RECT  23.065 24.0275 23.2 24.1625 ;
      RECT  22.36 45.5475 22.495 45.6825 ;
      RECT  20.245 32.0975 20.38 32.2325 ;
      RECT  20.245 21.3375 20.38 21.4725 ;
      RECT  23.065 29.4075 23.2 29.5425 ;
      RECT  19.8975 41.5125 20.0325 41.6475 ;
      RECT  23.6175 20.165 23.7525 20.235 ;
      RECT  22.7175 28.0625 22.8525 28.1975 ;
      RECT  22.7175 19.9925 22.8525 20.1275 ;
      RECT  19.8975 19.9925 20.0325 20.1275 ;
      RECT  23.6175 44.375 23.7525 44.445 ;
      RECT  19.7025 20.165 19.8375 20.235 ;
      RECT  22.7175 38.8225 22.8525 38.9575 ;
      RECT  19.8975 22.6825 20.0325 22.8175 ;
      RECT  22.7175 41.5125 22.8525 41.6475 ;
      RECT  22.0125 19.9925 22.1475 20.1275 ;
      RECT  21.3075 44.2025 21.4425 44.3375 ;
      RECT  19.8975 36.1325 20.0325 36.2675 ;
      RECT  22.7175 25.3725 22.8525 25.5075 ;
      RECT  19.8975 30.7525 20.0325 30.8875 ;
      RECT  19.8975 38.8225 20.0325 38.9575 ;
      RECT  22.7175 22.6825 22.8525 22.8175 ;
      RECT  19.8975 33.4425 20.0325 33.5775 ;
      RECT  19.8975 44.2025 20.0325 44.3375 ;
      RECT  22.7175 30.7525 22.8525 30.8875 ;
      RECT  19.8975 25.3725 20.0325 25.5075 ;
      RECT  21.3075 19.9925 21.4425 20.1275 ;
      RECT  19.8975 28.0625 20.0325 28.1975 ;
      RECT  22.7175 44.2025 22.8525 44.3375 ;
      RECT  20.6025 19.9925 20.7375 20.1275 ;
      RECT  22.7175 33.4425 22.8525 33.5775 ;
      RECT  20.6025 44.2025 20.7375 44.3375 ;
      RECT  22.7175 36.1325 22.8525 36.2675 ;
      RECT  19.7025 44.375 19.8375 44.445 ;
      RECT  22.0125 44.2025 22.1475 44.3375 ;
      RECT  21.0075 19.3325 21.0775 19.4675 ;
      RECT  21.7125 19.3325 21.7825 19.4675 ;
      RECT  22.4175 19.3325 22.4875 19.4675 ;
      RECT  21.0075 19.3325 21.0775 19.4675 ;
      RECT  22.4175 19.3325 22.4875 19.4675 ;
      RECT  21.7125 19.3325 21.7825 19.4675 ;
      RECT  21.6925 13.2925 21.7625 13.4275 ;
      RECT  22.3975 13.2925 22.4675 13.4275 ;
      RECT  22.75 17.3275 22.82 17.4625 ;
      RECT  22.045 17.3275 22.115 17.4625 ;
      RECT  21.5125 8.5075 21.5825 8.6425 ;
      RECT  22.2175 8.5075 22.2875 8.6425 ;
      RECT  22.045 10.5575 22.115 10.6925 ;
      RECT  21.34 10.5575 21.41 10.6925 ;
      RECT  22.2175 8.6425 22.2875 8.5075 ;
      RECT  21.5125 8.6425 21.5825 8.5075 ;
      RECT  22.3975 13.4275 22.4675 13.2925 ;
      RECT  21.6925 13.4275 21.7625 13.2925 ;
      RECT  22.4175 19.4675 22.4875 19.3325 ;
      RECT  21.0075 19.4675 21.0775 19.3325 ;
      RECT  21.7125 19.4675 21.7825 19.3325 ;
      RECT  22.75 17.4625 22.82 17.3275 ;
      RECT  21.34 10.6925 21.41 10.5575 ;
      RECT  22.045 10.6925 22.115 10.5575 ;
      RECT  22.045 17.4625 22.115 17.3275 ;
      RECT  12.56 24.0275 12.695 24.1625 ;
      RECT  11.0325 26.7175 11.1675 26.8525 ;
      RECT  11.0325 24.0275 11.1675 24.1625 ;
      RECT  12.56 26.7175 12.695 26.8525 ;
      RECT  12.56 25.3725 12.695 25.5075 ;
      RECT  11.0325 22.6825 11.1675 22.8175 ;
      RECT  11.0325 25.3725 11.1675 25.5075 ;
      RECT  12.56 22.6825 12.695 22.8175 ;
      RECT  11.0325 28.0625 11.1675 28.1975 ;
      RECT  12.56 28.0625 12.695 28.1975 ;
      RECT  12.56 32.0975 12.695 32.2325 ;
      RECT  11.0325 34.7875 11.1675 34.9225 ;
      RECT  11.0325 32.0975 11.1675 32.2325 ;
      RECT  12.56 34.7875 12.695 34.9225 ;
      RECT  12.56 33.4425 12.695 33.5775 ;
      RECT  11.0325 30.7525 11.1675 30.8875 ;
      RECT  11.0325 33.4425 11.1675 33.5775 ;
      RECT  12.56 30.7525 12.695 30.8875 ;
      RECT  11.0325 36.1325 11.1675 36.2675 ;
      RECT  12.56 36.1325 12.695 36.2675 ;
      RECT  12.56 32.0975 12.695 32.2325 ;
      RECT  11.0325 26.7175 11.1675 26.8525 ;
      RECT  11.0325 34.7875 11.1675 34.9225 ;
      RECT  11.0325 32.0975 11.1675 32.2325 ;
      RECT  17.1025 40.1675 17.2375 40.3025 ;
      RECT  17.1025 26.7175 17.2375 26.8525 ;
      RECT  11.0325 24.0275 11.1675 24.1625 ;
      RECT  12.56 26.7175 12.695 26.8525 ;
      RECT  17.1025 29.4075 17.2375 29.5425 ;
      RECT  17.1025 29.4075 17.2375 29.5425 ;
      RECT  12.56 24.0275 12.695 24.1625 ;
      RECT  17.1025 32.0975 17.2375 32.2325 ;
      RECT  17.1025 37.4775 17.2375 37.6125 ;
      RECT  17.1025 34.7875 17.2375 34.9225 ;
      RECT  12.56 34.7875 12.695 34.9225 ;
      RECT  17.1025 24.0275 17.2375 24.1625 ;
      RECT  17.1025 42.8575 17.2375 42.9925 ;
      RECT  17.1025 42.8575 17.2375 42.9925 ;
      RECT  17.1025 36.1325 17.2375 36.2675 ;
      RECT  11.0325 25.3725 11.1675 25.5075 ;
      RECT  12.56 36.1325 12.695 36.2675 ;
      RECT  11.0325 22.6825 11.1675 22.8175 ;
      RECT  17.1025 28.0625 17.2375 28.1975 ;
      RECT  17.1025 33.4425 17.2375 33.5775 ;
      RECT  12.56 33.4425 12.695 33.5775 ;
      RECT  17.1025 22.6825 17.2375 22.8175 ;
      RECT  17.1025 41.5125 17.2375 41.6475 ;
      RECT  11.0325 33.4425 11.1675 33.5775 ;
      RECT  11.0325 28.0625 11.1675 28.1975 ;
      RECT  11.0325 30.7525 11.1675 30.8875 ;
      RECT  17.1025 38.8225 17.2375 38.9575 ;
      RECT  17.1025 44.2025 17.2375 44.3375 ;
      RECT  17.1025 25.3725 17.2375 25.5075 ;
      RECT  12.56 30.7525 12.695 30.8875 ;
      RECT  12.56 25.3725 12.695 25.5075 ;
      RECT  17.1025 30.7525 17.2375 30.8875 ;
      RECT  12.56 28.0625 12.695 28.1975 ;
      RECT  11.0325 36.1325 11.1675 36.2675 ;
      RECT  12.56 22.6825 12.695 22.8175 ;
      RECT  18.6925 29.4075 18.8275 29.5425 ;
      RECT  18.6925 29.4075 18.8275 29.5425 ;
      RECT  18.6925 34.7875 18.8275 34.9225 ;
      RECT  18.6925 42.8575 18.8275 42.9925 ;
      RECT  18.6925 42.8575 18.8275 42.9925 ;
      RECT  18.6925 37.4775 18.8275 37.6125 ;
      RECT  18.6925 24.0275 18.8275 24.1625 ;
      RECT  18.6925 26.7175 18.8275 26.8525 ;
      RECT  18.6925 32.0975 18.8275 32.2325 ;
      RECT  18.6925 40.1675 18.8275 40.3025 ;
      RECT  18.6925 38.8225 18.8275 38.9575 ;
      RECT  18.6925 33.4425 18.8275 33.5775 ;
      RECT  18.6925 28.0625 18.8275 28.1975 ;
      RECT  18.6925 25.3725 18.8275 25.5075 ;
      RECT  18.6925 44.2025 18.8275 44.3375 ;
      RECT  18.6925 36.1325 18.8275 36.2675 ;
      RECT  18.6925 22.6825 18.8275 22.8175 ;
      RECT  18.6925 30.7525 18.8275 30.8875 ;
      RECT  18.6925 41.5125 18.8275 41.6475 ;
      RECT  11.0325 34.7875 11.1675 34.9225 ;
      RECT  18.6925 42.8575 18.8275 42.9925 ;
      RECT  18.6925 29.4075 18.8275 29.5425 ;
      RECT  18.6925 24.0275 18.8275 24.1625 ;
      RECT  12.56 34.7875 12.695 34.9225 ;
      RECT  18.6925 37.4775 18.8275 37.6125 ;
      RECT  17.1025 34.7875 17.2375 34.9225 ;
      RECT  12.56 24.0275 12.695 24.1625 ;
      RECT  11.0325 26.7175 11.1675 26.8525 ;
      RECT  18.6925 34.7875 18.8275 34.9225 ;
      RECT  18.6925 32.0975 18.8275 32.2325 ;
      RECT  18.6925 40.1675 18.8275 40.3025 ;
      RECT  12.56 26.7175 12.695 26.8525 ;
      RECT  12.56 32.0975 12.695 32.2325 ;
      RECT  17.1025 42.8575 17.2375 42.9925 ;
      RECT  17.1025 29.4075 17.2375 29.5425 ;
      RECT  18.6925 26.7175 18.8275 26.8525 ;
      RECT  17.915 21.3375 18.05 21.4725 ;
      RECT  17.1025 37.4775 17.2375 37.6125 ;
      RECT  17.1025 26.7175 17.2375 26.8525 ;
      RECT  17.1025 32.0975 17.2375 32.2325 ;
      RECT  17.1025 24.0275 17.2375 24.1625 ;
      RECT  17.1025 40.1675 17.2375 40.3025 ;
      RECT  11.0325 24.0275 11.1675 24.1625 ;
      RECT  11.0325 32.0975 11.1675 32.2325 ;
      RECT  12.56 22.6825 12.695 22.8175 ;
      RECT  12.56 36.1325 12.695 36.2675 ;
      RECT  11.0325 33.4425 11.1675 33.5775 ;
      RECT  18.6925 44.2025 18.8275 44.3375 ;
      RECT  17.1025 41.5125 17.2375 41.6475 ;
      RECT  17.1025 44.2025 17.2375 44.3375 ;
      RECT  11.0325 30.7525 11.1675 30.8875 ;
      RECT  18.6925 22.6825 18.8275 22.8175 ;
      RECT  18.6925 33.4425 18.8275 33.5775 ;
      RECT  12.56 25.3725 12.695 25.5075 ;
      RECT  12.56 33.4425 12.695 33.5775 ;
      RECT  12.56 28.0625 12.695 28.1975 ;
      RECT  17.1025 30.7525 17.2375 30.8875 ;
      RECT  18.6925 30.7525 18.8275 30.8875 ;
      RECT  12.56 30.7525 12.695 30.8875 ;
      RECT  11.0325 25.3725 11.1675 25.5075 ;
      RECT  18.6925 38.8225 18.8275 38.9575 ;
      RECT  17.1025 33.4425 17.2375 33.5775 ;
      RECT  17.1025 28.0625 17.2375 28.1975 ;
      RECT  17.1025 38.8225 17.2375 38.9575 ;
      RECT  11.0325 22.6825 11.1675 22.8175 ;
      RECT  18.6925 25.3725 18.8275 25.5075 ;
      RECT  17.1025 36.1325 17.2375 36.2675 ;
      RECT  11.0325 36.1325 11.1675 36.2675 ;
      RECT  18.6925 41.5125 18.8275 41.6475 ;
      RECT  17.1025 22.6825 17.2375 22.8175 ;
      RECT  17.1025 25.3725 17.2375 25.5075 ;
      RECT  11.0325 28.0625 11.1675 28.1975 ;
      RECT  18.6925 36.1325 18.8275 36.2675 ;
      RECT  18.6925 28.0625 18.8275 28.1975 ;
      RECT  9.9475 18.04 20.81 18.11 ;
      RECT  21.7125 19.3325 21.7825 19.4675 ;
      RECT  20.245 26.7175 20.38 26.8525 ;
      RECT  20.245 45.5475 20.38 45.6825 ;
      RECT  17.1025 32.0975 17.2375 32.2325 ;
      RECT  18.6925 26.7175 18.8275 26.8525 ;
      RECT  23.065 37.4775 23.2 37.6125 ;
      RECT  21.655 21.3375 21.79 21.4725 ;
      RECT  21.6925 13.2925 21.7625 13.4275 ;
      RECT  12.56 32.0975 12.695 32.2325 ;
      RECT  17.1025 29.4075 17.2375 29.5425 ;
      RECT  20.245 40.1675 20.38 40.3025 ;
      RECT  22.4175 19.3325 22.4875 19.4675 ;
      RECT  21.0075 19.3325 21.0775 19.4675 ;
      RECT  18.6925 32.0975 18.8275 32.2325 ;
      RECT  11.0325 34.7875 11.1675 34.9225 ;
      RECT  23.065 42.8575 23.2 42.9925 ;
      RECT  11.0325 32.0975 11.1675 32.2325 ;
      RECT  18.6925 40.1675 18.8275 40.3025 ;
      RECT  12.56 24.0275 12.695 24.1625 ;
      RECT  17.915 21.3375 18.05 21.4725 ;
      RECT  22.36 21.3375 22.495 21.4725 ;
      RECT  22.3975 13.2925 22.4675 13.4275 ;
      RECT  17.1025 34.7875 17.2375 34.9225 ;
      RECT  23.065 40.1675 23.2 40.3025 ;
      RECT  17.1025 40.1675 17.2375 40.3025 ;
      RECT  20.245 24.0275 20.38 24.1625 ;
      RECT  20.245 34.7875 20.38 34.9225 ;
      RECT  21.655 45.5475 21.79 45.6825 ;
      RECT  11.0325 24.0275 11.1675 24.1625 ;
      RECT  18.6925 37.4775 18.8275 37.6125 ;
      RECT  23.065 45.5475 23.2 45.6825 ;
      RECT  23.065 34.7875 23.2 34.9225 ;
      RECT  20.245 29.4075 20.38 29.5425 ;
      RECT  20.245 42.8575 20.38 42.9925 ;
      RECT  20.95 45.5475 21.085 45.6825 ;
      RECT  18.6925 42.8575 18.8275 42.9925 ;
      RECT  22.2175 8.5075 22.2875 8.6425 ;
      RECT  18.6925 24.0275 18.8275 24.1625 ;
      RECT  23.065 21.3375 23.2 21.4725 ;
      RECT  11.0325 26.7175 11.1675 26.8525 ;
      RECT  12.56 26.7175 12.695 26.8525 ;
      RECT  20.245 21.3375 20.38 21.4725 ;
      RECT  20.245 37.4775 20.38 37.6125 ;
      RECT  21.5125 8.5075 21.5825 8.6425 ;
      RECT  23.065 32.0975 23.2 32.2325 ;
      RECT  20.95 21.3375 21.085 21.4725 ;
      RECT  18.6925 29.4075 18.8275 29.5425 ;
      RECT  12.56 34.7875 12.695 34.9225 ;
      RECT  23.065 26.7175 23.2 26.8525 ;
      RECT  23.065 24.0275 23.2 24.1625 ;
      RECT  17.1025 26.7175 17.2375 26.8525 ;
      RECT  17.1025 24.0275 17.2375 24.1625 ;
      RECT  17.1025 37.4775 17.2375 37.6125 ;
      RECT  20.245 32.0975 20.38 32.2325 ;
      RECT  17.1025 42.8575 17.2375 42.9925 ;
      RECT  18.6925 34.7875 18.8275 34.9225 ;
      RECT  22.36 45.5475 22.495 45.6825 ;
      RECT  23.065 29.4075 23.2 29.5425 ;
      RECT  18.6925 44.2025 18.8275 44.3375 ;
      RECT  11.0325 30.7525 11.1675 30.8875 ;
      RECT  19.8975 41.5125 20.0325 41.6475 ;
      RECT  23.6175 20.165 23.7525 20.235 ;
      RECT  22.7175 28.0625 22.8525 28.1975 ;
      RECT  22.7175 19.9925 22.8525 20.1275 ;
      RECT  19.8975 19.9925 20.0325 20.1275 ;
      RECT  17.1025 30.7525 17.2375 30.8875 ;
      RECT  18.6925 36.1325 18.8275 36.2675 ;
      RECT  12.56 33.4425 12.695 33.5775 ;
      RECT  23.6175 44.375 23.7525 44.445 ;
      RECT  19.7025 20.165 19.8375 20.235 ;
      RECT  18.6925 30.7525 18.8275 30.8875 ;
      RECT  17.1025 28.0625 17.2375 28.1975 ;
      RECT  17.1025 25.3725 17.2375 25.5075 ;
      RECT  22.7175 38.8225 22.8525 38.9575 ;
      RECT  19.8975 22.6825 20.0325 22.8175 ;
      RECT  12.56 28.0625 12.695 28.1975 ;
      RECT  11.0325 28.0625 11.1675 28.1975 ;
      RECT  22.7175 41.5125 22.8525 41.6475 ;
      RECT  22.0125 19.9925 22.1475 20.1275 ;
      RECT  21.3075 44.2025 21.4425 44.3375 ;
      RECT  19.8975 36.1325 20.0325 36.2675 ;
      RECT  18.6925 28.0625 18.8275 28.1975 ;
      RECT  18.6925 25.3725 18.8275 25.5075 ;
      RECT  22.7175 25.3725 22.8525 25.5075 ;
      RECT  17.1025 36.1325 17.2375 36.2675 ;
      RECT  11.0325 36.1325 11.1675 36.2675 ;
      RECT  19.8975 30.7525 20.0325 30.8875 ;
      RECT  18.6925 22.6825 18.8275 22.8175 ;
      RECT  17.1025 44.2025 17.2375 44.3375 ;
      RECT  19.8975 38.8225 20.0325 38.9575 ;
      RECT  11.0325 22.6825 11.1675 22.8175 ;
      RECT  22.75 17.3275 22.82 17.4625 ;
      RECT  22.7175 22.6825 22.8525 22.8175 ;
      RECT  12.56 36.1325 12.695 36.2675 ;
      RECT  19.8975 33.4425 20.0325 33.5775 ;
      RECT  17.1025 22.6825 17.2375 22.8175 ;
      RECT  19.8975 44.2025 20.0325 44.3375 ;
      RECT  22.7175 30.7525 22.8525 30.8875 ;
      RECT  19.8975 25.3725 20.0325 25.5075 ;
      RECT  21.3075 19.9925 21.4425 20.1275 ;
      RECT  11.0325 25.3725 11.1675 25.5075 ;
      RECT  18.6925 33.4425 18.8275 33.5775 ;
      RECT  17.1025 38.8225 17.2375 38.9575 ;
      RECT  19.8975 28.0625 20.0325 28.1975 ;
      RECT  18.6925 41.5125 18.8275 41.6475 ;
      RECT  22.7175 44.2025 22.8525 44.3375 ;
      RECT  12.56 30.7525 12.695 30.8875 ;
      RECT  20.6025 19.9925 20.7375 20.1275 ;
      RECT  22.045 10.5575 22.115 10.6925 ;
      RECT  11.0325 33.4425 11.1675 33.5775 ;
      RECT  22.7175 33.4425 22.8525 33.5775 ;
      RECT  20.6025 44.2025 20.7375 44.3375 ;
      RECT  18.6925 38.8225 18.8275 38.9575 ;
      RECT  17.1025 33.4425 17.2375 33.5775 ;
      RECT  22.7175 36.1325 22.8525 36.2675 ;
      RECT  19.7025 44.375 19.8375 44.445 ;
      RECT  22.045 17.3275 22.115 17.4625 ;
      RECT  22.0125 44.2025 22.1475 44.3375 ;
      RECT  17.1025 41.5125 17.2375 41.6475 ;
      RECT  12.56 22.6825 12.695 22.8175 ;
      RECT  12.56 25.3725 12.695 25.5075 ;
      RECT  21.34 10.5575 21.41 10.6925 ;
      RECT  -0.0675 2.4125 0.0675 2.5475 ;
      RECT  -0.0675 2.4025 0.0675 2.5375 ;
      RECT  -0.0675 -0.0675 0.0675 0.0675 ;
      RECT  -0.0675 4.8825 0.0675 5.0175 ;
      RECT  2.26 29.0925 2.125 29.2275 ;
      RECT  2.26 25.4525 2.125 25.5875 ;
      RECT  2.26 29.0925 2.125 29.2275 ;
      RECT  2.26 36.3725 2.125 36.5075 ;
      RECT  0.885 36.3725 0.75 36.5075 ;
      RECT  0.885 21.8125 0.75 21.9475 ;
      RECT  2.26 32.7325 2.125 32.8675 ;
      RECT  2.26 21.8125 2.125 21.9475 ;
      RECT  0.885 29.0925 0.75 29.2275 ;
      RECT  0.885 29.0925 0.75 29.2275 ;
      RECT  0.885 32.7325 0.75 32.8675 ;
      RECT  0.885 25.4525 0.75 25.5875 ;
      RECT  2.26 23.6325 2.125 23.7675 ;
      RECT  0.885 27.2725 0.75 27.4075 ;
      RECT  0.885 19.9925 0.75 20.1275 ;
      RECT  2.26 27.2725 2.125 27.4075 ;
      RECT  0.885 34.5525 0.75 34.6875 ;
      RECT  0.885 23.6325 0.75 23.7675 ;
      RECT  2.26 19.9925 2.125 20.1275 ;
      RECT  0.885 30.9125 0.75 31.0475 ;
      RECT  2.26 30.9125 2.125 31.0475 ;
      RECT  2.26 34.5525 2.125 34.6875 ;
      RECT  0.75 25.4525 0.885 25.5875 ;
      RECT  9.46 7.3575 9.595 7.4925 ;
      RECT  9.46 2.4075 9.595 2.5425 ;
      RECT  9.46 7.3575 9.595 7.4925 ;
      RECT  9.46 2.4075 9.595 2.5425 ;
      RECT  2.125 36.3725 2.26 36.5075 ;
      RECT  0.75 32.7325 0.885 32.8675 ;
      RECT  -0.0675 2.4125 0.0675 2.5475 ;
      RECT  2.125 25.4525 2.26 25.5875 ;
      RECT  2.125 32.7325 2.26 32.8675 ;
      RECT  9.46 17.2575 9.595 17.3925 ;
      RECT  9.46 17.2575 9.595 17.3925 ;
      RECT  2.125 29.0925 2.26 29.2275 ;
      RECT  0.75 21.8125 0.885 21.9475 ;
      RECT  9.46 12.3075 9.595 12.4425 ;
      RECT  0.75 29.0925 0.885 29.2275 ;
      RECT  0.75 36.3725 0.885 36.5075 ;
      RECT  2.125 21.8125 2.26 21.9475 ;
      RECT  -0.0675 2.4025 0.0675 2.5375 ;
      RECT  9.46 -0.0675 9.595 0.0675 ;
      RECT  9.46 14.7825 9.595 14.9175 ;
      RECT  -0.0675 -0.0675 0.0675 0.0675 ;
      RECT  2.125 34.5525 2.26 34.6875 ;
      RECT  0.75 19.9925 0.885 20.1275 ;
      RECT  -0.0675 4.8825 0.0675 5.0175 ;
      RECT  9.46 4.8825 9.595 5.0175 ;
      RECT  0.75 23.6325 0.885 23.7675 ;
      RECT  2.125 23.6325 2.26 23.7675 ;
      RECT  0.75 27.2725 0.885 27.4075 ;
      RECT  9.46 9.8325 9.595 9.9675 ;
      RECT  2.125 19.9925 2.26 20.1275 ;
      RECT  0.75 30.9125 0.885 31.0475 ;
      RECT  2.125 27.2725 2.26 27.4075 ;
      RECT  2.125 30.9125 2.26 31.0475 ;
      RECT  9.46 19.7325 9.595 19.8675 ;
      RECT  0.75 34.5525 0.885 34.6875 ;
      RECT  6.8075 37.015 9.6675 37.085 ;
      RECT  8.12 39.1125 8.255 39.2475 ;
      RECT  8.12 44.0625 8.255 44.1975 ;
      RECT  8.12 39.1025 8.255 39.2375 ;
      RECT  8.12 44.0525 8.255 44.1875 ;
      RECT  8.17 41.5825 8.305 41.7175 ;
      RECT  8.17 46.5325 8.305 46.6675 ;
      RECT  8.17 36.6325 8.305 36.7675 ;
      RECT  12.5275 0.315 18.2475 0.385 ;
      RECT  16.7 2.4025 16.835 2.5375 ;
      RECT  13.84 2.4025 13.975 2.5375 ;
      RECT  16.75 -0.0675 16.885 0.0675 ;
      RECT  13.89 -0.0675 14.025 0.0675 ;
   LAYER  metal4 ;
   END
   END    sram_2_16_1_freepdk45
END    LIBRARY
