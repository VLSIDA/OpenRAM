magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1260 -1260 1326 1334
<< metal2 >>
rect 5 65 61 74
rect 5 0 61 9
<< via2 >>
rect 5 9 61 65
<< metal3 >>
rect 0 65 66 70
rect 0 9 5 65
rect 61 9 66 65
rect 0 4 66 9
<< properties >>
string FIXED_BBOX 0 0 66 74
<< end >>
