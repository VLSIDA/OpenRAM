VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 533700.0 by 1216800.0 ;
END  MacroSite
MACRO sram_1rw_8b_256w_1bank_scn3me_subm
   CLASS BLOCK ;
   SIZE 533700.0 BY 1216800.0 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN DATA[0]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  204600.0 600.0 205500.0 2400.0 ;
      END
   END DATA[0]
   PIN DATA[1]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  245400.0 600.0 246300.0 2400.0 ;
      END
   END DATA[1]
   PIN DATA[2]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  286200.0 600.0 287100.0 2400.0 ;
      END
   END DATA[2]
   PIN DATA[3]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  327000.0 600.0 327900.0 2400.0 ;
      END
   END DATA[3]
   PIN DATA[4]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  367800.0 600.0 368700.0 2400.0 ;
      END
   END DATA[4]
   PIN DATA[5]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  408600.0 600.0 409500.0 2400.0 ;
      END
   END DATA[5]
   PIN DATA[6]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  449400.0 600.0 450300.0 2400.0 ;
      END
   END DATA[6]
   PIN DATA[7]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  490200.0 600.0 491100.0 2400.0 ;
      END
   END DATA[7]
   PIN ADDR[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 136800.0 60000.0 138300.0 ;
      END
   END ADDR[0]
   PIN ADDR[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 126600.0 60000.0 128100.0 ;
      END
   END ADDR[1]
   PIN ADDR[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 116400.0 60000.0 117900.0 ;
      END
   END ADDR[2]
   PIN ADDR[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 106200.0 60000.0 107700.0 ;
      END
   END ADDR[3]
   PIN ADDR[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 96000.0 60000.0 97500.0 ;
      END
   END ADDR[4]
   PIN ADDR[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 85800.0 60000.0 87300.0 ;
      END
   END ADDR[5]
   PIN ADDR[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 75600.0 60000.0 77100.0 ;
      END
   END ADDR[6]
   PIN ADDR[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 65400.0 60000.0 66900.0 ;
      END
   END ADDR[7]
   PIN CSb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  14400.0 317700.0 16200.0 319500.0 ;
      END
   END CSb
   PIN WEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  24600.0 317700.0 26400.0 319500.0 ;
      END
   END WEb
   PIN OEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4200.0 317700.0 6000.0 319500.0 ;
      END
   END OEb
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER metal1 ;
         RECT  42600.0 316800.0 43800.0 320400.0 ;
      END
   END clk
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal1 ;
         RECT  529200.0 600.0 533700.0 1217400.0 ;
         LAYER metal1 ;
         RECT  52800.0 600.0 57300.0 1217400.0 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal2 ;
         RECT  172650.0 600.0 177150.0 1217400.0 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  54600.0 410250.0 55500.0 412950.0 ;
      RECT  107100.0 319950.0 108000.0 320850.0 ;
      RECT  107100.0 317550.0 108000.0 318450.0 ;
      RECT  105750.0 319950.0 107550.0 320850.0 ;
      RECT  107100.0 318000.0 108000.0 320400.0 ;
      RECT  107550.0 317550.0 109500.0 318450.0 ;
      RECT  172050.0 319950.0 172950.0 320850.0 ;
      RECT  172050.0 315450.0 172950.0 316350.0 ;
      RECT  145650.0 319950.0 172500.0 320850.0 ;
      RECT  172050.0 315900.0 172950.0 320400.0 ;
      RECT  172500.0 315450.0 199500.0 316350.0 ;
      RECT  107100.0 334350.0 108000.0 335250.0 ;
      RECT  107100.0 336750.0 108000.0 337650.0 ;
      RECT  105750.0 334350.0 107550.0 335250.0 ;
      RECT  107100.0 334800.0 108000.0 337200.0 ;
      RECT  107550.0 336750.0 109500.0 337650.0 ;
      RECT  172050.0 334350.0 172950.0 335250.0 ;
      RECT  172050.0 338850.0 172950.0 339750.0 ;
      RECT  145650.0 334350.0 172500.0 335250.0 ;
      RECT  172050.0 334800.0 172950.0 339300.0 ;
      RECT  172500.0 338850.0 199500.0 339750.0 ;
      RECT  107100.0 347550.0 108000.0 348450.0 ;
      RECT  107100.0 345150.0 108000.0 346050.0 ;
      RECT  105750.0 347550.0 107550.0 348450.0 ;
      RECT  107100.0 345600.0 108000.0 348000.0 ;
      RECT  107550.0 345150.0 109500.0 346050.0 ;
      RECT  172050.0 347550.0 172950.0 348450.0 ;
      RECT  172050.0 343050.0 172950.0 343950.0 ;
      RECT  145650.0 347550.0 172500.0 348450.0 ;
      RECT  172050.0 343500.0 172950.0 348000.0 ;
      RECT  172500.0 343050.0 199500.0 343950.0 ;
      RECT  107100.0 361950.0 108000.0 362850.0 ;
      RECT  107100.0 364350.0 108000.0 365250.0 ;
      RECT  105750.0 361950.0 107550.0 362850.0 ;
      RECT  107100.0 362400.0 108000.0 364800.0 ;
      RECT  107550.0 364350.0 109500.0 365250.0 ;
      RECT  172050.0 361950.0 172950.0 362850.0 ;
      RECT  172050.0 366450.0 172950.0 367350.0 ;
      RECT  145650.0 361950.0 172500.0 362850.0 ;
      RECT  172050.0 362400.0 172950.0 366900.0 ;
      RECT  172500.0 366450.0 199500.0 367350.0 ;
      RECT  107100.0 375150.0 108000.0 376050.0 ;
      RECT  107100.0 372750.0 108000.0 373650.0 ;
      RECT  105750.0 375150.0 107550.0 376050.0 ;
      RECT  107100.0 373200.0 108000.0 375600.0 ;
      RECT  107550.0 372750.0 109500.0 373650.0 ;
      RECT  172050.0 375150.0 172950.0 376050.0 ;
      RECT  172050.0 370650.0 172950.0 371550.0 ;
      RECT  145650.0 375150.0 172500.0 376050.0 ;
      RECT  172050.0 371100.0 172950.0 375600.0 ;
      RECT  172500.0 370650.0 199500.0 371550.0 ;
      RECT  107100.0 389550.0 108000.0 390450.0 ;
      RECT  107100.0 391950.0 108000.0 392850.0 ;
      RECT  105750.0 389550.0 107550.0 390450.0 ;
      RECT  107100.0 390000.0 108000.0 392400.0 ;
      RECT  107550.0 391950.0 109500.0 392850.0 ;
      RECT  172050.0 389550.0 172950.0 390450.0 ;
      RECT  172050.0 394050.0 172950.0 394950.0 ;
      RECT  145650.0 389550.0 172500.0 390450.0 ;
      RECT  172050.0 390000.0 172950.0 394500.0 ;
      RECT  172500.0 394050.0 199500.0 394950.0 ;
      RECT  107100.0 402750.0 108000.0 403650.0 ;
      RECT  107100.0 400350.0 108000.0 401250.0 ;
      RECT  105750.0 402750.0 107550.0 403650.0 ;
      RECT  107100.0 400800.0 108000.0 403200.0 ;
      RECT  107550.0 400350.0 109500.0 401250.0 ;
      RECT  172050.0 402750.0 172950.0 403650.0 ;
      RECT  172050.0 398250.0 172950.0 399150.0 ;
      RECT  145650.0 402750.0 172500.0 403650.0 ;
      RECT  172050.0 398700.0 172950.0 403200.0 ;
      RECT  172500.0 398250.0 199500.0 399150.0 ;
      RECT  107100.0 417150.0 108000.0 418050.0 ;
      RECT  107100.0 419550.0 108000.0 420450.0 ;
      RECT  105750.0 417150.0 107550.0 418050.0 ;
      RECT  107100.0 417600.0 108000.0 420000.0 ;
      RECT  107550.0 419550.0 109500.0 420450.0 ;
      RECT  172050.0 417150.0 172950.0 418050.0 ;
      RECT  172050.0 421650.0 172950.0 422550.0 ;
      RECT  145650.0 417150.0 172500.0 418050.0 ;
      RECT  172050.0 417600.0 172950.0 422100.0 ;
      RECT  172500.0 421650.0 199500.0 422550.0 ;
      RECT  107100.0 430350.0 108000.0 431250.0 ;
      RECT  107100.0 427950.0 108000.0 428850.0 ;
      RECT  105750.0 430350.0 107550.0 431250.0 ;
      RECT  107100.0 428400.0 108000.0 430800.0 ;
      RECT  107550.0 427950.0 109500.0 428850.0 ;
      RECT  172050.0 430350.0 172950.0 431250.0 ;
      RECT  172050.0 425850.0 172950.0 426750.0 ;
      RECT  145650.0 430350.0 172500.0 431250.0 ;
      RECT  172050.0 426300.0 172950.0 430800.0 ;
      RECT  172500.0 425850.0 199500.0 426750.0 ;
      RECT  107100.0 444750.0 108000.0 445650.0 ;
      RECT  107100.0 447150.0 108000.0 448050.0 ;
      RECT  105750.0 444750.0 107550.0 445650.0 ;
      RECT  107100.0 445200.0 108000.0 447600.0 ;
      RECT  107550.0 447150.0 109500.0 448050.0 ;
      RECT  172050.0 444750.0 172950.0 445650.0 ;
      RECT  172050.0 449250.0 172950.0 450150.0 ;
      RECT  145650.0 444750.0 172500.0 445650.0 ;
      RECT  172050.0 445200.0 172950.0 449700.0 ;
      RECT  172500.0 449250.0 199500.0 450150.0 ;
      RECT  107100.0 457950.0 108000.0 458850.0 ;
      RECT  107100.0 455550.0 108000.0 456450.0 ;
      RECT  105750.0 457950.0 107550.0 458850.0 ;
      RECT  107100.0 456000.0 108000.0 458400.0 ;
      RECT  107550.0 455550.0 109500.0 456450.0 ;
      RECT  172050.0 457950.0 172950.0 458850.0 ;
      RECT  172050.0 453450.0 172950.0 454350.0 ;
      RECT  145650.0 457950.0 172500.0 458850.0 ;
      RECT  172050.0 453900.0 172950.0 458400.0 ;
      RECT  172500.0 453450.0 199500.0 454350.0 ;
      RECT  107100.0 472350.0 108000.0 473250.0 ;
      RECT  107100.0 474750.0 108000.0 475650.0 ;
      RECT  105750.0 472350.0 107550.0 473250.0 ;
      RECT  107100.0 472800.0 108000.0 475200.0 ;
      RECT  107550.0 474750.0 109500.0 475650.0 ;
      RECT  172050.0 472350.0 172950.0 473250.0 ;
      RECT  172050.0 476850.0 172950.0 477750.0 ;
      RECT  145650.0 472350.0 172500.0 473250.0 ;
      RECT  172050.0 472800.0 172950.0 477300.0 ;
      RECT  172500.0 476850.0 199500.0 477750.0 ;
      RECT  107100.0 485550.0 108000.0 486450.0 ;
      RECT  107100.0 483150.0 108000.0 484050.0 ;
      RECT  105750.0 485550.0 107550.0 486450.0 ;
      RECT  107100.0 483600.0 108000.0 486000.0 ;
      RECT  107550.0 483150.0 109500.0 484050.0 ;
      RECT  172050.0 485550.0 172950.0 486450.0 ;
      RECT  172050.0 481050.0 172950.0 481950.0 ;
      RECT  145650.0 485550.0 172500.0 486450.0 ;
      RECT  172050.0 481500.0 172950.0 486000.0 ;
      RECT  172500.0 481050.0 199500.0 481950.0 ;
      RECT  107100.0 499950.0 108000.0 500850.0 ;
      RECT  107100.0 502350.0 108000.0 503250.0 ;
      RECT  105750.0 499950.0 107550.0 500850.0 ;
      RECT  107100.0 500400.0 108000.0 502800.0 ;
      RECT  107550.0 502350.0 109500.0 503250.0 ;
      RECT  172050.0 499950.0 172950.0 500850.0 ;
      RECT  172050.0 504450.0 172950.0 505350.0 ;
      RECT  145650.0 499950.0 172500.0 500850.0 ;
      RECT  172050.0 500400.0 172950.0 504900.0 ;
      RECT  172500.0 504450.0 199500.0 505350.0 ;
      RECT  107100.0 513150.0 108000.0 514050.0 ;
      RECT  107100.0 510750.0 108000.0 511650.0 ;
      RECT  105750.0 513150.0 107550.0 514050.0 ;
      RECT  107100.0 511200.0 108000.0 513600.0 ;
      RECT  107550.0 510750.0 109500.0 511650.0 ;
      RECT  172050.0 513150.0 172950.0 514050.0 ;
      RECT  172050.0 508650.0 172950.0 509550.0 ;
      RECT  145650.0 513150.0 172500.0 514050.0 ;
      RECT  172050.0 509100.0 172950.0 513600.0 ;
      RECT  172500.0 508650.0 199500.0 509550.0 ;
      RECT  107100.0 527550.0 108000.0 528450.0 ;
      RECT  107100.0 529950.0 108000.0 530850.0 ;
      RECT  105750.0 527550.0 107550.0 528450.0 ;
      RECT  107100.0 528000.0 108000.0 530400.0 ;
      RECT  107550.0 529950.0 109500.0 530850.0 ;
      RECT  172050.0 527550.0 172950.0 528450.0 ;
      RECT  172050.0 532050.0 172950.0 532950.0 ;
      RECT  145650.0 527550.0 172500.0 528450.0 ;
      RECT  172050.0 528000.0 172950.0 532500.0 ;
      RECT  172500.0 532050.0 199500.0 532950.0 ;
      RECT  107100.0 540750.0 108000.0 541650.0 ;
      RECT  107100.0 538350.0 108000.0 539250.0 ;
      RECT  105750.0 540750.0 107550.0 541650.0 ;
      RECT  107100.0 538800.0 108000.0 541200.0 ;
      RECT  107550.0 538350.0 109500.0 539250.0 ;
      RECT  172050.0 540750.0 172950.0 541650.0 ;
      RECT  172050.0 536250.0 172950.0 537150.0 ;
      RECT  145650.0 540750.0 172500.0 541650.0 ;
      RECT  172050.0 536700.0 172950.0 541200.0 ;
      RECT  172500.0 536250.0 199500.0 537150.0 ;
      RECT  107100.0 555150.0 108000.0 556050.0 ;
      RECT  107100.0 557550.0 108000.0 558450.0 ;
      RECT  105750.0 555150.0 107550.0 556050.0 ;
      RECT  107100.0 555600.0 108000.0 558000.0 ;
      RECT  107550.0 557550.0 109500.0 558450.0 ;
      RECT  172050.0 555150.0 172950.0 556050.0 ;
      RECT  172050.0 559650.0 172950.0 560550.0 ;
      RECT  145650.0 555150.0 172500.0 556050.0 ;
      RECT  172050.0 555600.0 172950.0 560100.0 ;
      RECT  172500.0 559650.0 199500.0 560550.0 ;
      RECT  107100.0 568350.0 108000.0 569250.0 ;
      RECT  107100.0 565950.0 108000.0 566850.0 ;
      RECT  105750.0 568350.0 107550.0 569250.0 ;
      RECT  107100.0 566400.0 108000.0 568800.0 ;
      RECT  107550.0 565950.0 109500.0 566850.0 ;
      RECT  172050.0 568350.0 172950.0 569250.0 ;
      RECT  172050.0 563850.0 172950.0 564750.0 ;
      RECT  145650.0 568350.0 172500.0 569250.0 ;
      RECT  172050.0 564300.0 172950.0 568800.0 ;
      RECT  172500.0 563850.0 199500.0 564750.0 ;
      RECT  107100.0 582750.0 108000.0 583650.0 ;
      RECT  107100.0 585150.0 108000.0 586050.0 ;
      RECT  105750.0 582750.0 107550.0 583650.0 ;
      RECT  107100.0 583200.0 108000.0 585600.0 ;
      RECT  107550.0 585150.0 109500.0 586050.0 ;
      RECT  172050.0 582750.0 172950.0 583650.0 ;
      RECT  172050.0 587250.0 172950.0 588150.0 ;
      RECT  145650.0 582750.0 172500.0 583650.0 ;
      RECT  172050.0 583200.0 172950.0 587700.0 ;
      RECT  172500.0 587250.0 199500.0 588150.0 ;
      RECT  107100.0 595950.0 108000.0 596850.0 ;
      RECT  107100.0 593550.0 108000.0 594450.0 ;
      RECT  105750.0 595950.0 107550.0 596850.0 ;
      RECT  107100.0 594000.0 108000.0 596400.0 ;
      RECT  107550.0 593550.0 109500.0 594450.0 ;
      RECT  172050.0 595950.0 172950.0 596850.0 ;
      RECT  172050.0 591450.0 172950.0 592350.0 ;
      RECT  145650.0 595950.0 172500.0 596850.0 ;
      RECT  172050.0 591900.0 172950.0 596400.0 ;
      RECT  172500.0 591450.0 199500.0 592350.0 ;
      RECT  107100.0 610350.0 108000.0 611250.0 ;
      RECT  107100.0 612750.0 108000.0 613650.0 ;
      RECT  105750.0 610350.0 107550.0 611250.0 ;
      RECT  107100.0 610800.0 108000.0 613200.0 ;
      RECT  107550.0 612750.0 109500.0 613650.0 ;
      RECT  172050.0 610350.0 172950.0 611250.0 ;
      RECT  172050.0 614850.0 172950.0 615750.0 ;
      RECT  145650.0 610350.0 172500.0 611250.0 ;
      RECT  172050.0 610800.0 172950.0 615300.0 ;
      RECT  172500.0 614850.0 199500.0 615750.0 ;
      RECT  107100.0 623550.0 108000.0 624450.0 ;
      RECT  107100.0 621150.0 108000.0 622050.0 ;
      RECT  105750.0 623550.0 107550.0 624450.0 ;
      RECT  107100.0 621600.0 108000.0 624000.0 ;
      RECT  107550.0 621150.0 109500.0 622050.0 ;
      RECT  172050.0 623550.0 172950.0 624450.0 ;
      RECT  172050.0 619050.0 172950.0 619950.0 ;
      RECT  145650.0 623550.0 172500.0 624450.0 ;
      RECT  172050.0 619500.0 172950.0 624000.0 ;
      RECT  172500.0 619050.0 199500.0 619950.0 ;
      RECT  107100.0 637950.0 108000.0 638850.0 ;
      RECT  107100.0 640350.0 108000.0 641250.0 ;
      RECT  105750.0 637950.0 107550.0 638850.0 ;
      RECT  107100.0 638400.0 108000.0 640800.0 ;
      RECT  107550.0 640350.0 109500.0 641250.0 ;
      RECT  172050.0 637950.0 172950.0 638850.0 ;
      RECT  172050.0 642450.0 172950.0 643350.0 ;
      RECT  145650.0 637950.0 172500.0 638850.0 ;
      RECT  172050.0 638400.0 172950.0 642900.0 ;
      RECT  172500.0 642450.0 199500.0 643350.0 ;
      RECT  107100.0 651150.0 108000.0 652050.0 ;
      RECT  107100.0 648750.0 108000.0 649650.0 ;
      RECT  105750.0 651150.0 107550.0 652050.0 ;
      RECT  107100.0 649200.0 108000.0 651600.0 ;
      RECT  107550.0 648750.0 109500.0 649650.0 ;
      RECT  172050.0 651150.0 172950.0 652050.0 ;
      RECT  172050.0 646650.0 172950.0 647550.0 ;
      RECT  145650.0 651150.0 172500.0 652050.0 ;
      RECT  172050.0 647100.0 172950.0 651600.0 ;
      RECT  172500.0 646650.0 199500.0 647550.0 ;
      RECT  107100.0 665550.0 108000.0 666450.0 ;
      RECT  107100.0 667950.0 108000.0 668850.0 ;
      RECT  105750.0 665550.0 107550.0 666450.0 ;
      RECT  107100.0 666000.0 108000.0 668400.0 ;
      RECT  107550.0 667950.0 109500.0 668850.0 ;
      RECT  172050.0 665550.0 172950.0 666450.0 ;
      RECT  172050.0 670050.0 172950.0 670950.0 ;
      RECT  145650.0 665550.0 172500.0 666450.0 ;
      RECT  172050.0 666000.0 172950.0 670500.0 ;
      RECT  172500.0 670050.0 199500.0 670950.0 ;
      RECT  107100.0 678750.0 108000.0 679650.0 ;
      RECT  107100.0 676350.0 108000.0 677250.0 ;
      RECT  105750.0 678750.0 107550.0 679650.0 ;
      RECT  107100.0 676800.0 108000.0 679200.0 ;
      RECT  107550.0 676350.0 109500.0 677250.0 ;
      RECT  172050.0 678750.0 172950.0 679650.0 ;
      RECT  172050.0 674250.0 172950.0 675150.0 ;
      RECT  145650.0 678750.0 172500.0 679650.0 ;
      RECT  172050.0 674700.0 172950.0 679200.0 ;
      RECT  172500.0 674250.0 199500.0 675150.0 ;
      RECT  107100.0 693150.0 108000.0 694050.0 ;
      RECT  107100.0 695550.0 108000.0 696450.0 ;
      RECT  105750.0 693150.0 107550.0 694050.0 ;
      RECT  107100.0 693600.0 108000.0 696000.0 ;
      RECT  107550.0 695550.0 109500.0 696450.0 ;
      RECT  172050.0 693150.0 172950.0 694050.0 ;
      RECT  172050.0 697650.0 172950.0 698550.0 ;
      RECT  145650.0 693150.0 172500.0 694050.0 ;
      RECT  172050.0 693600.0 172950.0 698100.0 ;
      RECT  172500.0 697650.0 199500.0 698550.0 ;
      RECT  107100.0 706350.0 108000.0 707250.0 ;
      RECT  107100.0 703950.0 108000.0 704850.0 ;
      RECT  105750.0 706350.0 107550.0 707250.0 ;
      RECT  107100.0 704400.0 108000.0 706800.0 ;
      RECT  107550.0 703950.0 109500.0 704850.0 ;
      RECT  172050.0 706350.0 172950.0 707250.0 ;
      RECT  172050.0 701850.0 172950.0 702750.0 ;
      RECT  145650.0 706350.0 172500.0 707250.0 ;
      RECT  172050.0 702300.0 172950.0 706800.0 ;
      RECT  172500.0 701850.0 199500.0 702750.0 ;
      RECT  107100.0 720750.0 108000.0 721650.0 ;
      RECT  107100.0 723150.0 108000.0 724050.0 ;
      RECT  105750.0 720750.0 107550.0 721650.0 ;
      RECT  107100.0 721200.0 108000.0 723600.0 ;
      RECT  107550.0 723150.0 109500.0 724050.0 ;
      RECT  172050.0 720750.0 172950.0 721650.0 ;
      RECT  172050.0 725250.0 172950.0 726150.0 ;
      RECT  145650.0 720750.0 172500.0 721650.0 ;
      RECT  172050.0 721200.0 172950.0 725700.0 ;
      RECT  172500.0 725250.0 199500.0 726150.0 ;
      RECT  107100.0 733950.0 108000.0 734850.0 ;
      RECT  107100.0 731550.0 108000.0 732450.0 ;
      RECT  105750.0 733950.0 107550.0 734850.0 ;
      RECT  107100.0 732000.0 108000.0 734400.0 ;
      RECT  107550.0 731550.0 109500.0 732450.0 ;
      RECT  172050.0 733950.0 172950.0 734850.0 ;
      RECT  172050.0 729450.0 172950.0 730350.0 ;
      RECT  145650.0 733950.0 172500.0 734850.0 ;
      RECT  172050.0 729900.0 172950.0 734400.0 ;
      RECT  172500.0 729450.0 199500.0 730350.0 ;
      RECT  107100.0 748350.0 108000.0 749250.0 ;
      RECT  107100.0 750750.0 108000.0 751650.0 ;
      RECT  105750.0 748350.0 107550.0 749250.0 ;
      RECT  107100.0 748800.0 108000.0 751200.0 ;
      RECT  107550.0 750750.0 109500.0 751650.0 ;
      RECT  172050.0 748350.0 172950.0 749250.0 ;
      RECT  172050.0 752850.0 172950.0 753750.0 ;
      RECT  145650.0 748350.0 172500.0 749250.0 ;
      RECT  172050.0 748800.0 172950.0 753300.0 ;
      RECT  172500.0 752850.0 199500.0 753750.0 ;
      RECT  107100.0 761550.0 108000.0 762450.0 ;
      RECT  107100.0 759150.0 108000.0 760050.0 ;
      RECT  105750.0 761550.0 107550.0 762450.0 ;
      RECT  107100.0 759600.0 108000.0 762000.0 ;
      RECT  107550.0 759150.0 109500.0 760050.0 ;
      RECT  172050.0 761550.0 172950.0 762450.0 ;
      RECT  172050.0 757050.0 172950.0 757950.0 ;
      RECT  145650.0 761550.0 172500.0 762450.0 ;
      RECT  172050.0 757500.0 172950.0 762000.0 ;
      RECT  172500.0 757050.0 199500.0 757950.0 ;
      RECT  107100.0 775950.0 108000.0 776850.0 ;
      RECT  107100.0 778350.0 108000.0 779250.0 ;
      RECT  105750.0 775950.0 107550.0 776850.0 ;
      RECT  107100.0 776400.0 108000.0 778800.0 ;
      RECT  107550.0 778350.0 109500.0 779250.0 ;
      RECT  172050.0 775950.0 172950.0 776850.0 ;
      RECT  172050.0 780450.0 172950.0 781350.0 ;
      RECT  145650.0 775950.0 172500.0 776850.0 ;
      RECT  172050.0 776400.0 172950.0 780900.0 ;
      RECT  172500.0 780450.0 199500.0 781350.0 ;
      RECT  107100.0 789150.0 108000.0 790050.0 ;
      RECT  107100.0 786750.0 108000.0 787650.0 ;
      RECT  105750.0 789150.0 107550.0 790050.0 ;
      RECT  107100.0 787200.0 108000.0 789600.0 ;
      RECT  107550.0 786750.0 109500.0 787650.0 ;
      RECT  172050.0 789150.0 172950.0 790050.0 ;
      RECT  172050.0 784650.0 172950.0 785550.0 ;
      RECT  145650.0 789150.0 172500.0 790050.0 ;
      RECT  172050.0 785100.0 172950.0 789600.0 ;
      RECT  172500.0 784650.0 199500.0 785550.0 ;
      RECT  107100.0 803550.0 108000.0 804450.0 ;
      RECT  107100.0 805950.0 108000.0 806850.0 ;
      RECT  105750.0 803550.0 107550.0 804450.0 ;
      RECT  107100.0 804000.0 108000.0 806400.0 ;
      RECT  107550.0 805950.0 109500.0 806850.0 ;
      RECT  172050.0 803550.0 172950.0 804450.0 ;
      RECT  172050.0 808050.0 172950.0 808950.0 ;
      RECT  145650.0 803550.0 172500.0 804450.0 ;
      RECT  172050.0 804000.0 172950.0 808500.0 ;
      RECT  172500.0 808050.0 199500.0 808950.0 ;
      RECT  107100.0 816750.0 108000.0 817650.0 ;
      RECT  107100.0 814350.0 108000.0 815250.0 ;
      RECT  105750.0 816750.0 107550.0 817650.0 ;
      RECT  107100.0 814800.0 108000.0 817200.0 ;
      RECT  107550.0 814350.0 109500.0 815250.0 ;
      RECT  172050.0 816750.0 172950.0 817650.0 ;
      RECT  172050.0 812250.0 172950.0 813150.0 ;
      RECT  145650.0 816750.0 172500.0 817650.0 ;
      RECT  172050.0 812700.0 172950.0 817200.0 ;
      RECT  172500.0 812250.0 199500.0 813150.0 ;
      RECT  107100.0 831150.0 108000.0 832050.0 ;
      RECT  107100.0 833550.0 108000.0 834450.0 ;
      RECT  105750.0 831150.0 107550.0 832050.0 ;
      RECT  107100.0 831600.0 108000.0 834000.0 ;
      RECT  107550.0 833550.0 109500.0 834450.0 ;
      RECT  172050.0 831150.0 172950.0 832050.0 ;
      RECT  172050.0 835650.0 172950.0 836550.0 ;
      RECT  145650.0 831150.0 172500.0 832050.0 ;
      RECT  172050.0 831600.0 172950.0 836100.0 ;
      RECT  172500.0 835650.0 199500.0 836550.0 ;
      RECT  107100.0 844350.0 108000.0 845250.0 ;
      RECT  107100.0 841950.0 108000.0 842850.0 ;
      RECT  105750.0 844350.0 107550.0 845250.0 ;
      RECT  107100.0 842400.0 108000.0 844800.0 ;
      RECT  107550.0 841950.0 109500.0 842850.0 ;
      RECT  172050.0 844350.0 172950.0 845250.0 ;
      RECT  172050.0 839850.0 172950.0 840750.0 ;
      RECT  145650.0 844350.0 172500.0 845250.0 ;
      RECT  172050.0 840300.0 172950.0 844800.0 ;
      RECT  172500.0 839850.0 199500.0 840750.0 ;
      RECT  107100.0 858750.0 108000.0 859650.0 ;
      RECT  107100.0 861150.0 108000.0 862050.0 ;
      RECT  105750.0 858750.0 107550.0 859650.0 ;
      RECT  107100.0 859200.0 108000.0 861600.0 ;
      RECT  107550.0 861150.0 109500.0 862050.0 ;
      RECT  172050.0 858750.0 172950.0 859650.0 ;
      RECT  172050.0 863250.0 172950.0 864150.0 ;
      RECT  145650.0 858750.0 172500.0 859650.0 ;
      RECT  172050.0 859200.0 172950.0 863700.0 ;
      RECT  172500.0 863250.0 199500.0 864150.0 ;
      RECT  107100.0 871950.0 108000.0 872850.0 ;
      RECT  107100.0 869550.0 108000.0 870450.0 ;
      RECT  105750.0 871950.0 107550.0 872850.0 ;
      RECT  107100.0 870000.0 108000.0 872400.0 ;
      RECT  107550.0 869550.0 109500.0 870450.0 ;
      RECT  172050.0 871950.0 172950.0 872850.0 ;
      RECT  172050.0 867450.0 172950.0 868350.0 ;
      RECT  145650.0 871950.0 172500.0 872850.0 ;
      RECT  172050.0 867900.0 172950.0 872400.0 ;
      RECT  172500.0 867450.0 199500.0 868350.0 ;
      RECT  107100.0 886350.0 108000.0 887250.0 ;
      RECT  107100.0 888750.0 108000.0 889650.0 ;
      RECT  105750.0 886350.0 107550.0 887250.0 ;
      RECT  107100.0 886800.0 108000.0 889200.0 ;
      RECT  107550.0 888750.0 109500.0 889650.0 ;
      RECT  172050.0 886350.0 172950.0 887250.0 ;
      RECT  172050.0 890850.0 172950.0 891750.0 ;
      RECT  145650.0 886350.0 172500.0 887250.0 ;
      RECT  172050.0 886800.0 172950.0 891300.0 ;
      RECT  172500.0 890850.0 199500.0 891750.0 ;
      RECT  107100.0 899550.0 108000.0 900450.0 ;
      RECT  107100.0 897150.0 108000.0 898050.0 ;
      RECT  105750.0 899550.0 107550.0 900450.0 ;
      RECT  107100.0 897600.0 108000.0 900000.0 ;
      RECT  107550.0 897150.0 109500.0 898050.0 ;
      RECT  172050.0 899550.0 172950.0 900450.0 ;
      RECT  172050.0 895050.0 172950.0 895950.0 ;
      RECT  145650.0 899550.0 172500.0 900450.0 ;
      RECT  172050.0 895500.0 172950.0 900000.0 ;
      RECT  172500.0 895050.0 199500.0 895950.0 ;
      RECT  107100.0 913950.0 108000.0 914850.0 ;
      RECT  107100.0 916350.0 108000.0 917250.0 ;
      RECT  105750.0 913950.0 107550.0 914850.0 ;
      RECT  107100.0 914400.0 108000.0 916800.0 ;
      RECT  107550.0 916350.0 109500.0 917250.0 ;
      RECT  172050.0 913950.0 172950.0 914850.0 ;
      RECT  172050.0 918450.0 172950.0 919350.0 ;
      RECT  145650.0 913950.0 172500.0 914850.0 ;
      RECT  172050.0 914400.0 172950.0 918900.0 ;
      RECT  172500.0 918450.0 199500.0 919350.0 ;
      RECT  107100.0 927150.0 108000.0 928050.0 ;
      RECT  107100.0 924750.0 108000.0 925650.0 ;
      RECT  105750.0 927150.0 107550.0 928050.0 ;
      RECT  107100.0 925200.0 108000.0 927600.0 ;
      RECT  107550.0 924750.0 109500.0 925650.0 ;
      RECT  172050.0 927150.0 172950.0 928050.0 ;
      RECT  172050.0 922650.0 172950.0 923550.0 ;
      RECT  145650.0 927150.0 172500.0 928050.0 ;
      RECT  172050.0 923100.0 172950.0 927600.0 ;
      RECT  172500.0 922650.0 199500.0 923550.0 ;
      RECT  107100.0 941550.0 108000.0 942450.0 ;
      RECT  107100.0 943950.0 108000.0 944850.0 ;
      RECT  105750.0 941550.0 107550.0 942450.0 ;
      RECT  107100.0 942000.0 108000.0 944400.0 ;
      RECT  107550.0 943950.0 109500.0 944850.0 ;
      RECT  172050.0 941550.0 172950.0 942450.0 ;
      RECT  172050.0 946050.0 172950.0 946950.0 ;
      RECT  145650.0 941550.0 172500.0 942450.0 ;
      RECT  172050.0 942000.0 172950.0 946500.0 ;
      RECT  172500.0 946050.0 199500.0 946950.0 ;
      RECT  107100.0 954750.0 108000.0 955650.0 ;
      RECT  107100.0 952350.0 108000.0 953250.0 ;
      RECT  105750.0 954750.0 107550.0 955650.0 ;
      RECT  107100.0 952800.0 108000.0 955200.0 ;
      RECT  107550.0 952350.0 109500.0 953250.0 ;
      RECT  172050.0 954750.0 172950.0 955650.0 ;
      RECT  172050.0 950250.0 172950.0 951150.0 ;
      RECT  145650.0 954750.0 172500.0 955650.0 ;
      RECT  172050.0 950700.0 172950.0 955200.0 ;
      RECT  172500.0 950250.0 199500.0 951150.0 ;
      RECT  107100.0 969150.0 108000.0 970050.0 ;
      RECT  107100.0 971550.0 108000.0 972450.0 ;
      RECT  105750.0 969150.0 107550.0 970050.0 ;
      RECT  107100.0 969600.0 108000.0 972000.0 ;
      RECT  107550.0 971550.0 109500.0 972450.0 ;
      RECT  172050.0 969150.0 172950.0 970050.0 ;
      RECT  172050.0 973650.0 172950.0 974550.0 ;
      RECT  145650.0 969150.0 172500.0 970050.0 ;
      RECT  172050.0 969600.0 172950.0 974100.0 ;
      RECT  172500.0 973650.0 199500.0 974550.0 ;
      RECT  107100.0 982350.0 108000.0 983250.0 ;
      RECT  107100.0 979950.0 108000.0 980850.0 ;
      RECT  105750.0 982350.0 107550.0 983250.0 ;
      RECT  107100.0 980400.0 108000.0 982800.0 ;
      RECT  107550.0 979950.0 109500.0 980850.0 ;
      RECT  172050.0 982350.0 172950.0 983250.0 ;
      RECT  172050.0 977850.0 172950.0 978750.0 ;
      RECT  145650.0 982350.0 172500.0 983250.0 ;
      RECT  172050.0 978300.0 172950.0 982800.0 ;
      RECT  172500.0 977850.0 199500.0 978750.0 ;
      RECT  107100.0 996750.0 108000.0 997650.0 ;
      RECT  107100.0 999150.0 108000.0 1000050.0 ;
      RECT  105750.0 996750.0 107550.0 997650.0 ;
      RECT  107100.0 997200.0 108000.0 999600.0 ;
      RECT  107550.0 999150.0 109500.0 1000050.0 ;
      RECT  172050.0 996750.0 172950.0 997650.0 ;
      RECT  172050.0 1001250.0 172950.0 1002150.0 ;
      RECT  145650.0 996750.0 172500.0 997650.0 ;
      RECT  172050.0 997200.0 172950.0 1001700.0 ;
      RECT  172500.0 1001250.0 199500.0 1002150.0 ;
      RECT  107100.0 1009950.0 108000.0 1010850.0 ;
      RECT  107100.0 1007550.0 108000.0 1008450.0 ;
      RECT  105750.0 1009950.0 107550.0 1010850.0 ;
      RECT  107100.0 1008000.0 108000.0 1010400.0 ;
      RECT  107550.0 1007550.0 109500.0 1008450.0 ;
      RECT  172050.0 1009950.0 172950.0 1010850.0 ;
      RECT  172050.0 1005450.0 172950.0 1006350.0 ;
      RECT  145650.0 1009950.0 172500.0 1010850.0 ;
      RECT  172050.0 1005900.0 172950.0 1010400.0 ;
      RECT  172500.0 1005450.0 199500.0 1006350.0 ;
      RECT  107100.0 1024350.0 108000.0 1025250.0 ;
      RECT  107100.0 1026750.0 108000.0 1027650.0 ;
      RECT  105750.0 1024350.0 107550.0 1025250.0 ;
      RECT  107100.0 1024800.0 108000.0 1027200.0 ;
      RECT  107550.0 1026750.0 109500.0 1027650.0 ;
      RECT  172050.0 1024350.0 172950.0 1025250.0 ;
      RECT  172050.0 1028850.0 172950.0 1029750.0 ;
      RECT  145650.0 1024350.0 172500.0 1025250.0 ;
      RECT  172050.0 1024800.0 172950.0 1029300.0 ;
      RECT  172500.0 1028850.0 199500.0 1029750.0 ;
      RECT  107100.0 1037550.0 108000.0 1038450.0 ;
      RECT  107100.0 1035150.0 108000.0 1036050.0 ;
      RECT  105750.0 1037550.0 107550.0 1038450.0 ;
      RECT  107100.0 1035600.0 108000.0 1038000.0 ;
      RECT  107550.0 1035150.0 109500.0 1036050.0 ;
      RECT  172050.0 1037550.0 172950.0 1038450.0 ;
      RECT  172050.0 1033050.0 172950.0 1033950.0 ;
      RECT  145650.0 1037550.0 172500.0 1038450.0 ;
      RECT  172050.0 1033500.0 172950.0 1038000.0 ;
      RECT  172500.0 1033050.0 199500.0 1033950.0 ;
      RECT  107100.0 1051950.0 108000.0 1052850.0 ;
      RECT  107100.0 1054350.0 108000.0 1055250.0 ;
      RECT  105750.0 1051950.0 107550.0 1052850.0 ;
      RECT  107100.0 1052400.0 108000.0 1054800.0 ;
      RECT  107550.0 1054350.0 109500.0 1055250.0 ;
      RECT  172050.0 1051950.0 172950.0 1052850.0 ;
      RECT  172050.0 1056450.0 172950.0 1057350.0 ;
      RECT  145650.0 1051950.0 172500.0 1052850.0 ;
      RECT  172050.0 1052400.0 172950.0 1056900.0 ;
      RECT  172500.0 1056450.0 199500.0 1057350.0 ;
      RECT  107100.0 1065150.0 108000.0 1066050.0 ;
      RECT  107100.0 1062750.0 108000.0 1063650.0 ;
      RECT  105750.0 1065150.0 107550.0 1066050.0 ;
      RECT  107100.0 1063200.0 108000.0 1065600.0 ;
      RECT  107550.0 1062750.0 109500.0 1063650.0 ;
      RECT  172050.0 1065150.0 172950.0 1066050.0 ;
      RECT  172050.0 1060650.0 172950.0 1061550.0 ;
      RECT  145650.0 1065150.0 172500.0 1066050.0 ;
      RECT  172050.0 1061100.0 172950.0 1065600.0 ;
      RECT  172500.0 1060650.0 199500.0 1061550.0 ;
      RECT  107100.0 1079550.0 108000.0 1080450.0 ;
      RECT  107100.0 1081950.0 108000.0 1082850.0 ;
      RECT  105750.0 1079550.0 107550.0 1080450.0 ;
      RECT  107100.0 1080000.0 108000.0 1082400.0 ;
      RECT  107550.0 1081950.0 109500.0 1082850.0 ;
      RECT  172050.0 1079550.0 172950.0 1080450.0 ;
      RECT  172050.0 1084050.0 172950.0 1084950.0 ;
      RECT  145650.0 1079550.0 172500.0 1080450.0 ;
      RECT  172050.0 1080000.0 172950.0 1084500.0 ;
      RECT  172500.0 1084050.0 199500.0 1084950.0 ;
      RECT  107100.0 1092750.0 108000.0 1093650.0 ;
      RECT  107100.0 1090350.0 108000.0 1091250.0 ;
      RECT  105750.0 1092750.0 107550.0 1093650.0 ;
      RECT  107100.0 1090800.0 108000.0 1093200.0 ;
      RECT  107550.0 1090350.0 109500.0 1091250.0 ;
      RECT  172050.0 1092750.0 172950.0 1093650.0 ;
      RECT  172050.0 1088250.0 172950.0 1089150.0 ;
      RECT  145650.0 1092750.0 172500.0 1093650.0 ;
      RECT  172050.0 1088700.0 172950.0 1093200.0 ;
      RECT  172500.0 1088250.0 199500.0 1089150.0 ;
      RECT  107100.0 1107150.0 108000.0 1108050.0 ;
      RECT  107100.0 1109550.0 108000.0 1110450.0 ;
      RECT  105750.0 1107150.0 107550.0 1108050.0 ;
      RECT  107100.0 1107600.0 108000.0 1110000.0 ;
      RECT  107550.0 1109550.0 109500.0 1110450.0 ;
      RECT  172050.0 1107150.0 172950.0 1108050.0 ;
      RECT  172050.0 1111650.0 172950.0 1112550.0 ;
      RECT  145650.0 1107150.0 172500.0 1108050.0 ;
      RECT  172050.0 1107600.0 172950.0 1112100.0 ;
      RECT  172500.0 1111650.0 199500.0 1112550.0 ;
      RECT  107100.0 1120350.0 108000.0 1121250.0 ;
      RECT  107100.0 1117950.0 108000.0 1118850.0 ;
      RECT  105750.0 1120350.0 107550.0 1121250.0 ;
      RECT  107100.0 1118400.0 108000.0 1120800.0 ;
      RECT  107550.0 1117950.0 109500.0 1118850.0 ;
      RECT  172050.0 1120350.0 172950.0 1121250.0 ;
      RECT  172050.0 1115850.0 172950.0 1116750.0 ;
      RECT  145650.0 1120350.0 172500.0 1121250.0 ;
      RECT  172050.0 1116300.0 172950.0 1120800.0 ;
      RECT  172500.0 1115850.0 199500.0 1116750.0 ;
      RECT  107100.0 1134750.0 108000.0 1135650.0 ;
      RECT  107100.0 1137150.0 108000.0 1138050.0 ;
      RECT  105750.0 1134750.0 107550.0 1135650.0 ;
      RECT  107100.0 1135200.0 108000.0 1137600.0 ;
      RECT  107550.0 1137150.0 109500.0 1138050.0 ;
      RECT  172050.0 1134750.0 172950.0 1135650.0 ;
      RECT  172050.0 1139250.0 172950.0 1140150.0 ;
      RECT  145650.0 1134750.0 172500.0 1135650.0 ;
      RECT  172050.0 1135200.0 172950.0 1139700.0 ;
      RECT  172500.0 1139250.0 199500.0 1140150.0 ;
      RECT  107100.0 1147950.0 108000.0 1148850.0 ;
      RECT  107100.0 1145550.0 108000.0 1146450.0 ;
      RECT  105750.0 1147950.0 107550.0 1148850.0 ;
      RECT  107100.0 1146000.0 108000.0 1148400.0 ;
      RECT  107550.0 1145550.0 109500.0 1146450.0 ;
      RECT  172050.0 1147950.0 172950.0 1148850.0 ;
      RECT  172050.0 1143450.0 172950.0 1144350.0 ;
      RECT  145650.0 1147950.0 172500.0 1148850.0 ;
      RECT  172050.0 1143900.0 172950.0 1148400.0 ;
      RECT  172500.0 1143450.0 199500.0 1144350.0 ;
      RECT  107100.0 1162350.0 108000.0 1163250.0 ;
      RECT  107100.0 1164750.0 108000.0 1165650.0 ;
      RECT  105750.0 1162350.0 107550.0 1163250.0 ;
      RECT  107100.0 1162800.0 108000.0 1165200.0 ;
      RECT  107550.0 1164750.0 109500.0 1165650.0 ;
      RECT  172050.0 1162350.0 172950.0 1163250.0 ;
      RECT  172050.0 1166850.0 172950.0 1167750.0 ;
      RECT  145650.0 1162350.0 172500.0 1163250.0 ;
      RECT  172050.0 1162800.0 172950.0 1167300.0 ;
      RECT  172500.0 1166850.0 199500.0 1167750.0 ;
      RECT  107100.0 1175550.0 108000.0 1176450.0 ;
      RECT  107100.0 1173150.0 108000.0 1174050.0 ;
      RECT  105750.0 1175550.0 107550.0 1176450.0 ;
      RECT  107100.0 1173600.0 108000.0 1176000.0 ;
      RECT  107550.0 1173150.0 109500.0 1174050.0 ;
      RECT  172050.0 1175550.0 172950.0 1176450.0 ;
      RECT  172050.0 1171050.0 172950.0 1171950.0 ;
      RECT  145650.0 1175550.0 172500.0 1176450.0 ;
      RECT  172050.0 1171500.0 172950.0 1176000.0 ;
      RECT  172500.0 1171050.0 199500.0 1171950.0 ;
      RECT  107100.0 1189950.0 108000.0 1190850.0 ;
      RECT  107100.0 1192350.0 108000.0 1193250.0 ;
      RECT  105750.0 1189950.0 107550.0 1190850.0 ;
      RECT  107100.0 1190400.0 108000.0 1192800.0 ;
      RECT  107550.0 1192350.0 109500.0 1193250.0 ;
      RECT  172050.0 1189950.0 172950.0 1190850.0 ;
      RECT  172050.0 1194450.0 172950.0 1195350.0 ;
      RECT  145650.0 1189950.0 172500.0 1190850.0 ;
      RECT  172050.0 1190400.0 172950.0 1194900.0 ;
      RECT  172500.0 1194450.0 199500.0 1195350.0 ;
      RECT  115800.0 313350.0 200100.0 314250.0 ;
      RECT  115800.0 340950.0 200100.0 341850.0 ;
      RECT  115800.0 368550.0 200100.0 369450.0 ;
      RECT  115800.0 396150.0 200100.0 397050.0 ;
      RECT  115800.0 423750.0 200100.0 424650.0 ;
      RECT  115800.0 451350.0 200100.0 452250.0 ;
      RECT  115800.0 478950.0 200100.0 479850.0 ;
      RECT  115800.0 506550.0 200100.0 507450.0 ;
      RECT  115800.0 534150.0 200100.0 535050.0 ;
      RECT  115800.0 561750.0 200100.0 562650.0 ;
      RECT  115800.0 589350.0 200100.0 590250.0 ;
      RECT  115800.0 616950.0 200100.0 617850.0 ;
      RECT  115800.0 644550.0 200100.0 645450.0 ;
      RECT  115800.0 672150.0 200100.0 673050.0 ;
      RECT  115800.0 699750.0 200100.0 700650.0 ;
      RECT  115800.0 727350.0 200100.0 728250.0 ;
      RECT  115800.0 754950.0 200100.0 755850.0 ;
      RECT  115800.0 782550.0 200100.0 783450.0 ;
      RECT  115800.0 810150.0 200100.0 811050.0 ;
      RECT  115800.0 837750.0 200100.0 838650.0 ;
      RECT  115800.0 865350.0 200100.0 866250.0 ;
      RECT  115800.0 892950.0 200100.0 893850.0 ;
      RECT  115800.0 920550.0 200100.0 921450.0 ;
      RECT  115800.0 948150.0 200100.0 949050.0 ;
      RECT  115800.0 975750.0 200100.0 976650.0 ;
      RECT  115800.0 1003350.0 200100.0 1004250.0 ;
      RECT  115800.0 1030950.0 200100.0 1031850.0 ;
      RECT  115800.0 1058550.0 200100.0 1059450.0 ;
      RECT  115800.0 1086150.0 200100.0 1087050.0 ;
      RECT  115800.0 1113750.0 200100.0 1114650.0 ;
      RECT  115800.0 1141350.0 200100.0 1142250.0 ;
      RECT  115800.0 1168950.0 200100.0 1169850.0 ;
      RECT  115800.0 1196550.0 200100.0 1197450.0 ;
      RECT  52800.0 327150.0 533700.0 328050.0 ;
      RECT  52800.0 354750.0 533700.0 355650.0 ;
      RECT  52800.0 382350.0 533700.0 383250.0 ;
      RECT  52800.0 409950.0 533700.0 410850.0 ;
      RECT  52800.0 437550.0 533700.0 438450.0 ;
      RECT  52800.0 465150.0 533700.0 466050.0 ;
      RECT  52800.0 492750.0 533700.0 493650.0 ;
      RECT  52800.0 520350.0 533700.0 521250.0 ;
      RECT  52800.0 547950.0 533700.0 548850.0 ;
      RECT  52800.0 575550.0 533700.0 576450.0 ;
      RECT  52800.0 603150.0 533700.0 604050.0 ;
      RECT  52800.0 630750.0 533700.0 631650.0 ;
      RECT  52800.0 658350.0 533700.0 659250.0 ;
      RECT  52800.0 685950.0 533700.0 686850.0 ;
      RECT  52800.0 713550.0 533700.0 714450.0 ;
      RECT  52800.0 741150.0 533700.0 742050.0 ;
      RECT  52800.0 768750.0 533700.0 769650.0 ;
      RECT  52800.0 796350.0 533700.0 797250.0 ;
      RECT  52800.0 823950.0 533700.0 824850.0 ;
      RECT  52800.0 851550.0 533700.0 852450.0 ;
      RECT  52800.0 879150.0 533700.0 880050.0 ;
      RECT  52800.0 906750.0 533700.0 907650.0 ;
      RECT  52800.0 934350.0 533700.0 935250.0 ;
      RECT  52800.0 961950.0 533700.0 962850.0 ;
      RECT  52800.0 989550.0 533700.0 990450.0 ;
      RECT  52800.0 1017150.0 533700.0 1018050.0 ;
      RECT  52800.0 1044750.0 533700.0 1045650.0 ;
      RECT  52800.0 1072350.0 533700.0 1073250.0 ;
      RECT  52800.0 1099950.0 533700.0 1100850.0 ;
      RECT  52800.0 1127550.0 533700.0 1128450.0 ;
      RECT  52800.0 1155150.0 533700.0 1156050.0 ;
      RECT  52800.0 1182750.0 533700.0 1183650.0 ;
      RECT  138900.0 150450.0 143400.0 151350.0 ;
      RECT  135900.0 164250.0 146100.0 165150.0 ;
      RECT  138900.0 205650.0 148800.0 206550.0 ;
      RECT  135900.0 219450.0 151500.0 220350.0 ;
      RECT  138900.0 260850.0 154200.0 261750.0 ;
      RECT  135900.0 274650.0 156900.0 275550.0 ;
      RECT  138900.0 147750.0 140400.0 148650.0 ;
      RECT  138900.0 175350.0 140400.0 176250.0 ;
      RECT  138900.0 202950.0 140400.0 203850.0 ;
      RECT  138900.0 230550.0 140400.0 231450.0 ;
      RECT  138900.0 258150.0 140400.0 259050.0 ;
      RECT  138900.0 285750.0 140400.0 286650.0 ;
      RECT  52800.0 161550.0 138900.0 162450.0 ;
      RECT  52800.0 189150.0 138900.0 190050.0 ;
      RECT  52800.0 216750.0 138900.0 217650.0 ;
      RECT  52800.0 244350.0 138900.0 245250.0 ;
      RECT  52800.0 271950.0 138900.0 272850.0 ;
      RECT  52800.0 299550.0 138900.0 300450.0 ;
      RECT  159600.0 285900.0 200100.0 286800.0 ;
      RECT  162300.0 283800.0 200100.0 284700.0 ;
      RECT  165000.0 281700.0 200100.0 282600.0 ;
      RECT  167700.0 279600.0 200100.0 280500.0 ;
      RECT  133500.0 6750.0 159600.0 7650.0 ;
      RECT  133500.0 21150.0 162300.0 22050.0 ;
      RECT  133500.0 34350.0 165000.0 35250.0 ;
      RECT  133500.0 48750.0 167700.0 49650.0 ;
      RECT  133500.0 150.0 172650.0 1050.0 ;
      RECT  133500.0 27750.0 172650.0 28650.0 ;
      RECT  133500.0 55350.0 172650.0 56250.0 ;
      RECT  52800.0 13950.0 172650.0 14850.0 ;
      RECT  52800.0 41550.0 172650.0 42450.0 ;
      RECT  117900.0 136500.0 143400.0 137400.0 ;
      RECT  117900.0 127800.0 146100.0 128700.0 ;
      RECT  117900.0 116100.0 148800.0 117000.0 ;
      RECT  117900.0 107400.0 151500.0 108300.0 ;
      RECT  117900.0 95700.0 154200.0 96600.0 ;
      RECT  117900.0 87000.0 156900.0 87900.0 ;
      RECT  119100.0 132150.0 173850.0 133050.0 ;
      RECT  119100.0 111750.0 173850.0 112650.0 ;
      RECT  119100.0 91350.0 173850.0 92250.0 ;
      RECT  119100.0 70950.0 173850.0 71850.0 ;
      RECT  115500.0 58650.0 116400.0 59550.0 ;
      RECT  115500.0 59100.0 116400.0 61200.0 ;
      RECT  52800.0 58650.0 115950.0 59550.0 ;
      RECT  188400.0 106050.0 200100.0 106950.0 ;
      RECT  183000.0 101550.0 200100.0 102450.0 ;
      RECT  185700.0 99150.0 200100.0 100050.0 ;
      RECT  188400.0 1205400.0 200100.0 1206300.0 ;
      RECT  191100.0 170850.0 200100.0 171750.0 ;
      RECT  193800.0 268950.0 200100.0 269850.0 ;
      RECT  61500.0 144450.0 62400.0 145350.0 ;
      RECT  61500.0 142800.0 62400.0 144900.0 ;
      RECT  61950.0 144450.0 180300.0 145350.0 ;
      RECT  112650.0 1198650.0 181200.0 1199550.0 ;
      RECT  200100.0 1216500.0 529200.0 1217400.0 ;
      RECT  200100.0 241650.0 529200.0 242550.0 ;
      RECT  200100.0 172950.0 529200.0 173850.0 ;
      RECT  200100.0 160050.0 529200.0 160950.0 ;
      RECT  200100.0 83250.0 529200.0 84150.0 ;
      RECT  177150.0 97050.0 200100.0 97950.0 ;
      RECT  177150.0 266850.0 200100.0 267750.0 ;
      RECT  177150.0 168750.0 200100.0 169650.0 ;
      RECT  200100.0 313800.0 210300.0 327600.0 ;
      RECT  200100.0 341400.0 210300.0 327600.0 ;
      RECT  200100.0 341400.0 210300.0 355200.0 ;
      RECT  200100.0 369000.0 210300.0 355200.0 ;
      RECT  200100.0 369000.0 210300.0 382800.0 ;
      RECT  200100.0 396600.0 210300.0 382800.0 ;
      RECT  200100.0 396600.0 210300.0 410400.0 ;
      RECT  200100.0 424200.0 210300.0 410400.0 ;
      RECT  200100.0 424200.0 210300.0 438000.0 ;
      RECT  200100.0 451800.0 210300.0 438000.0 ;
      RECT  200100.0 451800.0 210300.0 465600.0 ;
      RECT  200100.0 479400.0 210300.0 465600.0 ;
      RECT  200100.0 479400.0 210300.0 493200.0 ;
      RECT  200100.0 507000.0 210300.0 493200.0 ;
      RECT  200100.0 507000.0 210300.0 520800.0 ;
      RECT  200100.0 534600.0 210300.0 520800.0 ;
      RECT  200100.0 534600.0 210300.0 548400.0 ;
      RECT  200100.0 562200.0 210300.0 548400.0 ;
      RECT  200100.0 562200.0 210300.0 576000.0 ;
      RECT  200100.0 589800.0 210300.0 576000.0 ;
      RECT  200100.0 589800.0 210300.0 603600.0 ;
      RECT  200100.0 617400.0 210300.0 603600.0 ;
      RECT  200100.0 617400.0 210300.0 631200.0 ;
      RECT  200100.0 645000.0 210300.0 631200.0 ;
      RECT  200100.0 645000.0 210300.0 658800.0 ;
      RECT  200100.0 672600.0 210300.0 658800.0 ;
      RECT  200100.0 672600.0 210300.0 686400.0 ;
      RECT  200100.0 700200.0 210300.0 686400.0 ;
      RECT  200100.0 700200.0 210300.0 714000.0 ;
      RECT  200100.0 727800.0 210300.0 714000.0 ;
      RECT  200100.0 727800.0 210300.0 741600.0 ;
      RECT  200100.0 755400.0 210300.0 741600.0 ;
      RECT  200100.0 755400.0 210300.0 769200.0 ;
      RECT  200100.0 783000.0 210300.0 769200.0 ;
      RECT  200100.0 783000.0 210300.0 796800.0 ;
      RECT  200100.0 810600.0 210300.0 796800.0 ;
      RECT  200100.0 810600.0 210300.0 824400.0 ;
      RECT  200100.0 838200.0 210300.0 824400.0 ;
      RECT  200100.0 838200.0 210300.0 852000.0 ;
      RECT  200100.0 865800.0 210300.0 852000.0 ;
      RECT  200100.0 865800.0 210300.0 879600.0 ;
      RECT  200100.0 893400.0 210300.0 879600.0 ;
      RECT  200100.0 893400.0 210300.0 907200.0 ;
      RECT  200100.0 921000.0 210300.0 907200.0 ;
      RECT  200100.0 921000.0 210300.0 934800.0 ;
      RECT  200100.0 948600.0 210300.0 934800.0 ;
      RECT  200100.0 948600.0 210300.0 962400.0 ;
      RECT  200100.0 976200.0 210300.0 962400.0 ;
      RECT  200100.0 976200.0 210300.0 990000.0 ;
      RECT  200100.0 1003800.0 210300.0 990000.0 ;
      RECT  200100.0 1003800.0 210300.0 1017600.0 ;
      RECT  200100.0 1031400.0 210300.0 1017600.0 ;
      RECT  200100.0 1031400.0 210300.0 1045200.0 ;
      RECT  200100.0 1059000.0 210300.0 1045200.0 ;
      RECT  200100.0 1059000.0 210300.0 1072800.0 ;
      RECT  200100.0 1086600.0 210300.0 1072800.0 ;
      RECT  200100.0 1086600.0 210300.0 1100400.0 ;
      RECT  200100.0 1114200.0 210300.0 1100400.0 ;
      RECT  200100.0 1114200.0 210300.0 1128000.0 ;
      RECT  200100.0 1141800.0 210300.0 1128000.0 ;
      RECT  200100.0 1141800.0 210300.0 1155600.0 ;
      RECT  200100.0 1169400.0 210300.0 1155600.0 ;
      RECT  200100.0 1169400.0 210300.0 1183200.0 ;
      RECT  200100.0 1197000.0 210300.0 1183200.0 ;
      RECT  210300.0 313800.0 220500.0 327600.0 ;
      RECT  210300.0 341400.0 220500.0 327600.0 ;
      RECT  210300.0 341400.0 220500.0 355200.0 ;
      RECT  210300.0 369000.0 220500.0 355200.0 ;
      RECT  210300.0 369000.0 220500.0 382800.0 ;
      RECT  210300.0 396600.0 220500.0 382800.0 ;
      RECT  210300.0 396600.0 220500.0 410400.0 ;
      RECT  210300.0 424200.0 220500.0 410400.0 ;
      RECT  210300.0 424200.0 220500.0 438000.0 ;
      RECT  210300.0 451800.0 220500.0 438000.0 ;
      RECT  210300.0 451800.0 220500.0 465600.0 ;
      RECT  210300.0 479400.0 220500.0 465600.0 ;
      RECT  210300.0 479400.0 220500.0 493200.0 ;
      RECT  210300.0 507000.0 220500.0 493200.0 ;
      RECT  210300.0 507000.0 220500.0 520800.0 ;
      RECT  210300.0 534600.0 220500.0 520800.0 ;
      RECT  210300.0 534600.0 220500.0 548400.0 ;
      RECT  210300.0 562200.0 220500.0 548400.0 ;
      RECT  210300.0 562200.0 220500.0 576000.0 ;
      RECT  210300.0 589800.0 220500.0 576000.0 ;
      RECT  210300.0 589800.0 220500.0 603600.0 ;
      RECT  210300.0 617400.0 220500.0 603600.0 ;
      RECT  210300.0 617400.0 220500.0 631200.0 ;
      RECT  210300.0 645000.0 220500.0 631200.0 ;
      RECT  210300.0 645000.0 220500.0 658800.0 ;
      RECT  210300.0 672600.0 220500.0 658800.0 ;
      RECT  210300.0 672600.0 220500.0 686400.0 ;
      RECT  210300.0 700200.0 220500.0 686400.0 ;
      RECT  210300.0 700200.0 220500.0 714000.0 ;
      RECT  210300.0 727800.0 220500.0 714000.0 ;
      RECT  210300.0 727800.0 220500.0 741600.0 ;
      RECT  210300.0 755400.0 220500.0 741600.0 ;
      RECT  210300.0 755400.0 220500.0 769200.0 ;
      RECT  210300.0 783000.0 220500.0 769200.0 ;
      RECT  210300.0 783000.0 220500.0 796800.0 ;
      RECT  210300.0 810600.0 220500.0 796800.0 ;
      RECT  210300.0 810600.0 220500.0 824400.0 ;
      RECT  210300.0 838200.0 220500.0 824400.0 ;
      RECT  210300.0 838200.0 220500.0 852000.0 ;
      RECT  210300.0 865800.0 220500.0 852000.0 ;
      RECT  210300.0 865800.0 220500.0 879600.0 ;
      RECT  210300.0 893400.0 220500.0 879600.0 ;
      RECT  210300.0 893400.0 220500.0 907200.0 ;
      RECT  210300.0 921000.0 220500.0 907200.0 ;
      RECT  210300.0 921000.0 220500.0 934800.0 ;
      RECT  210300.0 948600.0 220500.0 934800.0 ;
      RECT  210300.0 948600.0 220500.0 962400.0 ;
      RECT  210300.0 976200.0 220500.0 962400.0 ;
      RECT  210300.0 976200.0 220500.0 990000.0 ;
      RECT  210300.0 1003800.0 220500.0 990000.0 ;
      RECT  210300.0 1003800.0 220500.0 1017600.0 ;
      RECT  210300.0 1031400.0 220500.0 1017600.0 ;
      RECT  210300.0 1031400.0 220500.0 1045200.0 ;
      RECT  210300.0 1059000.0 220500.0 1045200.0 ;
      RECT  210300.0 1059000.0 220500.0 1072800.0 ;
      RECT  210300.0 1086600.0 220500.0 1072800.0 ;
      RECT  210300.0 1086600.0 220500.0 1100400.0 ;
      RECT  210300.0 1114200.0 220500.0 1100400.0 ;
      RECT  210300.0 1114200.0 220500.0 1128000.0 ;
      RECT  210300.0 1141800.0 220500.0 1128000.0 ;
      RECT  210300.0 1141800.0 220500.0 1155600.0 ;
      RECT  210300.0 1169400.0 220500.0 1155600.0 ;
      RECT  210300.0 1169400.0 220500.0 1183200.0 ;
      RECT  210300.0 1197000.0 220500.0 1183200.0 ;
      RECT  220500.0 313800.0 230700.0 327600.0 ;
      RECT  220500.0 341400.0 230700.0 327600.0 ;
      RECT  220500.0 341400.0 230700.0 355200.0 ;
      RECT  220500.0 369000.0 230700.0 355200.0 ;
      RECT  220500.0 369000.0 230700.0 382800.0 ;
      RECT  220500.0 396600.0 230700.0 382800.0 ;
      RECT  220500.0 396600.0 230700.0 410400.0 ;
      RECT  220500.0 424200.0 230700.0 410400.0 ;
      RECT  220500.0 424200.0 230700.0 438000.0 ;
      RECT  220500.0 451800.0 230700.0 438000.0 ;
      RECT  220500.0 451800.0 230700.0 465600.0 ;
      RECT  220500.0 479400.0 230700.0 465600.0 ;
      RECT  220500.0 479400.0 230700.0 493200.0 ;
      RECT  220500.0 507000.0 230700.0 493200.0 ;
      RECT  220500.0 507000.0 230700.0 520800.0 ;
      RECT  220500.0 534600.0 230700.0 520800.0 ;
      RECT  220500.0 534600.0 230700.0 548400.0 ;
      RECT  220500.0 562200.0 230700.0 548400.0 ;
      RECT  220500.0 562200.0 230700.0 576000.0 ;
      RECT  220500.0 589800.0 230700.0 576000.0 ;
      RECT  220500.0 589800.0 230700.0 603600.0 ;
      RECT  220500.0 617400.0 230700.0 603600.0 ;
      RECT  220500.0 617400.0 230700.0 631200.0 ;
      RECT  220500.0 645000.0 230700.0 631200.0 ;
      RECT  220500.0 645000.0 230700.0 658800.0 ;
      RECT  220500.0 672600.0 230700.0 658800.0 ;
      RECT  220500.0 672600.0 230700.0 686400.0 ;
      RECT  220500.0 700200.0 230700.0 686400.0 ;
      RECT  220500.0 700200.0 230700.0 714000.0 ;
      RECT  220500.0 727800.0 230700.0 714000.0 ;
      RECT  220500.0 727800.0 230700.0 741600.0 ;
      RECT  220500.0 755400.0 230700.0 741600.0 ;
      RECT  220500.0 755400.0 230700.0 769200.0 ;
      RECT  220500.0 783000.0 230700.0 769200.0 ;
      RECT  220500.0 783000.0 230700.0 796800.0 ;
      RECT  220500.0 810600.0 230700.0 796800.0 ;
      RECT  220500.0 810600.0 230700.0 824400.0 ;
      RECT  220500.0 838200.0 230700.0 824400.0 ;
      RECT  220500.0 838200.0 230700.0 852000.0 ;
      RECT  220500.0 865800.0 230700.0 852000.0 ;
      RECT  220500.0 865800.0 230700.0 879600.0 ;
      RECT  220500.0 893400.0 230700.0 879600.0 ;
      RECT  220500.0 893400.0 230700.0 907200.0 ;
      RECT  220500.0 921000.0 230700.0 907200.0 ;
      RECT  220500.0 921000.0 230700.0 934800.0 ;
      RECT  220500.0 948600.0 230700.0 934800.0 ;
      RECT  220500.0 948600.0 230700.0 962400.0 ;
      RECT  220500.0 976200.0 230700.0 962400.0 ;
      RECT  220500.0 976200.0 230700.0 990000.0 ;
      RECT  220500.0 1003800.0 230700.0 990000.0 ;
      RECT  220500.0 1003800.0 230700.0 1017600.0 ;
      RECT  220500.0 1031400.0 230700.0 1017600.0 ;
      RECT  220500.0 1031400.0 230700.0 1045200.0 ;
      RECT  220500.0 1059000.0 230700.0 1045200.0 ;
      RECT  220500.0 1059000.0 230700.0 1072800.0 ;
      RECT  220500.0 1086600.0 230700.0 1072800.0 ;
      RECT  220500.0 1086600.0 230700.0 1100400.0 ;
      RECT  220500.0 1114200.0 230700.0 1100400.0 ;
      RECT  220500.0 1114200.0 230700.0 1128000.0 ;
      RECT  220500.0 1141800.0 230700.0 1128000.0 ;
      RECT  220500.0 1141800.0 230700.0 1155600.0 ;
      RECT  220500.0 1169400.0 230700.0 1155600.0 ;
      RECT  220500.0 1169400.0 230700.0 1183200.0 ;
      RECT  220500.0 1197000.0 230700.0 1183200.0 ;
      RECT  230700.0 313800.0 240900.0 327600.0 ;
      RECT  230700.0 341400.0 240900.0 327600.0 ;
      RECT  230700.0 341400.0 240900.0 355200.0 ;
      RECT  230700.0 369000.0 240900.0 355200.0 ;
      RECT  230700.0 369000.0 240900.0 382800.0 ;
      RECT  230700.0 396600.0 240900.0 382800.0 ;
      RECT  230700.0 396600.0 240900.0 410400.0 ;
      RECT  230700.0 424200.0 240900.0 410400.0 ;
      RECT  230700.0 424200.0 240900.0 438000.0 ;
      RECT  230700.0 451800.0 240900.0 438000.0 ;
      RECT  230700.0 451800.0 240900.0 465600.0 ;
      RECT  230700.0 479400.0 240900.0 465600.0 ;
      RECT  230700.0 479400.0 240900.0 493200.0 ;
      RECT  230700.0 507000.0 240900.0 493200.0 ;
      RECT  230700.0 507000.0 240900.0 520800.0 ;
      RECT  230700.0 534600.0 240900.0 520800.0 ;
      RECT  230700.0 534600.0 240900.0 548400.0 ;
      RECT  230700.0 562200.0 240900.0 548400.0 ;
      RECT  230700.0 562200.0 240900.0 576000.0 ;
      RECT  230700.0 589800.0 240900.0 576000.0 ;
      RECT  230700.0 589800.0 240900.0 603600.0 ;
      RECT  230700.0 617400.0 240900.0 603600.0 ;
      RECT  230700.0 617400.0 240900.0 631200.0 ;
      RECT  230700.0 645000.0 240900.0 631200.0 ;
      RECT  230700.0 645000.0 240900.0 658800.0 ;
      RECT  230700.0 672600.0 240900.0 658800.0 ;
      RECT  230700.0 672600.0 240900.0 686400.0 ;
      RECT  230700.0 700200.0 240900.0 686400.0 ;
      RECT  230700.0 700200.0 240900.0 714000.0 ;
      RECT  230700.0 727800.0 240900.0 714000.0 ;
      RECT  230700.0 727800.0 240900.0 741600.0 ;
      RECT  230700.0 755400.0 240900.0 741600.0 ;
      RECT  230700.0 755400.0 240900.0 769200.0 ;
      RECT  230700.0 783000.0 240900.0 769200.0 ;
      RECT  230700.0 783000.0 240900.0 796800.0 ;
      RECT  230700.0 810600.0 240900.0 796800.0 ;
      RECT  230700.0 810600.0 240900.0 824400.0 ;
      RECT  230700.0 838200.0 240900.0 824400.0 ;
      RECT  230700.0 838200.0 240900.0 852000.0 ;
      RECT  230700.0 865800.0 240900.0 852000.0 ;
      RECT  230700.0 865800.0 240900.0 879600.0 ;
      RECT  230700.0 893400.0 240900.0 879600.0 ;
      RECT  230700.0 893400.0 240900.0 907200.0 ;
      RECT  230700.0 921000.0 240900.0 907200.0 ;
      RECT  230700.0 921000.0 240900.0 934800.0 ;
      RECT  230700.0 948600.0 240900.0 934800.0 ;
      RECT  230700.0 948600.0 240900.0 962400.0 ;
      RECT  230700.0 976200.0 240900.0 962400.0 ;
      RECT  230700.0 976200.0 240900.0 990000.0 ;
      RECT  230700.0 1003800.0 240900.0 990000.0 ;
      RECT  230700.0 1003800.0 240900.0 1017600.0 ;
      RECT  230700.0 1031400.0 240900.0 1017600.0 ;
      RECT  230700.0 1031400.0 240900.0 1045200.0 ;
      RECT  230700.0 1059000.0 240900.0 1045200.0 ;
      RECT  230700.0 1059000.0 240900.0 1072800.0 ;
      RECT  230700.0 1086600.0 240900.0 1072800.0 ;
      RECT  230700.0 1086600.0 240900.0 1100400.0 ;
      RECT  230700.0 1114200.0 240900.0 1100400.0 ;
      RECT  230700.0 1114200.0 240900.0 1128000.0 ;
      RECT  230700.0 1141800.0 240900.0 1128000.0 ;
      RECT  230700.0 1141800.0 240900.0 1155600.0 ;
      RECT  230700.0 1169400.0 240900.0 1155600.0 ;
      RECT  230700.0 1169400.0 240900.0 1183200.0 ;
      RECT  230700.0 1197000.0 240900.0 1183200.0 ;
      RECT  240900.0 313800.0 251100.0 327600.0 ;
      RECT  240900.0 341400.0 251100.0 327600.0 ;
      RECT  240900.0 341400.0 251100.0 355200.0 ;
      RECT  240900.0 369000.0 251100.0 355200.0 ;
      RECT  240900.0 369000.0 251100.0 382800.0 ;
      RECT  240900.0 396600.0 251100.0 382800.0 ;
      RECT  240900.0 396600.0 251100.0 410400.0 ;
      RECT  240900.0 424200.0 251100.0 410400.0 ;
      RECT  240900.0 424200.0 251100.0 438000.0 ;
      RECT  240900.0 451800.0 251100.0 438000.0 ;
      RECT  240900.0 451800.0 251100.0 465600.0 ;
      RECT  240900.0 479400.0 251100.0 465600.0 ;
      RECT  240900.0 479400.0 251100.0 493200.0 ;
      RECT  240900.0 507000.0 251100.0 493200.0 ;
      RECT  240900.0 507000.0 251100.0 520800.0 ;
      RECT  240900.0 534600.0 251100.0 520800.0 ;
      RECT  240900.0 534600.0 251100.0 548400.0 ;
      RECT  240900.0 562200.0 251100.0 548400.0 ;
      RECT  240900.0 562200.0 251100.0 576000.0 ;
      RECT  240900.0 589800.0 251100.0 576000.0 ;
      RECT  240900.0 589800.0 251100.0 603600.0 ;
      RECT  240900.0 617400.0 251100.0 603600.0 ;
      RECT  240900.0 617400.0 251100.0 631200.0 ;
      RECT  240900.0 645000.0 251100.0 631200.0 ;
      RECT  240900.0 645000.0 251100.0 658800.0 ;
      RECT  240900.0 672600.0 251100.0 658800.0 ;
      RECT  240900.0 672600.0 251100.0 686400.0 ;
      RECT  240900.0 700200.0 251100.0 686400.0 ;
      RECT  240900.0 700200.0 251100.0 714000.0 ;
      RECT  240900.0 727800.0 251100.0 714000.0 ;
      RECT  240900.0 727800.0 251100.0 741600.0 ;
      RECT  240900.0 755400.0 251100.0 741600.0 ;
      RECT  240900.0 755400.0 251100.0 769200.0 ;
      RECT  240900.0 783000.0 251100.0 769200.0 ;
      RECT  240900.0 783000.0 251100.0 796800.0 ;
      RECT  240900.0 810600.0 251100.0 796800.0 ;
      RECT  240900.0 810600.0 251100.0 824400.0 ;
      RECT  240900.0 838200.0 251100.0 824400.0 ;
      RECT  240900.0 838200.0 251100.0 852000.0 ;
      RECT  240900.0 865800.0 251100.0 852000.0 ;
      RECT  240900.0 865800.0 251100.0 879600.0 ;
      RECT  240900.0 893400.0 251100.0 879600.0 ;
      RECT  240900.0 893400.0 251100.0 907200.0 ;
      RECT  240900.0 921000.0 251100.0 907200.0 ;
      RECT  240900.0 921000.0 251100.0 934800.0 ;
      RECT  240900.0 948600.0 251100.0 934800.0 ;
      RECT  240900.0 948600.0 251100.0 962400.0 ;
      RECT  240900.0 976200.0 251100.0 962400.0 ;
      RECT  240900.0 976200.0 251100.0 990000.0 ;
      RECT  240900.0 1003800.0 251100.0 990000.0 ;
      RECT  240900.0 1003800.0 251100.0 1017600.0 ;
      RECT  240900.0 1031400.0 251100.0 1017600.0 ;
      RECT  240900.0 1031400.0 251100.0 1045200.0 ;
      RECT  240900.0 1059000.0 251100.0 1045200.0 ;
      RECT  240900.0 1059000.0 251100.0 1072800.0 ;
      RECT  240900.0 1086600.0 251100.0 1072800.0 ;
      RECT  240900.0 1086600.0 251100.0 1100400.0 ;
      RECT  240900.0 1114200.0 251100.0 1100400.0 ;
      RECT  240900.0 1114200.0 251100.0 1128000.0 ;
      RECT  240900.0 1141800.0 251100.0 1128000.0 ;
      RECT  240900.0 1141800.0 251100.0 1155600.0 ;
      RECT  240900.0 1169400.0 251100.0 1155600.0 ;
      RECT  240900.0 1169400.0 251100.0 1183200.0 ;
      RECT  240900.0 1197000.0 251100.0 1183200.0 ;
      RECT  251100.0 313800.0 261300.0 327600.0 ;
      RECT  251100.0 341400.0 261300.0 327600.0 ;
      RECT  251100.0 341400.0 261300.0 355200.0 ;
      RECT  251100.0 369000.0 261300.0 355200.0 ;
      RECT  251100.0 369000.0 261300.0 382800.0 ;
      RECT  251100.0 396600.0 261300.0 382800.0 ;
      RECT  251100.0 396600.0 261300.0 410400.0 ;
      RECT  251100.0 424200.0 261300.0 410400.0 ;
      RECT  251100.0 424200.0 261300.0 438000.0 ;
      RECT  251100.0 451800.0 261300.0 438000.0 ;
      RECT  251100.0 451800.0 261300.0 465600.0 ;
      RECT  251100.0 479400.0 261300.0 465600.0 ;
      RECT  251100.0 479400.0 261300.0 493200.0 ;
      RECT  251100.0 507000.0 261300.0 493200.0 ;
      RECT  251100.0 507000.0 261300.0 520800.0 ;
      RECT  251100.0 534600.0 261300.0 520800.0 ;
      RECT  251100.0 534600.0 261300.0 548400.0 ;
      RECT  251100.0 562200.0 261300.0 548400.0 ;
      RECT  251100.0 562200.0 261300.0 576000.0 ;
      RECT  251100.0 589800.0 261300.0 576000.0 ;
      RECT  251100.0 589800.0 261300.0 603600.0 ;
      RECT  251100.0 617400.0 261300.0 603600.0 ;
      RECT  251100.0 617400.0 261300.0 631200.0 ;
      RECT  251100.0 645000.0 261300.0 631200.0 ;
      RECT  251100.0 645000.0 261300.0 658800.0 ;
      RECT  251100.0 672600.0 261300.0 658800.0 ;
      RECT  251100.0 672600.0 261300.0 686400.0 ;
      RECT  251100.0 700200.0 261300.0 686400.0 ;
      RECT  251100.0 700200.0 261300.0 714000.0 ;
      RECT  251100.0 727800.0 261300.0 714000.0 ;
      RECT  251100.0 727800.0 261300.0 741600.0 ;
      RECT  251100.0 755400.0 261300.0 741600.0 ;
      RECT  251100.0 755400.0 261300.0 769200.0 ;
      RECT  251100.0 783000.0 261300.0 769200.0 ;
      RECT  251100.0 783000.0 261300.0 796800.0 ;
      RECT  251100.0 810600.0 261300.0 796800.0 ;
      RECT  251100.0 810600.0 261300.0 824400.0 ;
      RECT  251100.0 838200.0 261300.0 824400.0 ;
      RECT  251100.0 838200.0 261300.0 852000.0 ;
      RECT  251100.0 865800.0 261300.0 852000.0 ;
      RECT  251100.0 865800.0 261300.0 879600.0 ;
      RECT  251100.0 893400.0 261300.0 879600.0 ;
      RECT  251100.0 893400.0 261300.0 907200.0 ;
      RECT  251100.0 921000.0 261300.0 907200.0 ;
      RECT  251100.0 921000.0 261300.0 934800.0 ;
      RECT  251100.0 948600.0 261300.0 934800.0 ;
      RECT  251100.0 948600.0 261300.0 962400.0 ;
      RECT  251100.0 976200.0 261300.0 962400.0 ;
      RECT  251100.0 976200.0 261300.0 990000.0 ;
      RECT  251100.0 1003800.0 261300.0 990000.0 ;
      RECT  251100.0 1003800.0 261300.0 1017600.0 ;
      RECT  251100.0 1031400.0 261300.0 1017600.0 ;
      RECT  251100.0 1031400.0 261300.0 1045200.0 ;
      RECT  251100.0 1059000.0 261300.0 1045200.0 ;
      RECT  251100.0 1059000.0 261300.0 1072800.0 ;
      RECT  251100.0 1086600.0 261300.0 1072800.0 ;
      RECT  251100.0 1086600.0 261300.0 1100400.0 ;
      RECT  251100.0 1114200.0 261300.0 1100400.0 ;
      RECT  251100.0 1114200.0 261300.0 1128000.0 ;
      RECT  251100.0 1141800.0 261300.0 1128000.0 ;
      RECT  251100.0 1141800.0 261300.0 1155600.0 ;
      RECT  251100.0 1169400.0 261300.0 1155600.0 ;
      RECT  251100.0 1169400.0 261300.0 1183200.0 ;
      RECT  251100.0 1197000.0 261300.0 1183200.0 ;
      RECT  261300.0 313800.0 271500.0 327600.0 ;
      RECT  261300.0 341400.0 271500.0 327600.0 ;
      RECT  261300.0 341400.0 271500.0 355200.0 ;
      RECT  261300.0 369000.0 271500.0 355200.0 ;
      RECT  261300.0 369000.0 271500.0 382800.0 ;
      RECT  261300.0 396600.0 271500.0 382800.0 ;
      RECT  261300.0 396600.0 271500.0 410400.0 ;
      RECT  261300.0 424200.0 271500.0 410400.0 ;
      RECT  261300.0 424200.0 271500.0 438000.0 ;
      RECT  261300.0 451800.0 271500.0 438000.0 ;
      RECT  261300.0 451800.0 271500.0 465600.0 ;
      RECT  261300.0 479400.0 271500.0 465600.0 ;
      RECT  261300.0 479400.0 271500.0 493200.0 ;
      RECT  261300.0 507000.0 271500.0 493200.0 ;
      RECT  261300.0 507000.0 271500.0 520800.0 ;
      RECT  261300.0 534600.0 271500.0 520800.0 ;
      RECT  261300.0 534600.0 271500.0 548400.0 ;
      RECT  261300.0 562200.0 271500.0 548400.0 ;
      RECT  261300.0 562200.0 271500.0 576000.0 ;
      RECT  261300.0 589800.0 271500.0 576000.0 ;
      RECT  261300.0 589800.0 271500.0 603600.0 ;
      RECT  261300.0 617400.0 271500.0 603600.0 ;
      RECT  261300.0 617400.0 271500.0 631200.0 ;
      RECT  261300.0 645000.0 271500.0 631200.0 ;
      RECT  261300.0 645000.0 271500.0 658800.0 ;
      RECT  261300.0 672600.0 271500.0 658800.0 ;
      RECT  261300.0 672600.0 271500.0 686400.0 ;
      RECT  261300.0 700200.0 271500.0 686400.0 ;
      RECT  261300.0 700200.0 271500.0 714000.0 ;
      RECT  261300.0 727800.0 271500.0 714000.0 ;
      RECT  261300.0 727800.0 271500.0 741600.0 ;
      RECT  261300.0 755400.0 271500.0 741600.0 ;
      RECT  261300.0 755400.0 271500.0 769200.0 ;
      RECT  261300.0 783000.0 271500.0 769200.0 ;
      RECT  261300.0 783000.0 271500.0 796800.0 ;
      RECT  261300.0 810600.0 271500.0 796800.0 ;
      RECT  261300.0 810600.0 271500.0 824400.0 ;
      RECT  261300.0 838200.0 271500.0 824400.0 ;
      RECT  261300.0 838200.0 271500.0 852000.0 ;
      RECT  261300.0 865800.0 271500.0 852000.0 ;
      RECT  261300.0 865800.0 271500.0 879600.0 ;
      RECT  261300.0 893400.0 271500.0 879600.0 ;
      RECT  261300.0 893400.0 271500.0 907200.0 ;
      RECT  261300.0 921000.0 271500.0 907200.0 ;
      RECT  261300.0 921000.0 271500.0 934800.0 ;
      RECT  261300.0 948600.0 271500.0 934800.0 ;
      RECT  261300.0 948600.0 271500.0 962400.0 ;
      RECT  261300.0 976200.0 271500.0 962400.0 ;
      RECT  261300.0 976200.0 271500.0 990000.0 ;
      RECT  261300.0 1003800.0 271500.0 990000.0 ;
      RECT  261300.0 1003800.0 271500.0 1017600.0 ;
      RECT  261300.0 1031400.0 271500.0 1017600.0 ;
      RECT  261300.0 1031400.0 271500.0 1045200.0 ;
      RECT  261300.0 1059000.0 271500.0 1045200.0 ;
      RECT  261300.0 1059000.0 271500.0 1072800.0 ;
      RECT  261300.0 1086600.0 271500.0 1072800.0 ;
      RECT  261300.0 1086600.0 271500.0 1100400.0 ;
      RECT  261300.0 1114200.0 271500.0 1100400.0 ;
      RECT  261300.0 1114200.0 271500.0 1128000.0 ;
      RECT  261300.0 1141800.0 271500.0 1128000.0 ;
      RECT  261300.0 1141800.0 271500.0 1155600.0 ;
      RECT  261300.0 1169400.0 271500.0 1155600.0 ;
      RECT  261300.0 1169400.0 271500.0 1183200.0 ;
      RECT  261300.0 1197000.0 271500.0 1183200.0 ;
      RECT  271500.0 313800.0 281700.0 327600.0 ;
      RECT  271500.0 341400.0 281700.0 327600.0 ;
      RECT  271500.0 341400.0 281700.0 355200.0 ;
      RECT  271500.0 369000.0 281700.0 355200.0 ;
      RECT  271500.0 369000.0 281700.0 382800.0 ;
      RECT  271500.0 396600.0 281700.0 382800.0 ;
      RECT  271500.0 396600.0 281700.0 410400.0 ;
      RECT  271500.0 424200.0 281700.0 410400.0 ;
      RECT  271500.0 424200.0 281700.0 438000.0 ;
      RECT  271500.0 451800.0 281700.0 438000.0 ;
      RECT  271500.0 451800.0 281700.0 465600.0 ;
      RECT  271500.0 479400.0 281700.0 465600.0 ;
      RECT  271500.0 479400.0 281700.0 493200.0 ;
      RECT  271500.0 507000.0 281700.0 493200.0 ;
      RECT  271500.0 507000.0 281700.0 520800.0 ;
      RECT  271500.0 534600.0 281700.0 520800.0 ;
      RECT  271500.0 534600.0 281700.0 548400.0 ;
      RECT  271500.0 562200.0 281700.0 548400.0 ;
      RECT  271500.0 562200.0 281700.0 576000.0 ;
      RECT  271500.0 589800.0 281700.0 576000.0 ;
      RECT  271500.0 589800.0 281700.0 603600.0 ;
      RECT  271500.0 617400.0 281700.0 603600.0 ;
      RECT  271500.0 617400.0 281700.0 631200.0 ;
      RECT  271500.0 645000.0 281700.0 631200.0 ;
      RECT  271500.0 645000.0 281700.0 658800.0 ;
      RECT  271500.0 672600.0 281700.0 658800.0 ;
      RECT  271500.0 672600.0 281700.0 686400.0 ;
      RECT  271500.0 700200.0 281700.0 686400.0 ;
      RECT  271500.0 700200.0 281700.0 714000.0 ;
      RECT  271500.0 727800.0 281700.0 714000.0 ;
      RECT  271500.0 727800.0 281700.0 741600.0 ;
      RECT  271500.0 755400.0 281700.0 741600.0 ;
      RECT  271500.0 755400.0 281700.0 769200.0 ;
      RECT  271500.0 783000.0 281700.0 769200.0 ;
      RECT  271500.0 783000.0 281700.0 796800.0 ;
      RECT  271500.0 810600.0 281700.0 796800.0 ;
      RECT  271500.0 810600.0 281700.0 824400.0 ;
      RECT  271500.0 838200.0 281700.0 824400.0 ;
      RECT  271500.0 838200.0 281700.0 852000.0 ;
      RECT  271500.0 865800.0 281700.0 852000.0 ;
      RECT  271500.0 865800.0 281700.0 879600.0 ;
      RECT  271500.0 893400.0 281700.0 879600.0 ;
      RECT  271500.0 893400.0 281700.0 907200.0 ;
      RECT  271500.0 921000.0 281700.0 907200.0 ;
      RECT  271500.0 921000.0 281700.0 934800.0 ;
      RECT  271500.0 948600.0 281700.0 934800.0 ;
      RECT  271500.0 948600.0 281700.0 962400.0 ;
      RECT  271500.0 976200.0 281700.0 962400.0 ;
      RECT  271500.0 976200.0 281700.0 990000.0 ;
      RECT  271500.0 1003800.0 281700.0 990000.0 ;
      RECT  271500.0 1003800.0 281700.0 1017600.0 ;
      RECT  271500.0 1031400.0 281700.0 1017600.0 ;
      RECT  271500.0 1031400.0 281700.0 1045200.0 ;
      RECT  271500.0 1059000.0 281700.0 1045200.0 ;
      RECT  271500.0 1059000.0 281700.0 1072800.0 ;
      RECT  271500.0 1086600.0 281700.0 1072800.0 ;
      RECT  271500.0 1086600.0 281700.0 1100400.0 ;
      RECT  271500.0 1114200.0 281700.0 1100400.0 ;
      RECT  271500.0 1114200.0 281700.0 1128000.0 ;
      RECT  271500.0 1141800.0 281700.0 1128000.0 ;
      RECT  271500.0 1141800.0 281700.0 1155600.0 ;
      RECT  271500.0 1169400.0 281700.0 1155600.0 ;
      RECT  271500.0 1169400.0 281700.0 1183200.0 ;
      RECT  271500.0 1197000.0 281700.0 1183200.0 ;
      RECT  281700.0 313800.0 291900.0 327600.0 ;
      RECT  281700.0 341400.0 291900.0 327600.0 ;
      RECT  281700.0 341400.0 291900.0 355200.0 ;
      RECT  281700.0 369000.0 291900.0 355200.0 ;
      RECT  281700.0 369000.0 291900.0 382800.0 ;
      RECT  281700.0 396600.0 291900.0 382800.0 ;
      RECT  281700.0 396600.0 291900.0 410400.0 ;
      RECT  281700.0 424200.0 291900.0 410400.0 ;
      RECT  281700.0 424200.0 291900.0 438000.0 ;
      RECT  281700.0 451800.0 291900.0 438000.0 ;
      RECT  281700.0 451800.0 291900.0 465600.0 ;
      RECT  281700.0 479400.0 291900.0 465600.0 ;
      RECT  281700.0 479400.0 291900.0 493200.0 ;
      RECT  281700.0 507000.0 291900.0 493200.0 ;
      RECT  281700.0 507000.0 291900.0 520800.0 ;
      RECT  281700.0 534600.0 291900.0 520800.0 ;
      RECT  281700.0 534600.0 291900.0 548400.0 ;
      RECT  281700.0 562200.0 291900.0 548400.0 ;
      RECT  281700.0 562200.0 291900.0 576000.0 ;
      RECT  281700.0 589800.0 291900.0 576000.0 ;
      RECT  281700.0 589800.0 291900.0 603600.0 ;
      RECT  281700.0 617400.0 291900.0 603600.0 ;
      RECT  281700.0 617400.0 291900.0 631200.0 ;
      RECT  281700.0 645000.0 291900.0 631200.0 ;
      RECT  281700.0 645000.0 291900.0 658800.0 ;
      RECT  281700.0 672600.0 291900.0 658800.0 ;
      RECT  281700.0 672600.0 291900.0 686400.0 ;
      RECT  281700.0 700200.0 291900.0 686400.0 ;
      RECT  281700.0 700200.0 291900.0 714000.0 ;
      RECT  281700.0 727800.0 291900.0 714000.0 ;
      RECT  281700.0 727800.0 291900.0 741600.0 ;
      RECT  281700.0 755400.0 291900.0 741600.0 ;
      RECT  281700.0 755400.0 291900.0 769200.0 ;
      RECT  281700.0 783000.0 291900.0 769200.0 ;
      RECT  281700.0 783000.0 291900.0 796800.0 ;
      RECT  281700.0 810600.0 291900.0 796800.0 ;
      RECT  281700.0 810600.0 291900.0 824400.0 ;
      RECT  281700.0 838200.0 291900.0 824400.0 ;
      RECT  281700.0 838200.0 291900.0 852000.0 ;
      RECT  281700.0 865800.0 291900.0 852000.0 ;
      RECT  281700.0 865800.0 291900.0 879600.0 ;
      RECT  281700.0 893400.0 291900.0 879600.0 ;
      RECT  281700.0 893400.0 291900.0 907200.0 ;
      RECT  281700.0 921000.0 291900.0 907200.0 ;
      RECT  281700.0 921000.0 291900.0 934800.0 ;
      RECT  281700.0 948600.0 291900.0 934800.0 ;
      RECT  281700.0 948600.0 291900.0 962400.0 ;
      RECT  281700.0 976200.0 291900.0 962400.0 ;
      RECT  281700.0 976200.0 291900.0 990000.0 ;
      RECT  281700.0 1003800.0 291900.0 990000.0 ;
      RECT  281700.0 1003800.0 291900.0 1017600.0 ;
      RECT  281700.0 1031400.0 291900.0 1017600.0 ;
      RECT  281700.0 1031400.0 291900.0 1045200.0 ;
      RECT  281700.0 1059000.0 291900.0 1045200.0 ;
      RECT  281700.0 1059000.0 291900.0 1072800.0 ;
      RECT  281700.0 1086600.0 291900.0 1072800.0 ;
      RECT  281700.0 1086600.0 291900.0 1100400.0 ;
      RECT  281700.0 1114200.0 291900.0 1100400.0 ;
      RECT  281700.0 1114200.0 291900.0 1128000.0 ;
      RECT  281700.0 1141800.0 291900.0 1128000.0 ;
      RECT  281700.0 1141800.0 291900.0 1155600.0 ;
      RECT  281700.0 1169400.0 291900.0 1155600.0 ;
      RECT  281700.0 1169400.0 291900.0 1183200.0 ;
      RECT  281700.0 1197000.0 291900.0 1183200.0 ;
      RECT  291900.0 313800.0 302100.0 327600.0 ;
      RECT  291900.0 341400.0 302100.0 327600.0 ;
      RECT  291900.0 341400.0 302100.0 355200.0 ;
      RECT  291900.0 369000.0 302100.0 355200.0 ;
      RECT  291900.0 369000.0 302100.0 382800.0 ;
      RECT  291900.0 396600.0 302100.0 382800.0 ;
      RECT  291900.0 396600.0 302100.0 410400.0 ;
      RECT  291900.0 424200.0 302100.0 410400.0 ;
      RECT  291900.0 424200.0 302100.0 438000.0 ;
      RECT  291900.0 451800.0 302100.0 438000.0 ;
      RECT  291900.0 451800.0 302100.0 465600.0 ;
      RECT  291900.0 479400.0 302100.0 465600.0 ;
      RECT  291900.0 479400.0 302100.0 493200.0 ;
      RECT  291900.0 507000.0 302100.0 493200.0 ;
      RECT  291900.0 507000.0 302100.0 520800.0 ;
      RECT  291900.0 534600.0 302100.0 520800.0 ;
      RECT  291900.0 534600.0 302100.0 548400.0 ;
      RECT  291900.0 562200.0 302100.0 548400.0 ;
      RECT  291900.0 562200.0 302100.0 576000.0 ;
      RECT  291900.0 589800.0 302100.0 576000.0 ;
      RECT  291900.0 589800.0 302100.0 603600.0 ;
      RECT  291900.0 617400.0 302100.0 603600.0 ;
      RECT  291900.0 617400.0 302100.0 631200.0 ;
      RECT  291900.0 645000.0 302100.0 631200.0 ;
      RECT  291900.0 645000.0 302100.0 658800.0 ;
      RECT  291900.0 672600.0 302100.0 658800.0 ;
      RECT  291900.0 672600.0 302100.0 686400.0 ;
      RECT  291900.0 700200.0 302100.0 686400.0 ;
      RECT  291900.0 700200.0 302100.0 714000.0 ;
      RECT  291900.0 727800.0 302100.0 714000.0 ;
      RECT  291900.0 727800.0 302100.0 741600.0 ;
      RECT  291900.0 755400.0 302100.0 741600.0 ;
      RECT  291900.0 755400.0 302100.0 769200.0 ;
      RECT  291900.0 783000.0 302100.0 769200.0 ;
      RECT  291900.0 783000.0 302100.0 796800.0 ;
      RECT  291900.0 810600.0 302100.0 796800.0 ;
      RECT  291900.0 810600.0 302100.0 824400.0 ;
      RECT  291900.0 838200.0 302100.0 824400.0 ;
      RECT  291900.0 838200.0 302100.0 852000.0 ;
      RECT  291900.0 865800.0 302100.0 852000.0 ;
      RECT  291900.0 865800.0 302100.0 879600.0 ;
      RECT  291900.0 893400.0 302100.0 879600.0 ;
      RECT  291900.0 893400.0 302100.0 907200.0 ;
      RECT  291900.0 921000.0 302100.0 907200.0 ;
      RECT  291900.0 921000.0 302100.0 934800.0 ;
      RECT  291900.0 948600.0 302100.0 934800.0 ;
      RECT  291900.0 948600.0 302100.0 962400.0 ;
      RECT  291900.0 976200.0 302100.0 962400.0 ;
      RECT  291900.0 976200.0 302100.0 990000.0 ;
      RECT  291900.0 1003800.0 302100.0 990000.0 ;
      RECT  291900.0 1003800.0 302100.0 1017600.0 ;
      RECT  291900.0 1031400.0 302100.0 1017600.0 ;
      RECT  291900.0 1031400.0 302100.0 1045200.0 ;
      RECT  291900.0 1059000.0 302100.0 1045200.0 ;
      RECT  291900.0 1059000.0 302100.0 1072800.0 ;
      RECT  291900.0 1086600.0 302100.0 1072800.0 ;
      RECT  291900.0 1086600.0 302100.0 1100400.0 ;
      RECT  291900.0 1114200.0 302100.0 1100400.0 ;
      RECT  291900.0 1114200.0 302100.0 1128000.0 ;
      RECT  291900.0 1141800.0 302100.0 1128000.0 ;
      RECT  291900.0 1141800.0 302100.0 1155600.0 ;
      RECT  291900.0 1169400.0 302100.0 1155600.0 ;
      RECT  291900.0 1169400.0 302100.0 1183200.0 ;
      RECT  291900.0 1197000.0 302100.0 1183200.0 ;
      RECT  302100.0 313800.0 312300.0 327600.0 ;
      RECT  302100.0 341400.0 312300.0 327600.0 ;
      RECT  302100.0 341400.0 312300.0 355200.0 ;
      RECT  302100.0 369000.0 312300.0 355200.0 ;
      RECT  302100.0 369000.0 312300.0 382800.0 ;
      RECT  302100.0 396600.0 312300.0 382800.0 ;
      RECT  302100.0 396600.0 312300.0 410400.0 ;
      RECT  302100.0 424200.0 312300.0 410400.0 ;
      RECT  302100.0 424200.0 312300.0 438000.0 ;
      RECT  302100.0 451800.0 312300.0 438000.0 ;
      RECT  302100.0 451800.0 312300.0 465600.0 ;
      RECT  302100.0 479400.0 312300.0 465600.0 ;
      RECT  302100.0 479400.0 312300.0 493200.0 ;
      RECT  302100.0 507000.0 312300.0 493200.0 ;
      RECT  302100.0 507000.0 312300.0 520800.0 ;
      RECT  302100.0 534600.0 312300.0 520800.0 ;
      RECT  302100.0 534600.0 312300.0 548400.0 ;
      RECT  302100.0 562200.0 312300.0 548400.0 ;
      RECT  302100.0 562200.0 312300.0 576000.0 ;
      RECT  302100.0 589800.0 312300.0 576000.0 ;
      RECT  302100.0 589800.0 312300.0 603600.0 ;
      RECT  302100.0 617400.0 312300.0 603600.0 ;
      RECT  302100.0 617400.0 312300.0 631200.0 ;
      RECT  302100.0 645000.0 312300.0 631200.0 ;
      RECT  302100.0 645000.0 312300.0 658800.0 ;
      RECT  302100.0 672600.0 312300.0 658800.0 ;
      RECT  302100.0 672600.0 312300.0 686400.0 ;
      RECT  302100.0 700200.0 312300.0 686400.0 ;
      RECT  302100.0 700200.0 312300.0 714000.0 ;
      RECT  302100.0 727800.0 312300.0 714000.0 ;
      RECT  302100.0 727800.0 312300.0 741600.0 ;
      RECT  302100.0 755400.0 312300.0 741600.0 ;
      RECT  302100.0 755400.0 312300.0 769200.0 ;
      RECT  302100.0 783000.0 312300.0 769200.0 ;
      RECT  302100.0 783000.0 312300.0 796800.0 ;
      RECT  302100.0 810600.0 312300.0 796800.0 ;
      RECT  302100.0 810600.0 312300.0 824400.0 ;
      RECT  302100.0 838200.0 312300.0 824400.0 ;
      RECT  302100.0 838200.0 312300.0 852000.0 ;
      RECT  302100.0 865800.0 312300.0 852000.0 ;
      RECT  302100.0 865800.0 312300.0 879600.0 ;
      RECT  302100.0 893400.0 312300.0 879600.0 ;
      RECT  302100.0 893400.0 312300.0 907200.0 ;
      RECT  302100.0 921000.0 312300.0 907200.0 ;
      RECT  302100.0 921000.0 312300.0 934800.0 ;
      RECT  302100.0 948600.0 312300.0 934800.0 ;
      RECT  302100.0 948600.0 312300.0 962400.0 ;
      RECT  302100.0 976200.0 312300.0 962400.0 ;
      RECT  302100.0 976200.0 312300.0 990000.0 ;
      RECT  302100.0 1003800.0 312300.0 990000.0 ;
      RECT  302100.0 1003800.0 312300.0 1017600.0 ;
      RECT  302100.0 1031400.0 312300.0 1017600.0 ;
      RECT  302100.0 1031400.0 312300.0 1045200.0 ;
      RECT  302100.0 1059000.0 312300.0 1045200.0 ;
      RECT  302100.0 1059000.0 312300.0 1072800.0 ;
      RECT  302100.0 1086600.0 312300.0 1072800.0 ;
      RECT  302100.0 1086600.0 312300.0 1100400.0 ;
      RECT  302100.0 1114200.0 312300.0 1100400.0 ;
      RECT  302100.0 1114200.0 312300.0 1128000.0 ;
      RECT  302100.0 1141800.0 312300.0 1128000.0 ;
      RECT  302100.0 1141800.0 312300.0 1155600.0 ;
      RECT  302100.0 1169400.0 312300.0 1155600.0 ;
      RECT  302100.0 1169400.0 312300.0 1183200.0 ;
      RECT  302100.0 1197000.0 312300.0 1183200.0 ;
      RECT  312300.0 313800.0 322500.0 327600.0 ;
      RECT  312300.0 341400.0 322500.0 327600.0 ;
      RECT  312300.0 341400.0 322500.0 355200.0 ;
      RECT  312300.0 369000.0 322500.0 355200.0 ;
      RECT  312300.0 369000.0 322500.0 382800.0 ;
      RECT  312300.0 396600.0 322500.0 382800.0 ;
      RECT  312300.0 396600.0 322500.0 410400.0 ;
      RECT  312300.0 424200.0 322500.0 410400.0 ;
      RECT  312300.0 424200.0 322500.0 438000.0 ;
      RECT  312300.0 451800.0 322500.0 438000.0 ;
      RECT  312300.0 451800.0 322500.0 465600.0 ;
      RECT  312300.0 479400.0 322500.0 465600.0 ;
      RECT  312300.0 479400.0 322500.0 493200.0 ;
      RECT  312300.0 507000.0 322500.0 493200.0 ;
      RECT  312300.0 507000.0 322500.0 520800.0 ;
      RECT  312300.0 534600.0 322500.0 520800.0 ;
      RECT  312300.0 534600.0 322500.0 548400.0 ;
      RECT  312300.0 562200.0 322500.0 548400.0 ;
      RECT  312300.0 562200.0 322500.0 576000.0 ;
      RECT  312300.0 589800.0 322500.0 576000.0 ;
      RECT  312300.0 589800.0 322500.0 603600.0 ;
      RECT  312300.0 617400.0 322500.0 603600.0 ;
      RECT  312300.0 617400.0 322500.0 631200.0 ;
      RECT  312300.0 645000.0 322500.0 631200.0 ;
      RECT  312300.0 645000.0 322500.0 658800.0 ;
      RECT  312300.0 672600.0 322500.0 658800.0 ;
      RECT  312300.0 672600.0 322500.0 686400.0 ;
      RECT  312300.0 700200.0 322500.0 686400.0 ;
      RECT  312300.0 700200.0 322500.0 714000.0 ;
      RECT  312300.0 727800.0 322500.0 714000.0 ;
      RECT  312300.0 727800.0 322500.0 741600.0 ;
      RECT  312300.0 755400.0 322500.0 741600.0 ;
      RECT  312300.0 755400.0 322500.0 769200.0 ;
      RECT  312300.0 783000.0 322500.0 769200.0 ;
      RECT  312300.0 783000.0 322500.0 796800.0 ;
      RECT  312300.0 810600.0 322500.0 796800.0 ;
      RECT  312300.0 810600.0 322500.0 824400.0 ;
      RECT  312300.0 838200.0 322500.0 824400.0 ;
      RECT  312300.0 838200.0 322500.0 852000.0 ;
      RECT  312300.0 865800.0 322500.0 852000.0 ;
      RECT  312300.0 865800.0 322500.0 879600.0 ;
      RECT  312300.0 893400.0 322500.0 879600.0 ;
      RECT  312300.0 893400.0 322500.0 907200.0 ;
      RECT  312300.0 921000.0 322500.0 907200.0 ;
      RECT  312300.0 921000.0 322500.0 934800.0 ;
      RECT  312300.0 948600.0 322500.0 934800.0 ;
      RECT  312300.0 948600.0 322500.0 962400.0 ;
      RECT  312300.0 976200.0 322500.0 962400.0 ;
      RECT  312300.0 976200.0 322500.0 990000.0 ;
      RECT  312300.0 1003800.0 322500.0 990000.0 ;
      RECT  312300.0 1003800.0 322500.0 1017600.0 ;
      RECT  312300.0 1031400.0 322500.0 1017600.0 ;
      RECT  312300.0 1031400.0 322500.0 1045200.0 ;
      RECT  312300.0 1059000.0 322500.0 1045200.0 ;
      RECT  312300.0 1059000.0 322500.0 1072800.0 ;
      RECT  312300.0 1086600.0 322500.0 1072800.0 ;
      RECT  312300.0 1086600.0 322500.0 1100400.0 ;
      RECT  312300.0 1114200.0 322500.0 1100400.0 ;
      RECT  312300.0 1114200.0 322500.0 1128000.0 ;
      RECT  312300.0 1141800.0 322500.0 1128000.0 ;
      RECT  312300.0 1141800.0 322500.0 1155600.0 ;
      RECT  312300.0 1169400.0 322500.0 1155600.0 ;
      RECT  312300.0 1169400.0 322500.0 1183200.0 ;
      RECT  312300.0 1197000.0 322500.0 1183200.0 ;
      RECT  322500.0 313800.0 332700.0 327600.0 ;
      RECT  322500.0 341400.0 332700.0 327600.0 ;
      RECT  322500.0 341400.0 332700.0 355200.0 ;
      RECT  322500.0 369000.0 332700.0 355200.0 ;
      RECT  322500.0 369000.0 332700.0 382800.0 ;
      RECT  322500.0 396600.0 332700.0 382800.0 ;
      RECT  322500.0 396600.0 332700.0 410400.0 ;
      RECT  322500.0 424200.0 332700.0 410400.0 ;
      RECT  322500.0 424200.0 332700.0 438000.0 ;
      RECT  322500.0 451800.0 332700.0 438000.0 ;
      RECT  322500.0 451800.0 332700.0 465600.0 ;
      RECT  322500.0 479400.0 332700.0 465600.0 ;
      RECT  322500.0 479400.0 332700.0 493200.0 ;
      RECT  322500.0 507000.0 332700.0 493200.0 ;
      RECT  322500.0 507000.0 332700.0 520800.0 ;
      RECT  322500.0 534600.0 332700.0 520800.0 ;
      RECT  322500.0 534600.0 332700.0 548400.0 ;
      RECT  322500.0 562200.0 332700.0 548400.0 ;
      RECT  322500.0 562200.0 332700.0 576000.0 ;
      RECT  322500.0 589800.0 332700.0 576000.0 ;
      RECT  322500.0 589800.0 332700.0 603600.0 ;
      RECT  322500.0 617400.0 332700.0 603600.0 ;
      RECT  322500.0 617400.0 332700.0 631200.0 ;
      RECT  322500.0 645000.0 332700.0 631200.0 ;
      RECT  322500.0 645000.0 332700.0 658800.0 ;
      RECT  322500.0 672600.0 332700.0 658800.0 ;
      RECT  322500.0 672600.0 332700.0 686400.0 ;
      RECT  322500.0 700200.0 332700.0 686400.0 ;
      RECT  322500.0 700200.0 332700.0 714000.0 ;
      RECT  322500.0 727800.0 332700.0 714000.0 ;
      RECT  322500.0 727800.0 332700.0 741600.0 ;
      RECT  322500.0 755400.0 332700.0 741600.0 ;
      RECT  322500.0 755400.0 332700.0 769200.0 ;
      RECT  322500.0 783000.0 332700.0 769200.0 ;
      RECT  322500.0 783000.0 332700.0 796800.0 ;
      RECT  322500.0 810600.0 332700.0 796800.0 ;
      RECT  322500.0 810600.0 332700.0 824400.0 ;
      RECT  322500.0 838200.0 332700.0 824400.0 ;
      RECT  322500.0 838200.0 332700.0 852000.0 ;
      RECT  322500.0 865800.0 332700.0 852000.0 ;
      RECT  322500.0 865800.0 332700.0 879600.0 ;
      RECT  322500.0 893400.0 332700.0 879600.0 ;
      RECT  322500.0 893400.0 332700.0 907200.0 ;
      RECT  322500.0 921000.0 332700.0 907200.0 ;
      RECT  322500.0 921000.0 332700.0 934800.0 ;
      RECT  322500.0 948600.0 332700.0 934800.0 ;
      RECT  322500.0 948600.0 332700.0 962400.0 ;
      RECT  322500.0 976200.0 332700.0 962400.0 ;
      RECT  322500.0 976200.0 332700.0 990000.0 ;
      RECT  322500.0 1003800.0 332700.0 990000.0 ;
      RECT  322500.0 1003800.0 332700.0 1017600.0 ;
      RECT  322500.0 1031400.0 332700.0 1017600.0 ;
      RECT  322500.0 1031400.0 332700.0 1045200.0 ;
      RECT  322500.0 1059000.0 332700.0 1045200.0 ;
      RECT  322500.0 1059000.0 332700.0 1072800.0 ;
      RECT  322500.0 1086600.0 332700.0 1072800.0 ;
      RECT  322500.0 1086600.0 332700.0 1100400.0 ;
      RECT  322500.0 1114200.0 332700.0 1100400.0 ;
      RECT  322500.0 1114200.0 332700.0 1128000.0 ;
      RECT  322500.0 1141800.0 332700.0 1128000.0 ;
      RECT  322500.0 1141800.0 332700.0 1155600.0 ;
      RECT  322500.0 1169400.0 332700.0 1155600.0 ;
      RECT  322500.0 1169400.0 332700.0 1183200.0 ;
      RECT  322500.0 1197000.0 332700.0 1183200.0 ;
      RECT  332700.0 313800.0 342900.0 327600.0 ;
      RECT  332700.0 341400.0 342900.0 327600.0 ;
      RECT  332700.0 341400.0 342900.0 355200.0 ;
      RECT  332700.0 369000.0 342900.0 355200.0 ;
      RECT  332700.0 369000.0 342900.0 382800.0 ;
      RECT  332700.0 396600.0 342900.0 382800.0 ;
      RECT  332700.0 396600.0 342900.0 410400.0 ;
      RECT  332700.0 424200.0 342900.0 410400.0 ;
      RECT  332700.0 424200.0 342900.0 438000.0 ;
      RECT  332700.0 451800.0 342900.0 438000.0 ;
      RECT  332700.0 451800.0 342900.0 465600.0 ;
      RECT  332700.0 479400.0 342900.0 465600.0 ;
      RECT  332700.0 479400.0 342900.0 493200.0 ;
      RECT  332700.0 507000.0 342900.0 493200.0 ;
      RECT  332700.0 507000.0 342900.0 520800.0 ;
      RECT  332700.0 534600.0 342900.0 520800.0 ;
      RECT  332700.0 534600.0 342900.0 548400.0 ;
      RECT  332700.0 562200.0 342900.0 548400.0 ;
      RECT  332700.0 562200.0 342900.0 576000.0 ;
      RECT  332700.0 589800.0 342900.0 576000.0 ;
      RECT  332700.0 589800.0 342900.0 603600.0 ;
      RECT  332700.0 617400.0 342900.0 603600.0 ;
      RECT  332700.0 617400.0 342900.0 631200.0 ;
      RECT  332700.0 645000.0 342900.0 631200.0 ;
      RECT  332700.0 645000.0 342900.0 658800.0 ;
      RECT  332700.0 672600.0 342900.0 658800.0 ;
      RECT  332700.0 672600.0 342900.0 686400.0 ;
      RECT  332700.0 700200.0 342900.0 686400.0 ;
      RECT  332700.0 700200.0 342900.0 714000.0 ;
      RECT  332700.0 727800.0 342900.0 714000.0 ;
      RECT  332700.0 727800.0 342900.0 741600.0 ;
      RECT  332700.0 755400.0 342900.0 741600.0 ;
      RECT  332700.0 755400.0 342900.0 769200.0 ;
      RECT  332700.0 783000.0 342900.0 769200.0 ;
      RECT  332700.0 783000.0 342900.0 796800.0 ;
      RECT  332700.0 810600.0 342900.0 796800.0 ;
      RECT  332700.0 810600.0 342900.0 824400.0 ;
      RECT  332700.0 838200.0 342900.0 824400.0 ;
      RECT  332700.0 838200.0 342900.0 852000.0 ;
      RECT  332700.0 865800.0 342900.0 852000.0 ;
      RECT  332700.0 865800.0 342900.0 879600.0 ;
      RECT  332700.0 893400.0 342900.0 879600.0 ;
      RECT  332700.0 893400.0 342900.0 907200.0 ;
      RECT  332700.0 921000.0 342900.0 907200.0 ;
      RECT  332700.0 921000.0 342900.0 934800.0 ;
      RECT  332700.0 948600.0 342900.0 934800.0 ;
      RECT  332700.0 948600.0 342900.0 962400.0 ;
      RECT  332700.0 976200.0 342900.0 962400.0 ;
      RECT  332700.0 976200.0 342900.0 990000.0 ;
      RECT  332700.0 1003800.0 342900.0 990000.0 ;
      RECT  332700.0 1003800.0 342900.0 1017600.0 ;
      RECT  332700.0 1031400.0 342900.0 1017600.0 ;
      RECT  332700.0 1031400.0 342900.0 1045200.0 ;
      RECT  332700.0 1059000.0 342900.0 1045200.0 ;
      RECT  332700.0 1059000.0 342900.0 1072800.0 ;
      RECT  332700.0 1086600.0 342900.0 1072800.0 ;
      RECT  332700.0 1086600.0 342900.0 1100400.0 ;
      RECT  332700.0 1114200.0 342900.0 1100400.0 ;
      RECT  332700.0 1114200.0 342900.0 1128000.0 ;
      RECT  332700.0 1141800.0 342900.0 1128000.0 ;
      RECT  332700.0 1141800.0 342900.0 1155600.0 ;
      RECT  332700.0 1169400.0 342900.0 1155600.0 ;
      RECT  332700.0 1169400.0 342900.0 1183200.0 ;
      RECT  332700.0 1197000.0 342900.0 1183200.0 ;
      RECT  342900.0 313800.0 353100.0 327600.0 ;
      RECT  342900.0 341400.0 353100.0 327600.0 ;
      RECT  342900.0 341400.0 353100.0 355200.0 ;
      RECT  342900.0 369000.0 353100.0 355200.0 ;
      RECT  342900.0 369000.0 353100.0 382800.0 ;
      RECT  342900.0 396600.0 353100.0 382800.0 ;
      RECT  342900.0 396600.0 353100.0 410400.0 ;
      RECT  342900.0 424200.0 353100.0 410400.0 ;
      RECT  342900.0 424200.0 353100.0 438000.0 ;
      RECT  342900.0 451800.0 353100.0 438000.0 ;
      RECT  342900.0 451800.0 353100.0 465600.0 ;
      RECT  342900.0 479400.0 353100.0 465600.0 ;
      RECT  342900.0 479400.0 353100.0 493200.0 ;
      RECT  342900.0 507000.0 353100.0 493200.0 ;
      RECT  342900.0 507000.0 353100.0 520800.0 ;
      RECT  342900.0 534600.0 353100.0 520800.0 ;
      RECT  342900.0 534600.0 353100.0 548400.0 ;
      RECT  342900.0 562200.0 353100.0 548400.0 ;
      RECT  342900.0 562200.0 353100.0 576000.0 ;
      RECT  342900.0 589800.0 353100.0 576000.0 ;
      RECT  342900.0 589800.0 353100.0 603600.0 ;
      RECT  342900.0 617400.0 353100.0 603600.0 ;
      RECT  342900.0 617400.0 353100.0 631200.0 ;
      RECT  342900.0 645000.0 353100.0 631200.0 ;
      RECT  342900.0 645000.0 353100.0 658800.0 ;
      RECT  342900.0 672600.0 353100.0 658800.0 ;
      RECT  342900.0 672600.0 353100.0 686400.0 ;
      RECT  342900.0 700200.0 353100.0 686400.0 ;
      RECT  342900.0 700200.0 353100.0 714000.0 ;
      RECT  342900.0 727800.0 353100.0 714000.0 ;
      RECT  342900.0 727800.0 353100.0 741600.0 ;
      RECT  342900.0 755400.0 353100.0 741600.0 ;
      RECT  342900.0 755400.0 353100.0 769200.0 ;
      RECT  342900.0 783000.0 353100.0 769200.0 ;
      RECT  342900.0 783000.0 353100.0 796800.0 ;
      RECT  342900.0 810600.0 353100.0 796800.0 ;
      RECT  342900.0 810600.0 353100.0 824400.0 ;
      RECT  342900.0 838200.0 353100.0 824400.0 ;
      RECT  342900.0 838200.0 353100.0 852000.0 ;
      RECT  342900.0 865800.0 353100.0 852000.0 ;
      RECT  342900.0 865800.0 353100.0 879600.0 ;
      RECT  342900.0 893400.0 353100.0 879600.0 ;
      RECT  342900.0 893400.0 353100.0 907200.0 ;
      RECT  342900.0 921000.0 353100.0 907200.0 ;
      RECT  342900.0 921000.0 353100.0 934800.0 ;
      RECT  342900.0 948600.0 353100.0 934800.0 ;
      RECT  342900.0 948600.0 353100.0 962400.0 ;
      RECT  342900.0 976200.0 353100.0 962400.0 ;
      RECT  342900.0 976200.0 353100.0 990000.0 ;
      RECT  342900.0 1003800.0 353100.0 990000.0 ;
      RECT  342900.0 1003800.0 353100.0 1017600.0 ;
      RECT  342900.0 1031400.0 353100.0 1017600.0 ;
      RECT  342900.0 1031400.0 353100.0 1045200.0 ;
      RECT  342900.0 1059000.0 353100.0 1045200.0 ;
      RECT  342900.0 1059000.0 353100.0 1072800.0 ;
      RECT  342900.0 1086600.0 353100.0 1072800.0 ;
      RECT  342900.0 1086600.0 353100.0 1100400.0 ;
      RECT  342900.0 1114200.0 353100.0 1100400.0 ;
      RECT  342900.0 1114200.0 353100.0 1128000.0 ;
      RECT  342900.0 1141800.0 353100.0 1128000.0 ;
      RECT  342900.0 1141800.0 353100.0 1155600.0 ;
      RECT  342900.0 1169400.0 353100.0 1155600.0 ;
      RECT  342900.0 1169400.0 353100.0 1183200.0 ;
      RECT  342900.0 1197000.0 353100.0 1183200.0 ;
      RECT  353100.0 313800.0 363300.0 327600.0 ;
      RECT  353100.0 341400.0 363300.0 327600.0 ;
      RECT  353100.0 341400.0 363300.0 355200.0 ;
      RECT  353100.0 369000.0 363300.0 355200.0 ;
      RECT  353100.0 369000.0 363300.0 382800.0 ;
      RECT  353100.0 396600.0 363300.0 382800.0 ;
      RECT  353100.0 396600.0 363300.0 410400.0 ;
      RECT  353100.0 424200.0 363300.0 410400.0 ;
      RECT  353100.0 424200.0 363300.0 438000.0 ;
      RECT  353100.0 451800.0 363300.0 438000.0 ;
      RECT  353100.0 451800.0 363300.0 465600.0 ;
      RECT  353100.0 479400.0 363300.0 465600.0 ;
      RECT  353100.0 479400.0 363300.0 493200.0 ;
      RECT  353100.0 507000.0 363300.0 493200.0 ;
      RECT  353100.0 507000.0 363300.0 520800.0 ;
      RECT  353100.0 534600.0 363300.0 520800.0 ;
      RECT  353100.0 534600.0 363300.0 548400.0 ;
      RECT  353100.0 562200.0 363300.0 548400.0 ;
      RECT  353100.0 562200.0 363300.0 576000.0 ;
      RECT  353100.0 589800.0 363300.0 576000.0 ;
      RECT  353100.0 589800.0 363300.0 603600.0 ;
      RECT  353100.0 617400.0 363300.0 603600.0 ;
      RECT  353100.0 617400.0 363300.0 631200.0 ;
      RECT  353100.0 645000.0 363300.0 631200.0 ;
      RECT  353100.0 645000.0 363300.0 658800.0 ;
      RECT  353100.0 672600.0 363300.0 658800.0 ;
      RECT  353100.0 672600.0 363300.0 686400.0 ;
      RECT  353100.0 700200.0 363300.0 686400.0 ;
      RECT  353100.0 700200.0 363300.0 714000.0 ;
      RECT  353100.0 727800.0 363300.0 714000.0 ;
      RECT  353100.0 727800.0 363300.0 741600.0 ;
      RECT  353100.0 755400.0 363300.0 741600.0 ;
      RECT  353100.0 755400.0 363300.0 769200.0 ;
      RECT  353100.0 783000.0 363300.0 769200.0 ;
      RECT  353100.0 783000.0 363300.0 796800.0 ;
      RECT  353100.0 810600.0 363300.0 796800.0 ;
      RECT  353100.0 810600.0 363300.0 824400.0 ;
      RECT  353100.0 838200.0 363300.0 824400.0 ;
      RECT  353100.0 838200.0 363300.0 852000.0 ;
      RECT  353100.0 865800.0 363300.0 852000.0 ;
      RECT  353100.0 865800.0 363300.0 879600.0 ;
      RECT  353100.0 893400.0 363300.0 879600.0 ;
      RECT  353100.0 893400.0 363300.0 907200.0 ;
      RECT  353100.0 921000.0 363300.0 907200.0 ;
      RECT  353100.0 921000.0 363300.0 934800.0 ;
      RECT  353100.0 948600.0 363300.0 934800.0 ;
      RECT  353100.0 948600.0 363300.0 962400.0 ;
      RECT  353100.0 976200.0 363300.0 962400.0 ;
      RECT  353100.0 976200.0 363300.0 990000.0 ;
      RECT  353100.0 1003800.0 363300.0 990000.0 ;
      RECT  353100.0 1003800.0 363300.0 1017600.0 ;
      RECT  353100.0 1031400.0 363300.0 1017600.0 ;
      RECT  353100.0 1031400.0 363300.0 1045200.0 ;
      RECT  353100.0 1059000.0 363300.0 1045200.0 ;
      RECT  353100.0 1059000.0 363300.0 1072800.0 ;
      RECT  353100.0 1086600.0 363300.0 1072800.0 ;
      RECT  353100.0 1086600.0 363300.0 1100400.0 ;
      RECT  353100.0 1114200.0 363300.0 1100400.0 ;
      RECT  353100.0 1114200.0 363300.0 1128000.0 ;
      RECT  353100.0 1141800.0 363300.0 1128000.0 ;
      RECT  353100.0 1141800.0 363300.0 1155600.0 ;
      RECT  353100.0 1169400.0 363300.0 1155600.0 ;
      RECT  353100.0 1169400.0 363300.0 1183200.0 ;
      RECT  353100.0 1197000.0 363300.0 1183200.0 ;
      RECT  363300.0 313800.0 373500.0 327600.0 ;
      RECT  363300.0 341400.0 373500.0 327600.0 ;
      RECT  363300.0 341400.0 373500.0 355200.0 ;
      RECT  363300.0 369000.0 373500.0 355200.0 ;
      RECT  363300.0 369000.0 373500.0 382800.0 ;
      RECT  363300.0 396600.0 373500.0 382800.0 ;
      RECT  363300.0 396600.0 373500.0 410400.0 ;
      RECT  363300.0 424200.0 373500.0 410400.0 ;
      RECT  363300.0 424200.0 373500.0 438000.0 ;
      RECT  363300.0 451800.0 373500.0 438000.0 ;
      RECT  363300.0 451800.0 373500.0 465600.0 ;
      RECT  363300.0 479400.0 373500.0 465600.0 ;
      RECT  363300.0 479400.0 373500.0 493200.0 ;
      RECT  363300.0 507000.0 373500.0 493200.0 ;
      RECT  363300.0 507000.0 373500.0 520800.0 ;
      RECT  363300.0 534600.0 373500.0 520800.0 ;
      RECT  363300.0 534600.0 373500.0 548400.0 ;
      RECT  363300.0 562200.0 373500.0 548400.0 ;
      RECT  363300.0 562200.0 373500.0 576000.0 ;
      RECT  363300.0 589800.0 373500.0 576000.0 ;
      RECT  363300.0 589800.0 373500.0 603600.0 ;
      RECT  363300.0 617400.0 373500.0 603600.0 ;
      RECT  363300.0 617400.0 373500.0 631200.0 ;
      RECT  363300.0 645000.0 373500.0 631200.0 ;
      RECT  363300.0 645000.0 373500.0 658800.0 ;
      RECT  363300.0 672600.0 373500.0 658800.0 ;
      RECT  363300.0 672600.0 373500.0 686400.0 ;
      RECT  363300.0 700200.0 373500.0 686400.0 ;
      RECT  363300.0 700200.0 373500.0 714000.0 ;
      RECT  363300.0 727800.0 373500.0 714000.0 ;
      RECT  363300.0 727800.0 373500.0 741600.0 ;
      RECT  363300.0 755400.0 373500.0 741600.0 ;
      RECT  363300.0 755400.0 373500.0 769200.0 ;
      RECT  363300.0 783000.0 373500.0 769200.0 ;
      RECT  363300.0 783000.0 373500.0 796800.0 ;
      RECT  363300.0 810600.0 373500.0 796800.0 ;
      RECT  363300.0 810600.0 373500.0 824400.0 ;
      RECT  363300.0 838200.0 373500.0 824400.0 ;
      RECT  363300.0 838200.0 373500.0 852000.0 ;
      RECT  363300.0 865800.0 373500.0 852000.0 ;
      RECT  363300.0 865800.0 373500.0 879600.0 ;
      RECT  363300.0 893400.0 373500.0 879600.0 ;
      RECT  363300.0 893400.0 373500.0 907200.0 ;
      RECT  363300.0 921000.0 373500.0 907200.0 ;
      RECT  363300.0 921000.0 373500.0 934800.0 ;
      RECT  363300.0 948600.0 373500.0 934800.0 ;
      RECT  363300.0 948600.0 373500.0 962400.0 ;
      RECT  363300.0 976200.0 373500.0 962400.0 ;
      RECT  363300.0 976200.0 373500.0 990000.0 ;
      RECT  363300.0 1003800.0 373500.0 990000.0 ;
      RECT  363300.0 1003800.0 373500.0 1017600.0 ;
      RECT  363300.0 1031400.0 373500.0 1017600.0 ;
      RECT  363300.0 1031400.0 373500.0 1045200.0 ;
      RECT  363300.0 1059000.0 373500.0 1045200.0 ;
      RECT  363300.0 1059000.0 373500.0 1072800.0 ;
      RECT  363300.0 1086600.0 373500.0 1072800.0 ;
      RECT  363300.0 1086600.0 373500.0 1100400.0 ;
      RECT  363300.0 1114200.0 373500.0 1100400.0 ;
      RECT  363300.0 1114200.0 373500.0 1128000.0 ;
      RECT  363300.0 1141800.0 373500.0 1128000.0 ;
      RECT  363300.0 1141800.0 373500.0 1155600.0 ;
      RECT  363300.0 1169400.0 373500.0 1155600.0 ;
      RECT  363300.0 1169400.0 373500.0 1183200.0 ;
      RECT  363300.0 1197000.0 373500.0 1183200.0 ;
      RECT  373500.0 313800.0 383700.0 327600.0 ;
      RECT  373500.0 341400.0 383700.0 327600.0 ;
      RECT  373500.0 341400.0 383700.0 355200.0 ;
      RECT  373500.0 369000.0 383700.0 355200.0 ;
      RECT  373500.0 369000.0 383700.0 382800.0 ;
      RECT  373500.0 396600.0 383700.0 382800.0 ;
      RECT  373500.0 396600.0 383700.0 410400.0 ;
      RECT  373500.0 424200.0 383700.0 410400.0 ;
      RECT  373500.0 424200.0 383700.0 438000.0 ;
      RECT  373500.0 451800.0 383700.0 438000.0 ;
      RECT  373500.0 451800.0 383700.0 465600.0 ;
      RECT  373500.0 479400.0 383700.0 465600.0 ;
      RECT  373500.0 479400.0 383700.0 493200.0 ;
      RECT  373500.0 507000.0 383700.0 493200.0 ;
      RECT  373500.0 507000.0 383700.0 520800.0 ;
      RECT  373500.0 534600.0 383700.0 520800.0 ;
      RECT  373500.0 534600.0 383700.0 548400.0 ;
      RECT  373500.0 562200.0 383700.0 548400.0 ;
      RECT  373500.0 562200.0 383700.0 576000.0 ;
      RECT  373500.0 589800.0 383700.0 576000.0 ;
      RECT  373500.0 589800.0 383700.0 603600.0 ;
      RECT  373500.0 617400.0 383700.0 603600.0 ;
      RECT  373500.0 617400.0 383700.0 631200.0 ;
      RECT  373500.0 645000.0 383700.0 631200.0 ;
      RECT  373500.0 645000.0 383700.0 658800.0 ;
      RECT  373500.0 672600.0 383700.0 658800.0 ;
      RECT  373500.0 672600.0 383700.0 686400.0 ;
      RECT  373500.0 700200.0 383700.0 686400.0 ;
      RECT  373500.0 700200.0 383700.0 714000.0 ;
      RECT  373500.0 727800.0 383700.0 714000.0 ;
      RECT  373500.0 727800.0 383700.0 741600.0 ;
      RECT  373500.0 755400.0 383700.0 741600.0 ;
      RECT  373500.0 755400.0 383700.0 769200.0 ;
      RECT  373500.0 783000.0 383700.0 769200.0 ;
      RECT  373500.0 783000.0 383700.0 796800.0 ;
      RECT  373500.0 810600.0 383700.0 796800.0 ;
      RECT  373500.0 810600.0 383700.0 824400.0 ;
      RECT  373500.0 838200.0 383700.0 824400.0 ;
      RECT  373500.0 838200.0 383700.0 852000.0 ;
      RECT  373500.0 865800.0 383700.0 852000.0 ;
      RECT  373500.0 865800.0 383700.0 879600.0 ;
      RECT  373500.0 893400.0 383700.0 879600.0 ;
      RECT  373500.0 893400.0 383700.0 907200.0 ;
      RECT  373500.0 921000.0 383700.0 907200.0 ;
      RECT  373500.0 921000.0 383700.0 934800.0 ;
      RECT  373500.0 948600.0 383700.0 934800.0 ;
      RECT  373500.0 948600.0 383700.0 962400.0 ;
      RECT  373500.0 976200.0 383700.0 962400.0 ;
      RECT  373500.0 976200.0 383700.0 990000.0 ;
      RECT  373500.0 1003800.0 383700.0 990000.0 ;
      RECT  373500.0 1003800.0 383700.0 1017600.0 ;
      RECT  373500.0 1031400.0 383700.0 1017600.0 ;
      RECT  373500.0 1031400.0 383700.0 1045200.0 ;
      RECT  373500.0 1059000.0 383700.0 1045200.0 ;
      RECT  373500.0 1059000.0 383700.0 1072800.0 ;
      RECT  373500.0 1086600.0 383700.0 1072800.0 ;
      RECT  373500.0 1086600.0 383700.0 1100400.0 ;
      RECT  373500.0 1114200.0 383700.0 1100400.0 ;
      RECT  373500.0 1114200.0 383700.0 1128000.0 ;
      RECT  373500.0 1141800.0 383700.0 1128000.0 ;
      RECT  373500.0 1141800.0 383700.0 1155600.0 ;
      RECT  373500.0 1169400.0 383700.0 1155600.0 ;
      RECT  373500.0 1169400.0 383700.0 1183200.0 ;
      RECT  373500.0 1197000.0 383700.0 1183200.0 ;
      RECT  383700.0 313800.0 393900.0 327600.0 ;
      RECT  383700.0 341400.0 393900.0 327600.0 ;
      RECT  383700.0 341400.0 393900.0 355200.0 ;
      RECT  383700.0 369000.0 393900.0 355200.0 ;
      RECT  383700.0 369000.0 393900.0 382800.0 ;
      RECT  383700.0 396600.0 393900.0 382800.0 ;
      RECT  383700.0 396600.0 393900.0 410400.0 ;
      RECT  383700.0 424200.0 393900.0 410400.0 ;
      RECT  383700.0 424200.0 393900.0 438000.0 ;
      RECT  383700.0 451800.0 393900.0 438000.0 ;
      RECT  383700.0 451800.0 393900.0 465600.0 ;
      RECT  383700.0 479400.0 393900.0 465600.0 ;
      RECT  383700.0 479400.0 393900.0 493200.0 ;
      RECT  383700.0 507000.0 393900.0 493200.0 ;
      RECT  383700.0 507000.0 393900.0 520800.0 ;
      RECT  383700.0 534600.0 393900.0 520800.0 ;
      RECT  383700.0 534600.0 393900.0 548400.0 ;
      RECT  383700.0 562200.0 393900.0 548400.0 ;
      RECT  383700.0 562200.0 393900.0 576000.0 ;
      RECT  383700.0 589800.0 393900.0 576000.0 ;
      RECT  383700.0 589800.0 393900.0 603600.0 ;
      RECT  383700.0 617400.0 393900.0 603600.0 ;
      RECT  383700.0 617400.0 393900.0 631200.0 ;
      RECT  383700.0 645000.0 393900.0 631200.0 ;
      RECT  383700.0 645000.0 393900.0 658800.0 ;
      RECT  383700.0 672600.0 393900.0 658800.0 ;
      RECT  383700.0 672600.0 393900.0 686400.0 ;
      RECT  383700.0 700200.0 393900.0 686400.0 ;
      RECT  383700.0 700200.0 393900.0 714000.0 ;
      RECT  383700.0 727800.0 393900.0 714000.0 ;
      RECT  383700.0 727800.0 393900.0 741600.0 ;
      RECT  383700.0 755400.0 393900.0 741600.0 ;
      RECT  383700.0 755400.0 393900.0 769200.0 ;
      RECT  383700.0 783000.0 393900.0 769200.0 ;
      RECT  383700.0 783000.0 393900.0 796800.0 ;
      RECT  383700.0 810600.0 393900.0 796800.0 ;
      RECT  383700.0 810600.0 393900.0 824400.0 ;
      RECT  383700.0 838200.0 393900.0 824400.0 ;
      RECT  383700.0 838200.0 393900.0 852000.0 ;
      RECT  383700.0 865800.0 393900.0 852000.0 ;
      RECT  383700.0 865800.0 393900.0 879600.0 ;
      RECT  383700.0 893400.0 393900.0 879600.0 ;
      RECT  383700.0 893400.0 393900.0 907200.0 ;
      RECT  383700.0 921000.0 393900.0 907200.0 ;
      RECT  383700.0 921000.0 393900.0 934800.0 ;
      RECT  383700.0 948600.0 393900.0 934800.0 ;
      RECT  383700.0 948600.0 393900.0 962400.0 ;
      RECT  383700.0 976200.0 393900.0 962400.0 ;
      RECT  383700.0 976200.0 393900.0 990000.0 ;
      RECT  383700.0 1003800.0 393900.0 990000.0 ;
      RECT  383700.0 1003800.0 393900.0 1017600.0 ;
      RECT  383700.0 1031400.0 393900.0 1017600.0 ;
      RECT  383700.0 1031400.0 393900.0 1045200.0 ;
      RECT  383700.0 1059000.0 393900.0 1045200.0 ;
      RECT  383700.0 1059000.0 393900.0 1072800.0 ;
      RECT  383700.0 1086600.0 393900.0 1072800.0 ;
      RECT  383700.0 1086600.0 393900.0 1100400.0 ;
      RECT  383700.0 1114200.0 393900.0 1100400.0 ;
      RECT  383700.0 1114200.0 393900.0 1128000.0 ;
      RECT  383700.0 1141800.0 393900.0 1128000.0 ;
      RECT  383700.0 1141800.0 393900.0 1155600.0 ;
      RECT  383700.0 1169400.0 393900.0 1155600.0 ;
      RECT  383700.0 1169400.0 393900.0 1183200.0 ;
      RECT  383700.0 1197000.0 393900.0 1183200.0 ;
      RECT  393900.0 313800.0 404100.0 327600.0 ;
      RECT  393900.0 341400.0 404100.0 327600.0 ;
      RECT  393900.0 341400.0 404100.0 355200.0 ;
      RECT  393900.0 369000.0 404100.0 355200.0 ;
      RECT  393900.0 369000.0 404100.0 382800.0 ;
      RECT  393900.0 396600.0 404100.0 382800.0 ;
      RECT  393900.0 396600.0 404100.0 410400.0 ;
      RECT  393900.0 424200.0 404100.0 410400.0 ;
      RECT  393900.0 424200.0 404100.0 438000.0 ;
      RECT  393900.0 451800.0 404100.0 438000.0 ;
      RECT  393900.0 451800.0 404100.0 465600.0 ;
      RECT  393900.0 479400.0 404100.0 465600.0 ;
      RECT  393900.0 479400.0 404100.0 493200.0 ;
      RECT  393900.0 507000.0 404100.0 493200.0 ;
      RECT  393900.0 507000.0 404100.0 520800.0 ;
      RECT  393900.0 534600.0 404100.0 520800.0 ;
      RECT  393900.0 534600.0 404100.0 548400.0 ;
      RECT  393900.0 562200.0 404100.0 548400.0 ;
      RECT  393900.0 562200.0 404100.0 576000.0 ;
      RECT  393900.0 589800.0 404100.0 576000.0 ;
      RECT  393900.0 589800.0 404100.0 603600.0 ;
      RECT  393900.0 617400.0 404100.0 603600.0 ;
      RECT  393900.0 617400.0 404100.0 631200.0 ;
      RECT  393900.0 645000.0 404100.0 631200.0 ;
      RECT  393900.0 645000.0 404100.0 658800.0 ;
      RECT  393900.0 672600.0 404100.0 658800.0 ;
      RECT  393900.0 672600.0 404100.0 686400.0 ;
      RECT  393900.0 700200.0 404100.0 686400.0 ;
      RECT  393900.0 700200.0 404100.0 714000.0 ;
      RECT  393900.0 727800.0 404100.0 714000.0 ;
      RECT  393900.0 727800.0 404100.0 741600.0 ;
      RECT  393900.0 755400.0 404100.0 741600.0 ;
      RECT  393900.0 755400.0 404100.0 769200.0 ;
      RECT  393900.0 783000.0 404100.0 769200.0 ;
      RECT  393900.0 783000.0 404100.0 796800.0 ;
      RECT  393900.0 810600.0 404100.0 796800.0 ;
      RECT  393900.0 810600.0 404100.0 824400.0 ;
      RECT  393900.0 838200.0 404100.0 824400.0 ;
      RECT  393900.0 838200.0 404100.0 852000.0 ;
      RECT  393900.0 865800.0 404100.0 852000.0 ;
      RECT  393900.0 865800.0 404100.0 879600.0 ;
      RECT  393900.0 893400.0 404100.0 879600.0 ;
      RECT  393900.0 893400.0 404100.0 907200.0 ;
      RECT  393900.0 921000.0 404100.0 907200.0 ;
      RECT  393900.0 921000.0 404100.0 934800.0 ;
      RECT  393900.0 948600.0 404100.0 934800.0 ;
      RECT  393900.0 948600.0 404100.0 962400.0 ;
      RECT  393900.0 976200.0 404100.0 962400.0 ;
      RECT  393900.0 976200.0 404100.0 990000.0 ;
      RECT  393900.0 1003800.0 404100.0 990000.0 ;
      RECT  393900.0 1003800.0 404100.0 1017600.0 ;
      RECT  393900.0 1031400.0 404100.0 1017600.0 ;
      RECT  393900.0 1031400.0 404100.0 1045200.0 ;
      RECT  393900.0 1059000.0 404100.0 1045200.0 ;
      RECT  393900.0 1059000.0 404100.0 1072800.0 ;
      RECT  393900.0 1086600.0 404100.0 1072800.0 ;
      RECT  393900.0 1086600.0 404100.0 1100400.0 ;
      RECT  393900.0 1114200.0 404100.0 1100400.0 ;
      RECT  393900.0 1114200.0 404100.0 1128000.0 ;
      RECT  393900.0 1141800.0 404100.0 1128000.0 ;
      RECT  393900.0 1141800.0 404100.0 1155600.0 ;
      RECT  393900.0 1169400.0 404100.0 1155600.0 ;
      RECT  393900.0 1169400.0 404100.0 1183200.0 ;
      RECT  393900.0 1197000.0 404100.0 1183200.0 ;
      RECT  404100.0 313800.0 414300.0 327600.0 ;
      RECT  404100.0 341400.0 414300.0 327600.0 ;
      RECT  404100.0 341400.0 414300.0 355200.0 ;
      RECT  404100.0 369000.0 414300.0 355200.0 ;
      RECT  404100.0 369000.0 414300.0 382800.0 ;
      RECT  404100.0 396600.0 414300.0 382800.0 ;
      RECT  404100.0 396600.0 414300.0 410400.0 ;
      RECT  404100.0 424200.0 414300.0 410400.0 ;
      RECT  404100.0 424200.0 414300.0 438000.0 ;
      RECT  404100.0 451800.0 414300.0 438000.0 ;
      RECT  404100.0 451800.0 414300.0 465600.0 ;
      RECT  404100.0 479400.0 414300.0 465600.0 ;
      RECT  404100.0 479400.0 414300.0 493200.0 ;
      RECT  404100.0 507000.0 414300.0 493200.0 ;
      RECT  404100.0 507000.0 414300.0 520800.0 ;
      RECT  404100.0 534600.0 414300.0 520800.0 ;
      RECT  404100.0 534600.0 414300.0 548400.0 ;
      RECT  404100.0 562200.0 414300.0 548400.0 ;
      RECT  404100.0 562200.0 414300.0 576000.0 ;
      RECT  404100.0 589800.0 414300.0 576000.0 ;
      RECT  404100.0 589800.0 414300.0 603600.0 ;
      RECT  404100.0 617400.0 414300.0 603600.0 ;
      RECT  404100.0 617400.0 414300.0 631200.0 ;
      RECT  404100.0 645000.0 414300.0 631200.0 ;
      RECT  404100.0 645000.0 414300.0 658800.0 ;
      RECT  404100.0 672600.0 414300.0 658800.0 ;
      RECT  404100.0 672600.0 414300.0 686400.0 ;
      RECT  404100.0 700200.0 414300.0 686400.0 ;
      RECT  404100.0 700200.0 414300.0 714000.0 ;
      RECT  404100.0 727800.0 414300.0 714000.0 ;
      RECT  404100.0 727800.0 414300.0 741600.0 ;
      RECT  404100.0 755400.0 414300.0 741600.0 ;
      RECT  404100.0 755400.0 414300.0 769200.0 ;
      RECT  404100.0 783000.0 414300.0 769200.0 ;
      RECT  404100.0 783000.0 414300.0 796800.0 ;
      RECT  404100.0 810600.0 414300.0 796800.0 ;
      RECT  404100.0 810600.0 414300.0 824400.0 ;
      RECT  404100.0 838200.0 414300.0 824400.0 ;
      RECT  404100.0 838200.0 414300.0 852000.0 ;
      RECT  404100.0 865800.0 414300.0 852000.0 ;
      RECT  404100.0 865800.0 414300.0 879600.0 ;
      RECT  404100.0 893400.0 414300.0 879600.0 ;
      RECT  404100.0 893400.0 414300.0 907200.0 ;
      RECT  404100.0 921000.0 414300.0 907200.0 ;
      RECT  404100.0 921000.0 414300.0 934800.0 ;
      RECT  404100.0 948600.0 414300.0 934800.0 ;
      RECT  404100.0 948600.0 414300.0 962400.0 ;
      RECT  404100.0 976200.0 414300.0 962400.0 ;
      RECT  404100.0 976200.0 414300.0 990000.0 ;
      RECT  404100.0 1003800.0 414300.0 990000.0 ;
      RECT  404100.0 1003800.0 414300.0 1017600.0 ;
      RECT  404100.0 1031400.0 414300.0 1017600.0 ;
      RECT  404100.0 1031400.0 414300.0 1045200.0 ;
      RECT  404100.0 1059000.0 414300.0 1045200.0 ;
      RECT  404100.0 1059000.0 414300.0 1072800.0 ;
      RECT  404100.0 1086600.0 414300.0 1072800.0 ;
      RECT  404100.0 1086600.0 414300.0 1100400.0 ;
      RECT  404100.0 1114200.0 414300.0 1100400.0 ;
      RECT  404100.0 1114200.0 414300.0 1128000.0 ;
      RECT  404100.0 1141800.0 414300.0 1128000.0 ;
      RECT  404100.0 1141800.0 414300.0 1155600.0 ;
      RECT  404100.0 1169400.0 414300.0 1155600.0 ;
      RECT  404100.0 1169400.0 414300.0 1183200.0 ;
      RECT  404100.0 1197000.0 414300.0 1183200.0 ;
      RECT  414300.0 313800.0 424500.0 327600.0 ;
      RECT  414300.0 341400.0 424500.0 327600.0 ;
      RECT  414300.0 341400.0 424500.0 355200.0 ;
      RECT  414300.0 369000.0 424500.0 355200.0 ;
      RECT  414300.0 369000.0 424500.0 382800.0 ;
      RECT  414300.0 396600.0 424500.0 382800.0 ;
      RECT  414300.0 396600.0 424500.0 410400.0 ;
      RECT  414300.0 424200.0 424500.0 410400.0 ;
      RECT  414300.0 424200.0 424500.0 438000.0 ;
      RECT  414300.0 451800.0 424500.0 438000.0 ;
      RECT  414300.0 451800.0 424500.0 465600.0 ;
      RECT  414300.0 479400.0 424500.0 465600.0 ;
      RECT  414300.0 479400.0 424500.0 493200.0 ;
      RECT  414300.0 507000.0 424500.0 493200.0 ;
      RECT  414300.0 507000.0 424500.0 520800.0 ;
      RECT  414300.0 534600.0 424500.0 520800.0 ;
      RECT  414300.0 534600.0 424500.0 548400.0 ;
      RECT  414300.0 562200.0 424500.0 548400.0 ;
      RECT  414300.0 562200.0 424500.0 576000.0 ;
      RECT  414300.0 589800.0 424500.0 576000.0 ;
      RECT  414300.0 589800.0 424500.0 603600.0 ;
      RECT  414300.0 617400.0 424500.0 603600.0 ;
      RECT  414300.0 617400.0 424500.0 631200.0 ;
      RECT  414300.0 645000.0 424500.0 631200.0 ;
      RECT  414300.0 645000.0 424500.0 658800.0 ;
      RECT  414300.0 672600.0 424500.0 658800.0 ;
      RECT  414300.0 672600.0 424500.0 686400.0 ;
      RECT  414300.0 700200.0 424500.0 686400.0 ;
      RECT  414300.0 700200.0 424500.0 714000.0 ;
      RECT  414300.0 727800.0 424500.0 714000.0 ;
      RECT  414300.0 727800.0 424500.0 741600.0 ;
      RECT  414300.0 755400.0 424500.0 741600.0 ;
      RECT  414300.0 755400.0 424500.0 769200.0 ;
      RECT  414300.0 783000.0 424500.0 769200.0 ;
      RECT  414300.0 783000.0 424500.0 796800.0 ;
      RECT  414300.0 810600.0 424500.0 796800.0 ;
      RECT  414300.0 810600.0 424500.0 824400.0 ;
      RECT  414300.0 838200.0 424500.0 824400.0 ;
      RECT  414300.0 838200.0 424500.0 852000.0 ;
      RECT  414300.0 865800.0 424500.0 852000.0 ;
      RECT  414300.0 865800.0 424500.0 879600.0 ;
      RECT  414300.0 893400.0 424500.0 879600.0 ;
      RECT  414300.0 893400.0 424500.0 907200.0 ;
      RECT  414300.0 921000.0 424500.0 907200.0 ;
      RECT  414300.0 921000.0 424500.0 934800.0 ;
      RECT  414300.0 948600.0 424500.0 934800.0 ;
      RECT  414300.0 948600.0 424500.0 962400.0 ;
      RECT  414300.0 976200.0 424500.0 962400.0 ;
      RECT  414300.0 976200.0 424500.0 990000.0 ;
      RECT  414300.0 1003800.0 424500.0 990000.0 ;
      RECT  414300.0 1003800.0 424500.0 1017600.0 ;
      RECT  414300.0 1031400.0 424500.0 1017600.0 ;
      RECT  414300.0 1031400.0 424500.0 1045200.0 ;
      RECT  414300.0 1059000.0 424500.0 1045200.0 ;
      RECT  414300.0 1059000.0 424500.0 1072800.0 ;
      RECT  414300.0 1086600.0 424500.0 1072800.0 ;
      RECT  414300.0 1086600.0 424500.0 1100400.0 ;
      RECT  414300.0 1114200.0 424500.0 1100400.0 ;
      RECT  414300.0 1114200.0 424500.0 1128000.0 ;
      RECT  414300.0 1141800.0 424500.0 1128000.0 ;
      RECT  414300.0 1141800.0 424500.0 1155600.0 ;
      RECT  414300.0 1169400.0 424500.0 1155600.0 ;
      RECT  414300.0 1169400.0 424500.0 1183200.0 ;
      RECT  414300.0 1197000.0 424500.0 1183200.0 ;
      RECT  424500.0 313800.0 434700.0 327600.0 ;
      RECT  424500.0 341400.0 434700.0 327600.0 ;
      RECT  424500.0 341400.0 434700.0 355200.0 ;
      RECT  424500.0 369000.0 434700.0 355200.0 ;
      RECT  424500.0 369000.0 434700.0 382800.0 ;
      RECT  424500.0 396600.0 434700.0 382800.0 ;
      RECT  424500.0 396600.0 434700.0 410400.0 ;
      RECT  424500.0 424200.0 434700.0 410400.0 ;
      RECT  424500.0 424200.0 434700.0 438000.0 ;
      RECT  424500.0 451800.0 434700.0 438000.0 ;
      RECT  424500.0 451800.0 434700.0 465600.0 ;
      RECT  424500.0 479400.0 434700.0 465600.0 ;
      RECT  424500.0 479400.0 434700.0 493200.0 ;
      RECT  424500.0 507000.0 434700.0 493200.0 ;
      RECT  424500.0 507000.0 434700.0 520800.0 ;
      RECT  424500.0 534600.0 434700.0 520800.0 ;
      RECT  424500.0 534600.0 434700.0 548400.0 ;
      RECT  424500.0 562200.0 434700.0 548400.0 ;
      RECT  424500.0 562200.0 434700.0 576000.0 ;
      RECT  424500.0 589800.0 434700.0 576000.0 ;
      RECT  424500.0 589800.0 434700.0 603600.0 ;
      RECT  424500.0 617400.0 434700.0 603600.0 ;
      RECT  424500.0 617400.0 434700.0 631200.0 ;
      RECT  424500.0 645000.0 434700.0 631200.0 ;
      RECT  424500.0 645000.0 434700.0 658800.0 ;
      RECT  424500.0 672600.0 434700.0 658800.0 ;
      RECT  424500.0 672600.0 434700.0 686400.0 ;
      RECT  424500.0 700200.0 434700.0 686400.0 ;
      RECT  424500.0 700200.0 434700.0 714000.0 ;
      RECT  424500.0 727800.0 434700.0 714000.0 ;
      RECT  424500.0 727800.0 434700.0 741600.0 ;
      RECT  424500.0 755400.0 434700.0 741600.0 ;
      RECT  424500.0 755400.0 434700.0 769200.0 ;
      RECT  424500.0 783000.0 434700.0 769200.0 ;
      RECT  424500.0 783000.0 434700.0 796800.0 ;
      RECT  424500.0 810600.0 434700.0 796800.0 ;
      RECT  424500.0 810600.0 434700.0 824400.0 ;
      RECT  424500.0 838200.0 434700.0 824400.0 ;
      RECT  424500.0 838200.0 434700.0 852000.0 ;
      RECT  424500.0 865800.0 434700.0 852000.0 ;
      RECT  424500.0 865800.0 434700.0 879600.0 ;
      RECT  424500.0 893400.0 434700.0 879600.0 ;
      RECT  424500.0 893400.0 434700.0 907200.0 ;
      RECT  424500.0 921000.0 434700.0 907200.0 ;
      RECT  424500.0 921000.0 434700.0 934800.0 ;
      RECT  424500.0 948600.0 434700.0 934800.0 ;
      RECT  424500.0 948600.0 434700.0 962400.0 ;
      RECT  424500.0 976200.0 434700.0 962400.0 ;
      RECT  424500.0 976200.0 434700.0 990000.0 ;
      RECT  424500.0 1003800.0 434700.0 990000.0 ;
      RECT  424500.0 1003800.0 434700.0 1017600.0 ;
      RECT  424500.0 1031400.0 434700.0 1017600.0 ;
      RECT  424500.0 1031400.0 434700.0 1045200.0 ;
      RECT  424500.0 1059000.0 434700.0 1045200.0 ;
      RECT  424500.0 1059000.0 434700.0 1072800.0 ;
      RECT  424500.0 1086600.0 434700.0 1072800.0 ;
      RECT  424500.0 1086600.0 434700.0 1100400.0 ;
      RECT  424500.0 1114200.0 434700.0 1100400.0 ;
      RECT  424500.0 1114200.0 434700.0 1128000.0 ;
      RECT  424500.0 1141800.0 434700.0 1128000.0 ;
      RECT  424500.0 1141800.0 434700.0 1155600.0 ;
      RECT  424500.0 1169400.0 434700.0 1155600.0 ;
      RECT  424500.0 1169400.0 434700.0 1183200.0 ;
      RECT  424500.0 1197000.0 434700.0 1183200.0 ;
      RECT  434700.0 313800.0 444900.0 327600.0 ;
      RECT  434700.0 341400.0 444900.0 327600.0 ;
      RECT  434700.0 341400.0 444900.0 355200.0 ;
      RECT  434700.0 369000.0 444900.0 355200.0 ;
      RECT  434700.0 369000.0 444900.0 382800.0 ;
      RECT  434700.0 396600.0 444900.0 382800.0 ;
      RECT  434700.0 396600.0 444900.0 410400.0 ;
      RECT  434700.0 424200.0 444900.0 410400.0 ;
      RECT  434700.0 424200.0 444900.0 438000.0 ;
      RECT  434700.0 451800.0 444900.0 438000.0 ;
      RECT  434700.0 451800.0 444900.0 465600.0 ;
      RECT  434700.0 479400.0 444900.0 465600.0 ;
      RECT  434700.0 479400.0 444900.0 493200.0 ;
      RECT  434700.0 507000.0 444900.0 493200.0 ;
      RECT  434700.0 507000.0 444900.0 520800.0 ;
      RECT  434700.0 534600.0 444900.0 520800.0 ;
      RECT  434700.0 534600.0 444900.0 548400.0 ;
      RECT  434700.0 562200.0 444900.0 548400.0 ;
      RECT  434700.0 562200.0 444900.0 576000.0 ;
      RECT  434700.0 589800.0 444900.0 576000.0 ;
      RECT  434700.0 589800.0 444900.0 603600.0 ;
      RECT  434700.0 617400.0 444900.0 603600.0 ;
      RECT  434700.0 617400.0 444900.0 631200.0 ;
      RECT  434700.0 645000.0 444900.0 631200.0 ;
      RECT  434700.0 645000.0 444900.0 658800.0 ;
      RECT  434700.0 672600.0 444900.0 658800.0 ;
      RECT  434700.0 672600.0 444900.0 686400.0 ;
      RECT  434700.0 700200.0 444900.0 686400.0 ;
      RECT  434700.0 700200.0 444900.0 714000.0 ;
      RECT  434700.0 727800.0 444900.0 714000.0 ;
      RECT  434700.0 727800.0 444900.0 741600.0 ;
      RECT  434700.0 755400.0 444900.0 741600.0 ;
      RECT  434700.0 755400.0 444900.0 769200.0 ;
      RECT  434700.0 783000.0 444900.0 769200.0 ;
      RECT  434700.0 783000.0 444900.0 796800.0 ;
      RECT  434700.0 810600.0 444900.0 796800.0 ;
      RECT  434700.0 810600.0 444900.0 824400.0 ;
      RECT  434700.0 838200.0 444900.0 824400.0 ;
      RECT  434700.0 838200.0 444900.0 852000.0 ;
      RECT  434700.0 865800.0 444900.0 852000.0 ;
      RECT  434700.0 865800.0 444900.0 879600.0 ;
      RECT  434700.0 893400.0 444900.0 879600.0 ;
      RECT  434700.0 893400.0 444900.0 907200.0 ;
      RECT  434700.0 921000.0 444900.0 907200.0 ;
      RECT  434700.0 921000.0 444900.0 934800.0 ;
      RECT  434700.0 948600.0 444900.0 934800.0 ;
      RECT  434700.0 948600.0 444900.0 962400.0 ;
      RECT  434700.0 976200.0 444900.0 962400.0 ;
      RECT  434700.0 976200.0 444900.0 990000.0 ;
      RECT  434700.0 1003800.0 444900.0 990000.0 ;
      RECT  434700.0 1003800.0 444900.0 1017600.0 ;
      RECT  434700.0 1031400.0 444900.0 1017600.0 ;
      RECT  434700.0 1031400.0 444900.0 1045200.0 ;
      RECT  434700.0 1059000.0 444900.0 1045200.0 ;
      RECT  434700.0 1059000.0 444900.0 1072800.0 ;
      RECT  434700.0 1086600.0 444900.0 1072800.0 ;
      RECT  434700.0 1086600.0 444900.0 1100400.0 ;
      RECT  434700.0 1114200.0 444900.0 1100400.0 ;
      RECT  434700.0 1114200.0 444900.0 1128000.0 ;
      RECT  434700.0 1141800.0 444900.0 1128000.0 ;
      RECT  434700.0 1141800.0 444900.0 1155600.0 ;
      RECT  434700.0 1169400.0 444900.0 1155600.0 ;
      RECT  434700.0 1169400.0 444900.0 1183200.0 ;
      RECT  434700.0 1197000.0 444900.0 1183200.0 ;
      RECT  444900.0 313800.0 455100.0 327600.0 ;
      RECT  444900.0 341400.0 455100.0 327600.0 ;
      RECT  444900.0 341400.0 455100.0 355200.0 ;
      RECT  444900.0 369000.0 455100.0 355200.0 ;
      RECT  444900.0 369000.0 455100.0 382800.0 ;
      RECT  444900.0 396600.0 455100.0 382800.0 ;
      RECT  444900.0 396600.0 455100.0 410400.0 ;
      RECT  444900.0 424200.0 455100.0 410400.0 ;
      RECT  444900.0 424200.0 455100.0 438000.0 ;
      RECT  444900.0 451800.0 455100.0 438000.0 ;
      RECT  444900.0 451800.0 455100.0 465600.0 ;
      RECT  444900.0 479400.0 455100.0 465600.0 ;
      RECT  444900.0 479400.0 455100.0 493200.0 ;
      RECT  444900.0 507000.0 455100.0 493200.0 ;
      RECT  444900.0 507000.0 455100.0 520800.0 ;
      RECT  444900.0 534600.0 455100.0 520800.0 ;
      RECT  444900.0 534600.0 455100.0 548400.0 ;
      RECT  444900.0 562200.0 455100.0 548400.0 ;
      RECT  444900.0 562200.0 455100.0 576000.0 ;
      RECT  444900.0 589800.0 455100.0 576000.0 ;
      RECT  444900.0 589800.0 455100.0 603600.0 ;
      RECT  444900.0 617400.0 455100.0 603600.0 ;
      RECT  444900.0 617400.0 455100.0 631200.0 ;
      RECT  444900.0 645000.0 455100.0 631200.0 ;
      RECT  444900.0 645000.0 455100.0 658800.0 ;
      RECT  444900.0 672600.0 455100.0 658800.0 ;
      RECT  444900.0 672600.0 455100.0 686400.0 ;
      RECT  444900.0 700200.0 455100.0 686400.0 ;
      RECT  444900.0 700200.0 455100.0 714000.0 ;
      RECT  444900.0 727800.0 455100.0 714000.0 ;
      RECT  444900.0 727800.0 455100.0 741600.0 ;
      RECT  444900.0 755400.0 455100.0 741600.0 ;
      RECT  444900.0 755400.0 455100.0 769200.0 ;
      RECT  444900.0 783000.0 455100.0 769200.0 ;
      RECT  444900.0 783000.0 455100.0 796800.0 ;
      RECT  444900.0 810600.0 455100.0 796800.0 ;
      RECT  444900.0 810600.0 455100.0 824400.0 ;
      RECT  444900.0 838200.0 455100.0 824400.0 ;
      RECT  444900.0 838200.0 455100.0 852000.0 ;
      RECT  444900.0 865800.0 455100.0 852000.0 ;
      RECT  444900.0 865800.0 455100.0 879600.0 ;
      RECT  444900.0 893400.0 455100.0 879600.0 ;
      RECT  444900.0 893400.0 455100.0 907200.0 ;
      RECT  444900.0 921000.0 455100.0 907200.0 ;
      RECT  444900.0 921000.0 455100.0 934800.0 ;
      RECT  444900.0 948600.0 455100.0 934800.0 ;
      RECT  444900.0 948600.0 455100.0 962400.0 ;
      RECT  444900.0 976200.0 455100.0 962400.0 ;
      RECT  444900.0 976200.0 455100.0 990000.0 ;
      RECT  444900.0 1003800.0 455100.0 990000.0 ;
      RECT  444900.0 1003800.0 455100.0 1017600.0 ;
      RECT  444900.0 1031400.0 455100.0 1017600.0 ;
      RECT  444900.0 1031400.0 455100.0 1045200.0 ;
      RECT  444900.0 1059000.0 455100.0 1045200.0 ;
      RECT  444900.0 1059000.0 455100.0 1072800.0 ;
      RECT  444900.0 1086600.0 455100.0 1072800.0 ;
      RECT  444900.0 1086600.0 455100.0 1100400.0 ;
      RECT  444900.0 1114200.0 455100.0 1100400.0 ;
      RECT  444900.0 1114200.0 455100.0 1128000.0 ;
      RECT  444900.0 1141800.0 455100.0 1128000.0 ;
      RECT  444900.0 1141800.0 455100.0 1155600.0 ;
      RECT  444900.0 1169400.0 455100.0 1155600.0 ;
      RECT  444900.0 1169400.0 455100.0 1183200.0 ;
      RECT  444900.0 1197000.0 455100.0 1183200.0 ;
      RECT  455100.0 313800.0 465300.0 327600.0 ;
      RECT  455100.0 341400.0 465300.0 327600.0 ;
      RECT  455100.0 341400.0 465300.0 355200.0 ;
      RECT  455100.0 369000.0 465300.0 355200.0 ;
      RECT  455100.0 369000.0 465300.0 382800.0 ;
      RECT  455100.0 396600.0 465300.0 382800.0 ;
      RECT  455100.0 396600.0 465300.0 410400.0 ;
      RECT  455100.0 424200.0 465300.0 410400.0 ;
      RECT  455100.0 424200.0 465300.0 438000.0 ;
      RECT  455100.0 451800.0 465300.0 438000.0 ;
      RECT  455100.0 451800.0 465300.0 465600.0 ;
      RECT  455100.0 479400.0 465300.0 465600.0 ;
      RECT  455100.0 479400.0 465300.0 493200.0 ;
      RECT  455100.0 507000.0 465300.0 493200.0 ;
      RECT  455100.0 507000.0 465300.0 520800.0 ;
      RECT  455100.0 534600.0 465300.0 520800.0 ;
      RECT  455100.0 534600.0 465300.0 548400.0 ;
      RECT  455100.0 562200.0 465300.0 548400.0 ;
      RECT  455100.0 562200.0 465300.0 576000.0 ;
      RECT  455100.0 589800.0 465300.0 576000.0 ;
      RECT  455100.0 589800.0 465300.0 603600.0 ;
      RECT  455100.0 617400.0 465300.0 603600.0 ;
      RECT  455100.0 617400.0 465300.0 631200.0 ;
      RECT  455100.0 645000.0 465300.0 631200.0 ;
      RECT  455100.0 645000.0 465300.0 658800.0 ;
      RECT  455100.0 672600.0 465300.0 658800.0 ;
      RECT  455100.0 672600.0 465300.0 686400.0 ;
      RECT  455100.0 700200.0 465300.0 686400.0 ;
      RECT  455100.0 700200.0 465300.0 714000.0 ;
      RECT  455100.0 727800.0 465300.0 714000.0 ;
      RECT  455100.0 727800.0 465300.0 741600.0 ;
      RECT  455100.0 755400.0 465300.0 741600.0 ;
      RECT  455100.0 755400.0 465300.0 769200.0 ;
      RECT  455100.0 783000.0 465300.0 769200.0 ;
      RECT  455100.0 783000.0 465300.0 796800.0 ;
      RECT  455100.0 810600.0 465300.0 796800.0 ;
      RECT  455100.0 810600.0 465300.0 824400.0 ;
      RECT  455100.0 838200.0 465300.0 824400.0 ;
      RECT  455100.0 838200.0 465300.0 852000.0 ;
      RECT  455100.0 865800.0 465300.0 852000.0 ;
      RECT  455100.0 865800.0 465300.0 879600.0 ;
      RECT  455100.0 893400.0 465300.0 879600.0 ;
      RECT  455100.0 893400.0 465300.0 907200.0 ;
      RECT  455100.0 921000.0 465300.0 907200.0 ;
      RECT  455100.0 921000.0 465300.0 934800.0 ;
      RECT  455100.0 948600.0 465300.0 934800.0 ;
      RECT  455100.0 948600.0 465300.0 962400.0 ;
      RECT  455100.0 976200.0 465300.0 962400.0 ;
      RECT  455100.0 976200.0 465300.0 990000.0 ;
      RECT  455100.0 1003800.0 465300.0 990000.0 ;
      RECT  455100.0 1003800.0 465300.0 1017600.0 ;
      RECT  455100.0 1031400.0 465300.0 1017600.0 ;
      RECT  455100.0 1031400.0 465300.0 1045200.0 ;
      RECT  455100.0 1059000.0 465300.0 1045200.0 ;
      RECT  455100.0 1059000.0 465300.0 1072800.0 ;
      RECT  455100.0 1086600.0 465300.0 1072800.0 ;
      RECT  455100.0 1086600.0 465300.0 1100400.0 ;
      RECT  455100.0 1114200.0 465300.0 1100400.0 ;
      RECT  455100.0 1114200.0 465300.0 1128000.0 ;
      RECT  455100.0 1141800.0 465300.0 1128000.0 ;
      RECT  455100.0 1141800.0 465300.0 1155600.0 ;
      RECT  455100.0 1169400.0 465300.0 1155600.0 ;
      RECT  455100.0 1169400.0 465300.0 1183200.0 ;
      RECT  455100.0 1197000.0 465300.0 1183200.0 ;
      RECT  465300.0 313800.0 475500.0 327600.0 ;
      RECT  465300.0 341400.0 475500.0 327600.0 ;
      RECT  465300.0 341400.0 475500.0 355200.0 ;
      RECT  465300.0 369000.0 475500.0 355200.0 ;
      RECT  465300.0 369000.0 475500.0 382800.0 ;
      RECT  465300.0 396600.0 475500.0 382800.0 ;
      RECT  465300.0 396600.0 475500.0 410400.0 ;
      RECT  465300.0 424200.0 475500.0 410400.0 ;
      RECT  465300.0 424200.0 475500.0 438000.0 ;
      RECT  465300.0 451800.0 475500.0 438000.0 ;
      RECT  465300.0 451800.0 475500.0 465600.0 ;
      RECT  465300.0 479400.0 475500.0 465600.0 ;
      RECT  465300.0 479400.0 475500.0 493200.0 ;
      RECT  465300.0 507000.0 475500.0 493200.0 ;
      RECT  465300.0 507000.0 475500.0 520800.0 ;
      RECT  465300.0 534600.0 475500.0 520800.0 ;
      RECT  465300.0 534600.0 475500.0 548400.0 ;
      RECT  465300.0 562200.0 475500.0 548400.0 ;
      RECT  465300.0 562200.0 475500.0 576000.0 ;
      RECT  465300.0 589800.0 475500.0 576000.0 ;
      RECT  465300.0 589800.0 475500.0 603600.0 ;
      RECT  465300.0 617400.0 475500.0 603600.0 ;
      RECT  465300.0 617400.0 475500.0 631200.0 ;
      RECT  465300.0 645000.0 475500.0 631200.0 ;
      RECT  465300.0 645000.0 475500.0 658800.0 ;
      RECT  465300.0 672600.0 475500.0 658800.0 ;
      RECT  465300.0 672600.0 475500.0 686400.0 ;
      RECT  465300.0 700200.0 475500.0 686400.0 ;
      RECT  465300.0 700200.0 475500.0 714000.0 ;
      RECT  465300.0 727800.0 475500.0 714000.0 ;
      RECT  465300.0 727800.0 475500.0 741600.0 ;
      RECT  465300.0 755400.0 475500.0 741600.0 ;
      RECT  465300.0 755400.0 475500.0 769200.0 ;
      RECT  465300.0 783000.0 475500.0 769200.0 ;
      RECT  465300.0 783000.0 475500.0 796800.0 ;
      RECT  465300.0 810600.0 475500.0 796800.0 ;
      RECT  465300.0 810600.0 475500.0 824400.0 ;
      RECT  465300.0 838200.0 475500.0 824400.0 ;
      RECT  465300.0 838200.0 475500.0 852000.0 ;
      RECT  465300.0 865800.0 475500.0 852000.0 ;
      RECT  465300.0 865800.0 475500.0 879600.0 ;
      RECT  465300.0 893400.0 475500.0 879600.0 ;
      RECT  465300.0 893400.0 475500.0 907200.0 ;
      RECT  465300.0 921000.0 475500.0 907200.0 ;
      RECT  465300.0 921000.0 475500.0 934800.0 ;
      RECT  465300.0 948600.0 475500.0 934800.0 ;
      RECT  465300.0 948600.0 475500.0 962400.0 ;
      RECT  465300.0 976200.0 475500.0 962400.0 ;
      RECT  465300.0 976200.0 475500.0 990000.0 ;
      RECT  465300.0 1003800.0 475500.0 990000.0 ;
      RECT  465300.0 1003800.0 475500.0 1017600.0 ;
      RECT  465300.0 1031400.0 475500.0 1017600.0 ;
      RECT  465300.0 1031400.0 475500.0 1045200.0 ;
      RECT  465300.0 1059000.0 475500.0 1045200.0 ;
      RECT  465300.0 1059000.0 475500.0 1072800.0 ;
      RECT  465300.0 1086600.0 475500.0 1072800.0 ;
      RECT  465300.0 1086600.0 475500.0 1100400.0 ;
      RECT  465300.0 1114200.0 475500.0 1100400.0 ;
      RECT  465300.0 1114200.0 475500.0 1128000.0 ;
      RECT  465300.0 1141800.0 475500.0 1128000.0 ;
      RECT  465300.0 1141800.0 475500.0 1155600.0 ;
      RECT  465300.0 1169400.0 475500.0 1155600.0 ;
      RECT  465300.0 1169400.0 475500.0 1183200.0 ;
      RECT  465300.0 1197000.0 475500.0 1183200.0 ;
      RECT  475500.0 313800.0 485700.0 327600.0 ;
      RECT  475500.0 341400.0 485700.0 327600.0 ;
      RECT  475500.0 341400.0 485700.0 355200.0 ;
      RECT  475500.0 369000.0 485700.0 355200.0 ;
      RECT  475500.0 369000.0 485700.0 382800.0 ;
      RECT  475500.0 396600.0 485700.0 382800.0 ;
      RECT  475500.0 396600.0 485700.0 410400.0 ;
      RECT  475500.0 424200.0 485700.0 410400.0 ;
      RECT  475500.0 424200.0 485700.0 438000.0 ;
      RECT  475500.0 451800.0 485700.0 438000.0 ;
      RECT  475500.0 451800.0 485700.0 465600.0 ;
      RECT  475500.0 479400.0 485700.0 465600.0 ;
      RECT  475500.0 479400.0 485700.0 493200.0 ;
      RECT  475500.0 507000.0 485700.0 493200.0 ;
      RECT  475500.0 507000.0 485700.0 520800.0 ;
      RECT  475500.0 534600.0 485700.0 520800.0 ;
      RECT  475500.0 534600.0 485700.0 548400.0 ;
      RECT  475500.0 562200.0 485700.0 548400.0 ;
      RECT  475500.0 562200.0 485700.0 576000.0 ;
      RECT  475500.0 589800.0 485700.0 576000.0 ;
      RECT  475500.0 589800.0 485700.0 603600.0 ;
      RECT  475500.0 617400.0 485700.0 603600.0 ;
      RECT  475500.0 617400.0 485700.0 631200.0 ;
      RECT  475500.0 645000.0 485700.0 631200.0 ;
      RECT  475500.0 645000.0 485700.0 658800.0 ;
      RECT  475500.0 672600.0 485700.0 658800.0 ;
      RECT  475500.0 672600.0 485700.0 686400.0 ;
      RECT  475500.0 700200.0 485700.0 686400.0 ;
      RECT  475500.0 700200.0 485700.0 714000.0 ;
      RECT  475500.0 727800.0 485700.0 714000.0 ;
      RECT  475500.0 727800.0 485700.0 741600.0 ;
      RECT  475500.0 755400.0 485700.0 741600.0 ;
      RECT  475500.0 755400.0 485700.0 769200.0 ;
      RECT  475500.0 783000.0 485700.0 769200.0 ;
      RECT  475500.0 783000.0 485700.0 796800.0 ;
      RECT  475500.0 810600.0 485700.0 796800.0 ;
      RECT  475500.0 810600.0 485700.0 824400.0 ;
      RECT  475500.0 838200.0 485700.0 824400.0 ;
      RECT  475500.0 838200.0 485700.0 852000.0 ;
      RECT  475500.0 865800.0 485700.0 852000.0 ;
      RECT  475500.0 865800.0 485700.0 879600.0 ;
      RECT  475500.0 893400.0 485700.0 879600.0 ;
      RECT  475500.0 893400.0 485700.0 907200.0 ;
      RECT  475500.0 921000.0 485700.0 907200.0 ;
      RECT  475500.0 921000.0 485700.0 934800.0 ;
      RECT  475500.0 948600.0 485700.0 934800.0 ;
      RECT  475500.0 948600.0 485700.0 962400.0 ;
      RECT  475500.0 976200.0 485700.0 962400.0 ;
      RECT  475500.0 976200.0 485700.0 990000.0 ;
      RECT  475500.0 1003800.0 485700.0 990000.0 ;
      RECT  475500.0 1003800.0 485700.0 1017600.0 ;
      RECT  475500.0 1031400.0 485700.0 1017600.0 ;
      RECT  475500.0 1031400.0 485700.0 1045200.0 ;
      RECT  475500.0 1059000.0 485700.0 1045200.0 ;
      RECT  475500.0 1059000.0 485700.0 1072800.0 ;
      RECT  475500.0 1086600.0 485700.0 1072800.0 ;
      RECT  475500.0 1086600.0 485700.0 1100400.0 ;
      RECT  475500.0 1114200.0 485700.0 1100400.0 ;
      RECT  475500.0 1114200.0 485700.0 1128000.0 ;
      RECT  475500.0 1141800.0 485700.0 1128000.0 ;
      RECT  475500.0 1141800.0 485700.0 1155600.0 ;
      RECT  475500.0 1169400.0 485700.0 1155600.0 ;
      RECT  475500.0 1169400.0 485700.0 1183200.0 ;
      RECT  475500.0 1197000.0 485700.0 1183200.0 ;
      RECT  485700.0 313800.0 495900.0 327600.0 ;
      RECT  485700.0 341400.0 495900.0 327600.0 ;
      RECT  485700.0 341400.0 495900.0 355200.0 ;
      RECT  485700.0 369000.0 495900.0 355200.0 ;
      RECT  485700.0 369000.0 495900.0 382800.0 ;
      RECT  485700.0 396600.0 495900.0 382800.0 ;
      RECT  485700.0 396600.0 495900.0 410400.0 ;
      RECT  485700.0 424200.0 495900.0 410400.0 ;
      RECT  485700.0 424200.0 495900.0 438000.0 ;
      RECT  485700.0 451800.0 495900.0 438000.0 ;
      RECT  485700.0 451800.0 495900.0 465600.0 ;
      RECT  485700.0 479400.0 495900.0 465600.0 ;
      RECT  485700.0 479400.0 495900.0 493200.0 ;
      RECT  485700.0 507000.0 495900.0 493200.0 ;
      RECT  485700.0 507000.0 495900.0 520800.0 ;
      RECT  485700.0 534600.0 495900.0 520800.0 ;
      RECT  485700.0 534600.0 495900.0 548400.0 ;
      RECT  485700.0 562200.0 495900.0 548400.0 ;
      RECT  485700.0 562200.0 495900.0 576000.0 ;
      RECT  485700.0 589800.0 495900.0 576000.0 ;
      RECT  485700.0 589800.0 495900.0 603600.0 ;
      RECT  485700.0 617400.0 495900.0 603600.0 ;
      RECT  485700.0 617400.0 495900.0 631200.0 ;
      RECT  485700.0 645000.0 495900.0 631200.0 ;
      RECT  485700.0 645000.0 495900.0 658800.0 ;
      RECT  485700.0 672600.0 495900.0 658800.0 ;
      RECT  485700.0 672600.0 495900.0 686400.0 ;
      RECT  485700.0 700200.0 495900.0 686400.0 ;
      RECT  485700.0 700200.0 495900.0 714000.0 ;
      RECT  485700.0 727800.0 495900.0 714000.0 ;
      RECT  485700.0 727800.0 495900.0 741600.0 ;
      RECT  485700.0 755400.0 495900.0 741600.0 ;
      RECT  485700.0 755400.0 495900.0 769200.0 ;
      RECT  485700.0 783000.0 495900.0 769200.0 ;
      RECT  485700.0 783000.0 495900.0 796800.0 ;
      RECT  485700.0 810600.0 495900.0 796800.0 ;
      RECT  485700.0 810600.0 495900.0 824400.0 ;
      RECT  485700.0 838200.0 495900.0 824400.0 ;
      RECT  485700.0 838200.0 495900.0 852000.0 ;
      RECT  485700.0 865800.0 495900.0 852000.0 ;
      RECT  485700.0 865800.0 495900.0 879600.0 ;
      RECT  485700.0 893400.0 495900.0 879600.0 ;
      RECT  485700.0 893400.0 495900.0 907200.0 ;
      RECT  485700.0 921000.0 495900.0 907200.0 ;
      RECT  485700.0 921000.0 495900.0 934800.0 ;
      RECT  485700.0 948600.0 495900.0 934800.0 ;
      RECT  485700.0 948600.0 495900.0 962400.0 ;
      RECT  485700.0 976200.0 495900.0 962400.0 ;
      RECT  485700.0 976200.0 495900.0 990000.0 ;
      RECT  485700.0 1003800.0 495900.0 990000.0 ;
      RECT  485700.0 1003800.0 495900.0 1017600.0 ;
      RECT  485700.0 1031400.0 495900.0 1017600.0 ;
      RECT  485700.0 1031400.0 495900.0 1045200.0 ;
      RECT  485700.0 1059000.0 495900.0 1045200.0 ;
      RECT  485700.0 1059000.0 495900.0 1072800.0 ;
      RECT  485700.0 1086600.0 495900.0 1072800.0 ;
      RECT  485700.0 1086600.0 495900.0 1100400.0 ;
      RECT  485700.0 1114200.0 495900.0 1100400.0 ;
      RECT  485700.0 1114200.0 495900.0 1128000.0 ;
      RECT  485700.0 1141800.0 495900.0 1128000.0 ;
      RECT  485700.0 1141800.0 495900.0 1155600.0 ;
      RECT  485700.0 1169400.0 495900.0 1155600.0 ;
      RECT  485700.0 1169400.0 495900.0 1183200.0 ;
      RECT  485700.0 1197000.0 495900.0 1183200.0 ;
      RECT  495900.0 313800.0 506100.0 327600.0 ;
      RECT  495900.0 341400.0 506100.0 327600.0 ;
      RECT  495900.0 341400.0 506100.0 355200.0 ;
      RECT  495900.0 369000.0 506100.0 355200.0 ;
      RECT  495900.0 369000.0 506100.0 382800.0 ;
      RECT  495900.0 396600.0 506100.0 382800.0 ;
      RECT  495900.0 396600.0 506100.0 410400.0 ;
      RECT  495900.0 424200.0 506100.0 410400.0 ;
      RECT  495900.0 424200.0 506100.0 438000.0 ;
      RECT  495900.0 451800.0 506100.0 438000.0 ;
      RECT  495900.0 451800.0 506100.0 465600.0 ;
      RECT  495900.0 479400.0 506100.0 465600.0 ;
      RECT  495900.0 479400.0 506100.0 493200.0 ;
      RECT  495900.0 507000.0 506100.0 493200.0 ;
      RECT  495900.0 507000.0 506100.0 520800.0 ;
      RECT  495900.0 534600.0 506100.0 520800.0 ;
      RECT  495900.0 534600.0 506100.0 548400.0 ;
      RECT  495900.0 562200.0 506100.0 548400.0 ;
      RECT  495900.0 562200.0 506100.0 576000.0 ;
      RECT  495900.0 589800.0 506100.0 576000.0 ;
      RECT  495900.0 589800.0 506100.0 603600.0 ;
      RECT  495900.0 617400.0 506100.0 603600.0 ;
      RECT  495900.0 617400.0 506100.0 631200.0 ;
      RECT  495900.0 645000.0 506100.0 631200.0 ;
      RECT  495900.0 645000.0 506100.0 658800.0 ;
      RECT  495900.0 672600.0 506100.0 658800.0 ;
      RECT  495900.0 672600.0 506100.0 686400.0 ;
      RECT  495900.0 700200.0 506100.0 686400.0 ;
      RECT  495900.0 700200.0 506100.0 714000.0 ;
      RECT  495900.0 727800.0 506100.0 714000.0 ;
      RECT  495900.0 727800.0 506100.0 741600.0 ;
      RECT  495900.0 755400.0 506100.0 741600.0 ;
      RECT  495900.0 755400.0 506100.0 769200.0 ;
      RECT  495900.0 783000.0 506100.0 769200.0 ;
      RECT  495900.0 783000.0 506100.0 796800.0 ;
      RECT  495900.0 810600.0 506100.0 796800.0 ;
      RECT  495900.0 810600.0 506100.0 824400.0 ;
      RECT  495900.0 838200.0 506100.0 824400.0 ;
      RECT  495900.0 838200.0 506100.0 852000.0 ;
      RECT  495900.0 865800.0 506100.0 852000.0 ;
      RECT  495900.0 865800.0 506100.0 879600.0 ;
      RECT  495900.0 893400.0 506100.0 879600.0 ;
      RECT  495900.0 893400.0 506100.0 907200.0 ;
      RECT  495900.0 921000.0 506100.0 907200.0 ;
      RECT  495900.0 921000.0 506100.0 934800.0 ;
      RECT  495900.0 948600.0 506100.0 934800.0 ;
      RECT  495900.0 948600.0 506100.0 962400.0 ;
      RECT  495900.0 976200.0 506100.0 962400.0 ;
      RECT  495900.0 976200.0 506100.0 990000.0 ;
      RECT  495900.0 1003800.0 506100.0 990000.0 ;
      RECT  495900.0 1003800.0 506100.0 1017600.0 ;
      RECT  495900.0 1031400.0 506100.0 1017600.0 ;
      RECT  495900.0 1031400.0 506100.0 1045200.0 ;
      RECT  495900.0 1059000.0 506100.0 1045200.0 ;
      RECT  495900.0 1059000.0 506100.0 1072800.0 ;
      RECT  495900.0 1086600.0 506100.0 1072800.0 ;
      RECT  495900.0 1086600.0 506100.0 1100400.0 ;
      RECT  495900.0 1114200.0 506100.0 1100400.0 ;
      RECT  495900.0 1114200.0 506100.0 1128000.0 ;
      RECT  495900.0 1141800.0 506100.0 1128000.0 ;
      RECT  495900.0 1141800.0 506100.0 1155600.0 ;
      RECT  495900.0 1169400.0 506100.0 1155600.0 ;
      RECT  495900.0 1169400.0 506100.0 1183200.0 ;
      RECT  495900.0 1197000.0 506100.0 1183200.0 ;
      RECT  506100.0 313800.0 516300.0 327600.0 ;
      RECT  506100.0 341400.0 516300.0 327600.0 ;
      RECT  506100.0 341400.0 516300.0 355200.0 ;
      RECT  506100.0 369000.0 516300.0 355200.0 ;
      RECT  506100.0 369000.0 516300.0 382800.0 ;
      RECT  506100.0 396600.0 516300.0 382800.0 ;
      RECT  506100.0 396600.0 516300.0 410400.0 ;
      RECT  506100.0 424200.0 516300.0 410400.0 ;
      RECT  506100.0 424200.0 516300.0 438000.0 ;
      RECT  506100.0 451800.0 516300.0 438000.0 ;
      RECT  506100.0 451800.0 516300.0 465600.0 ;
      RECT  506100.0 479400.0 516300.0 465600.0 ;
      RECT  506100.0 479400.0 516300.0 493200.0 ;
      RECT  506100.0 507000.0 516300.0 493200.0 ;
      RECT  506100.0 507000.0 516300.0 520800.0 ;
      RECT  506100.0 534600.0 516300.0 520800.0 ;
      RECT  506100.0 534600.0 516300.0 548400.0 ;
      RECT  506100.0 562200.0 516300.0 548400.0 ;
      RECT  506100.0 562200.0 516300.0 576000.0 ;
      RECT  506100.0 589800.0 516300.0 576000.0 ;
      RECT  506100.0 589800.0 516300.0 603600.0 ;
      RECT  506100.0 617400.0 516300.0 603600.0 ;
      RECT  506100.0 617400.0 516300.0 631200.0 ;
      RECT  506100.0 645000.0 516300.0 631200.0 ;
      RECT  506100.0 645000.0 516300.0 658800.0 ;
      RECT  506100.0 672600.0 516300.0 658800.0 ;
      RECT  506100.0 672600.0 516300.0 686400.0 ;
      RECT  506100.0 700200.0 516300.0 686400.0 ;
      RECT  506100.0 700200.0 516300.0 714000.0 ;
      RECT  506100.0 727800.0 516300.0 714000.0 ;
      RECT  506100.0 727800.0 516300.0 741600.0 ;
      RECT  506100.0 755400.0 516300.0 741600.0 ;
      RECT  506100.0 755400.0 516300.0 769200.0 ;
      RECT  506100.0 783000.0 516300.0 769200.0 ;
      RECT  506100.0 783000.0 516300.0 796800.0 ;
      RECT  506100.0 810600.0 516300.0 796800.0 ;
      RECT  506100.0 810600.0 516300.0 824400.0 ;
      RECT  506100.0 838200.0 516300.0 824400.0 ;
      RECT  506100.0 838200.0 516300.0 852000.0 ;
      RECT  506100.0 865800.0 516300.0 852000.0 ;
      RECT  506100.0 865800.0 516300.0 879600.0 ;
      RECT  506100.0 893400.0 516300.0 879600.0 ;
      RECT  506100.0 893400.0 516300.0 907200.0 ;
      RECT  506100.0 921000.0 516300.0 907200.0 ;
      RECT  506100.0 921000.0 516300.0 934800.0 ;
      RECT  506100.0 948600.0 516300.0 934800.0 ;
      RECT  506100.0 948600.0 516300.0 962400.0 ;
      RECT  506100.0 976200.0 516300.0 962400.0 ;
      RECT  506100.0 976200.0 516300.0 990000.0 ;
      RECT  506100.0 1003800.0 516300.0 990000.0 ;
      RECT  506100.0 1003800.0 516300.0 1017600.0 ;
      RECT  506100.0 1031400.0 516300.0 1017600.0 ;
      RECT  506100.0 1031400.0 516300.0 1045200.0 ;
      RECT  506100.0 1059000.0 516300.0 1045200.0 ;
      RECT  506100.0 1059000.0 516300.0 1072800.0 ;
      RECT  506100.0 1086600.0 516300.0 1072800.0 ;
      RECT  506100.0 1086600.0 516300.0 1100400.0 ;
      RECT  506100.0 1114200.0 516300.0 1100400.0 ;
      RECT  506100.0 1114200.0 516300.0 1128000.0 ;
      RECT  506100.0 1141800.0 516300.0 1128000.0 ;
      RECT  506100.0 1141800.0 516300.0 1155600.0 ;
      RECT  506100.0 1169400.0 516300.0 1155600.0 ;
      RECT  506100.0 1169400.0 516300.0 1183200.0 ;
      RECT  506100.0 1197000.0 516300.0 1183200.0 ;
      RECT  516300.0 313800.0 526500.0 327600.0 ;
      RECT  516300.0 341400.0 526500.0 327600.0 ;
      RECT  516300.0 341400.0 526500.0 355200.0 ;
      RECT  516300.0 369000.0 526500.0 355200.0 ;
      RECT  516300.0 369000.0 526500.0 382800.0 ;
      RECT  516300.0 396600.0 526500.0 382800.0 ;
      RECT  516300.0 396600.0 526500.0 410400.0 ;
      RECT  516300.0 424200.0 526500.0 410400.0 ;
      RECT  516300.0 424200.0 526500.0 438000.0 ;
      RECT  516300.0 451800.0 526500.0 438000.0 ;
      RECT  516300.0 451800.0 526500.0 465600.0 ;
      RECT  516300.0 479400.0 526500.0 465600.0 ;
      RECT  516300.0 479400.0 526500.0 493200.0 ;
      RECT  516300.0 507000.0 526500.0 493200.0 ;
      RECT  516300.0 507000.0 526500.0 520800.0 ;
      RECT  516300.0 534600.0 526500.0 520800.0 ;
      RECT  516300.0 534600.0 526500.0 548400.0 ;
      RECT  516300.0 562200.0 526500.0 548400.0 ;
      RECT  516300.0 562200.0 526500.0 576000.0 ;
      RECT  516300.0 589800.0 526500.0 576000.0 ;
      RECT  516300.0 589800.0 526500.0 603600.0 ;
      RECT  516300.0 617400.0 526500.0 603600.0 ;
      RECT  516300.0 617400.0 526500.0 631200.0 ;
      RECT  516300.0 645000.0 526500.0 631200.0 ;
      RECT  516300.0 645000.0 526500.0 658800.0 ;
      RECT  516300.0 672600.0 526500.0 658800.0 ;
      RECT  516300.0 672600.0 526500.0 686400.0 ;
      RECT  516300.0 700200.0 526500.0 686400.0 ;
      RECT  516300.0 700200.0 526500.0 714000.0 ;
      RECT  516300.0 727800.0 526500.0 714000.0 ;
      RECT  516300.0 727800.0 526500.0 741600.0 ;
      RECT  516300.0 755400.0 526500.0 741600.0 ;
      RECT  516300.0 755400.0 526500.0 769200.0 ;
      RECT  516300.0 783000.0 526500.0 769200.0 ;
      RECT  516300.0 783000.0 526500.0 796800.0 ;
      RECT  516300.0 810600.0 526500.0 796800.0 ;
      RECT  516300.0 810600.0 526500.0 824400.0 ;
      RECT  516300.0 838200.0 526500.0 824400.0 ;
      RECT  516300.0 838200.0 526500.0 852000.0 ;
      RECT  516300.0 865800.0 526500.0 852000.0 ;
      RECT  516300.0 865800.0 526500.0 879600.0 ;
      RECT  516300.0 893400.0 526500.0 879600.0 ;
      RECT  516300.0 893400.0 526500.0 907200.0 ;
      RECT  516300.0 921000.0 526500.0 907200.0 ;
      RECT  516300.0 921000.0 526500.0 934800.0 ;
      RECT  516300.0 948600.0 526500.0 934800.0 ;
      RECT  516300.0 948600.0 526500.0 962400.0 ;
      RECT  516300.0 976200.0 526500.0 962400.0 ;
      RECT  516300.0 976200.0 526500.0 990000.0 ;
      RECT  516300.0 1003800.0 526500.0 990000.0 ;
      RECT  516300.0 1003800.0 526500.0 1017600.0 ;
      RECT  516300.0 1031400.0 526500.0 1017600.0 ;
      RECT  516300.0 1031400.0 526500.0 1045200.0 ;
      RECT  516300.0 1059000.0 526500.0 1045200.0 ;
      RECT  516300.0 1059000.0 526500.0 1072800.0 ;
      RECT  516300.0 1086600.0 526500.0 1072800.0 ;
      RECT  516300.0 1086600.0 526500.0 1100400.0 ;
      RECT  516300.0 1114200.0 526500.0 1100400.0 ;
      RECT  516300.0 1114200.0 526500.0 1128000.0 ;
      RECT  516300.0 1141800.0 526500.0 1128000.0 ;
      RECT  516300.0 1141800.0 526500.0 1155600.0 ;
      RECT  516300.0 1169400.0 526500.0 1155600.0 ;
      RECT  516300.0 1169400.0 526500.0 1183200.0 ;
      RECT  516300.0 1197000.0 526500.0 1183200.0 ;
      RECT  199500.0 315300.0 527100.0 316500.0 ;
      RECT  199500.0 338700.0 527100.0 339900.0 ;
      RECT  199500.0 342900.0 527100.0 344100.0 ;
      RECT  199500.0 366300.0 527100.0 367500.0 ;
      RECT  199500.0 370500.0 527100.0 371700.0 ;
      RECT  199500.0 393900.0 527100.0 395100.0 ;
      RECT  199500.0 398100.0 527100.0 399300.0 ;
      RECT  199500.0 421500.0 527100.0 422700.0 ;
      RECT  199500.0 425700.0 527100.0 426900.0 ;
      RECT  199500.0 449100.0 527100.0 450300.0 ;
      RECT  199500.0 453300.0 527100.0 454500.0 ;
      RECT  199500.0 476700.0 527100.0 477900.0 ;
      RECT  199500.0 480900.0 527100.0 482100.0 ;
      RECT  199500.0 504300.0 527100.0 505500.0 ;
      RECT  199500.0 508500.0 527100.0 509700.0 ;
      RECT  199500.0 531900.0 527100.0 533100.0 ;
      RECT  199500.0 536100.0 527100.0 537300.0 ;
      RECT  199500.0 559500.0 527100.0 560700.0 ;
      RECT  199500.0 563700.0 527100.0 564900.0 ;
      RECT  199500.0 587100.0 527100.0 588300.0 ;
      RECT  199500.0 591300.0 527100.0 592500.0 ;
      RECT  199500.0 614700.0 527100.0 615900.0 ;
      RECT  199500.0 618900.0 527100.0 620100.0 ;
      RECT  199500.0 642300.0 527100.0 643500.0 ;
      RECT  199500.0 646500.0 527100.0 647700.0 ;
      RECT  199500.0 669900.0 527100.0 671100.0 ;
      RECT  199500.0 674100.0 527100.0 675300.0 ;
      RECT  199500.0 697500.0 527100.0 698700.0 ;
      RECT  199500.0 701700.0 527100.0 702900.0 ;
      RECT  199500.0 725100.0 527100.0 726300.0 ;
      RECT  199500.0 729300.0 527100.0 730500.0 ;
      RECT  199500.0 752700.0 527100.0 753900.0 ;
      RECT  199500.0 756900.0 527100.0 758100.0 ;
      RECT  199500.0 780300.0 527100.0 781500.0 ;
      RECT  199500.0 784500.0 527100.0 785700.0 ;
      RECT  199500.0 807900.0 527100.0 809100.0 ;
      RECT  199500.0 812100.0 527100.0 813300.0 ;
      RECT  199500.0 835500.0 527100.0 836700.0 ;
      RECT  199500.0 839700.0 527100.0 840900.0 ;
      RECT  199500.0 863100.0 527100.0 864300.0 ;
      RECT  199500.0 867300.0 527100.0 868500.0 ;
      RECT  199500.0 890700.0 527100.0 891900.0 ;
      RECT  199500.0 894900.0 527100.0 896100.0 ;
      RECT  199500.0 918300.0 527100.0 919500.0 ;
      RECT  199500.0 922500.0 527100.0 923700.0 ;
      RECT  199500.0 945900.0 527100.0 947100.0 ;
      RECT  199500.0 950100.0 527100.0 951300.0 ;
      RECT  199500.0 973500.0 527100.0 974700.0 ;
      RECT  199500.0 977700.0 527100.0 978900.0 ;
      RECT  199500.0 1001100.0 527100.0 1002300.0 ;
      RECT  199500.0 1005300.0 527100.0 1006500.0 ;
      RECT  199500.0 1028700.0 527100.0 1029900.0 ;
      RECT  199500.0 1032900.0 527100.0 1034100.0 ;
      RECT  199500.0 1056300.0 527100.0 1057500.0 ;
      RECT  199500.0 1060500.0 527100.0 1061700.0 ;
      RECT  199500.0 1083900.0 527100.0 1085100.0 ;
      RECT  199500.0 1088100.0 527100.0 1089300.0 ;
      RECT  199500.0 1111500.0 527100.0 1112700.0 ;
      RECT  199500.0 1115700.0 527100.0 1116900.0 ;
      RECT  199500.0 1139100.0 527100.0 1140300.0 ;
      RECT  199500.0 1143300.0 527100.0 1144500.0 ;
      RECT  199500.0 1166700.0 527100.0 1167900.0 ;
      RECT  199500.0 1170900.0 527100.0 1172100.0 ;
      RECT  199500.0 1194300.0 527100.0 1195500.0 ;
      RECT  199500.0 327000.0 527100.0 327900.0 ;
      RECT  199500.0 354600.0 527100.0 355500.0 ;
      RECT  199500.0 382200.0 527100.0 383100.0 ;
      RECT  199500.0 409800.0 527100.0 410700.0 ;
      RECT  199500.0 437400.0 527100.0 438300.0 ;
      RECT  199500.0 465000.0 527100.0 465900.0 ;
      RECT  199500.0 492600.0 527100.0 493500.0 ;
      RECT  199500.0 520200.0 527100.0 521100.0 ;
      RECT  199500.0 547800.0 527100.0 548700.0 ;
      RECT  199500.0 575400.0 527100.0 576300.0 ;
      RECT  199500.0 603000.0 527100.0 603900.0 ;
      RECT  199500.0 630600.0 527100.0 631500.0 ;
      RECT  199500.0 658200.0 527100.0 659100.0 ;
      RECT  199500.0 685800.0 527100.0 686700.0 ;
      RECT  199500.0 713400.0 527100.0 714300.0 ;
      RECT  199500.0 741000.0 527100.0 741900.0 ;
      RECT  199500.0 768600.0 527100.0 769500.0 ;
      RECT  199500.0 796200.0 527100.0 797100.0 ;
      RECT  199500.0 823800.0 527100.0 824700.0 ;
      RECT  199500.0 851400.0 527100.0 852300.0 ;
      RECT  199500.0 879000.0 527100.0 879900.0 ;
      RECT  199500.0 906600.0 527100.0 907500.0 ;
      RECT  199500.0 934200.0 527100.0 935100.0 ;
      RECT  199500.0 961800.0 527100.0 962700.0 ;
      RECT  199500.0 989400.0 527100.0 990300.0 ;
      RECT  199500.0 1017000.0 527100.0 1017900.0 ;
      RECT  199500.0 1044600.0 527100.0 1045500.0 ;
      RECT  199500.0 1072200.0 527100.0 1073100.0 ;
      RECT  199500.0 1099800.0 527100.0 1100700.0 ;
      RECT  199500.0 1127400.0 527100.0 1128300.0 ;
      RECT  199500.0 1155000.0 527100.0 1155900.0 ;
      RECT  199500.0 1182600.0 527100.0 1183500.0 ;
      RECT  205500.0 1210200.0 206700.0 1217400.0 ;
      RECT  203100.0 1203000.0 204300.0 1204200.0 ;
      RECT  205500.0 1203000.0 206700.0 1204200.0 ;
      RECT  205500.0 1203000.0 206700.0 1204200.0 ;
      RECT  203100.0 1203000.0 204300.0 1204200.0 ;
      RECT  203100.0 1210200.0 204300.0 1211400.0 ;
      RECT  205500.0 1210200.0 206700.0 1211400.0 ;
      RECT  205500.0 1210200.0 206700.0 1211400.0 ;
      RECT  203100.0 1210200.0 204300.0 1211400.0 ;
      RECT  205500.0 1210200.0 206700.0 1211400.0 ;
      RECT  207900.0 1210200.0 209100.0 1211400.0 ;
      RECT  207900.0 1210200.0 209100.0 1211400.0 ;
      RECT  205500.0 1210200.0 206700.0 1211400.0 ;
      RECT  205200.0 1205250.0 204000.0 1206450.0 ;
      RECT  205500.0 1215600.0 206700.0 1216800.0 ;
      RECT  203100.0 1203000.0 204300.0 1204200.0 ;
      RECT  205500.0 1203000.0 206700.0 1204200.0 ;
      RECT  203100.0 1210200.0 204300.0 1211400.0 ;
      RECT  207900.0 1210200.0 209100.0 1211400.0 ;
      RECT  200100.0 1205400.0 210300.0 1206300.0 ;
      RECT  200100.0 1216500.0 210300.0 1217400.0 ;
      RECT  215700.0 1210200.0 216900.0 1217400.0 ;
      RECT  213300.0 1203000.0 214500.0 1204200.0 ;
      RECT  215700.0 1203000.0 216900.0 1204200.0 ;
      RECT  215700.0 1203000.0 216900.0 1204200.0 ;
      RECT  213300.0 1203000.0 214500.0 1204200.0 ;
      RECT  213300.0 1210200.0 214500.0 1211400.0 ;
      RECT  215700.0 1210200.0 216900.0 1211400.0 ;
      RECT  215700.0 1210200.0 216900.0 1211400.0 ;
      RECT  213300.0 1210200.0 214500.0 1211400.0 ;
      RECT  215700.0 1210200.0 216900.0 1211400.0 ;
      RECT  218100.0 1210200.0 219300.0 1211400.0 ;
      RECT  218100.0 1210200.0 219300.0 1211400.0 ;
      RECT  215700.0 1210200.0 216900.0 1211400.0 ;
      RECT  215400.0 1205250.0 214200.0 1206450.0 ;
      RECT  215700.0 1215600.0 216900.0 1216800.0 ;
      RECT  213300.0 1203000.0 214500.0 1204200.0 ;
      RECT  215700.0 1203000.0 216900.0 1204200.0 ;
      RECT  213300.0 1210200.0 214500.0 1211400.0 ;
      RECT  218100.0 1210200.0 219300.0 1211400.0 ;
      RECT  210300.0 1205400.0 220500.0 1206300.0 ;
      RECT  210300.0 1216500.0 220500.0 1217400.0 ;
      RECT  225900.0 1210200.0 227100.0 1217400.0 ;
      RECT  223500.0 1203000.0 224700.0 1204200.0 ;
      RECT  225900.0 1203000.0 227100.0 1204200.0 ;
      RECT  225900.0 1203000.0 227100.0 1204200.0 ;
      RECT  223500.0 1203000.0 224700.0 1204200.0 ;
      RECT  223500.0 1210200.0 224700.0 1211400.0 ;
      RECT  225900.0 1210200.0 227100.0 1211400.0 ;
      RECT  225900.0 1210200.0 227100.0 1211400.0 ;
      RECT  223500.0 1210200.0 224700.0 1211400.0 ;
      RECT  225900.0 1210200.0 227100.0 1211400.0 ;
      RECT  228300.0 1210200.0 229500.0 1211400.0 ;
      RECT  228300.0 1210200.0 229500.0 1211400.0 ;
      RECT  225900.0 1210200.0 227100.0 1211400.0 ;
      RECT  225600.0 1205250.0 224400.0 1206450.0 ;
      RECT  225900.0 1215600.0 227100.0 1216800.0 ;
      RECT  223500.0 1203000.0 224700.0 1204200.0 ;
      RECT  225900.0 1203000.0 227100.0 1204200.0 ;
      RECT  223500.0 1210200.0 224700.0 1211400.0 ;
      RECT  228300.0 1210200.0 229500.0 1211400.0 ;
      RECT  220500.0 1205400.0 230700.0 1206300.0 ;
      RECT  220500.0 1216500.0 230700.0 1217400.0 ;
      RECT  236100.0 1210200.0 237300.0 1217400.0 ;
      RECT  233700.0 1203000.0 234900.0 1204200.0 ;
      RECT  236100.0 1203000.0 237300.0 1204200.0 ;
      RECT  236100.0 1203000.0 237300.0 1204200.0 ;
      RECT  233700.0 1203000.0 234900.0 1204200.0 ;
      RECT  233700.0 1210200.0 234900.0 1211400.0 ;
      RECT  236100.0 1210200.0 237300.0 1211400.0 ;
      RECT  236100.0 1210200.0 237300.0 1211400.0 ;
      RECT  233700.0 1210200.0 234900.0 1211400.0 ;
      RECT  236100.0 1210200.0 237300.0 1211400.0 ;
      RECT  238500.0 1210200.0 239700.0 1211400.0 ;
      RECT  238500.0 1210200.0 239700.0 1211400.0 ;
      RECT  236100.0 1210200.0 237300.0 1211400.0 ;
      RECT  235800.0 1205250.0 234600.0 1206450.0 ;
      RECT  236100.0 1215600.0 237300.0 1216800.0 ;
      RECT  233700.0 1203000.0 234900.0 1204200.0 ;
      RECT  236100.0 1203000.0 237300.0 1204200.0 ;
      RECT  233700.0 1210200.0 234900.0 1211400.0 ;
      RECT  238500.0 1210200.0 239700.0 1211400.0 ;
      RECT  230700.0 1205400.0 240900.0 1206300.0 ;
      RECT  230700.0 1216500.0 240900.0 1217400.0 ;
      RECT  246300.0 1210200.0 247500.0 1217400.0 ;
      RECT  243900.0 1203000.0 245100.0 1204200.0 ;
      RECT  246300.0 1203000.0 247500.0 1204200.0 ;
      RECT  246300.0 1203000.0 247500.0 1204200.0 ;
      RECT  243900.0 1203000.0 245100.0 1204200.0 ;
      RECT  243900.0 1210200.0 245100.0 1211400.0 ;
      RECT  246300.0 1210200.0 247500.0 1211400.0 ;
      RECT  246300.0 1210200.0 247500.0 1211400.0 ;
      RECT  243900.0 1210200.0 245100.0 1211400.0 ;
      RECT  246300.0 1210200.0 247500.0 1211400.0 ;
      RECT  248700.0 1210200.0 249900.0 1211400.0 ;
      RECT  248700.0 1210200.0 249900.0 1211400.0 ;
      RECT  246300.0 1210200.0 247500.0 1211400.0 ;
      RECT  246000.0 1205250.0 244800.0 1206450.0 ;
      RECT  246300.0 1215600.0 247500.0 1216800.0 ;
      RECT  243900.0 1203000.0 245100.0 1204200.0 ;
      RECT  246300.0 1203000.0 247500.0 1204200.0 ;
      RECT  243900.0 1210200.0 245100.0 1211400.0 ;
      RECT  248700.0 1210200.0 249900.0 1211400.0 ;
      RECT  240900.0 1205400.0 251100.0 1206300.0 ;
      RECT  240900.0 1216500.0 251100.0 1217400.0 ;
      RECT  256500.0 1210200.0 257700.0 1217400.0 ;
      RECT  254100.0 1203000.0 255300.0 1204200.0 ;
      RECT  256500.0 1203000.0 257700.0 1204200.0 ;
      RECT  256500.0 1203000.0 257700.0 1204200.0 ;
      RECT  254100.0 1203000.0 255300.0 1204200.0 ;
      RECT  254100.0 1210200.0 255300.0 1211400.0 ;
      RECT  256500.0 1210200.0 257700.0 1211400.0 ;
      RECT  256500.0 1210200.0 257700.0 1211400.0 ;
      RECT  254100.0 1210200.0 255300.0 1211400.0 ;
      RECT  256500.0 1210200.0 257700.0 1211400.0 ;
      RECT  258900.0 1210200.0 260100.0 1211400.0 ;
      RECT  258900.0 1210200.0 260100.0 1211400.0 ;
      RECT  256500.0 1210200.0 257700.0 1211400.0 ;
      RECT  256200.0 1205250.0 255000.0 1206450.0 ;
      RECT  256500.0 1215600.0 257700.0 1216800.0 ;
      RECT  254100.0 1203000.0 255300.0 1204200.0 ;
      RECT  256500.0 1203000.0 257700.0 1204200.0 ;
      RECT  254100.0 1210200.0 255300.0 1211400.0 ;
      RECT  258900.0 1210200.0 260100.0 1211400.0 ;
      RECT  251100.0 1205400.0 261300.0 1206300.0 ;
      RECT  251100.0 1216500.0 261300.0 1217400.0 ;
      RECT  266700.0 1210200.0 267900.0 1217400.0 ;
      RECT  264300.0 1203000.0 265500.0 1204200.0 ;
      RECT  266700.0 1203000.0 267900.0 1204200.0 ;
      RECT  266700.0 1203000.0 267900.0 1204200.0 ;
      RECT  264300.0 1203000.0 265500.0 1204200.0 ;
      RECT  264300.0 1210200.0 265500.0 1211400.0 ;
      RECT  266700.0 1210200.0 267900.0 1211400.0 ;
      RECT  266700.0 1210200.0 267900.0 1211400.0 ;
      RECT  264300.0 1210200.0 265500.0 1211400.0 ;
      RECT  266700.0 1210200.0 267900.0 1211400.0 ;
      RECT  269100.0 1210200.0 270300.0 1211400.0 ;
      RECT  269100.0 1210200.0 270300.0 1211400.0 ;
      RECT  266700.0 1210200.0 267900.0 1211400.0 ;
      RECT  266400.0 1205250.0 265200.0 1206450.0 ;
      RECT  266700.0 1215600.0 267900.0 1216800.0 ;
      RECT  264300.0 1203000.0 265500.0 1204200.0 ;
      RECT  266700.0 1203000.0 267900.0 1204200.0 ;
      RECT  264300.0 1210200.0 265500.0 1211400.0 ;
      RECT  269100.0 1210200.0 270300.0 1211400.0 ;
      RECT  261300.0 1205400.0 271500.0 1206300.0 ;
      RECT  261300.0 1216500.0 271500.0 1217400.0 ;
      RECT  276900.0 1210200.0 278100.0 1217400.0 ;
      RECT  274500.0 1203000.0 275700.0 1204200.0 ;
      RECT  276900.0 1203000.0 278100.0 1204200.0 ;
      RECT  276900.0 1203000.0 278100.0 1204200.0 ;
      RECT  274500.0 1203000.0 275700.0 1204200.0 ;
      RECT  274500.0 1210200.0 275700.0 1211400.0 ;
      RECT  276900.0 1210200.0 278100.0 1211400.0 ;
      RECT  276900.0 1210200.0 278100.0 1211400.0 ;
      RECT  274500.0 1210200.0 275700.0 1211400.0 ;
      RECT  276900.0 1210200.0 278100.0 1211400.0 ;
      RECT  279300.0 1210200.0 280500.0 1211400.0 ;
      RECT  279300.0 1210200.0 280500.0 1211400.0 ;
      RECT  276900.0 1210200.0 278100.0 1211400.0 ;
      RECT  276600.0 1205250.0 275400.0 1206450.0 ;
      RECT  276900.0 1215600.0 278100.0 1216800.0 ;
      RECT  274500.0 1203000.0 275700.0 1204200.0 ;
      RECT  276900.0 1203000.0 278100.0 1204200.0 ;
      RECT  274500.0 1210200.0 275700.0 1211400.0 ;
      RECT  279300.0 1210200.0 280500.0 1211400.0 ;
      RECT  271500.0 1205400.0 281700.0 1206300.0 ;
      RECT  271500.0 1216500.0 281700.0 1217400.0 ;
      RECT  287100.0 1210200.0 288300.0 1217400.0 ;
      RECT  284700.0 1203000.0 285900.0 1204200.0 ;
      RECT  287100.0 1203000.0 288300.0 1204200.0 ;
      RECT  287100.0 1203000.0 288300.0 1204200.0 ;
      RECT  284700.0 1203000.0 285900.0 1204200.0 ;
      RECT  284700.0 1210200.0 285900.0 1211400.0 ;
      RECT  287100.0 1210200.0 288300.0 1211400.0 ;
      RECT  287100.0 1210200.0 288300.0 1211400.0 ;
      RECT  284700.0 1210200.0 285900.0 1211400.0 ;
      RECT  287100.0 1210200.0 288300.0 1211400.0 ;
      RECT  289500.0 1210200.0 290700.0 1211400.0 ;
      RECT  289500.0 1210200.0 290700.0 1211400.0 ;
      RECT  287100.0 1210200.0 288300.0 1211400.0 ;
      RECT  286800.0 1205250.0 285600.0 1206450.0 ;
      RECT  287100.0 1215600.0 288300.0 1216800.0 ;
      RECT  284700.0 1203000.0 285900.0 1204200.0 ;
      RECT  287100.0 1203000.0 288300.0 1204200.0 ;
      RECT  284700.0 1210200.0 285900.0 1211400.0 ;
      RECT  289500.0 1210200.0 290700.0 1211400.0 ;
      RECT  281700.0 1205400.0 291900.0 1206300.0 ;
      RECT  281700.0 1216500.0 291900.0 1217400.0 ;
      RECT  297300.0 1210200.0 298500.0 1217400.0 ;
      RECT  294900.0 1203000.0 296100.0 1204200.0 ;
      RECT  297300.0 1203000.0 298500.0 1204200.0 ;
      RECT  297300.0 1203000.0 298500.0 1204200.0 ;
      RECT  294900.0 1203000.0 296100.0 1204200.0 ;
      RECT  294900.0 1210200.0 296100.0 1211400.0 ;
      RECT  297300.0 1210200.0 298500.0 1211400.0 ;
      RECT  297300.0 1210200.0 298500.0 1211400.0 ;
      RECT  294900.0 1210200.0 296100.0 1211400.0 ;
      RECT  297300.0 1210200.0 298500.0 1211400.0 ;
      RECT  299700.0 1210200.0 300900.0 1211400.0 ;
      RECT  299700.0 1210200.0 300900.0 1211400.0 ;
      RECT  297300.0 1210200.0 298500.0 1211400.0 ;
      RECT  297000.0 1205250.0 295800.0 1206450.0 ;
      RECT  297300.0 1215600.0 298500.0 1216800.0 ;
      RECT  294900.0 1203000.0 296100.0 1204200.0 ;
      RECT  297300.0 1203000.0 298500.0 1204200.0 ;
      RECT  294900.0 1210200.0 296100.0 1211400.0 ;
      RECT  299700.0 1210200.0 300900.0 1211400.0 ;
      RECT  291900.0 1205400.0 302100.0 1206300.0 ;
      RECT  291900.0 1216500.0 302100.0 1217400.0 ;
      RECT  307500.0 1210200.0 308700.0 1217400.0 ;
      RECT  305100.0 1203000.0 306300.0 1204200.0 ;
      RECT  307500.0 1203000.0 308700.0 1204200.0 ;
      RECT  307500.0 1203000.0 308700.0 1204200.0 ;
      RECT  305100.0 1203000.0 306300.0 1204200.0 ;
      RECT  305100.0 1210200.0 306300.0 1211400.0 ;
      RECT  307500.0 1210200.0 308700.0 1211400.0 ;
      RECT  307500.0 1210200.0 308700.0 1211400.0 ;
      RECT  305100.0 1210200.0 306300.0 1211400.0 ;
      RECT  307500.0 1210200.0 308700.0 1211400.0 ;
      RECT  309900.0 1210200.0 311100.0 1211400.0 ;
      RECT  309900.0 1210200.0 311100.0 1211400.0 ;
      RECT  307500.0 1210200.0 308700.0 1211400.0 ;
      RECT  307200.0 1205250.0 306000.0 1206450.0 ;
      RECT  307500.0 1215600.0 308700.0 1216800.0 ;
      RECT  305100.0 1203000.0 306300.0 1204200.0 ;
      RECT  307500.0 1203000.0 308700.0 1204200.0 ;
      RECT  305100.0 1210200.0 306300.0 1211400.0 ;
      RECT  309900.0 1210200.0 311100.0 1211400.0 ;
      RECT  302100.0 1205400.0 312300.0 1206300.0 ;
      RECT  302100.0 1216500.0 312300.0 1217400.0 ;
      RECT  317700.0 1210200.0 318900.0 1217400.0 ;
      RECT  315300.0 1203000.0 316500.0 1204200.0 ;
      RECT  317700.0 1203000.0 318900.0 1204200.0 ;
      RECT  317700.0 1203000.0 318900.0 1204200.0 ;
      RECT  315300.0 1203000.0 316500.0 1204200.0 ;
      RECT  315300.0 1210200.0 316500.0 1211400.0 ;
      RECT  317700.0 1210200.0 318900.0 1211400.0 ;
      RECT  317700.0 1210200.0 318900.0 1211400.0 ;
      RECT  315300.0 1210200.0 316500.0 1211400.0 ;
      RECT  317700.0 1210200.0 318900.0 1211400.0 ;
      RECT  320100.0 1210200.0 321300.0 1211400.0 ;
      RECT  320100.0 1210200.0 321300.0 1211400.0 ;
      RECT  317700.0 1210200.0 318900.0 1211400.0 ;
      RECT  317400.0 1205250.0 316200.0 1206450.0 ;
      RECT  317700.0 1215600.0 318900.0 1216800.0 ;
      RECT  315300.0 1203000.0 316500.0 1204200.0 ;
      RECT  317700.0 1203000.0 318900.0 1204200.0 ;
      RECT  315300.0 1210200.0 316500.0 1211400.0 ;
      RECT  320100.0 1210200.0 321300.0 1211400.0 ;
      RECT  312300.0 1205400.0 322500.0 1206300.0 ;
      RECT  312300.0 1216500.0 322500.0 1217400.0 ;
      RECT  327900.0 1210200.0 329100.0 1217400.0 ;
      RECT  325500.0 1203000.0 326700.0 1204200.0 ;
      RECT  327900.0 1203000.0 329100.0 1204200.0 ;
      RECT  327900.0 1203000.0 329100.0 1204200.0 ;
      RECT  325500.0 1203000.0 326700.0 1204200.0 ;
      RECT  325500.0 1210200.0 326700.0 1211400.0 ;
      RECT  327900.0 1210200.0 329100.0 1211400.0 ;
      RECT  327900.0 1210200.0 329100.0 1211400.0 ;
      RECT  325500.0 1210200.0 326700.0 1211400.0 ;
      RECT  327900.0 1210200.0 329100.0 1211400.0 ;
      RECT  330300.0 1210200.0 331500.0 1211400.0 ;
      RECT  330300.0 1210200.0 331500.0 1211400.0 ;
      RECT  327900.0 1210200.0 329100.0 1211400.0 ;
      RECT  327600.0 1205250.0 326400.0 1206450.0 ;
      RECT  327900.0 1215600.0 329100.0 1216800.0 ;
      RECT  325500.0 1203000.0 326700.0 1204200.0 ;
      RECT  327900.0 1203000.0 329100.0 1204200.0 ;
      RECT  325500.0 1210200.0 326700.0 1211400.0 ;
      RECT  330300.0 1210200.0 331500.0 1211400.0 ;
      RECT  322500.0 1205400.0 332700.0 1206300.0 ;
      RECT  322500.0 1216500.0 332700.0 1217400.0 ;
      RECT  338100.0 1210200.0 339300.0 1217400.0 ;
      RECT  335700.0 1203000.0 336900.0 1204200.0 ;
      RECT  338100.0 1203000.0 339300.0 1204200.0 ;
      RECT  338100.0 1203000.0 339300.0 1204200.0 ;
      RECT  335700.0 1203000.0 336900.0 1204200.0 ;
      RECT  335700.0 1210200.0 336900.0 1211400.0 ;
      RECT  338100.0 1210200.0 339300.0 1211400.0 ;
      RECT  338100.0 1210200.0 339300.0 1211400.0 ;
      RECT  335700.0 1210200.0 336900.0 1211400.0 ;
      RECT  338100.0 1210200.0 339300.0 1211400.0 ;
      RECT  340500.0 1210200.0 341700.0 1211400.0 ;
      RECT  340500.0 1210200.0 341700.0 1211400.0 ;
      RECT  338100.0 1210200.0 339300.0 1211400.0 ;
      RECT  337800.0 1205250.0 336600.0 1206450.0 ;
      RECT  338100.0 1215600.0 339300.0 1216800.0 ;
      RECT  335700.0 1203000.0 336900.0 1204200.0 ;
      RECT  338100.0 1203000.0 339300.0 1204200.0 ;
      RECT  335700.0 1210200.0 336900.0 1211400.0 ;
      RECT  340500.0 1210200.0 341700.0 1211400.0 ;
      RECT  332700.0 1205400.0 342900.0 1206300.0 ;
      RECT  332700.0 1216500.0 342900.0 1217400.0 ;
      RECT  348300.0 1210200.0 349500.0 1217400.0 ;
      RECT  345900.0 1203000.0 347100.0 1204200.0 ;
      RECT  348300.0 1203000.0 349500.0 1204200.0 ;
      RECT  348300.0 1203000.0 349500.0 1204200.0 ;
      RECT  345900.0 1203000.0 347100.0 1204200.0 ;
      RECT  345900.0 1210200.0 347100.0 1211400.0 ;
      RECT  348300.0 1210200.0 349500.0 1211400.0 ;
      RECT  348300.0 1210200.0 349500.0 1211400.0 ;
      RECT  345900.0 1210200.0 347100.0 1211400.0 ;
      RECT  348300.0 1210200.0 349500.0 1211400.0 ;
      RECT  350700.0 1210200.0 351900.0 1211400.0 ;
      RECT  350700.0 1210200.0 351900.0 1211400.0 ;
      RECT  348300.0 1210200.0 349500.0 1211400.0 ;
      RECT  348000.0 1205250.0 346800.0 1206450.0 ;
      RECT  348300.0 1215600.0 349500.0 1216800.0 ;
      RECT  345900.0 1203000.0 347100.0 1204200.0 ;
      RECT  348300.0 1203000.0 349500.0 1204200.0 ;
      RECT  345900.0 1210200.0 347100.0 1211400.0 ;
      RECT  350700.0 1210200.0 351900.0 1211400.0 ;
      RECT  342900.0 1205400.0 353100.0 1206300.0 ;
      RECT  342900.0 1216500.0 353100.0 1217400.0 ;
      RECT  358500.0 1210200.0 359700.0 1217400.0 ;
      RECT  356100.0 1203000.0 357300.0 1204200.0 ;
      RECT  358500.0 1203000.0 359700.0 1204200.0 ;
      RECT  358500.0 1203000.0 359700.0 1204200.0 ;
      RECT  356100.0 1203000.0 357300.0 1204200.0 ;
      RECT  356100.0 1210200.0 357300.0 1211400.0 ;
      RECT  358500.0 1210200.0 359700.0 1211400.0 ;
      RECT  358500.0 1210200.0 359700.0 1211400.0 ;
      RECT  356100.0 1210200.0 357300.0 1211400.0 ;
      RECT  358500.0 1210200.0 359700.0 1211400.0 ;
      RECT  360900.0 1210200.0 362100.0 1211400.0 ;
      RECT  360900.0 1210200.0 362100.0 1211400.0 ;
      RECT  358500.0 1210200.0 359700.0 1211400.0 ;
      RECT  358200.0 1205250.0 357000.0 1206450.0 ;
      RECT  358500.0 1215600.0 359700.0 1216800.0 ;
      RECT  356100.0 1203000.0 357300.0 1204200.0 ;
      RECT  358500.0 1203000.0 359700.0 1204200.0 ;
      RECT  356100.0 1210200.0 357300.0 1211400.0 ;
      RECT  360900.0 1210200.0 362100.0 1211400.0 ;
      RECT  353100.0 1205400.0 363300.0 1206300.0 ;
      RECT  353100.0 1216500.0 363300.0 1217400.0 ;
      RECT  368700.0 1210200.0 369900.0 1217400.0 ;
      RECT  366300.0 1203000.0 367500.0 1204200.0 ;
      RECT  368700.0 1203000.0 369900.0 1204200.0 ;
      RECT  368700.0 1203000.0 369900.0 1204200.0 ;
      RECT  366300.0 1203000.0 367500.0 1204200.0 ;
      RECT  366300.0 1210200.0 367500.0 1211400.0 ;
      RECT  368700.0 1210200.0 369900.0 1211400.0 ;
      RECT  368700.0 1210200.0 369900.0 1211400.0 ;
      RECT  366300.0 1210200.0 367500.0 1211400.0 ;
      RECT  368700.0 1210200.0 369900.0 1211400.0 ;
      RECT  371100.0 1210200.0 372300.0 1211400.0 ;
      RECT  371100.0 1210200.0 372300.0 1211400.0 ;
      RECT  368700.0 1210200.0 369900.0 1211400.0 ;
      RECT  368400.0 1205250.0 367200.0 1206450.0 ;
      RECT  368700.0 1215600.0 369900.0 1216800.0 ;
      RECT  366300.0 1203000.0 367500.0 1204200.0 ;
      RECT  368700.0 1203000.0 369900.0 1204200.0 ;
      RECT  366300.0 1210200.0 367500.0 1211400.0 ;
      RECT  371100.0 1210200.0 372300.0 1211400.0 ;
      RECT  363300.0 1205400.0 373500.0 1206300.0 ;
      RECT  363300.0 1216500.0 373500.0 1217400.0 ;
      RECT  378900.0 1210200.0 380100.0 1217400.0 ;
      RECT  376500.0 1203000.0 377700.0 1204200.0 ;
      RECT  378900.0 1203000.0 380100.0 1204200.0 ;
      RECT  378900.0 1203000.0 380100.0 1204200.0 ;
      RECT  376500.0 1203000.0 377700.0 1204200.0 ;
      RECT  376500.0 1210200.0 377700.0 1211400.0 ;
      RECT  378900.0 1210200.0 380100.0 1211400.0 ;
      RECT  378900.0 1210200.0 380100.0 1211400.0 ;
      RECT  376500.0 1210200.0 377700.0 1211400.0 ;
      RECT  378900.0 1210200.0 380100.0 1211400.0 ;
      RECT  381300.0 1210200.0 382500.0 1211400.0 ;
      RECT  381300.0 1210200.0 382500.0 1211400.0 ;
      RECT  378900.0 1210200.0 380100.0 1211400.0 ;
      RECT  378600.0 1205250.0 377400.0 1206450.0 ;
      RECT  378900.0 1215600.0 380100.0 1216800.0 ;
      RECT  376500.0 1203000.0 377700.0 1204200.0 ;
      RECT  378900.0 1203000.0 380100.0 1204200.0 ;
      RECT  376500.0 1210200.0 377700.0 1211400.0 ;
      RECT  381300.0 1210200.0 382500.0 1211400.0 ;
      RECT  373500.0 1205400.0 383700.0 1206300.0 ;
      RECT  373500.0 1216500.0 383700.0 1217400.0 ;
      RECT  389100.0 1210200.0 390300.0 1217400.0 ;
      RECT  386700.0 1203000.0 387900.0 1204200.0 ;
      RECT  389100.0 1203000.0 390300.0 1204200.0 ;
      RECT  389100.0 1203000.0 390300.0 1204200.0 ;
      RECT  386700.0 1203000.0 387900.0 1204200.0 ;
      RECT  386700.0 1210200.0 387900.0 1211400.0 ;
      RECT  389100.0 1210200.0 390300.0 1211400.0 ;
      RECT  389100.0 1210200.0 390300.0 1211400.0 ;
      RECT  386700.0 1210200.0 387900.0 1211400.0 ;
      RECT  389100.0 1210200.0 390300.0 1211400.0 ;
      RECT  391500.0 1210200.0 392700.0 1211400.0 ;
      RECT  391500.0 1210200.0 392700.0 1211400.0 ;
      RECT  389100.0 1210200.0 390300.0 1211400.0 ;
      RECT  388800.0 1205250.0 387600.0 1206450.0 ;
      RECT  389100.0 1215600.0 390300.0 1216800.0 ;
      RECT  386700.0 1203000.0 387900.0 1204200.0 ;
      RECT  389100.0 1203000.0 390300.0 1204200.0 ;
      RECT  386700.0 1210200.0 387900.0 1211400.0 ;
      RECT  391500.0 1210200.0 392700.0 1211400.0 ;
      RECT  383700.0 1205400.0 393900.0 1206300.0 ;
      RECT  383700.0 1216500.0 393900.0 1217400.0 ;
      RECT  399300.0 1210200.0 400500.0 1217400.0 ;
      RECT  396900.0 1203000.0 398100.0 1204200.0 ;
      RECT  399300.0 1203000.0 400500.0 1204200.0 ;
      RECT  399300.0 1203000.0 400500.0 1204200.0 ;
      RECT  396900.0 1203000.0 398100.0 1204200.0 ;
      RECT  396900.0 1210200.0 398100.0 1211400.0 ;
      RECT  399300.0 1210200.0 400500.0 1211400.0 ;
      RECT  399300.0 1210200.0 400500.0 1211400.0 ;
      RECT  396900.0 1210200.0 398100.0 1211400.0 ;
      RECT  399300.0 1210200.0 400500.0 1211400.0 ;
      RECT  401700.0 1210200.0 402900.0 1211400.0 ;
      RECT  401700.0 1210200.0 402900.0 1211400.0 ;
      RECT  399300.0 1210200.0 400500.0 1211400.0 ;
      RECT  399000.0 1205250.0 397800.0 1206450.0 ;
      RECT  399300.0 1215600.0 400500.0 1216800.0 ;
      RECT  396900.0 1203000.0 398100.0 1204200.0 ;
      RECT  399300.0 1203000.0 400500.0 1204200.0 ;
      RECT  396900.0 1210200.0 398100.0 1211400.0 ;
      RECT  401700.0 1210200.0 402900.0 1211400.0 ;
      RECT  393900.0 1205400.0 404100.0 1206300.0 ;
      RECT  393900.0 1216500.0 404100.0 1217400.0 ;
      RECT  409500.0 1210200.0 410700.0 1217400.0 ;
      RECT  407100.0 1203000.0 408300.0 1204200.0 ;
      RECT  409500.0 1203000.0 410700.0 1204200.0 ;
      RECT  409500.0 1203000.0 410700.0 1204200.0 ;
      RECT  407100.0 1203000.0 408300.0 1204200.0 ;
      RECT  407100.0 1210200.0 408300.0 1211400.0 ;
      RECT  409500.0 1210200.0 410700.0 1211400.0 ;
      RECT  409500.0 1210200.0 410700.0 1211400.0 ;
      RECT  407100.0 1210200.0 408300.0 1211400.0 ;
      RECT  409500.0 1210200.0 410700.0 1211400.0 ;
      RECT  411900.0 1210200.0 413100.0 1211400.0 ;
      RECT  411900.0 1210200.0 413100.0 1211400.0 ;
      RECT  409500.0 1210200.0 410700.0 1211400.0 ;
      RECT  409200.0 1205250.0 408000.0 1206450.0 ;
      RECT  409500.0 1215600.0 410700.0 1216800.0 ;
      RECT  407100.0 1203000.0 408300.0 1204200.0 ;
      RECT  409500.0 1203000.0 410700.0 1204200.0 ;
      RECT  407100.0 1210200.0 408300.0 1211400.0 ;
      RECT  411900.0 1210200.0 413100.0 1211400.0 ;
      RECT  404100.0 1205400.0 414300.0 1206300.0 ;
      RECT  404100.0 1216500.0 414300.0 1217400.0 ;
      RECT  419700.0 1210200.0 420900.0 1217400.0 ;
      RECT  417300.0 1203000.0 418500.0 1204200.0 ;
      RECT  419700.0 1203000.0 420900.0 1204200.0 ;
      RECT  419700.0 1203000.0 420900.0 1204200.0 ;
      RECT  417300.0 1203000.0 418500.0 1204200.0 ;
      RECT  417300.0 1210200.0 418500.0 1211400.0 ;
      RECT  419700.0 1210200.0 420900.0 1211400.0 ;
      RECT  419700.0 1210200.0 420900.0 1211400.0 ;
      RECT  417300.0 1210200.0 418500.0 1211400.0 ;
      RECT  419700.0 1210200.0 420900.0 1211400.0 ;
      RECT  422100.0 1210200.0 423300.0 1211400.0 ;
      RECT  422100.0 1210200.0 423300.0 1211400.0 ;
      RECT  419700.0 1210200.0 420900.0 1211400.0 ;
      RECT  419400.0 1205250.0 418200.0 1206450.0 ;
      RECT  419700.0 1215600.0 420900.0 1216800.0 ;
      RECT  417300.0 1203000.0 418500.0 1204200.0 ;
      RECT  419700.0 1203000.0 420900.0 1204200.0 ;
      RECT  417300.0 1210200.0 418500.0 1211400.0 ;
      RECT  422100.0 1210200.0 423300.0 1211400.0 ;
      RECT  414300.0 1205400.0 424500.0 1206300.0 ;
      RECT  414300.0 1216500.0 424500.0 1217400.0 ;
      RECT  429900.0 1210200.0 431100.0 1217400.0 ;
      RECT  427500.0 1203000.0 428700.0 1204200.0 ;
      RECT  429900.0 1203000.0 431100.0 1204200.0 ;
      RECT  429900.0 1203000.0 431100.0 1204200.0 ;
      RECT  427500.0 1203000.0 428700.0 1204200.0 ;
      RECT  427500.0 1210200.0 428700.0 1211400.0 ;
      RECT  429900.0 1210200.0 431100.0 1211400.0 ;
      RECT  429900.0 1210200.0 431100.0 1211400.0 ;
      RECT  427500.0 1210200.0 428700.0 1211400.0 ;
      RECT  429900.0 1210200.0 431100.0 1211400.0 ;
      RECT  432300.0 1210200.0 433500.0 1211400.0 ;
      RECT  432300.0 1210200.0 433500.0 1211400.0 ;
      RECT  429900.0 1210200.0 431100.0 1211400.0 ;
      RECT  429600.0 1205250.0 428400.0 1206450.0 ;
      RECT  429900.0 1215600.0 431100.0 1216800.0 ;
      RECT  427500.0 1203000.0 428700.0 1204200.0 ;
      RECT  429900.0 1203000.0 431100.0 1204200.0 ;
      RECT  427500.0 1210200.0 428700.0 1211400.0 ;
      RECT  432300.0 1210200.0 433500.0 1211400.0 ;
      RECT  424500.0 1205400.0 434700.0 1206300.0 ;
      RECT  424500.0 1216500.0 434700.0 1217400.0 ;
      RECT  440100.0 1210200.0 441300.0 1217400.0 ;
      RECT  437700.0 1203000.0 438900.0 1204200.0 ;
      RECT  440100.0 1203000.0 441300.0 1204200.0 ;
      RECT  440100.0 1203000.0 441300.0 1204200.0 ;
      RECT  437700.0 1203000.0 438900.0 1204200.0 ;
      RECT  437700.0 1210200.0 438900.0 1211400.0 ;
      RECT  440100.0 1210200.0 441300.0 1211400.0 ;
      RECT  440100.0 1210200.0 441300.0 1211400.0 ;
      RECT  437700.0 1210200.0 438900.0 1211400.0 ;
      RECT  440100.0 1210200.0 441300.0 1211400.0 ;
      RECT  442500.0 1210200.0 443700.0 1211400.0 ;
      RECT  442500.0 1210200.0 443700.0 1211400.0 ;
      RECT  440100.0 1210200.0 441300.0 1211400.0 ;
      RECT  439800.0 1205250.0 438600.0 1206450.0 ;
      RECT  440100.0 1215600.0 441300.0 1216800.0 ;
      RECT  437700.0 1203000.0 438900.0 1204200.0 ;
      RECT  440100.0 1203000.0 441300.0 1204200.0 ;
      RECT  437700.0 1210200.0 438900.0 1211400.0 ;
      RECT  442500.0 1210200.0 443700.0 1211400.0 ;
      RECT  434700.0 1205400.0 444900.0 1206300.0 ;
      RECT  434700.0 1216500.0 444900.0 1217400.0 ;
      RECT  450300.0 1210200.0 451500.0 1217400.0 ;
      RECT  447900.0 1203000.0 449100.0 1204200.0 ;
      RECT  450300.0 1203000.0 451500.0 1204200.0 ;
      RECT  450300.0 1203000.0 451500.0 1204200.0 ;
      RECT  447900.0 1203000.0 449100.0 1204200.0 ;
      RECT  447900.0 1210200.0 449100.0 1211400.0 ;
      RECT  450300.0 1210200.0 451500.0 1211400.0 ;
      RECT  450300.0 1210200.0 451500.0 1211400.0 ;
      RECT  447900.0 1210200.0 449100.0 1211400.0 ;
      RECT  450300.0 1210200.0 451500.0 1211400.0 ;
      RECT  452700.0 1210200.0 453900.0 1211400.0 ;
      RECT  452700.0 1210200.0 453900.0 1211400.0 ;
      RECT  450300.0 1210200.0 451500.0 1211400.0 ;
      RECT  450000.0 1205250.0 448800.0 1206450.0 ;
      RECT  450300.0 1215600.0 451500.0 1216800.0 ;
      RECT  447900.0 1203000.0 449100.0 1204200.0 ;
      RECT  450300.0 1203000.0 451500.0 1204200.0 ;
      RECT  447900.0 1210200.0 449100.0 1211400.0 ;
      RECT  452700.0 1210200.0 453900.0 1211400.0 ;
      RECT  444900.0 1205400.0 455100.0 1206300.0 ;
      RECT  444900.0 1216500.0 455100.0 1217400.0 ;
      RECT  460500.0 1210200.0 461700.0 1217400.0 ;
      RECT  458100.0 1203000.0 459300.0 1204200.0 ;
      RECT  460500.0 1203000.0 461700.0 1204200.0 ;
      RECT  460500.0 1203000.0 461700.0 1204200.0 ;
      RECT  458100.0 1203000.0 459300.0 1204200.0 ;
      RECT  458100.0 1210200.0 459300.0 1211400.0 ;
      RECT  460500.0 1210200.0 461700.0 1211400.0 ;
      RECT  460500.0 1210200.0 461700.0 1211400.0 ;
      RECT  458100.0 1210200.0 459300.0 1211400.0 ;
      RECT  460500.0 1210200.0 461700.0 1211400.0 ;
      RECT  462900.0 1210200.0 464100.0 1211400.0 ;
      RECT  462900.0 1210200.0 464100.0 1211400.0 ;
      RECT  460500.0 1210200.0 461700.0 1211400.0 ;
      RECT  460200.0 1205250.0 459000.0 1206450.0 ;
      RECT  460500.0 1215600.0 461700.0 1216800.0 ;
      RECT  458100.0 1203000.0 459300.0 1204200.0 ;
      RECT  460500.0 1203000.0 461700.0 1204200.0 ;
      RECT  458100.0 1210200.0 459300.0 1211400.0 ;
      RECT  462900.0 1210200.0 464100.0 1211400.0 ;
      RECT  455100.0 1205400.0 465300.0 1206300.0 ;
      RECT  455100.0 1216500.0 465300.0 1217400.0 ;
      RECT  470700.0 1210200.0 471900.0 1217400.0 ;
      RECT  468300.0 1203000.0 469500.0 1204200.0 ;
      RECT  470700.0 1203000.0 471900.0 1204200.0 ;
      RECT  470700.0 1203000.0 471900.0 1204200.0 ;
      RECT  468300.0 1203000.0 469500.0 1204200.0 ;
      RECT  468300.0 1210200.0 469500.0 1211400.0 ;
      RECT  470700.0 1210200.0 471900.0 1211400.0 ;
      RECT  470700.0 1210200.0 471900.0 1211400.0 ;
      RECT  468300.0 1210200.0 469500.0 1211400.0 ;
      RECT  470700.0 1210200.0 471900.0 1211400.0 ;
      RECT  473100.0 1210200.0 474300.0 1211400.0 ;
      RECT  473100.0 1210200.0 474300.0 1211400.0 ;
      RECT  470700.0 1210200.0 471900.0 1211400.0 ;
      RECT  470400.0 1205250.0 469200.0 1206450.0 ;
      RECT  470700.0 1215600.0 471900.0 1216800.0 ;
      RECT  468300.0 1203000.0 469500.0 1204200.0 ;
      RECT  470700.0 1203000.0 471900.0 1204200.0 ;
      RECT  468300.0 1210200.0 469500.0 1211400.0 ;
      RECT  473100.0 1210200.0 474300.0 1211400.0 ;
      RECT  465300.0 1205400.0 475500.0 1206300.0 ;
      RECT  465300.0 1216500.0 475500.0 1217400.0 ;
      RECT  480900.0 1210200.0 482100.0 1217400.0 ;
      RECT  478500.0 1203000.0 479700.0 1204200.0 ;
      RECT  480900.0 1203000.0 482100.0 1204200.0 ;
      RECT  480900.0 1203000.0 482100.0 1204200.0 ;
      RECT  478500.0 1203000.0 479700.0 1204200.0 ;
      RECT  478500.0 1210200.0 479700.0 1211400.0 ;
      RECT  480900.0 1210200.0 482100.0 1211400.0 ;
      RECT  480900.0 1210200.0 482100.0 1211400.0 ;
      RECT  478500.0 1210200.0 479700.0 1211400.0 ;
      RECT  480900.0 1210200.0 482100.0 1211400.0 ;
      RECT  483300.0 1210200.0 484500.0 1211400.0 ;
      RECT  483300.0 1210200.0 484500.0 1211400.0 ;
      RECT  480900.0 1210200.0 482100.0 1211400.0 ;
      RECT  480600.0 1205250.0 479400.0 1206450.0 ;
      RECT  480900.0 1215600.0 482100.0 1216800.0 ;
      RECT  478500.0 1203000.0 479700.0 1204200.0 ;
      RECT  480900.0 1203000.0 482100.0 1204200.0 ;
      RECT  478500.0 1210200.0 479700.0 1211400.0 ;
      RECT  483300.0 1210200.0 484500.0 1211400.0 ;
      RECT  475500.0 1205400.0 485700.0 1206300.0 ;
      RECT  475500.0 1216500.0 485700.0 1217400.0 ;
      RECT  491100.0 1210200.0 492300.0 1217400.0 ;
      RECT  488700.0 1203000.0 489900.0 1204200.0 ;
      RECT  491100.0 1203000.0 492300.0 1204200.0 ;
      RECT  491100.0 1203000.0 492300.0 1204200.0 ;
      RECT  488700.0 1203000.0 489900.0 1204200.0 ;
      RECT  488700.0 1210200.0 489900.0 1211400.0 ;
      RECT  491100.0 1210200.0 492300.0 1211400.0 ;
      RECT  491100.0 1210200.0 492300.0 1211400.0 ;
      RECT  488700.0 1210200.0 489900.0 1211400.0 ;
      RECT  491100.0 1210200.0 492300.0 1211400.0 ;
      RECT  493500.0 1210200.0 494700.0 1211400.0 ;
      RECT  493500.0 1210200.0 494700.0 1211400.0 ;
      RECT  491100.0 1210200.0 492300.0 1211400.0 ;
      RECT  490800.0 1205250.0 489600.0 1206450.0 ;
      RECT  491100.0 1215600.0 492300.0 1216800.0 ;
      RECT  488700.0 1203000.0 489900.0 1204200.0 ;
      RECT  491100.0 1203000.0 492300.0 1204200.0 ;
      RECT  488700.0 1210200.0 489900.0 1211400.0 ;
      RECT  493500.0 1210200.0 494700.0 1211400.0 ;
      RECT  485700.0 1205400.0 495900.0 1206300.0 ;
      RECT  485700.0 1216500.0 495900.0 1217400.0 ;
      RECT  501300.0 1210200.0 502500.0 1217400.0 ;
      RECT  498900.0 1203000.0 500100.0 1204200.0 ;
      RECT  501300.0 1203000.0 502500.0 1204200.0 ;
      RECT  501300.0 1203000.0 502500.0 1204200.0 ;
      RECT  498900.0 1203000.0 500100.0 1204200.0 ;
      RECT  498900.0 1210200.0 500100.0 1211400.0 ;
      RECT  501300.0 1210200.0 502500.0 1211400.0 ;
      RECT  501300.0 1210200.0 502500.0 1211400.0 ;
      RECT  498900.0 1210200.0 500100.0 1211400.0 ;
      RECT  501300.0 1210200.0 502500.0 1211400.0 ;
      RECT  503700.0 1210200.0 504900.0 1211400.0 ;
      RECT  503700.0 1210200.0 504900.0 1211400.0 ;
      RECT  501300.0 1210200.0 502500.0 1211400.0 ;
      RECT  501000.0 1205250.0 499800.0 1206450.0 ;
      RECT  501300.0 1215600.0 502500.0 1216800.0 ;
      RECT  498900.0 1203000.0 500100.0 1204200.0 ;
      RECT  501300.0 1203000.0 502500.0 1204200.0 ;
      RECT  498900.0 1210200.0 500100.0 1211400.0 ;
      RECT  503700.0 1210200.0 504900.0 1211400.0 ;
      RECT  495900.0 1205400.0 506100.0 1206300.0 ;
      RECT  495900.0 1216500.0 506100.0 1217400.0 ;
      RECT  511500.0 1210200.0 512700.0 1217400.0 ;
      RECT  509100.0 1203000.0 510300.0 1204200.0 ;
      RECT  511500.0 1203000.0 512700.0 1204200.0 ;
      RECT  511500.0 1203000.0 512700.0 1204200.0 ;
      RECT  509100.0 1203000.0 510300.0 1204200.0 ;
      RECT  509100.0 1210200.0 510300.0 1211400.0 ;
      RECT  511500.0 1210200.0 512700.0 1211400.0 ;
      RECT  511500.0 1210200.0 512700.0 1211400.0 ;
      RECT  509100.0 1210200.0 510300.0 1211400.0 ;
      RECT  511500.0 1210200.0 512700.0 1211400.0 ;
      RECT  513900.0 1210200.0 515100.0 1211400.0 ;
      RECT  513900.0 1210200.0 515100.0 1211400.0 ;
      RECT  511500.0 1210200.0 512700.0 1211400.0 ;
      RECT  511200.0 1205250.0 510000.0 1206450.0 ;
      RECT  511500.0 1215600.0 512700.0 1216800.0 ;
      RECT  509100.0 1203000.0 510300.0 1204200.0 ;
      RECT  511500.0 1203000.0 512700.0 1204200.0 ;
      RECT  509100.0 1210200.0 510300.0 1211400.0 ;
      RECT  513900.0 1210200.0 515100.0 1211400.0 ;
      RECT  506100.0 1205400.0 516300.0 1206300.0 ;
      RECT  506100.0 1216500.0 516300.0 1217400.0 ;
      RECT  521700.0 1210200.0 522900.0 1217400.0 ;
      RECT  519300.0 1203000.0 520500.0 1204200.0 ;
      RECT  521700.0 1203000.0 522900.0 1204200.0 ;
      RECT  521700.0 1203000.0 522900.0 1204200.0 ;
      RECT  519300.0 1203000.0 520500.0 1204200.0 ;
      RECT  519300.0 1210200.0 520500.0 1211400.0 ;
      RECT  521700.0 1210200.0 522900.0 1211400.0 ;
      RECT  521700.0 1210200.0 522900.0 1211400.0 ;
      RECT  519300.0 1210200.0 520500.0 1211400.0 ;
      RECT  521700.0 1210200.0 522900.0 1211400.0 ;
      RECT  524100.0 1210200.0 525300.0 1211400.0 ;
      RECT  524100.0 1210200.0 525300.0 1211400.0 ;
      RECT  521700.0 1210200.0 522900.0 1211400.0 ;
      RECT  521400.0 1205250.0 520200.0 1206450.0 ;
      RECT  521700.0 1215600.0 522900.0 1216800.0 ;
      RECT  519300.0 1203000.0 520500.0 1204200.0 ;
      RECT  521700.0 1203000.0 522900.0 1204200.0 ;
      RECT  519300.0 1210200.0 520500.0 1211400.0 ;
      RECT  524100.0 1210200.0 525300.0 1211400.0 ;
      RECT  516300.0 1205400.0 526500.0 1206300.0 ;
      RECT  516300.0 1216500.0 526500.0 1217400.0 ;
      RECT  200100.0 1205400.0 526500.0 1206300.0 ;
      RECT  200100.0 1216500.0 526500.0 1217400.0 ;
      RECT  203100.0 277350.0 234900.0 278250.0 ;
      RECT  206100.0 275250.0 237900.0 276150.0 ;
      RECT  243900.0 277350.0 275700.0 278250.0 ;
      RECT  246900.0 275250.0 278700.0 276150.0 ;
      RECT  284700.0 277350.0 316500.0 278250.0 ;
      RECT  287700.0 275250.0 319500.0 276150.0 ;
      RECT  325500.0 277350.0 357300.0 278250.0 ;
      RECT  328500.0 275250.0 360300.0 276150.0 ;
      RECT  366300.0 277350.0 398100.0 278250.0 ;
      RECT  369300.0 275250.0 401100.0 276150.0 ;
      RECT  407100.0 277350.0 438900.0 278250.0 ;
      RECT  410100.0 275250.0 441900.0 276150.0 ;
      RECT  447900.0 277350.0 479700.0 278250.0 ;
      RECT  450900.0 275250.0 482700.0 276150.0 ;
      RECT  488700.0 277350.0 520500.0 278250.0 ;
      RECT  491700.0 275250.0 523500.0 276150.0 ;
      RECT  205950.0 311100.0 206850.0 312000.0 ;
      RECT  203100.0 311100.0 206400.0 312000.0 ;
      RECT  205950.0 304950.0 206850.0 311550.0 ;
      RECT  203550.0 289200.0 204450.0 290100.0 ;
      RECT  204000.0 289200.0 206550.0 290100.0 ;
      RECT  203550.0 289650.0 204450.0 294450.0 ;
      RECT  203400.0 293850.0 204600.0 295050.0 ;
      RECT  205800.0 293850.0 207000.0 295050.0 ;
      RECT  205800.0 293850.0 207000.0 295050.0 ;
      RECT  203400.0 293850.0 204600.0 295050.0 ;
      RECT  203400.0 304350.0 204600.0 305550.0 ;
      RECT  205800.0 304350.0 207000.0 305550.0 ;
      RECT  205800.0 304350.0 207000.0 305550.0 ;
      RECT  203400.0 304350.0 204600.0 305550.0 ;
      RECT  202950.0 310950.0 204150.0 312150.0 ;
      RECT  205950.0 289050.0 207150.0 290250.0 ;
      RECT  203400.0 304350.0 204600.0 305550.0 ;
      RECT  205800.0 293850.0 207000.0 295050.0 ;
      RECT  209700.0 292050.0 210900.0 293250.0 ;
      RECT  209700.0 292050.0 210900.0 293250.0 ;
      RECT  216150.0 311100.0 217050.0 312000.0 ;
      RECT  213300.0 311100.0 216600.0 312000.0 ;
      RECT  216150.0 304950.0 217050.0 311550.0 ;
      RECT  213750.0 289200.0 214650.0 290100.0 ;
      RECT  214200.0 289200.0 216750.0 290100.0 ;
      RECT  213750.0 289650.0 214650.0 294450.0 ;
      RECT  213600.0 293850.0 214800.0 295050.0 ;
      RECT  216000.0 293850.0 217200.0 295050.0 ;
      RECT  216000.0 293850.0 217200.0 295050.0 ;
      RECT  213600.0 293850.0 214800.0 295050.0 ;
      RECT  213600.0 304350.0 214800.0 305550.0 ;
      RECT  216000.0 304350.0 217200.0 305550.0 ;
      RECT  216000.0 304350.0 217200.0 305550.0 ;
      RECT  213600.0 304350.0 214800.0 305550.0 ;
      RECT  213150.0 310950.0 214350.0 312150.0 ;
      RECT  216150.0 289050.0 217350.0 290250.0 ;
      RECT  213600.0 304350.0 214800.0 305550.0 ;
      RECT  216000.0 293850.0 217200.0 295050.0 ;
      RECT  219900.0 292050.0 221100.0 293250.0 ;
      RECT  219900.0 292050.0 221100.0 293250.0 ;
      RECT  226350.0 311100.0 227250.0 312000.0 ;
      RECT  223500.0 311100.0 226800.0 312000.0 ;
      RECT  226350.0 304950.0 227250.0 311550.0 ;
      RECT  223950.0 289200.0 224850.0 290100.0 ;
      RECT  224400.0 289200.0 226950.0 290100.0 ;
      RECT  223950.0 289650.0 224850.0 294450.0 ;
      RECT  223800.0 293850.0 225000.0 295050.0 ;
      RECT  226200.0 293850.0 227400.0 295050.0 ;
      RECT  226200.0 293850.0 227400.0 295050.0 ;
      RECT  223800.0 293850.0 225000.0 295050.0 ;
      RECT  223800.0 304350.0 225000.0 305550.0 ;
      RECT  226200.0 304350.0 227400.0 305550.0 ;
      RECT  226200.0 304350.0 227400.0 305550.0 ;
      RECT  223800.0 304350.0 225000.0 305550.0 ;
      RECT  223350.0 310950.0 224550.0 312150.0 ;
      RECT  226350.0 289050.0 227550.0 290250.0 ;
      RECT  223800.0 304350.0 225000.0 305550.0 ;
      RECT  226200.0 293850.0 227400.0 295050.0 ;
      RECT  230100.0 292050.0 231300.0 293250.0 ;
      RECT  230100.0 292050.0 231300.0 293250.0 ;
      RECT  236550.0 311100.0 237450.0 312000.0 ;
      RECT  233700.0 311100.0 237000.0 312000.0 ;
      RECT  236550.0 304950.0 237450.0 311550.0 ;
      RECT  234150.0 289200.0 235050.0 290100.0 ;
      RECT  234600.0 289200.0 237150.0 290100.0 ;
      RECT  234150.0 289650.0 235050.0 294450.0 ;
      RECT  234000.0 293850.0 235200.0 295050.0 ;
      RECT  236400.0 293850.0 237600.0 295050.0 ;
      RECT  236400.0 293850.0 237600.0 295050.0 ;
      RECT  234000.0 293850.0 235200.0 295050.0 ;
      RECT  234000.0 304350.0 235200.0 305550.0 ;
      RECT  236400.0 304350.0 237600.0 305550.0 ;
      RECT  236400.0 304350.0 237600.0 305550.0 ;
      RECT  234000.0 304350.0 235200.0 305550.0 ;
      RECT  233550.0 310950.0 234750.0 312150.0 ;
      RECT  236550.0 289050.0 237750.0 290250.0 ;
      RECT  234000.0 304350.0 235200.0 305550.0 ;
      RECT  236400.0 293850.0 237600.0 295050.0 ;
      RECT  240300.0 292050.0 241500.0 293250.0 ;
      RECT  240300.0 292050.0 241500.0 293250.0 ;
      RECT  246750.0 311100.0 247650.0 312000.0 ;
      RECT  243900.0 311100.0 247200.0 312000.0 ;
      RECT  246750.0 304950.0 247650.0 311550.0 ;
      RECT  244350.0 289200.0 245250.0 290100.0 ;
      RECT  244800.0 289200.0 247350.0 290100.0 ;
      RECT  244350.0 289650.0 245250.0 294450.0 ;
      RECT  244200.0 293850.0 245400.0 295050.0 ;
      RECT  246600.0 293850.0 247800.0 295050.0 ;
      RECT  246600.0 293850.0 247800.0 295050.0 ;
      RECT  244200.0 293850.0 245400.0 295050.0 ;
      RECT  244200.0 304350.0 245400.0 305550.0 ;
      RECT  246600.0 304350.0 247800.0 305550.0 ;
      RECT  246600.0 304350.0 247800.0 305550.0 ;
      RECT  244200.0 304350.0 245400.0 305550.0 ;
      RECT  243750.0 310950.0 244950.0 312150.0 ;
      RECT  246750.0 289050.0 247950.0 290250.0 ;
      RECT  244200.0 304350.0 245400.0 305550.0 ;
      RECT  246600.0 293850.0 247800.0 295050.0 ;
      RECT  250500.0 292050.0 251700.0 293250.0 ;
      RECT  250500.0 292050.0 251700.0 293250.0 ;
      RECT  256950.0 311100.0 257850.0 312000.0 ;
      RECT  254100.0 311100.0 257400.0 312000.0 ;
      RECT  256950.0 304950.0 257850.0 311550.0 ;
      RECT  254550.0 289200.0 255450.0 290100.0 ;
      RECT  255000.0 289200.0 257550.0 290100.0 ;
      RECT  254550.0 289650.0 255450.0 294450.0 ;
      RECT  254400.0 293850.0 255600.0 295050.0 ;
      RECT  256800.0 293850.0 258000.0 295050.0 ;
      RECT  256800.0 293850.0 258000.0 295050.0 ;
      RECT  254400.0 293850.0 255600.0 295050.0 ;
      RECT  254400.0 304350.0 255600.0 305550.0 ;
      RECT  256800.0 304350.0 258000.0 305550.0 ;
      RECT  256800.0 304350.0 258000.0 305550.0 ;
      RECT  254400.0 304350.0 255600.0 305550.0 ;
      RECT  253950.0 310950.0 255150.0 312150.0 ;
      RECT  256950.0 289050.0 258150.0 290250.0 ;
      RECT  254400.0 304350.0 255600.0 305550.0 ;
      RECT  256800.0 293850.0 258000.0 295050.0 ;
      RECT  260700.0 292050.0 261900.0 293250.0 ;
      RECT  260700.0 292050.0 261900.0 293250.0 ;
      RECT  267150.0 311100.0 268050.0 312000.0 ;
      RECT  264300.0 311100.0 267600.0 312000.0 ;
      RECT  267150.0 304950.0 268050.0 311550.0 ;
      RECT  264750.0 289200.0 265650.0 290100.0 ;
      RECT  265200.0 289200.0 267750.0 290100.0 ;
      RECT  264750.0 289650.0 265650.0 294450.0 ;
      RECT  264600.0 293850.0 265800.0 295050.0 ;
      RECT  267000.0 293850.0 268200.0 295050.0 ;
      RECT  267000.0 293850.0 268200.0 295050.0 ;
      RECT  264600.0 293850.0 265800.0 295050.0 ;
      RECT  264600.0 304350.0 265800.0 305550.0 ;
      RECT  267000.0 304350.0 268200.0 305550.0 ;
      RECT  267000.0 304350.0 268200.0 305550.0 ;
      RECT  264600.0 304350.0 265800.0 305550.0 ;
      RECT  264150.0 310950.0 265350.0 312150.0 ;
      RECT  267150.0 289050.0 268350.0 290250.0 ;
      RECT  264600.0 304350.0 265800.0 305550.0 ;
      RECT  267000.0 293850.0 268200.0 295050.0 ;
      RECT  270900.0 292050.0 272100.0 293250.0 ;
      RECT  270900.0 292050.0 272100.0 293250.0 ;
      RECT  277350.0 311100.0 278250.0 312000.0 ;
      RECT  274500.0 311100.0 277800.0 312000.0 ;
      RECT  277350.0 304950.0 278250.0 311550.0 ;
      RECT  274950.0 289200.0 275850.0 290100.0 ;
      RECT  275400.0 289200.0 277950.0 290100.0 ;
      RECT  274950.0 289650.0 275850.0 294450.0 ;
      RECT  274800.0 293850.0 276000.0 295050.0 ;
      RECT  277200.0 293850.0 278400.0 295050.0 ;
      RECT  277200.0 293850.0 278400.0 295050.0 ;
      RECT  274800.0 293850.0 276000.0 295050.0 ;
      RECT  274800.0 304350.0 276000.0 305550.0 ;
      RECT  277200.0 304350.0 278400.0 305550.0 ;
      RECT  277200.0 304350.0 278400.0 305550.0 ;
      RECT  274800.0 304350.0 276000.0 305550.0 ;
      RECT  274350.0 310950.0 275550.0 312150.0 ;
      RECT  277350.0 289050.0 278550.0 290250.0 ;
      RECT  274800.0 304350.0 276000.0 305550.0 ;
      RECT  277200.0 293850.0 278400.0 295050.0 ;
      RECT  281100.0 292050.0 282300.0 293250.0 ;
      RECT  281100.0 292050.0 282300.0 293250.0 ;
      RECT  287550.0 311100.0 288450.0 312000.0 ;
      RECT  284700.0 311100.0 288000.0 312000.0 ;
      RECT  287550.0 304950.0 288450.0 311550.0 ;
      RECT  285150.0 289200.0 286050.0 290100.0 ;
      RECT  285600.0 289200.0 288150.0 290100.0 ;
      RECT  285150.0 289650.0 286050.0 294450.0 ;
      RECT  285000.0 293850.0 286200.0 295050.0 ;
      RECT  287400.0 293850.0 288600.0 295050.0 ;
      RECT  287400.0 293850.0 288600.0 295050.0 ;
      RECT  285000.0 293850.0 286200.0 295050.0 ;
      RECT  285000.0 304350.0 286200.0 305550.0 ;
      RECT  287400.0 304350.0 288600.0 305550.0 ;
      RECT  287400.0 304350.0 288600.0 305550.0 ;
      RECT  285000.0 304350.0 286200.0 305550.0 ;
      RECT  284550.0 310950.0 285750.0 312150.0 ;
      RECT  287550.0 289050.0 288750.0 290250.0 ;
      RECT  285000.0 304350.0 286200.0 305550.0 ;
      RECT  287400.0 293850.0 288600.0 295050.0 ;
      RECT  291300.0 292050.0 292500.0 293250.0 ;
      RECT  291300.0 292050.0 292500.0 293250.0 ;
      RECT  297750.0 311100.0 298650.0 312000.0 ;
      RECT  294900.0 311100.0 298200.0 312000.0 ;
      RECT  297750.0 304950.0 298650.0 311550.0 ;
      RECT  295350.0 289200.0 296250.0 290100.0 ;
      RECT  295800.0 289200.0 298350.0 290100.0 ;
      RECT  295350.0 289650.0 296250.0 294450.0 ;
      RECT  295200.0 293850.0 296400.0 295050.0 ;
      RECT  297600.0 293850.0 298800.0 295050.0 ;
      RECT  297600.0 293850.0 298800.0 295050.0 ;
      RECT  295200.0 293850.0 296400.0 295050.0 ;
      RECT  295200.0 304350.0 296400.0 305550.0 ;
      RECT  297600.0 304350.0 298800.0 305550.0 ;
      RECT  297600.0 304350.0 298800.0 305550.0 ;
      RECT  295200.0 304350.0 296400.0 305550.0 ;
      RECT  294750.0 310950.0 295950.0 312150.0 ;
      RECT  297750.0 289050.0 298950.0 290250.0 ;
      RECT  295200.0 304350.0 296400.0 305550.0 ;
      RECT  297600.0 293850.0 298800.0 295050.0 ;
      RECT  301500.0 292050.0 302700.0 293250.0 ;
      RECT  301500.0 292050.0 302700.0 293250.0 ;
      RECT  307950.0 311100.0 308850.0 312000.0 ;
      RECT  305100.0 311100.0 308400.0 312000.0 ;
      RECT  307950.0 304950.0 308850.0 311550.0 ;
      RECT  305550.0 289200.0 306450.0 290100.0 ;
      RECT  306000.0 289200.0 308550.0 290100.0 ;
      RECT  305550.0 289650.0 306450.0 294450.0 ;
      RECT  305400.0 293850.0 306600.0 295050.0 ;
      RECT  307800.0 293850.0 309000.0 295050.0 ;
      RECT  307800.0 293850.0 309000.0 295050.0 ;
      RECT  305400.0 293850.0 306600.0 295050.0 ;
      RECT  305400.0 304350.0 306600.0 305550.0 ;
      RECT  307800.0 304350.0 309000.0 305550.0 ;
      RECT  307800.0 304350.0 309000.0 305550.0 ;
      RECT  305400.0 304350.0 306600.0 305550.0 ;
      RECT  304950.0 310950.0 306150.0 312150.0 ;
      RECT  307950.0 289050.0 309150.0 290250.0 ;
      RECT  305400.0 304350.0 306600.0 305550.0 ;
      RECT  307800.0 293850.0 309000.0 295050.0 ;
      RECT  311700.0 292050.0 312900.0 293250.0 ;
      RECT  311700.0 292050.0 312900.0 293250.0 ;
      RECT  318150.0 311100.0 319050.0 312000.0 ;
      RECT  315300.0 311100.0 318600.0 312000.0 ;
      RECT  318150.0 304950.0 319050.0 311550.0 ;
      RECT  315750.0 289200.0 316650.0 290100.0 ;
      RECT  316200.0 289200.0 318750.0 290100.0 ;
      RECT  315750.0 289650.0 316650.0 294450.0 ;
      RECT  315600.0 293850.0 316800.0 295050.0 ;
      RECT  318000.0 293850.0 319200.0 295050.0 ;
      RECT  318000.0 293850.0 319200.0 295050.0 ;
      RECT  315600.0 293850.0 316800.0 295050.0 ;
      RECT  315600.0 304350.0 316800.0 305550.0 ;
      RECT  318000.0 304350.0 319200.0 305550.0 ;
      RECT  318000.0 304350.0 319200.0 305550.0 ;
      RECT  315600.0 304350.0 316800.0 305550.0 ;
      RECT  315150.0 310950.0 316350.0 312150.0 ;
      RECT  318150.0 289050.0 319350.0 290250.0 ;
      RECT  315600.0 304350.0 316800.0 305550.0 ;
      RECT  318000.0 293850.0 319200.0 295050.0 ;
      RECT  321900.0 292050.0 323100.0 293250.0 ;
      RECT  321900.0 292050.0 323100.0 293250.0 ;
      RECT  328350.0 311100.0 329250.0 312000.0 ;
      RECT  325500.0 311100.0 328800.0 312000.0 ;
      RECT  328350.0 304950.0 329250.0 311550.0 ;
      RECT  325950.0 289200.0 326850.0 290100.0 ;
      RECT  326400.0 289200.0 328950.0 290100.0 ;
      RECT  325950.0 289650.0 326850.0 294450.0 ;
      RECT  325800.0 293850.0 327000.0 295050.0 ;
      RECT  328200.0 293850.0 329400.0 295050.0 ;
      RECT  328200.0 293850.0 329400.0 295050.0 ;
      RECT  325800.0 293850.0 327000.0 295050.0 ;
      RECT  325800.0 304350.0 327000.0 305550.0 ;
      RECT  328200.0 304350.0 329400.0 305550.0 ;
      RECT  328200.0 304350.0 329400.0 305550.0 ;
      RECT  325800.0 304350.0 327000.0 305550.0 ;
      RECT  325350.0 310950.0 326550.0 312150.0 ;
      RECT  328350.0 289050.0 329550.0 290250.0 ;
      RECT  325800.0 304350.0 327000.0 305550.0 ;
      RECT  328200.0 293850.0 329400.0 295050.0 ;
      RECT  332100.0 292050.0 333300.0 293250.0 ;
      RECT  332100.0 292050.0 333300.0 293250.0 ;
      RECT  338550.0 311100.0 339450.0 312000.0 ;
      RECT  335700.0 311100.0 339000.0 312000.0 ;
      RECT  338550.0 304950.0 339450.0 311550.0 ;
      RECT  336150.0 289200.0 337050.0 290100.0 ;
      RECT  336600.0 289200.0 339150.0 290100.0 ;
      RECT  336150.0 289650.0 337050.0 294450.0 ;
      RECT  336000.0 293850.0 337200.0 295050.0 ;
      RECT  338400.0 293850.0 339600.0 295050.0 ;
      RECT  338400.0 293850.0 339600.0 295050.0 ;
      RECT  336000.0 293850.0 337200.0 295050.0 ;
      RECT  336000.0 304350.0 337200.0 305550.0 ;
      RECT  338400.0 304350.0 339600.0 305550.0 ;
      RECT  338400.0 304350.0 339600.0 305550.0 ;
      RECT  336000.0 304350.0 337200.0 305550.0 ;
      RECT  335550.0 310950.0 336750.0 312150.0 ;
      RECT  338550.0 289050.0 339750.0 290250.0 ;
      RECT  336000.0 304350.0 337200.0 305550.0 ;
      RECT  338400.0 293850.0 339600.0 295050.0 ;
      RECT  342300.0 292050.0 343500.0 293250.0 ;
      RECT  342300.0 292050.0 343500.0 293250.0 ;
      RECT  348750.0 311100.0 349650.0 312000.0 ;
      RECT  345900.0 311100.0 349200.0 312000.0 ;
      RECT  348750.0 304950.0 349650.0 311550.0 ;
      RECT  346350.0 289200.0 347250.0 290100.0 ;
      RECT  346800.0 289200.0 349350.0 290100.0 ;
      RECT  346350.0 289650.0 347250.0 294450.0 ;
      RECT  346200.0 293850.0 347400.0 295050.0 ;
      RECT  348600.0 293850.0 349800.0 295050.0 ;
      RECT  348600.0 293850.0 349800.0 295050.0 ;
      RECT  346200.0 293850.0 347400.0 295050.0 ;
      RECT  346200.0 304350.0 347400.0 305550.0 ;
      RECT  348600.0 304350.0 349800.0 305550.0 ;
      RECT  348600.0 304350.0 349800.0 305550.0 ;
      RECT  346200.0 304350.0 347400.0 305550.0 ;
      RECT  345750.0 310950.0 346950.0 312150.0 ;
      RECT  348750.0 289050.0 349950.0 290250.0 ;
      RECT  346200.0 304350.0 347400.0 305550.0 ;
      RECT  348600.0 293850.0 349800.0 295050.0 ;
      RECT  352500.0 292050.0 353700.0 293250.0 ;
      RECT  352500.0 292050.0 353700.0 293250.0 ;
      RECT  358950.0 311100.0 359850.0 312000.0 ;
      RECT  356100.0 311100.0 359400.0 312000.0 ;
      RECT  358950.0 304950.0 359850.0 311550.0 ;
      RECT  356550.0 289200.0 357450.0 290100.0 ;
      RECT  357000.0 289200.0 359550.0 290100.0 ;
      RECT  356550.0 289650.0 357450.0 294450.0 ;
      RECT  356400.0 293850.0 357600.0 295050.0 ;
      RECT  358800.0 293850.0 360000.0 295050.0 ;
      RECT  358800.0 293850.0 360000.0 295050.0 ;
      RECT  356400.0 293850.0 357600.0 295050.0 ;
      RECT  356400.0 304350.0 357600.0 305550.0 ;
      RECT  358800.0 304350.0 360000.0 305550.0 ;
      RECT  358800.0 304350.0 360000.0 305550.0 ;
      RECT  356400.0 304350.0 357600.0 305550.0 ;
      RECT  355950.0 310950.0 357150.0 312150.0 ;
      RECT  358950.0 289050.0 360150.0 290250.0 ;
      RECT  356400.0 304350.0 357600.0 305550.0 ;
      RECT  358800.0 293850.0 360000.0 295050.0 ;
      RECT  362700.0 292050.0 363900.0 293250.0 ;
      RECT  362700.0 292050.0 363900.0 293250.0 ;
      RECT  369150.0 311100.0 370050.0 312000.0 ;
      RECT  366300.0 311100.0 369600.0 312000.0 ;
      RECT  369150.0 304950.0 370050.0 311550.0 ;
      RECT  366750.0 289200.0 367650.0 290100.0 ;
      RECT  367200.0 289200.0 369750.0 290100.0 ;
      RECT  366750.0 289650.0 367650.0 294450.0 ;
      RECT  366600.0 293850.0 367800.0 295050.0 ;
      RECT  369000.0 293850.0 370200.0 295050.0 ;
      RECT  369000.0 293850.0 370200.0 295050.0 ;
      RECT  366600.0 293850.0 367800.0 295050.0 ;
      RECT  366600.0 304350.0 367800.0 305550.0 ;
      RECT  369000.0 304350.0 370200.0 305550.0 ;
      RECT  369000.0 304350.0 370200.0 305550.0 ;
      RECT  366600.0 304350.0 367800.0 305550.0 ;
      RECT  366150.0 310950.0 367350.0 312150.0 ;
      RECT  369150.0 289050.0 370350.0 290250.0 ;
      RECT  366600.0 304350.0 367800.0 305550.0 ;
      RECT  369000.0 293850.0 370200.0 295050.0 ;
      RECT  372900.0 292050.0 374100.0 293250.0 ;
      RECT  372900.0 292050.0 374100.0 293250.0 ;
      RECT  379350.0 311100.0 380250.0 312000.0 ;
      RECT  376500.0 311100.0 379800.0 312000.0 ;
      RECT  379350.0 304950.0 380250.0 311550.0 ;
      RECT  376950.0 289200.0 377850.0 290100.0 ;
      RECT  377400.0 289200.0 379950.0 290100.0 ;
      RECT  376950.0 289650.0 377850.0 294450.0 ;
      RECT  376800.0 293850.0 378000.0 295050.0 ;
      RECT  379200.0 293850.0 380400.0 295050.0 ;
      RECT  379200.0 293850.0 380400.0 295050.0 ;
      RECT  376800.0 293850.0 378000.0 295050.0 ;
      RECT  376800.0 304350.0 378000.0 305550.0 ;
      RECT  379200.0 304350.0 380400.0 305550.0 ;
      RECT  379200.0 304350.0 380400.0 305550.0 ;
      RECT  376800.0 304350.0 378000.0 305550.0 ;
      RECT  376350.0 310950.0 377550.0 312150.0 ;
      RECT  379350.0 289050.0 380550.0 290250.0 ;
      RECT  376800.0 304350.0 378000.0 305550.0 ;
      RECT  379200.0 293850.0 380400.0 295050.0 ;
      RECT  383100.0 292050.0 384300.0 293250.0 ;
      RECT  383100.0 292050.0 384300.0 293250.0 ;
      RECT  389550.0 311100.0 390450.0 312000.0 ;
      RECT  386700.0 311100.0 390000.0 312000.0 ;
      RECT  389550.0 304950.0 390450.0 311550.0 ;
      RECT  387150.0 289200.0 388050.0 290100.0 ;
      RECT  387600.0 289200.0 390150.0 290100.0 ;
      RECT  387150.0 289650.0 388050.0 294450.0 ;
      RECT  387000.0 293850.0 388200.0 295050.0 ;
      RECT  389400.0 293850.0 390600.0 295050.0 ;
      RECT  389400.0 293850.0 390600.0 295050.0 ;
      RECT  387000.0 293850.0 388200.0 295050.0 ;
      RECT  387000.0 304350.0 388200.0 305550.0 ;
      RECT  389400.0 304350.0 390600.0 305550.0 ;
      RECT  389400.0 304350.0 390600.0 305550.0 ;
      RECT  387000.0 304350.0 388200.0 305550.0 ;
      RECT  386550.0 310950.0 387750.0 312150.0 ;
      RECT  389550.0 289050.0 390750.0 290250.0 ;
      RECT  387000.0 304350.0 388200.0 305550.0 ;
      RECT  389400.0 293850.0 390600.0 295050.0 ;
      RECT  393300.0 292050.0 394500.0 293250.0 ;
      RECT  393300.0 292050.0 394500.0 293250.0 ;
      RECT  399750.0 311100.0 400650.0 312000.0 ;
      RECT  396900.0 311100.0 400200.0 312000.0 ;
      RECT  399750.0 304950.0 400650.0 311550.0 ;
      RECT  397350.0 289200.0 398250.0 290100.0 ;
      RECT  397800.0 289200.0 400350.0 290100.0 ;
      RECT  397350.0 289650.0 398250.0 294450.0 ;
      RECT  397200.0 293850.0 398400.0 295050.0 ;
      RECT  399600.0 293850.0 400800.0 295050.0 ;
      RECT  399600.0 293850.0 400800.0 295050.0 ;
      RECT  397200.0 293850.0 398400.0 295050.0 ;
      RECT  397200.0 304350.0 398400.0 305550.0 ;
      RECT  399600.0 304350.0 400800.0 305550.0 ;
      RECT  399600.0 304350.0 400800.0 305550.0 ;
      RECT  397200.0 304350.0 398400.0 305550.0 ;
      RECT  396750.0 310950.0 397950.0 312150.0 ;
      RECT  399750.0 289050.0 400950.0 290250.0 ;
      RECT  397200.0 304350.0 398400.0 305550.0 ;
      RECT  399600.0 293850.0 400800.0 295050.0 ;
      RECT  403500.0 292050.0 404700.0 293250.0 ;
      RECT  403500.0 292050.0 404700.0 293250.0 ;
      RECT  409950.0 311100.0 410850.0 312000.0 ;
      RECT  407100.0 311100.0 410400.0 312000.0 ;
      RECT  409950.0 304950.0 410850.0 311550.0 ;
      RECT  407550.0 289200.0 408450.0 290100.0 ;
      RECT  408000.0 289200.0 410550.0 290100.0 ;
      RECT  407550.0 289650.0 408450.0 294450.0 ;
      RECT  407400.0 293850.0 408600.0 295050.0 ;
      RECT  409800.0 293850.0 411000.0 295050.0 ;
      RECT  409800.0 293850.0 411000.0 295050.0 ;
      RECT  407400.0 293850.0 408600.0 295050.0 ;
      RECT  407400.0 304350.0 408600.0 305550.0 ;
      RECT  409800.0 304350.0 411000.0 305550.0 ;
      RECT  409800.0 304350.0 411000.0 305550.0 ;
      RECT  407400.0 304350.0 408600.0 305550.0 ;
      RECT  406950.0 310950.0 408150.0 312150.0 ;
      RECT  409950.0 289050.0 411150.0 290250.0 ;
      RECT  407400.0 304350.0 408600.0 305550.0 ;
      RECT  409800.0 293850.0 411000.0 295050.0 ;
      RECT  413700.0 292050.0 414900.0 293250.0 ;
      RECT  413700.0 292050.0 414900.0 293250.0 ;
      RECT  420150.0 311100.0 421050.0 312000.0 ;
      RECT  417300.0 311100.0 420600.0 312000.0 ;
      RECT  420150.0 304950.0 421050.0 311550.0 ;
      RECT  417750.0 289200.0 418650.0 290100.0 ;
      RECT  418200.0 289200.0 420750.0 290100.0 ;
      RECT  417750.0 289650.0 418650.0 294450.0 ;
      RECT  417600.0 293850.0 418800.0 295050.0 ;
      RECT  420000.0 293850.0 421200.0 295050.0 ;
      RECT  420000.0 293850.0 421200.0 295050.0 ;
      RECT  417600.0 293850.0 418800.0 295050.0 ;
      RECT  417600.0 304350.0 418800.0 305550.0 ;
      RECT  420000.0 304350.0 421200.0 305550.0 ;
      RECT  420000.0 304350.0 421200.0 305550.0 ;
      RECT  417600.0 304350.0 418800.0 305550.0 ;
      RECT  417150.0 310950.0 418350.0 312150.0 ;
      RECT  420150.0 289050.0 421350.0 290250.0 ;
      RECT  417600.0 304350.0 418800.0 305550.0 ;
      RECT  420000.0 293850.0 421200.0 295050.0 ;
      RECT  423900.0 292050.0 425100.0 293250.0 ;
      RECT  423900.0 292050.0 425100.0 293250.0 ;
      RECT  430350.0 311100.0 431250.0 312000.0 ;
      RECT  427500.0 311100.0 430800.0 312000.0 ;
      RECT  430350.0 304950.0 431250.0 311550.0 ;
      RECT  427950.0 289200.0 428850.0 290100.0 ;
      RECT  428400.0 289200.0 430950.0 290100.0 ;
      RECT  427950.0 289650.0 428850.0 294450.0 ;
      RECT  427800.0 293850.0 429000.0 295050.0 ;
      RECT  430200.0 293850.0 431400.0 295050.0 ;
      RECT  430200.0 293850.0 431400.0 295050.0 ;
      RECT  427800.0 293850.0 429000.0 295050.0 ;
      RECT  427800.0 304350.0 429000.0 305550.0 ;
      RECT  430200.0 304350.0 431400.0 305550.0 ;
      RECT  430200.0 304350.0 431400.0 305550.0 ;
      RECT  427800.0 304350.0 429000.0 305550.0 ;
      RECT  427350.0 310950.0 428550.0 312150.0 ;
      RECT  430350.0 289050.0 431550.0 290250.0 ;
      RECT  427800.0 304350.0 429000.0 305550.0 ;
      RECT  430200.0 293850.0 431400.0 295050.0 ;
      RECT  434100.0 292050.0 435300.0 293250.0 ;
      RECT  434100.0 292050.0 435300.0 293250.0 ;
      RECT  440550.0 311100.0 441450.0 312000.0 ;
      RECT  437700.0 311100.0 441000.0 312000.0 ;
      RECT  440550.0 304950.0 441450.0 311550.0 ;
      RECT  438150.0 289200.0 439050.0 290100.0 ;
      RECT  438600.0 289200.0 441150.0 290100.0 ;
      RECT  438150.0 289650.0 439050.0 294450.0 ;
      RECT  438000.0 293850.0 439200.0 295050.0 ;
      RECT  440400.0 293850.0 441600.0 295050.0 ;
      RECT  440400.0 293850.0 441600.0 295050.0 ;
      RECT  438000.0 293850.0 439200.0 295050.0 ;
      RECT  438000.0 304350.0 439200.0 305550.0 ;
      RECT  440400.0 304350.0 441600.0 305550.0 ;
      RECT  440400.0 304350.0 441600.0 305550.0 ;
      RECT  438000.0 304350.0 439200.0 305550.0 ;
      RECT  437550.0 310950.0 438750.0 312150.0 ;
      RECT  440550.0 289050.0 441750.0 290250.0 ;
      RECT  438000.0 304350.0 439200.0 305550.0 ;
      RECT  440400.0 293850.0 441600.0 295050.0 ;
      RECT  444300.0 292050.0 445500.0 293250.0 ;
      RECT  444300.0 292050.0 445500.0 293250.0 ;
      RECT  450750.0 311100.0 451650.0 312000.0 ;
      RECT  447900.0 311100.0 451200.0 312000.0 ;
      RECT  450750.0 304950.0 451650.0 311550.0 ;
      RECT  448350.0 289200.0 449250.0 290100.0 ;
      RECT  448800.0 289200.0 451350.0 290100.0 ;
      RECT  448350.0 289650.0 449250.0 294450.0 ;
      RECT  448200.0 293850.0 449400.0 295050.0 ;
      RECT  450600.0 293850.0 451800.0 295050.0 ;
      RECT  450600.0 293850.0 451800.0 295050.0 ;
      RECT  448200.0 293850.0 449400.0 295050.0 ;
      RECT  448200.0 304350.0 449400.0 305550.0 ;
      RECT  450600.0 304350.0 451800.0 305550.0 ;
      RECT  450600.0 304350.0 451800.0 305550.0 ;
      RECT  448200.0 304350.0 449400.0 305550.0 ;
      RECT  447750.0 310950.0 448950.0 312150.0 ;
      RECT  450750.0 289050.0 451950.0 290250.0 ;
      RECT  448200.0 304350.0 449400.0 305550.0 ;
      RECT  450600.0 293850.0 451800.0 295050.0 ;
      RECT  454500.0 292050.0 455700.0 293250.0 ;
      RECT  454500.0 292050.0 455700.0 293250.0 ;
      RECT  460950.0 311100.0 461850.0 312000.0 ;
      RECT  458100.0 311100.0 461400.0 312000.0 ;
      RECT  460950.0 304950.0 461850.0 311550.0 ;
      RECT  458550.0 289200.0 459450.0 290100.0 ;
      RECT  459000.0 289200.0 461550.0 290100.0 ;
      RECT  458550.0 289650.0 459450.0 294450.0 ;
      RECT  458400.0 293850.0 459600.0 295050.0 ;
      RECT  460800.0 293850.0 462000.0 295050.0 ;
      RECT  460800.0 293850.0 462000.0 295050.0 ;
      RECT  458400.0 293850.0 459600.0 295050.0 ;
      RECT  458400.0 304350.0 459600.0 305550.0 ;
      RECT  460800.0 304350.0 462000.0 305550.0 ;
      RECT  460800.0 304350.0 462000.0 305550.0 ;
      RECT  458400.0 304350.0 459600.0 305550.0 ;
      RECT  457950.0 310950.0 459150.0 312150.0 ;
      RECT  460950.0 289050.0 462150.0 290250.0 ;
      RECT  458400.0 304350.0 459600.0 305550.0 ;
      RECT  460800.0 293850.0 462000.0 295050.0 ;
      RECT  464700.0 292050.0 465900.0 293250.0 ;
      RECT  464700.0 292050.0 465900.0 293250.0 ;
      RECT  471150.0 311100.0 472050.0 312000.0 ;
      RECT  468300.0 311100.0 471600.0 312000.0 ;
      RECT  471150.0 304950.0 472050.0 311550.0 ;
      RECT  468750.0 289200.0 469650.0 290100.0 ;
      RECT  469200.0 289200.0 471750.0 290100.0 ;
      RECT  468750.0 289650.0 469650.0 294450.0 ;
      RECT  468600.0 293850.0 469800.0 295050.0 ;
      RECT  471000.0 293850.0 472200.0 295050.0 ;
      RECT  471000.0 293850.0 472200.0 295050.0 ;
      RECT  468600.0 293850.0 469800.0 295050.0 ;
      RECT  468600.0 304350.0 469800.0 305550.0 ;
      RECT  471000.0 304350.0 472200.0 305550.0 ;
      RECT  471000.0 304350.0 472200.0 305550.0 ;
      RECT  468600.0 304350.0 469800.0 305550.0 ;
      RECT  468150.0 310950.0 469350.0 312150.0 ;
      RECT  471150.0 289050.0 472350.0 290250.0 ;
      RECT  468600.0 304350.0 469800.0 305550.0 ;
      RECT  471000.0 293850.0 472200.0 295050.0 ;
      RECT  474900.0 292050.0 476100.0 293250.0 ;
      RECT  474900.0 292050.0 476100.0 293250.0 ;
      RECT  481350.0 311100.0 482250.0 312000.0 ;
      RECT  478500.0 311100.0 481800.0 312000.0 ;
      RECT  481350.0 304950.0 482250.0 311550.0 ;
      RECT  478950.0 289200.0 479850.0 290100.0 ;
      RECT  479400.0 289200.0 481950.0 290100.0 ;
      RECT  478950.0 289650.0 479850.0 294450.0 ;
      RECT  478800.0 293850.0 480000.0 295050.0 ;
      RECT  481200.0 293850.0 482400.0 295050.0 ;
      RECT  481200.0 293850.0 482400.0 295050.0 ;
      RECT  478800.0 293850.0 480000.0 295050.0 ;
      RECT  478800.0 304350.0 480000.0 305550.0 ;
      RECT  481200.0 304350.0 482400.0 305550.0 ;
      RECT  481200.0 304350.0 482400.0 305550.0 ;
      RECT  478800.0 304350.0 480000.0 305550.0 ;
      RECT  478350.0 310950.0 479550.0 312150.0 ;
      RECT  481350.0 289050.0 482550.0 290250.0 ;
      RECT  478800.0 304350.0 480000.0 305550.0 ;
      RECT  481200.0 293850.0 482400.0 295050.0 ;
      RECT  485100.0 292050.0 486300.0 293250.0 ;
      RECT  485100.0 292050.0 486300.0 293250.0 ;
      RECT  491550.0 311100.0 492450.0 312000.0 ;
      RECT  488700.0 311100.0 492000.0 312000.0 ;
      RECT  491550.0 304950.0 492450.0 311550.0 ;
      RECT  489150.0 289200.0 490050.0 290100.0 ;
      RECT  489600.0 289200.0 492150.0 290100.0 ;
      RECT  489150.0 289650.0 490050.0 294450.0 ;
      RECT  489000.0 293850.0 490200.0 295050.0 ;
      RECT  491400.0 293850.0 492600.0 295050.0 ;
      RECT  491400.0 293850.0 492600.0 295050.0 ;
      RECT  489000.0 293850.0 490200.0 295050.0 ;
      RECT  489000.0 304350.0 490200.0 305550.0 ;
      RECT  491400.0 304350.0 492600.0 305550.0 ;
      RECT  491400.0 304350.0 492600.0 305550.0 ;
      RECT  489000.0 304350.0 490200.0 305550.0 ;
      RECT  488550.0 310950.0 489750.0 312150.0 ;
      RECT  491550.0 289050.0 492750.0 290250.0 ;
      RECT  489000.0 304350.0 490200.0 305550.0 ;
      RECT  491400.0 293850.0 492600.0 295050.0 ;
      RECT  495300.0 292050.0 496500.0 293250.0 ;
      RECT  495300.0 292050.0 496500.0 293250.0 ;
      RECT  501750.0 311100.0 502650.0 312000.0 ;
      RECT  498900.0 311100.0 502200.0 312000.0 ;
      RECT  501750.0 304950.0 502650.0 311550.0 ;
      RECT  499350.0 289200.0 500250.0 290100.0 ;
      RECT  499800.0 289200.0 502350.0 290100.0 ;
      RECT  499350.0 289650.0 500250.0 294450.0 ;
      RECT  499200.0 293850.0 500400.0 295050.0 ;
      RECT  501600.0 293850.0 502800.0 295050.0 ;
      RECT  501600.0 293850.0 502800.0 295050.0 ;
      RECT  499200.0 293850.0 500400.0 295050.0 ;
      RECT  499200.0 304350.0 500400.0 305550.0 ;
      RECT  501600.0 304350.0 502800.0 305550.0 ;
      RECT  501600.0 304350.0 502800.0 305550.0 ;
      RECT  499200.0 304350.0 500400.0 305550.0 ;
      RECT  498750.0 310950.0 499950.0 312150.0 ;
      RECT  501750.0 289050.0 502950.0 290250.0 ;
      RECT  499200.0 304350.0 500400.0 305550.0 ;
      RECT  501600.0 293850.0 502800.0 295050.0 ;
      RECT  505500.0 292050.0 506700.0 293250.0 ;
      RECT  505500.0 292050.0 506700.0 293250.0 ;
      RECT  511950.0 311100.0 512850.0 312000.0 ;
      RECT  509100.0 311100.0 512400.0 312000.0 ;
      RECT  511950.0 304950.0 512850.0 311550.0 ;
      RECT  509550.0 289200.0 510450.0 290100.0 ;
      RECT  510000.0 289200.0 512550.0 290100.0 ;
      RECT  509550.0 289650.0 510450.0 294450.0 ;
      RECT  509400.0 293850.0 510600.0 295050.0 ;
      RECT  511800.0 293850.0 513000.0 295050.0 ;
      RECT  511800.0 293850.0 513000.0 295050.0 ;
      RECT  509400.0 293850.0 510600.0 295050.0 ;
      RECT  509400.0 304350.0 510600.0 305550.0 ;
      RECT  511800.0 304350.0 513000.0 305550.0 ;
      RECT  511800.0 304350.0 513000.0 305550.0 ;
      RECT  509400.0 304350.0 510600.0 305550.0 ;
      RECT  508950.0 310950.0 510150.0 312150.0 ;
      RECT  511950.0 289050.0 513150.0 290250.0 ;
      RECT  509400.0 304350.0 510600.0 305550.0 ;
      RECT  511800.0 293850.0 513000.0 295050.0 ;
      RECT  515700.0 292050.0 516900.0 293250.0 ;
      RECT  515700.0 292050.0 516900.0 293250.0 ;
      RECT  522150.0 311100.0 523050.0 312000.0 ;
      RECT  519300.0 311100.0 522600.0 312000.0 ;
      RECT  522150.0 304950.0 523050.0 311550.0 ;
      RECT  519750.0 289200.0 520650.0 290100.0 ;
      RECT  520200.0 289200.0 522750.0 290100.0 ;
      RECT  519750.0 289650.0 520650.0 294450.0 ;
      RECT  519600.0 293850.0 520800.0 295050.0 ;
      RECT  522000.0 293850.0 523200.0 295050.0 ;
      RECT  522000.0 293850.0 523200.0 295050.0 ;
      RECT  519600.0 293850.0 520800.0 295050.0 ;
      RECT  519600.0 304350.0 520800.0 305550.0 ;
      RECT  522000.0 304350.0 523200.0 305550.0 ;
      RECT  522000.0 304350.0 523200.0 305550.0 ;
      RECT  519600.0 304350.0 520800.0 305550.0 ;
      RECT  519150.0 310950.0 520350.0 312150.0 ;
      RECT  522150.0 289050.0 523350.0 290250.0 ;
      RECT  519600.0 304350.0 520800.0 305550.0 ;
      RECT  522000.0 293850.0 523200.0 295050.0 ;
      RECT  525900.0 292050.0 527100.0 293250.0 ;
      RECT  525900.0 292050.0 527100.0 293250.0 ;
      RECT  205800.0 285750.0 204600.0 286950.0 ;
      RECT  216000.0 283650.0 214800.0 284850.0 ;
      RECT  226200.0 281550.0 225000.0 282750.0 ;
      RECT  236400.0 279450.0 235200.0 280650.0 ;
      RECT  246600.0 285750.0 245400.0 286950.0 ;
      RECT  256800.0 283650.0 255600.0 284850.0 ;
      RECT  267000.0 281550.0 265800.0 282750.0 ;
      RECT  277200.0 279450.0 276000.0 280650.0 ;
      RECT  287400.0 285750.0 286200.0 286950.0 ;
      RECT  297600.0 283650.0 296400.0 284850.0 ;
      RECT  307800.0 281550.0 306600.0 282750.0 ;
      RECT  318000.0 279450.0 316800.0 280650.0 ;
      RECT  328200.0 285750.0 327000.0 286950.0 ;
      RECT  338400.0 283650.0 337200.0 284850.0 ;
      RECT  348600.0 281550.0 347400.0 282750.0 ;
      RECT  358800.0 279450.0 357600.0 280650.0 ;
      RECT  369000.0 285750.0 367800.0 286950.0 ;
      RECT  379200.0 283650.0 378000.0 284850.0 ;
      RECT  389400.0 281550.0 388200.0 282750.0 ;
      RECT  399600.0 279450.0 398400.0 280650.0 ;
      RECT  409800.0 285750.0 408600.0 286950.0 ;
      RECT  420000.0 283650.0 418800.0 284850.0 ;
      RECT  430200.0 281550.0 429000.0 282750.0 ;
      RECT  440400.0 279450.0 439200.0 280650.0 ;
      RECT  450600.0 285750.0 449400.0 286950.0 ;
      RECT  460800.0 283650.0 459600.0 284850.0 ;
      RECT  471000.0 281550.0 469800.0 282750.0 ;
      RECT  481200.0 279450.0 480000.0 280650.0 ;
      RECT  491400.0 285750.0 490200.0 286950.0 ;
      RECT  501600.0 283650.0 500400.0 284850.0 ;
      RECT  511800.0 281550.0 510600.0 282750.0 ;
      RECT  522000.0 279450.0 520800.0 280650.0 ;
      RECT  204300.0 277350.0 203100.0 278550.0 ;
      RECT  206100.0 275250.0 204900.0 276450.0 ;
      RECT  214500.0 277350.0 213300.0 278550.0 ;
      RECT  216300.0 275250.0 215100.0 276450.0 ;
      RECT  224700.0 277350.0 223500.0 278550.0 ;
      RECT  226500.0 275250.0 225300.0 276450.0 ;
      RECT  234900.0 277350.0 233700.0 278550.0 ;
      RECT  236700.0 275250.0 235500.0 276450.0 ;
      RECT  245100.0 277350.0 243900.0 278550.0 ;
      RECT  246900.0 275250.0 245700.0 276450.0 ;
      RECT  255300.0 277350.0 254100.0 278550.0 ;
      RECT  257100.0 275250.0 255900.0 276450.0 ;
      RECT  265500.0 277350.0 264300.0 278550.0 ;
      RECT  267300.0 275250.0 266100.0 276450.0 ;
      RECT  275700.0 277350.0 274500.0 278550.0 ;
      RECT  277500.0 275250.0 276300.0 276450.0 ;
      RECT  285900.0 277350.0 284700.0 278550.0 ;
      RECT  287700.0 275250.0 286500.0 276450.0 ;
      RECT  296100.0 277350.0 294900.0 278550.0 ;
      RECT  297900.0 275250.0 296700.0 276450.0 ;
      RECT  306300.0 277350.0 305100.0 278550.0 ;
      RECT  308100.0 275250.0 306900.0 276450.0 ;
      RECT  316500.0 277350.0 315300.0 278550.0 ;
      RECT  318300.0 275250.0 317100.0 276450.0 ;
      RECT  326700.0 277350.0 325500.0 278550.0 ;
      RECT  328500.0 275250.0 327300.0 276450.0 ;
      RECT  336900.0 277350.0 335700.0 278550.0 ;
      RECT  338700.0 275250.0 337500.0 276450.0 ;
      RECT  347100.0 277350.0 345900.0 278550.0 ;
      RECT  348900.0 275250.0 347700.0 276450.0 ;
      RECT  357300.0 277350.0 356100.0 278550.0 ;
      RECT  359100.0 275250.0 357900.0 276450.0 ;
      RECT  367500.0 277350.0 366300.0 278550.0 ;
      RECT  369300.0 275250.0 368100.0 276450.0 ;
      RECT  377700.0 277350.0 376500.0 278550.0 ;
      RECT  379500.0 275250.0 378300.0 276450.0 ;
      RECT  387900.0 277350.0 386700.0 278550.0 ;
      RECT  389700.0 275250.0 388500.0 276450.0 ;
      RECT  398100.0 277350.0 396900.0 278550.0 ;
      RECT  399900.0 275250.0 398700.0 276450.0 ;
      RECT  408300.0 277350.0 407100.0 278550.0 ;
      RECT  410100.0 275250.0 408900.0 276450.0 ;
      RECT  418500.0 277350.0 417300.0 278550.0 ;
      RECT  420300.0 275250.0 419100.0 276450.0 ;
      RECT  428700.0 277350.0 427500.0 278550.0 ;
      RECT  430500.0 275250.0 429300.0 276450.0 ;
      RECT  438900.0 277350.0 437700.0 278550.0 ;
      RECT  440700.0 275250.0 439500.0 276450.0 ;
      RECT  449100.0 277350.0 447900.0 278550.0 ;
      RECT  450900.0 275250.0 449700.0 276450.0 ;
      RECT  459300.0 277350.0 458100.0 278550.0 ;
      RECT  461100.0 275250.0 459900.0 276450.0 ;
      RECT  469500.0 277350.0 468300.0 278550.0 ;
      RECT  471300.0 275250.0 470100.0 276450.0 ;
      RECT  479700.0 277350.0 478500.0 278550.0 ;
      RECT  481500.0 275250.0 480300.0 276450.0 ;
      RECT  489900.0 277350.0 488700.0 278550.0 ;
      RECT  491700.0 275250.0 490500.0 276450.0 ;
      RECT  500100.0 277350.0 498900.0 278550.0 ;
      RECT  501900.0 275250.0 500700.0 276450.0 ;
      RECT  510300.0 277350.0 509100.0 278550.0 ;
      RECT  512100.0 275250.0 510900.0 276450.0 ;
      RECT  520500.0 277350.0 519300.0 278550.0 ;
      RECT  522300.0 275250.0 521100.0 276450.0 ;
      RECT  200100.0 285750.0 526500.0 286950.0 ;
      RECT  200100.0 283650.0 526500.0 284850.0 ;
      RECT  200100.0 281550.0 526500.0 282750.0 ;
      RECT  200100.0 279450.0 526500.0 280650.0 ;
      RECT  94950.0 6750.0 95850.0 7650.0 ;
      RECT  94950.0 11250.0 95850.0 12150.0 ;
      RECT  90750.0 6750.0 95400.0 7650.0 ;
      RECT  94950.0 7200.0 95850.0 11700.0 ;
      RECT  95400.0 11250.0 97950.0 12150.0 ;
      RECT  79350.0 6750.0 87300.0 7650.0 ;
      RECT  94950.0 21150.0 95850.0 22050.0 ;
      RECT  94950.0 25050.0 95850.0 25950.0 ;
      RECT  90750.0 21150.0 95400.0 22050.0 ;
      RECT  94950.0 21600.0 95850.0 25500.0 ;
      RECT  95400.0 25050.0 100950.0 25950.0 ;
      RECT  82350.0 21150.0 87300.0 22050.0 ;
      RECT  79350.0 29850.0 103950.0 30750.0 ;
      RECT  82350.0 43650.0 106950.0 44550.0 ;
      RECT  97950.0 7950.0 111900.0 8850.0 ;
      RECT  100950.0 5250.0 114900.0 6150.0 ;
      RECT  103950.0 19950.0 111900.0 20850.0 ;
      RECT  100950.0 22650.0 114900.0 23550.0 ;
      RECT  97950.0 35550.0 111900.0 36450.0 ;
      RECT  106950.0 32850.0 114900.0 33750.0 ;
      RECT  103950.0 47550.0 111900.0 48450.0 ;
      RECT  106950.0 50250.0 114900.0 51150.0 ;
      RECT  121350.0 7950.0 122250.0 8850.0 ;
      RECT  121350.0 6750.0 122250.0 7650.0 ;
      RECT  117300.0 7950.0 121800.0 8850.0 ;
      RECT  121350.0 7200.0 122250.0 8400.0 ;
      RECT  121800.0 6750.0 126300.0 7650.0 ;
      RECT  121350.0 19950.0 122250.0 20850.0 ;
      RECT  121350.0 21150.0 122250.0 22050.0 ;
      RECT  117300.0 19950.0 121800.0 20850.0 ;
      RECT  121350.0 20400.0 122250.0 21600.0 ;
      RECT  121800.0 21150.0 126300.0 22050.0 ;
      RECT  121350.0 35550.0 122250.0 36450.0 ;
      RECT  121350.0 34350.0 122250.0 35250.0 ;
      RECT  117300.0 35550.0 121800.0 36450.0 ;
      RECT  121350.0 34800.0 122250.0 36000.0 ;
      RECT  121800.0 34350.0 126300.0 35250.0 ;
      RECT  121350.0 47550.0 122250.0 48450.0 ;
      RECT  121350.0 48750.0 122250.0 49650.0 ;
      RECT  117300.0 47550.0 121800.0 48450.0 ;
      RECT  121350.0 48000.0 122250.0 49200.0 ;
      RECT  121800.0 48750.0 126300.0 49650.0 ;
      RECT  91500.0 12450.0 92700.0 14400.0 ;
      RECT  91500.0 600.0 92700.0 2550.0 ;
      RECT  86700.0 1950.0 87900.0 150.0 ;
      RECT  86700.0 11250.0 87900.0 14850.0 ;
      RECT  89400.0 1950.0 90300.0 11250.0 ;
      RECT  86700.0 11250.0 87900.0 12450.0 ;
      RECT  89100.0 11250.0 90300.0 12450.0 ;
      RECT  89100.0 11250.0 90300.0 12450.0 ;
      RECT  86700.0 11250.0 87900.0 12450.0 ;
      RECT  86700.0 1950.0 87900.0 3150.0 ;
      RECT  89100.0 1950.0 90300.0 3150.0 ;
      RECT  89100.0 1950.0 90300.0 3150.0 ;
      RECT  86700.0 1950.0 87900.0 3150.0 ;
      RECT  91500.0 11850.0 92700.0 13050.0 ;
      RECT  91500.0 1950.0 92700.0 3150.0 ;
      RECT  87300.0 6600.0 88500.0 7800.0 ;
      RECT  87300.0 6600.0 88500.0 7800.0 ;
      RECT  89850.0 6750.0 90750.0 7650.0 ;
      RECT  84900.0 13950.0 94500.0 14850.0 ;
      RECT  84900.0 150.0 94500.0 1050.0 ;
      RECT  91500.0 16350.0 92700.0 14400.0 ;
      RECT  91500.0 28200.0 92700.0 26250.0 ;
      RECT  86700.0 26850.0 87900.0 28650.0 ;
      RECT  86700.0 17550.0 87900.0 13950.0 ;
      RECT  89400.0 26850.0 90300.0 17550.0 ;
      RECT  86700.0 17550.0 87900.0 16350.0 ;
      RECT  89100.0 17550.0 90300.0 16350.0 ;
      RECT  89100.0 17550.0 90300.0 16350.0 ;
      RECT  86700.0 17550.0 87900.0 16350.0 ;
      RECT  86700.0 26850.0 87900.0 25650.0 ;
      RECT  89100.0 26850.0 90300.0 25650.0 ;
      RECT  89100.0 26850.0 90300.0 25650.0 ;
      RECT  86700.0 26850.0 87900.0 25650.0 ;
      RECT  91500.0 16950.0 92700.0 15750.0 ;
      RECT  91500.0 26850.0 92700.0 25650.0 ;
      RECT  87300.0 22200.0 88500.0 21000.0 ;
      RECT  87300.0 22200.0 88500.0 21000.0 ;
      RECT  89850.0 22050.0 90750.0 21150.0 ;
      RECT  84900.0 14850.0 94500.0 13950.0 ;
      RECT  84900.0 28650.0 94500.0 27750.0 ;
      RECT  130500.0 12450.0 131700.0 14400.0 ;
      RECT  130500.0 600.0 131700.0 2550.0 ;
      RECT  125700.0 1950.0 126900.0 150.0 ;
      RECT  125700.0 11250.0 126900.0 14850.0 ;
      RECT  128400.0 1950.0 129300.0 11250.0 ;
      RECT  125700.0 11250.0 126900.0 12450.0 ;
      RECT  128100.0 11250.0 129300.0 12450.0 ;
      RECT  128100.0 11250.0 129300.0 12450.0 ;
      RECT  125700.0 11250.0 126900.0 12450.0 ;
      RECT  125700.0 1950.0 126900.0 3150.0 ;
      RECT  128100.0 1950.0 129300.0 3150.0 ;
      RECT  128100.0 1950.0 129300.0 3150.0 ;
      RECT  125700.0 1950.0 126900.0 3150.0 ;
      RECT  130500.0 11850.0 131700.0 13050.0 ;
      RECT  130500.0 1950.0 131700.0 3150.0 ;
      RECT  126300.0 6600.0 127500.0 7800.0 ;
      RECT  126300.0 6600.0 127500.0 7800.0 ;
      RECT  128850.0 6750.0 129750.0 7650.0 ;
      RECT  123900.0 13950.0 133500.0 14850.0 ;
      RECT  123900.0 150.0 133500.0 1050.0 ;
      RECT  130500.0 16350.0 131700.0 14400.0 ;
      RECT  130500.0 28200.0 131700.0 26250.0 ;
      RECT  125700.0 26850.0 126900.0 28650.0 ;
      RECT  125700.0 17550.0 126900.0 13950.0 ;
      RECT  128400.0 26850.0 129300.0 17550.0 ;
      RECT  125700.0 17550.0 126900.0 16350.0 ;
      RECT  128100.0 17550.0 129300.0 16350.0 ;
      RECT  128100.0 17550.0 129300.0 16350.0 ;
      RECT  125700.0 17550.0 126900.0 16350.0 ;
      RECT  125700.0 26850.0 126900.0 25650.0 ;
      RECT  128100.0 26850.0 129300.0 25650.0 ;
      RECT  128100.0 26850.0 129300.0 25650.0 ;
      RECT  125700.0 26850.0 126900.0 25650.0 ;
      RECT  130500.0 16950.0 131700.0 15750.0 ;
      RECT  130500.0 26850.0 131700.0 25650.0 ;
      RECT  126300.0 22200.0 127500.0 21000.0 ;
      RECT  126300.0 22200.0 127500.0 21000.0 ;
      RECT  128850.0 22050.0 129750.0 21150.0 ;
      RECT  123900.0 14850.0 133500.0 13950.0 ;
      RECT  123900.0 28650.0 133500.0 27750.0 ;
      RECT  130500.0 40050.0 131700.0 42000.0 ;
      RECT  130500.0 28200.0 131700.0 30150.0 ;
      RECT  125700.0 29550.0 126900.0 27750.0 ;
      RECT  125700.0 38850.0 126900.0 42450.0 ;
      RECT  128400.0 29550.0 129300.0 38850.0 ;
      RECT  125700.0 38850.0 126900.0 40050.0 ;
      RECT  128100.0 38850.0 129300.0 40050.0 ;
      RECT  128100.0 38850.0 129300.0 40050.0 ;
      RECT  125700.0 38850.0 126900.0 40050.0 ;
      RECT  125700.0 29550.0 126900.0 30750.0 ;
      RECT  128100.0 29550.0 129300.0 30750.0 ;
      RECT  128100.0 29550.0 129300.0 30750.0 ;
      RECT  125700.0 29550.0 126900.0 30750.0 ;
      RECT  130500.0 39450.0 131700.0 40650.0 ;
      RECT  130500.0 29550.0 131700.0 30750.0 ;
      RECT  126300.0 34200.0 127500.0 35400.0 ;
      RECT  126300.0 34200.0 127500.0 35400.0 ;
      RECT  128850.0 34350.0 129750.0 35250.0 ;
      RECT  123900.0 41550.0 133500.0 42450.0 ;
      RECT  123900.0 27750.0 133500.0 28650.0 ;
      RECT  130500.0 43950.0 131700.0 42000.0 ;
      RECT  130500.0 55800.0 131700.0 53850.0 ;
      RECT  125700.0 54450.0 126900.0 56250.0 ;
      RECT  125700.0 45150.0 126900.0 41550.0 ;
      RECT  128400.0 54450.0 129300.0 45150.0 ;
      RECT  125700.0 45150.0 126900.0 43950.0 ;
      RECT  128100.0 45150.0 129300.0 43950.0 ;
      RECT  128100.0 45150.0 129300.0 43950.0 ;
      RECT  125700.0 45150.0 126900.0 43950.0 ;
      RECT  125700.0 54450.0 126900.0 53250.0 ;
      RECT  128100.0 54450.0 129300.0 53250.0 ;
      RECT  128100.0 54450.0 129300.0 53250.0 ;
      RECT  125700.0 54450.0 126900.0 53250.0 ;
      RECT  130500.0 44550.0 131700.0 43350.0 ;
      RECT  130500.0 54450.0 131700.0 53250.0 ;
      RECT  126300.0 49800.0 127500.0 48600.0 ;
      RECT  126300.0 49800.0 127500.0 48600.0 ;
      RECT  128850.0 49650.0 129750.0 48750.0 ;
      RECT  123900.0 42450.0 133500.0 41550.0 ;
      RECT  123900.0 56250.0 133500.0 55350.0 ;
      RECT  111300.0 2550.0 112500.0 150.0 ;
      RECT  111300.0 11250.0 112500.0 14850.0 ;
      RECT  116100.0 11250.0 117300.0 14850.0 ;
      RECT  118500.0 12450.0 119700.0 14400.0 ;
      RECT  118500.0 600.0 119700.0 2550.0 ;
      RECT  111300.0 11250.0 112500.0 12450.0 ;
      RECT  113700.0 11250.0 114900.0 12450.0 ;
      RECT  113700.0 11250.0 114900.0 12450.0 ;
      RECT  111300.0 11250.0 112500.0 12450.0 ;
      RECT  113700.0 11250.0 114900.0 12450.0 ;
      RECT  116100.0 11250.0 117300.0 12450.0 ;
      RECT  116100.0 11250.0 117300.0 12450.0 ;
      RECT  113700.0 11250.0 114900.0 12450.0 ;
      RECT  111300.0 2550.0 112500.0 3750.0 ;
      RECT  113700.0 2550.0 114900.0 3750.0 ;
      RECT  113700.0 2550.0 114900.0 3750.0 ;
      RECT  111300.0 2550.0 112500.0 3750.0 ;
      RECT  113700.0 2550.0 114900.0 3750.0 ;
      RECT  116100.0 2550.0 117300.0 3750.0 ;
      RECT  116100.0 2550.0 117300.0 3750.0 ;
      RECT  113700.0 2550.0 114900.0 3750.0 ;
      RECT  118500.0 11850.0 119700.0 13050.0 ;
      RECT  118500.0 1950.0 119700.0 3150.0 ;
      RECT  116100.0 5100.0 114900.0 6300.0 ;
      RECT  113100.0 7800.0 111900.0 9000.0 ;
      RECT  113700.0 11250.0 114900.0 12450.0 ;
      RECT  116100.0 2550.0 117300.0 3750.0 ;
      RECT  117300.0 7800.0 116100.0 9000.0 ;
      RECT  111900.0 7800.0 113100.0 9000.0 ;
      RECT  114900.0 5100.0 116100.0 6300.0 ;
      RECT  116100.0 7800.0 117300.0 9000.0 ;
      RECT  109500.0 13950.0 123900.0 14850.0 ;
      RECT  109500.0 150.0 123900.0 1050.0 ;
      RECT  111300.0 26250.0 112500.0 28650.0 ;
      RECT  111300.0 17550.0 112500.0 13950.0 ;
      RECT  116100.0 17550.0 117300.0 13950.0 ;
      RECT  118500.0 16350.0 119700.0 14400.0 ;
      RECT  118500.0 28200.0 119700.0 26250.0 ;
      RECT  111300.0 17550.0 112500.0 16350.0 ;
      RECT  113700.0 17550.0 114900.0 16350.0 ;
      RECT  113700.0 17550.0 114900.0 16350.0 ;
      RECT  111300.0 17550.0 112500.0 16350.0 ;
      RECT  113700.0 17550.0 114900.0 16350.0 ;
      RECT  116100.0 17550.0 117300.0 16350.0 ;
      RECT  116100.0 17550.0 117300.0 16350.0 ;
      RECT  113700.0 17550.0 114900.0 16350.0 ;
      RECT  111300.0 26250.0 112500.0 25050.0 ;
      RECT  113700.0 26250.0 114900.0 25050.0 ;
      RECT  113700.0 26250.0 114900.0 25050.0 ;
      RECT  111300.0 26250.0 112500.0 25050.0 ;
      RECT  113700.0 26250.0 114900.0 25050.0 ;
      RECT  116100.0 26250.0 117300.0 25050.0 ;
      RECT  116100.0 26250.0 117300.0 25050.0 ;
      RECT  113700.0 26250.0 114900.0 25050.0 ;
      RECT  118500.0 16950.0 119700.0 15750.0 ;
      RECT  118500.0 26850.0 119700.0 25650.0 ;
      RECT  116100.0 23700.0 114900.0 22500.0 ;
      RECT  113100.0 21000.0 111900.0 19800.0 ;
      RECT  113700.0 17550.0 114900.0 16350.0 ;
      RECT  116100.0 26250.0 117300.0 25050.0 ;
      RECT  117300.0 21000.0 116100.0 19800.0 ;
      RECT  111900.0 21000.0 113100.0 19800.0 ;
      RECT  114900.0 23700.0 116100.0 22500.0 ;
      RECT  116100.0 21000.0 117300.0 19800.0 ;
      RECT  109500.0 14850.0 123900.0 13950.0 ;
      RECT  109500.0 28650.0 123900.0 27750.0 ;
      RECT  111300.0 30150.0 112500.0 27750.0 ;
      RECT  111300.0 38850.0 112500.0 42450.0 ;
      RECT  116100.0 38850.0 117300.0 42450.0 ;
      RECT  118500.0 40050.0 119700.0 42000.0 ;
      RECT  118500.0 28200.0 119700.0 30150.0 ;
      RECT  111300.0 38850.0 112500.0 40050.0 ;
      RECT  113700.0 38850.0 114900.0 40050.0 ;
      RECT  113700.0 38850.0 114900.0 40050.0 ;
      RECT  111300.0 38850.0 112500.0 40050.0 ;
      RECT  113700.0 38850.0 114900.0 40050.0 ;
      RECT  116100.0 38850.0 117300.0 40050.0 ;
      RECT  116100.0 38850.0 117300.0 40050.0 ;
      RECT  113700.0 38850.0 114900.0 40050.0 ;
      RECT  111300.0 30150.0 112500.0 31350.0 ;
      RECT  113700.0 30150.0 114900.0 31350.0 ;
      RECT  113700.0 30150.0 114900.0 31350.0 ;
      RECT  111300.0 30150.0 112500.0 31350.0 ;
      RECT  113700.0 30150.0 114900.0 31350.0 ;
      RECT  116100.0 30150.0 117300.0 31350.0 ;
      RECT  116100.0 30150.0 117300.0 31350.0 ;
      RECT  113700.0 30150.0 114900.0 31350.0 ;
      RECT  118500.0 39450.0 119700.0 40650.0 ;
      RECT  118500.0 29550.0 119700.0 30750.0 ;
      RECT  116100.0 32700.0 114900.0 33900.0 ;
      RECT  113100.0 35400.0 111900.0 36600.0 ;
      RECT  113700.0 38850.0 114900.0 40050.0 ;
      RECT  116100.0 30150.0 117300.0 31350.0 ;
      RECT  117300.0 35400.0 116100.0 36600.0 ;
      RECT  111900.0 35400.0 113100.0 36600.0 ;
      RECT  114900.0 32700.0 116100.0 33900.0 ;
      RECT  116100.0 35400.0 117300.0 36600.0 ;
      RECT  109500.0 41550.0 123900.0 42450.0 ;
      RECT  109500.0 27750.0 123900.0 28650.0 ;
      RECT  111300.0 53850.0 112500.0 56250.0 ;
      RECT  111300.0 45150.0 112500.0 41550.0 ;
      RECT  116100.0 45150.0 117300.0 41550.0 ;
      RECT  118500.0 43950.0 119700.0 42000.0 ;
      RECT  118500.0 55800.0 119700.0 53850.0 ;
      RECT  111300.0 45150.0 112500.0 43950.0 ;
      RECT  113700.0 45150.0 114900.0 43950.0 ;
      RECT  113700.0 45150.0 114900.0 43950.0 ;
      RECT  111300.0 45150.0 112500.0 43950.0 ;
      RECT  113700.0 45150.0 114900.0 43950.0 ;
      RECT  116100.0 45150.0 117300.0 43950.0 ;
      RECT  116100.0 45150.0 117300.0 43950.0 ;
      RECT  113700.0 45150.0 114900.0 43950.0 ;
      RECT  111300.0 53850.0 112500.0 52650.0 ;
      RECT  113700.0 53850.0 114900.0 52650.0 ;
      RECT  113700.0 53850.0 114900.0 52650.0 ;
      RECT  111300.0 53850.0 112500.0 52650.0 ;
      RECT  113700.0 53850.0 114900.0 52650.0 ;
      RECT  116100.0 53850.0 117300.0 52650.0 ;
      RECT  116100.0 53850.0 117300.0 52650.0 ;
      RECT  113700.0 53850.0 114900.0 52650.0 ;
      RECT  118500.0 44550.0 119700.0 43350.0 ;
      RECT  118500.0 54450.0 119700.0 53250.0 ;
      RECT  116100.0 51300.0 114900.0 50100.0 ;
      RECT  113100.0 48600.0 111900.0 47400.0 ;
      RECT  113700.0 45150.0 114900.0 43950.0 ;
      RECT  116100.0 53850.0 117300.0 52650.0 ;
      RECT  117300.0 48600.0 116100.0 47400.0 ;
      RECT  111900.0 48600.0 113100.0 47400.0 ;
      RECT  114900.0 51300.0 116100.0 50100.0 ;
      RECT  116100.0 48600.0 117300.0 47400.0 ;
      RECT  109500.0 42450.0 123900.0 41550.0 ;
      RECT  109500.0 56250.0 123900.0 55350.0 ;
      RECT  98550.0 11100.0 97350.0 12300.0 ;
      RECT  79950.0 6600.0 78750.0 7800.0 ;
      RECT  101550.0 24900.0 100350.0 26100.0 ;
      RECT  82950.0 21000.0 81750.0 22200.0 ;
      RECT  79950.0 29700.0 78750.0 30900.0 ;
      RECT  104550.0 29700.0 103350.0 30900.0 ;
      RECT  82950.0 43500.0 81750.0 44700.0 ;
      RECT  107550.0 43500.0 106350.0 44700.0 ;
      RECT  98550.0 7800.0 97350.0 9000.0 ;
      RECT  101550.0 5100.0 100350.0 6300.0 ;
      RECT  104550.0 19800.0 103350.0 21000.0 ;
      RECT  101550.0 22500.0 100350.0 23700.0 ;
      RECT  98550.0 35400.0 97350.0 36600.0 ;
      RECT  107550.0 32700.0 106350.0 33900.0 ;
      RECT  104550.0 47400.0 103350.0 48600.0 ;
      RECT  107550.0 50100.0 106350.0 51300.0 ;
      RECT  129750.0 6750.0 133500.0 7650.0 ;
      RECT  129750.0 21150.0 133500.0 22050.0 ;
      RECT  129750.0 34350.0 133500.0 35250.0 ;
      RECT  129750.0 48750.0 133500.0 49650.0 ;
      RECT  78900.0 13950.0 133500.0 14850.0 ;
      RECT  78900.0 41550.0 133500.0 42450.0 ;
      RECT  78900.0 150.0 133500.0 1050.0 ;
      RECT  78900.0 27750.0 133500.0 28650.0 ;
      RECT  78900.0 55350.0 133500.0 56250.0 ;
      RECT  200100.0 224250.0 210300.0 273150.0 ;
      RECT  240900.0 224250.0 251100.0 273150.0 ;
      RECT  281700.0 224250.0 291900.0 273150.0 ;
      RECT  322500.0 224250.0 332700.0 273150.0 ;
      RECT  363300.0 224250.0 373500.0 273150.0 ;
      RECT  404100.0 224250.0 414300.0 273150.0 ;
      RECT  444900.0 224250.0 455100.0 273150.0 ;
      RECT  485700.0 224250.0 495900.0 273150.0 ;
      RECT  200100.0 268950.0 526500.0 269850.0 ;
      RECT  200100.0 241650.0 526500.0 242550.0 ;
      RECT  200100.0 266850.0 526500.0 267750.0 ;
      RECT  200100.0 163650.0 210300.0 224250.0 ;
      RECT  240900.0 163650.0 251100.0 224250.0 ;
      RECT  281700.0 163650.0 291900.0 224250.0 ;
      RECT  322500.0 163650.0 332700.0 224250.0 ;
      RECT  363300.0 163650.0 373500.0 224250.0 ;
      RECT  404100.0 163650.0 414300.0 224250.0 ;
      RECT  444900.0 163650.0 455100.0 224250.0 ;
      RECT  485700.0 163650.0 495900.0 224250.0 ;
      RECT  200100.0 170850.0 526500.0 171750.0 ;
      RECT  200100.0 172950.0 526500.0 173850.0 ;
      RECT  200100.0 168750.0 526500.0 169650.0 ;
      RECT  200100.0 103650.0 210300.0 163650.0 ;
      RECT  240900.0 103650.0 251100.0 163650.0 ;
      RECT  281700.0 103650.0 291900.0 163650.0 ;
      RECT  322500.0 103650.0 332700.0 163650.0 ;
      RECT  363300.0 103650.0 373500.0 163650.0 ;
      RECT  404100.0 103650.0 414300.0 163650.0 ;
      RECT  444900.0 103650.0 455100.0 163650.0 ;
      RECT  485700.0 103650.0 495900.0 163650.0 ;
      RECT  200100.0 106050.0 526500.0 106950.0 ;
      RECT  200100.0 160050.0 526500.0 160950.0 ;
      RECT  200100.0 103650.0 210300.0 81750.0 ;
      RECT  240900.0 103650.0 251100.0 81750.0 ;
      RECT  281700.0 103650.0 291900.0 81750.0 ;
      RECT  322500.0 103650.0 332700.0 81750.0 ;
      RECT  363300.0 103650.0 373500.0 81750.0 ;
      RECT  404100.0 103650.0 414300.0 81750.0 ;
      RECT  444900.0 103650.0 455100.0 81750.0 ;
      RECT  485700.0 103650.0 495900.0 81750.0 ;
      RECT  200100.0 100050.0 495900.0 99150.0 ;
      RECT  200100.0 102450.0 495900.0 101550.0 ;
      RECT  200100.0 84150.0 495900.0 83250.0 ;
      RECT  200100.0 97950.0 495900.0 97050.0 ;
      RECT  97950.0 321900.0 98850.0 322800.0 ;
      RECT  97950.0 319950.0 98850.0 320850.0 ;
      RECT  94500.0 321900.0 98400.0 322800.0 ;
      RECT  97950.0 320400.0 98850.0 322350.0 ;
      RECT  98400.0 319950.0 102300.0 320850.0 ;
      RECT  97950.0 332400.0 98850.0 333300.0 ;
      RECT  97950.0 334350.0 98850.0 335250.0 ;
      RECT  94500.0 332400.0 98400.0 333300.0 ;
      RECT  97950.0 332850.0 98850.0 334800.0 ;
      RECT  98400.0 334350.0 102300.0 335250.0 ;
      RECT  97950.0 349500.0 98850.0 350400.0 ;
      RECT  97950.0 347550.0 98850.0 348450.0 ;
      RECT  94500.0 349500.0 98400.0 350400.0 ;
      RECT  97950.0 348000.0 98850.0 349950.0 ;
      RECT  98400.0 347550.0 102300.0 348450.0 ;
      RECT  97950.0 360000.0 98850.0 360900.0 ;
      RECT  97950.0 361950.0 98850.0 362850.0 ;
      RECT  94500.0 360000.0 98400.0 360900.0 ;
      RECT  97950.0 360450.0 98850.0 362400.0 ;
      RECT  98400.0 361950.0 102300.0 362850.0 ;
      RECT  97950.0 377100.0 98850.0 378000.0 ;
      RECT  97950.0 375150.0 98850.0 376050.0 ;
      RECT  94500.0 377100.0 98400.0 378000.0 ;
      RECT  97950.0 375600.0 98850.0 377550.0 ;
      RECT  98400.0 375150.0 102300.0 376050.0 ;
      RECT  97950.0 387600.0 98850.0 388500.0 ;
      RECT  97950.0 389550.0 98850.0 390450.0 ;
      RECT  94500.0 387600.0 98400.0 388500.0 ;
      RECT  97950.0 388050.0 98850.0 390000.0 ;
      RECT  98400.0 389550.0 102300.0 390450.0 ;
      RECT  97950.0 404700.0 98850.0 405600.0 ;
      RECT  97950.0 402750.0 98850.0 403650.0 ;
      RECT  94500.0 404700.0 98400.0 405600.0 ;
      RECT  97950.0 403200.0 98850.0 405150.0 ;
      RECT  98400.0 402750.0 102300.0 403650.0 ;
      RECT  97950.0 415200.0 98850.0 416100.0 ;
      RECT  97950.0 417150.0 98850.0 418050.0 ;
      RECT  94500.0 415200.0 98400.0 416100.0 ;
      RECT  97950.0 415650.0 98850.0 417600.0 ;
      RECT  98400.0 417150.0 102300.0 418050.0 ;
      RECT  97950.0 432300.0 98850.0 433200.0 ;
      RECT  97950.0 430350.0 98850.0 431250.0 ;
      RECT  94500.0 432300.0 98400.0 433200.0 ;
      RECT  97950.0 430800.0 98850.0 432750.0 ;
      RECT  98400.0 430350.0 102300.0 431250.0 ;
      RECT  97950.0 442800.0 98850.0 443700.0 ;
      RECT  97950.0 444750.0 98850.0 445650.0 ;
      RECT  94500.0 442800.0 98400.0 443700.0 ;
      RECT  97950.0 443250.0 98850.0 445200.0 ;
      RECT  98400.0 444750.0 102300.0 445650.0 ;
      RECT  97950.0 459900.0 98850.0 460800.0 ;
      RECT  97950.0 457950.0 98850.0 458850.0 ;
      RECT  94500.0 459900.0 98400.0 460800.0 ;
      RECT  97950.0 458400.0 98850.0 460350.0 ;
      RECT  98400.0 457950.0 102300.0 458850.0 ;
      RECT  97950.0 470400.0 98850.0 471300.0 ;
      RECT  97950.0 472350.0 98850.0 473250.0 ;
      RECT  94500.0 470400.0 98400.0 471300.0 ;
      RECT  97950.0 470850.0 98850.0 472800.0 ;
      RECT  98400.0 472350.0 102300.0 473250.0 ;
      RECT  97950.0 487500.0 98850.0 488400.0 ;
      RECT  97950.0 485550.0 98850.0 486450.0 ;
      RECT  94500.0 487500.0 98400.0 488400.0 ;
      RECT  97950.0 486000.0 98850.0 487950.0 ;
      RECT  98400.0 485550.0 102300.0 486450.0 ;
      RECT  97950.0 498000.0 98850.0 498900.0 ;
      RECT  97950.0 499950.0 98850.0 500850.0 ;
      RECT  94500.0 498000.0 98400.0 498900.0 ;
      RECT  97950.0 498450.0 98850.0 500400.0 ;
      RECT  98400.0 499950.0 102300.0 500850.0 ;
      RECT  97950.0 515100.0 98850.0 516000.0 ;
      RECT  97950.0 513150.0 98850.0 514050.0 ;
      RECT  94500.0 515100.0 98400.0 516000.0 ;
      RECT  97950.0 513600.0 98850.0 515550.0 ;
      RECT  98400.0 513150.0 102300.0 514050.0 ;
      RECT  97950.0 525600.0 98850.0 526500.0 ;
      RECT  97950.0 527550.0 98850.0 528450.0 ;
      RECT  94500.0 525600.0 98400.0 526500.0 ;
      RECT  97950.0 526050.0 98850.0 528000.0 ;
      RECT  98400.0 527550.0 102300.0 528450.0 ;
      RECT  97950.0 542700.0 98850.0 543600.0 ;
      RECT  97950.0 540750.0 98850.0 541650.0 ;
      RECT  94500.0 542700.0 98400.0 543600.0 ;
      RECT  97950.0 541200.0 98850.0 543150.0 ;
      RECT  98400.0 540750.0 102300.0 541650.0 ;
      RECT  97950.0 553200.0 98850.0 554100.0 ;
      RECT  97950.0 555150.0 98850.0 556050.0 ;
      RECT  94500.0 553200.0 98400.0 554100.0 ;
      RECT  97950.0 553650.0 98850.0 555600.0 ;
      RECT  98400.0 555150.0 102300.0 556050.0 ;
      RECT  97950.0 570300.0 98850.0 571200.0 ;
      RECT  97950.0 568350.0 98850.0 569250.0 ;
      RECT  94500.0 570300.0 98400.0 571200.0 ;
      RECT  97950.0 568800.0 98850.0 570750.0 ;
      RECT  98400.0 568350.0 102300.0 569250.0 ;
      RECT  97950.0 580800.0 98850.0 581700.0 ;
      RECT  97950.0 582750.0 98850.0 583650.0 ;
      RECT  94500.0 580800.0 98400.0 581700.0 ;
      RECT  97950.0 581250.0 98850.0 583200.0 ;
      RECT  98400.0 582750.0 102300.0 583650.0 ;
      RECT  97950.0 597900.0 98850.0 598800.0 ;
      RECT  97950.0 595950.0 98850.0 596850.0 ;
      RECT  94500.0 597900.0 98400.0 598800.0 ;
      RECT  97950.0 596400.0 98850.0 598350.0 ;
      RECT  98400.0 595950.0 102300.0 596850.0 ;
      RECT  97950.0 608400.0 98850.0 609300.0 ;
      RECT  97950.0 610350.0 98850.0 611250.0 ;
      RECT  94500.0 608400.0 98400.0 609300.0 ;
      RECT  97950.0 608850.0 98850.0 610800.0 ;
      RECT  98400.0 610350.0 102300.0 611250.0 ;
      RECT  97950.0 625500.0 98850.0 626400.0 ;
      RECT  97950.0 623550.0 98850.0 624450.0 ;
      RECT  94500.0 625500.0 98400.0 626400.0 ;
      RECT  97950.0 624000.0 98850.0 625950.0 ;
      RECT  98400.0 623550.0 102300.0 624450.0 ;
      RECT  97950.0 636000.0 98850.0 636900.0 ;
      RECT  97950.0 637950.0 98850.0 638850.0 ;
      RECT  94500.0 636000.0 98400.0 636900.0 ;
      RECT  97950.0 636450.0 98850.0 638400.0 ;
      RECT  98400.0 637950.0 102300.0 638850.0 ;
      RECT  97950.0 653100.0 98850.0 654000.0 ;
      RECT  97950.0 651150.0 98850.0 652050.0 ;
      RECT  94500.0 653100.0 98400.0 654000.0 ;
      RECT  97950.0 651600.0 98850.0 653550.0 ;
      RECT  98400.0 651150.0 102300.0 652050.0 ;
      RECT  97950.0 663600.0 98850.0 664500.0 ;
      RECT  97950.0 665550.0 98850.0 666450.0 ;
      RECT  94500.0 663600.0 98400.0 664500.0 ;
      RECT  97950.0 664050.0 98850.0 666000.0 ;
      RECT  98400.0 665550.0 102300.0 666450.0 ;
      RECT  97950.0 680700.0 98850.0 681600.0 ;
      RECT  97950.0 678750.0 98850.0 679650.0 ;
      RECT  94500.0 680700.0 98400.0 681600.0 ;
      RECT  97950.0 679200.0 98850.0 681150.0 ;
      RECT  98400.0 678750.0 102300.0 679650.0 ;
      RECT  97950.0 691200.0 98850.0 692100.0 ;
      RECT  97950.0 693150.0 98850.0 694050.0 ;
      RECT  94500.0 691200.0 98400.0 692100.0 ;
      RECT  97950.0 691650.0 98850.0 693600.0 ;
      RECT  98400.0 693150.0 102300.0 694050.0 ;
      RECT  97950.0 708300.0 98850.0 709200.0 ;
      RECT  97950.0 706350.0 98850.0 707250.0 ;
      RECT  94500.0 708300.0 98400.0 709200.0 ;
      RECT  97950.0 706800.0 98850.0 708750.0 ;
      RECT  98400.0 706350.0 102300.0 707250.0 ;
      RECT  97950.0 718800.0 98850.0 719700.0 ;
      RECT  97950.0 720750.0 98850.0 721650.0 ;
      RECT  94500.0 718800.0 98400.0 719700.0 ;
      RECT  97950.0 719250.0 98850.0 721200.0 ;
      RECT  98400.0 720750.0 102300.0 721650.0 ;
      RECT  97950.0 735900.0 98850.0 736800.0 ;
      RECT  97950.0 733950.0 98850.0 734850.0 ;
      RECT  94500.0 735900.0 98400.0 736800.0 ;
      RECT  97950.0 734400.0 98850.0 736350.0 ;
      RECT  98400.0 733950.0 102300.0 734850.0 ;
      RECT  97950.0 746400.0 98850.0 747300.0 ;
      RECT  97950.0 748350.0 98850.0 749250.0 ;
      RECT  94500.0 746400.0 98400.0 747300.0 ;
      RECT  97950.0 746850.0 98850.0 748800.0 ;
      RECT  98400.0 748350.0 102300.0 749250.0 ;
      RECT  97950.0 763500.0 98850.0 764400.0 ;
      RECT  97950.0 761550.0 98850.0 762450.0 ;
      RECT  94500.0 763500.0 98400.0 764400.0 ;
      RECT  97950.0 762000.0 98850.0 763950.0 ;
      RECT  98400.0 761550.0 102300.0 762450.0 ;
      RECT  97950.0 774000.0 98850.0 774900.0 ;
      RECT  97950.0 775950.0 98850.0 776850.0 ;
      RECT  94500.0 774000.0 98400.0 774900.0 ;
      RECT  97950.0 774450.0 98850.0 776400.0 ;
      RECT  98400.0 775950.0 102300.0 776850.0 ;
      RECT  97950.0 791100.0 98850.0 792000.0 ;
      RECT  97950.0 789150.0 98850.0 790050.0 ;
      RECT  94500.0 791100.0 98400.0 792000.0 ;
      RECT  97950.0 789600.0 98850.0 791550.0 ;
      RECT  98400.0 789150.0 102300.0 790050.0 ;
      RECT  97950.0 801600.0 98850.0 802500.0 ;
      RECT  97950.0 803550.0 98850.0 804450.0 ;
      RECT  94500.0 801600.0 98400.0 802500.0 ;
      RECT  97950.0 802050.0 98850.0 804000.0 ;
      RECT  98400.0 803550.0 102300.0 804450.0 ;
      RECT  97950.0 818700.0 98850.0 819600.0 ;
      RECT  97950.0 816750.0 98850.0 817650.0 ;
      RECT  94500.0 818700.0 98400.0 819600.0 ;
      RECT  97950.0 817200.0 98850.0 819150.0 ;
      RECT  98400.0 816750.0 102300.0 817650.0 ;
      RECT  97950.0 829200.0 98850.0 830100.0 ;
      RECT  97950.0 831150.0 98850.0 832050.0 ;
      RECT  94500.0 829200.0 98400.0 830100.0 ;
      RECT  97950.0 829650.0 98850.0 831600.0 ;
      RECT  98400.0 831150.0 102300.0 832050.0 ;
      RECT  97950.0 846300.0 98850.0 847200.0 ;
      RECT  97950.0 844350.0 98850.0 845250.0 ;
      RECT  94500.0 846300.0 98400.0 847200.0 ;
      RECT  97950.0 844800.0 98850.0 846750.0 ;
      RECT  98400.0 844350.0 102300.0 845250.0 ;
      RECT  97950.0 856800.0 98850.0 857700.0 ;
      RECT  97950.0 858750.0 98850.0 859650.0 ;
      RECT  94500.0 856800.0 98400.0 857700.0 ;
      RECT  97950.0 857250.0 98850.0 859200.0 ;
      RECT  98400.0 858750.0 102300.0 859650.0 ;
      RECT  97950.0 873900.0 98850.0 874800.0 ;
      RECT  97950.0 871950.0 98850.0 872850.0 ;
      RECT  94500.0 873900.0 98400.0 874800.0 ;
      RECT  97950.0 872400.0 98850.0 874350.0 ;
      RECT  98400.0 871950.0 102300.0 872850.0 ;
      RECT  97950.0 884400.0 98850.0 885300.0 ;
      RECT  97950.0 886350.0 98850.0 887250.0 ;
      RECT  94500.0 884400.0 98400.0 885300.0 ;
      RECT  97950.0 884850.0 98850.0 886800.0 ;
      RECT  98400.0 886350.0 102300.0 887250.0 ;
      RECT  97950.0 901500.0 98850.0 902400.0 ;
      RECT  97950.0 899550.0 98850.0 900450.0 ;
      RECT  94500.0 901500.0 98400.0 902400.0 ;
      RECT  97950.0 900000.0 98850.0 901950.0 ;
      RECT  98400.0 899550.0 102300.0 900450.0 ;
      RECT  97950.0 912000.0 98850.0 912900.0 ;
      RECT  97950.0 913950.0 98850.0 914850.0 ;
      RECT  94500.0 912000.0 98400.0 912900.0 ;
      RECT  97950.0 912450.0 98850.0 914400.0 ;
      RECT  98400.0 913950.0 102300.0 914850.0 ;
      RECT  97950.0 929100.0 98850.0 930000.0 ;
      RECT  97950.0 927150.0 98850.0 928050.0 ;
      RECT  94500.0 929100.0 98400.0 930000.0 ;
      RECT  97950.0 927600.0 98850.0 929550.0 ;
      RECT  98400.0 927150.0 102300.0 928050.0 ;
      RECT  97950.0 939600.0 98850.0 940500.0 ;
      RECT  97950.0 941550.0 98850.0 942450.0 ;
      RECT  94500.0 939600.0 98400.0 940500.0 ;
      RECT  97950.0 940050.0 98850.0 942000.0 ;
      RECT  98400.0 941550.0 102300.0 942450.0 ;
      RECT  97950.0 956700.0 98850.0 957600.0 ;
      RECT  97950.0 954750.0 98850.0 955650.0 ;
      RECT  94500.0 956700.0 98400.0 957600.0 ;
      RECT  97950.0 955200.0 98850.0 957150.0 ;
      RECT  98400.0 954750.0 102300.0 955650.0 ;
      RECT  97950.0 967200.0 98850.0 968100.0 ;
      RECT  97950.0 969150.0 98850.0 970050.0 ;
      RECT  94500.0 967200.0 98400.0 968100.0 ;
      RECT  97950.0 967650.0 98850.0 969600.0 ;
      RECT  98400.0 969150.0 102300.0 970050.0 ;
      RECT  97950.0 984300.0 98850.0 985200.0 ;
      RECT  97950.0 982350.0 98850.0 983250.0 ;
      RECT  94500.0 984300.0 98400.0 985200.0 ;
      RECT  97950.0 982800.0 98850.0 984750.0 ;
      RECT  98400.0 982350.0 102300.0 983250.0 ;
      RECT  97950.0 994800.0 98850.0 995700.0 ;
      RECT  97950.0 996750.0 98850.0 997650.0 ;
      RECT  94500.0 994800.0 98400.0 995700.0 ;
      RECT  97950.0 995250.0 98850.0 997200.0 ;
      RECT  98400.0 996750.0 102300.0 997650.0 ;
      RECT  97950.0 1011900.0 98850.0 1012800.0 ;
      RECT  97950.0 1009950.0 98850.0 1010850.0 ;
      RECT  94500.0 1011900.0 98400.0 1012800.0 ;
      RECT  97950.0 1010400.0 98850.0 1012350.0 ;
      RECT  98400.0 1009950.0 102300.0 1010850.0 ;
      RECT  97950.0 1022400.0 98850.0 1023300.0 ;
      RECT  97950.0 1024350.0 98850.0 1025250.0 ;
      RECT  94500.0 1022400.0 98400.0 1023300.0 ;
      RECT  97950.0 1022850.0 98850.0 1024800.0 ;
      RECT  98400.0 1024350.0 102300.0 1025250.0 ;
      RECT  97950.0 1039500.0 98850.0 1040400.0 ;
      RECT  97950.0 1037550.0 98850.0 1038450.0 ;
      RECT  94500.0 1039500.0 98400.0 1040400.0 ;
      RECT  97950.0 1038000.0 98850.0 1039950.0 ;
      RECT  98400.0 1037550.0 102300.0 1038450.0 ;
      RECT  97950.0 1050000.0 98850.0 1050900.0 ;
      RECT  97950.0 1051950.0 98850.0 1052850.0 ;
      RECT  94500.0 1050000.0 98400.0 1050900.0 ;
      RECT  97950.0 1050450.0 98850.0 1052400.0 ;
      RECT  98400.0 1051950.0 102300.0 1052850.0 ;
      RECT  97950.0 1067100.0 98850.0 1068000.0 ;
      RECT  97950.0 1065150.0 98850.0 1066050.0 ;
      RECT  94500.0 1067100.0 98400.0 1068000.0 ;
      RECT  97950.0 1065600.0 98850.0 1067550.0 ;
      RECT  98400.0 1065150.0 102300.0 1066050.0 ;
      RECT  97950.0 1077600.0 98850.0 1078500.0 ;
      RECT  97950.0 1079550.0 98850.0 1080450.0 ;
      RECT  94500.0 1077600.0 98400.0 1078500.0 ;
      RECT  97950.0 1078050.0 98850.0 1080000.0 ;
      RECT  98400.0 1079550.0 102300.0 1080450.0 ;
      RECT  97950.0 1094700.0 98850.0 1095600.0 ;
      RECT  97950.0 1092750.0 98850.0 1093650.0 ;
      RECT  94500.0 1094700.0 98400.0 1095600.0 ;
      RECT  97950.0 1093200.0 98850.0 1095150.0 ;
      RECT  98400.0 1092750.0 102300.0 1093650.0 ;
      RECT  97950.0 1105200.0 98850.0 1106100.0 ;
      RECT  97950.0 1107150.0 98850.0 1108050.0 ;
      RECT  94500.0 1105200.0 98400.0 1106100.0 ;
      RECT  97950.0 1105650.0 98850.0 1107600.0 ;
      RECT  98400.0 1107150.0 102300.0 1108050.0 ;
      RECT  97950.0 1122300.0 98850.0 1123200.0 ;
      RECT  97950.0 1120350.0 98850.0 1121250.0 ;
      RECT  94500.0 1122300.0 98400.0 1123200.0 ;
      RECT  97950.0 1120800.0 98850.0 1122750.0 ;
      RECT  98400.0 1120350.0 102300.0 1121250.0 ;
      RECT  97950.0 1132800.0 98850.0 1133700.0 ;
      RECT  97950.0 1134750.0 98850.0 1135650.0 ;
      RECT  94500.0 1132800.0 98400.0 1133700.0 ;
      RECT  97950.0 1133250.0 98850.0 1135200.0 ;
      RECT  98400.0 1134750.0 102300.0 1135650.0 ;
      RECT  97950.0 1149900.0 98850.0 1150800.0 ;
      RECT  97950.0 1147950.0 98850.0 1148850.0 ;
      RECT  94500.0 1149900.0 98400.0 1150800.0 ;
      RECT  97950.0 1148400.0 98850.0 1150350.0 ;
      RECT  98400.0 1147950.0 102300.0 1148850.0 ;
      RECT  97950.0 1160400.0 98850.0 1161300.0 ;
      RECT  97950.0 1162350.0 98850.0 1163250.0 ;
      RECT  94500.0 1160400.0 98400.0 1161300.0 ;
      RECT  97950.0 1160850.0 98850.0 1162800.0 ;
      RECT  98400.0 1162350.0 102300.0 1163250.0 ;
      RECT  97950.0 1177500.0 98850.0 1178400.0 ;
      RECT  97950.0 1175550.0 98850.0 1176450.0 ;
      RECT  94500.0 1177500.0 98400.0 1178400.0 ;
      RECT  97950.0 1176000.0 98850.0 1177950.0 ;
      RECT  98400.0 1175550.0 102300.0 1176450.0 ;
      RECT  97950.0 1188000.0 98850.0 1188900.0 ;
      RECT  97950.0 1189950.0 98850.0 1190850.0 ;
      RECT  94500.0 1188000.0 98400.0 1188900.0 ;
      RECT  97950.0 1188450.0 98850.0 1190400.0 ;
      RECT  98400.0 1189950.0 102300.0 1190850.0 ;
      RECT  59550.0 154350.0 84300.0 155250.0 ;
      RECT  61650.0 168750.0 84300.0 169650.0 ;
      RECT  63750.0 181950.0 84300.0 182850.0 ;
      RECT  65850.0 196350.0 84300.0 197250.0 ;
      RECT  67950.0 209550.0 84300.0 210450.0 ;
      RECT  70050.0 223950.0 84300.0 224850.0 ;
      RECT  72150.0 237150.0 84300.0 238050.0 ;
      RECT  74250.0 251550.0 84300.0 252450.0 ;
      RECT  76350.0 264750.0 84300.0 265650.0 ;
      RECT  78450.0 279150.0 84300.0 280050.0 ;
      RECT  80550.0 292350.0 84300.0 293250.0 ;
      RECT  82650.0 306750.0 84300.0 307650.0 ;
      RECT  59550.0 321900.0 87300.0 322800.0 ;
      RECT  67950.0 319950.0 89700.0 320850.0 ;
      RECT  76350.0 318000.0 92100.0 318900.0 ;
      RECT  59550.0 332400.0 87300.0 333300.0 ;
      RECT  67950.0 334350.0 89700.0 335250.0 ;
      RECT  78450.0 336300.0 92100.0 337200.0 ;
      RECT  59550.0 349500.0 87300.0 350400.0 ;
      RECT  67950.0 347550.0 89700.0 348450.0 ;
      RECT  80550.0 345600.0 92100.0 346500.0 ;
      RECT  59550.0 360000.0 87300.0 360900.0 ;
      RECT  67950.0 361950.0 89700.0 362850.0 ;
      RECT  82650.0 363900.0 92100.0 364800.0 ;
      RECT  59550.0 377100.0 87300.0 378000.0 ;
      RECT  70050.0 375150.0 89700.0 376050.0 ;
      RECT  76350.0 373200.0 92100.0 374100.0 ;
      RECT  59550.0 387600.0 87300.0 388500.0 ;
      RECT  70050.0 389550.0 89700.0 390450.0 ;
      RECT  78450.0 391500.0 92100.0 392400.0 ;
      RECT  59550.0 404700.0 87300.0 405600.0 ;
      RECT  70050.0 402750.0 89700.0 403650.0 ;
      RECT  80550.0 400800.0 92100.0 401700.0 ;
      RECT  59550.0 415200.0 87300.0 416100.0 ;
      RECT  70050.0 417150.0 89700.0 418050.0 ;
      RECT  82650.0 419100.0 92100.0 420000.0 ;
      RECT  59550.0 432300.0 87300.0 433200.0 ;
      RECT  72150.0 430350.0 89700.0 431250.0 ;
      RECT  76350.0 428400.0 92100.0 429300.0 ;
      RECT  59550.0 442800.0 87300.0 443700.0 ;
      RECT  72150.0 444750.0 89700.0 445650.0 ;
      RECT  78450.0 446700.0 92100.0 447600.0 ;
      RECT  59550.0 459900.0 87300.0 460800.0 ;
      RECT  72150.0 457950.0 89700.0 458850.0 ;
      RECT  80550.0 456000.0 92100.0 456900.0 ;
      RECT  59550.0 470400.0 87300.0 471300.0 ;
      RECT  72150.0 472350.0 89700.0 473250.0 ;
      RECT  82650.0 474300.0 92100.0 475200.0 ;
      RECT  59550.0 487500.0 87300.0 488400.0 ;
      RECT  74250.0 485550.0 89700.0 486450.0 ;
      RECT  76350.0 483600.0 92100.0 484500.0 ;
      RECT  59550.0 498000.0 87300.0 498900.0 ;
      RECT  74250.0 499950.0 89700.0 500850.0 ;
      RECT  78450.0 501900.0 92100.0 502800.0 ;
      RECT  59550.0 515100.0 87300.0 516000.0 ;
      RECT  74250.0 513150.0 89700.0 514050.0 ;
      RECT  80550.0 511200.0 92100.0 512100.0 ;
      RECT  59550.0 525600.0 87300.0 526500.0 ;
      RECT  74250.0 527550.0 89700.0 528450.0 ;
      RECT  82650.0 529500.0 92100.0 530400.0 ;
      RECT  61650.0 542700.0 87300.0 543600.0 ;
      RECT  67950.0 540750.0 89700.0 541650.0 ;
      RECT  76350.0 538800.0 92100.0 539700.0 ;
      RECT  61650.0 553200.0 87300.0 554100.0 ;
      RECT  67950.0 555150.0 89700.0 556050.0 ;
      RECT  78450.0 557100.0 92100.0 558000.0 ;
      RECT  61650.0 570300.0 87300.0 571200.0 ;
      RECT  67950.0 568350.0 89700.0 569250.0 ;
      RECT  80550.0 566400.0 92100.0 567300.0 ;
      RECT  61650.0 580800.0 87300.0 581700.0 ;
      RECT  67950.0 582750.0 89700.0 583650.0 ;
      RECT  82650.0 584700.0 92100.0 585600.0 ;
      RECT  61650.0 597900.0 87300.0 598800.0 ;
      RECT  70050.0 595950.0 89700.0 596850.0 ;
      RECT  76350.0 594000.0 92100.0 594900.0 ;
      RECT  61650.0 608400.0 87300.0 609300.0 ;
      RECT  70050.0 610350.0 89700.0 611250.0 ;
      RECT  78450.0 612300.0 92100.0 613200.0 ;
      RECT  61650.0 625500.0 87300.0 626400.0 ;
      RECT  70050.0 623550.0 89700.0 624450.0 ;
      RECT  80550.0 621600.0 92100.0 622500.0 ;
      RECT  61650.0 636000.0 87300.0 636900.0 ;
      RECT  70050.0 637950.0 89700.0 638850.0 ;
      RECT  82650.0 639900.0 92100.0 640800.0 ;
      RECT  61650.0 653100.0 87300.0 654000.0 ;
      RECT  72150.0 651150.0 89700.0 652050.0 ;
      RECT  76350.0 649200.0 92100.0 650100.0 ;
      RECT  61650.0 663600.0 87300.0 664500.0 ;
      RECT  72150.0 665550.0 89700.0 666450.0 ;
      RECT  78450.0 667500.0 92100.0 668400.0 ;
      RECT  61650.0 680700.0 87300.0 681600.0 ;
      RECT  72150.0 678750.0 89700.0 679650.0 ;
      RECT  80550.0 676800.0 92100.0 677700.0 ;
      RECT  61650.0 691200.0 87300.0 692100.0 ;
      RECT  72150.0 693150.0 89700.0 694050.0 ;
      RECT  82650.0 695100.0 92100.0 696000.0 ;
      RECT  61650.0 708300.0 87300.0 709200.0 ;
      RECT  74250.0 706350.0 89700.0 707250.0 ;
      RECT  76350.0 704400.0 92100.0 705300.0 ;
      RECT  61650.0 718800.0 87300.0 719700.0 ;
      RECT  74250.0 720750.0 89700.0 721650.0 ;
      RECT  78450.0 722700.0 92100.0 723600.0 ;
      RECT  61650.0 735900.0 87300.0 736800.0 ;
      RECT  74250.0 733950.0 89700.0 734850.0 ;
      RECT  80550.0 732000.0 92100.0 732900.0 ;
      RECT  61650.0 746400.0 87300.0 747300.0 ;
      RECT  74250.0 748350.0 89700.0 749250.0 ;
      RECT  82650.0 750300.0 92100.0 751200.0 ;
      RECT  63750.0 763500.0 87300.0 764400.0 ;
      RECT  67950.0 761550.0 89700.0 762450.0 ;
      RECT  76350.0 759600.0 92100.0 760500.0 ;
      RECT  63750.0 774000.0 87300.0 774900.0 ;
      RECT  67950.0 775950.0 89700.0 776850.0 ;
      RECT  78450.0 777900.0 92100.0 778800.0 ;
      RECT  63750.0 791100.0 87300.0 792000.0 ;
      RECT  67950.0 789150.0 89700.0 790050.0 ;
      RECT  80550.0 787200.0 92100.0 788100.0 ;
      RECT  63750.0 801600.0 87300.0 802500.0 ;
      RECT  67950.0 803550.0 89700.0 804450.0 ;
      RECT  82650.0 805500.0 92100.0 806400.0 ;
      RECT  63750.0 818700.0 87300.0 819600.0 ;
      RECT  70050.0 816750.0 89700.0 817650.0 ;
      RECT  76350.0 814800.0 92100.0 815700.0 ;
      RECT  63750.0 829200.0 87300.0 830100.0 ;
      RECT  70050.0 831150.0 89700.0 832050.0 ;
      RECT  78450.0 833100.0 92100.0 834000.0 ;
      RECT  63750.0 846300.0 87300.0 847200.0 ;
      RECT  70050.0 844350.0 89700.0 845250.0 ;
      RECT  80550.0 842400.0 92100.0 843300.0 ;
      RECT  63750.0 856800.0 87300.0 857700.0 ;
      RECT  70050.0 858750.0 89700.0 859650.0 ;
      RECT  82650.0 860700.0 92100.0 861600.0 ;
      RECT  63750.0 873900.0 87300.0 874800.0 ;
      RECT  72150.0 871950.0 89700.0 872850.0 ;
      RECT  76350.0 870000.0 92100.0 870900.0 ;
      RECT  63750.0 884400.0 87300.0 885300.0 ;
      RECT  72150.0 886350.0 89700.0 887250.0 ;
      RECT  78450.0 888300.0 92100.0 889200.0 ;
      RECT  63750.0 901500.0 87300.0 902400.0 ;
      RECT  72150.0 899550.0 89700.0 900450.0 ;
      RECT  80550.0 897600.0 92100.0 898500.0 ;
      RECT  63750.0 912000.0 87300.0 912900.0 ;
      RECT  72150.0 913950.0 89700.0 914850.0 ;
      RECT  82650.0 915900.0 92100.0 916800.0 ;
      RECT  63750.0 929100.0 87300.0 930000.0 ;
      RECT  74250.0 927150.0 89700.0 928050.0 ;
      RECT  76350.0 925200.0 92100.0 926100.0 ;
      RECT  63750.0 939600.0 87300.0 940500.0 ;
      RECT  74250.0 941550.0 89700.0 942450.0 ;
      RECT  78450.0 943500.0 92100.0 944400.0 ;
      RECT  63750.0 956700.0 87300.0 957600.0 ;
      RECT  74250.0 954750.0 89700.0 955650.0 ;
      RECT  80550.0 952800.0 92100.0 953700.0 ;
      RECT  63750.0 967200.0 87300.0 968100.0 ;
      RECT  74250.0 969150.0 89700.0 970050.0 ;
      RECT  82650.0 971100.0 92100.0 972000.0 ;
      RECT  65850.0 984300.0 87300.0 985200.0 ;
      RECT  67950.0 982350.0 89700.0 983250.0 ;
      RECT  76350.0 980400.0 92100.0 981300.0 ;
      RECT  65850.0 994800.0 87300.0 995700.0 ;
      RECT  67950.0 996750.0 89700.0 997650.0 ;
      RECT  78450.0 998700.0 92100.0 999600.0 ;
      RECT  65850.0 1011900.0 87300.0 1012800.0 ;
      RECT  67950.0 1009950.0 89700.0 1010850.0 ;
      RECT  80550.0 1008000.0 92100.0 1008900.0 ;
      RECT  65850.0 1022400.0 87300.0 1023300.0 ;
      RECT  67950.0 1024350.0 89700.0 1025250.0 ;
      RECT  82650.0 1026300.0 92100.0 1027200.0 ;
      RECT  65850.0 1039500.0 87300.0 1040400.0 ;
      RECT  70050.0 1037550.0 89700.0 1038450.0 ;
      RECT  76350.0 1035600.0 92100.0 1036500.0 ;
      RECT  65850.0 1050000.0 87300.0 1050900.0 ;
      RECT  70050.0 1051950.0 89700.0 1052850.0 ;
      RECT  78450.0 1053900.0 92100.0 1054800.0 ;
      RECT  65850.0 1067100.0 87300.0 1068000.0 ;
      RECT  70050.0 1065150.0 89700.0 1066050.0 ;
      RECT  80550.0 1063200.0 92100.0 1064100.0 ;
      RECT  65850.0 1077600.0 87300.0 1078500.0 ;
      RECT  70050.0 1079550.0 89700.0 1080450.0 ;
      RECT  82650.0 1081500.0 92100.0 1082400.0 ;
      RECT  65850.0 1094700.0 87300.0 1095600.0 ;
      RECT  72150.0 1092750.0 89700.0 1093650.0 ;
      RECT  76350.0 1090800.0 92100.0 1091700.0 ;
      RECT  65850.0 1105200.0 87300.0 1106100.0 ;
      RECT  72150.0 1107150.0 89700.0 1108050.0 ;
      RECT  78450.0 1109100.0 92100.0 1110000.0 ;
      RECT  65850.0 1122300.0 87300.0 1123200.0 ;
      RECT  72150.0 1120350.0 89700.0 1121250.0 ;
      RECT  80550.0 1118400.0 92100.0 1119300.0 ;
      RECT  65850.0 1132800.0 87300.0 1133700.0 ;
      RECT  72150.0 1134750.0 89700.0 1135650.0 ;
      RECT  82650.0 1136700.0 92100.0 1137600.0 ;
      RECT  65850.0 1149900.0 87300.0 1150800.0 ;
      RECT  74250.0 1147950.0 89700.0 1148850.0 ;
      RECT  76350.0 1146000.0 92100.0 1146900.0 ;
      RECT  65850.0 1160400.0 87300.0 1161300.0 ;
      RECT  74250.0 1162350.0 89700.0 1163250.0 ;
      RECT  78450.0 1164300.0 92100.0 1165200.0 ;
      RECT  65850.0 1177500.0 87300.0 1178400.0 ;
      RECT  74250.0 1175550.0 89700.0 1176450.0 ;
      RECT  80550.0 1173600.0 92100.0 1174500.0 ;
      RECT  65850.0 1188000.0 87300.0 1188900.0 ;
      RECT  74250.0 1189950.0 89700.0 1190850.0 ;
      RECT  82650.0 1191900.0 92100.0 1192800.0 ;
      RECT  122850.0 154350.0 121950.0 155250.0 ;
      RECT  122850.0 158850.0 121950.0 159750.0 ;
      RECT  127050.0 154350.0 122400.0 155250.0 ;
      RECT  122850.0 154800.0 121950.0 159300.0 ;
      RECT  122400.0 158850.0 119850.0 159750.0 ;
      RECT  138450.0 154350.0 130500.0 155250.0 ;
      RECT  122850.0 168750.0 121950.0 169650.0 ;
      RECT  122850.0 172650.0 121950.0 173550.0 ;
      RECT  127050.0 168750.0 122400.0 169650.0 ;
      RECT  122850.0 169200.0 121950.0 173100.0 ;
      RECT  122400.0 172650.0 116850.0 173550.0 ;
      RECT  135450.0 168750.0 130500.0 169650.0 ;
      RECT  138450.0 177450.0 113850.0 178350.0 ;
      RECT  135450.0 191250.0 110850.0 192150.0 ;
      RECT  119850.0 155550.0 105900.0 156450.0 ;
      RECT  116850.0 152850.0 102900.0 153750.0 ;
      RECT  113850.0 167550.0 105900.0 168450.0 ;
      RECT  116850.0 170250.0 102900.0 171150.0 ;
      RECT  119850.0 183150.0 105900.0 184050.0 ;
      RECT  110850.0 180450.0 102900.0 181350.0 ;
      RECT  113850.0 195150.0 105900.0 196050.0 ;
      RECT  110850.0 197850.0 102900.0 198750.0 ;
      RECT  96450.0 155550.0 95550.0 156450.0 ;
      RECT  96450.0 154350.0 95550.0 155250.0 ;
      RECT  100500.0 155550.0 96000.0 156450.0 ;
      RECT  96450.0 154800.0 95550.0 156000.0 ;
      RECT  96000.0 154350.0 91500.0 155250.0 ;
      RECT  96450.0 167550.0 95550.0 168450.0 ;
      RECT  96450.0 168750.0 95550.0 169650.0 ;
      RECT  100500.0 167550.0 96000.0 168450.0 ;
      RECT  96450.0 168000.0 95550.0 169200.0 ;
      RECT  96000.0 168750.0 91500.0 169650.0 ;
      RECT  96450.0 183150.0 95550.0 184050.0 ;
      RECT  96450.0 181950.0 95550.0 182850.0 ;
      RECT  100500.0 183150.0 96000.0 184050.0 ;
      RECT  96450.0 182400.0 95550.0 183600.0 ;
      RECT  96000.0 181950.0 91500.0 182850.0 ;
      RECT  96450.0 195150.0 95550.0 196050.0 ;
      RECT  96450.0 196350.0 95550.0 197250.0 ;
      RECT  100500.0 195150.0 96000.0 196050.0 ;
      RECT  96450.0 195600.0 95550.0 196800.0 ;
      RECT  96000.0 196350.0 91500.0 197250.0 ;
      RECT  126300.0 160050.0 125100.0 162000.0 ;
      RECT  126300.0 148200.0 125100.0 150150.0 ;
      RECT  131100.0 149550.0 129900.0 147750.0 ;
      RECT  131100.0 158850.0 129900.0 162450.0 ;
      RECT  128400.0 149550.0 127500.0 158850.0 ;
      RECT  131100.0 158850.0 129900.0 160050.0 ;
      RECT  128700.0 158850.0 127500.0 160050.0 ;
      RECT  128700.0 158850.0 127500.0 160050.0 ;
      RECT  131100.0 158850.0 129900.0 160050.0 ;
      RECT  131100.0 149550.0 129900.0 150750.0 ;
      RECT  128700.0 149550.0 127500.0 150750.0 ;
      RECT  128700.0 149550.0 127500.0 150750.0 ;
      RECT  131100.0 149550.0 129900.0 150750.0 ;
      RECT  126300.0 159450.0 125100.0 160650.0 ;
      RECT  126300.0 149550.0 125100.0 150750.0 ;
      RECT  130500.0 154200.0 129300.0 155400.0 ;
      RECT  130500.0 154200.0 129300.0 155400.0 ;
      RECT  127950.0 154350.0 127050.0 155250.0 ;
      RECT  132900.0 161550.0 123300.0 162450.0 ;
      RECT  132900.0 147750.0 123300.0 148650.0 ;
      RECT  126300.0 163950.0 125100.0 162000.0 ;
      RECT  126300.0 175800.0 125100.0 173850.0 ;
      RECT  131100.0 174450.0 129900.0 176250.0 ;
      RECT  131100.0 165150.0 129900.0 161550.0 ;
      RECT  128400.0 174450.0 127500.0 165150.0 ;
      RECT  131100.0 165150.0 129900.0 163950.0 ;
      RECT  128700.0 165150.0 127500.0 163950.0 ;
      RECT  128700.0 165150.0 127500.0 163950.0 ;
      RECT  131100.0 165150.0 129900.0 163950.0 ;
      RECT  131100.0 174450.0 129900.0 173250.0 ;
      RECT  128700.0 174450.0 127500.0 173250.0 ;
      RECT  128700.0 174450.0 127500.0 173250.0 ;
      RECT  131100.0 174450.0 129900.0 173250.0 ;
      RECT  126300.0 164550.0 125100.0 163350.0 ;
      RECT  126300.0 174450.0 125100.0 173250.0 ;
      RECT  130500.0 169800.0 129300.0 168600.0 ;
      RECT  130500.0 169800.0 129300.0 168600.0 ;
      RECT  127950.0 169650.0 127050.0 168750.0 ;
      RECT  132900.0 162450.0 123300.0 161550.0 ;
      RECT  132900.0 176250.0 123300.0 175350.0 ;
      RECT  87300.0 160050.0 86100.0 162000.0 ;
      RECT  87300.0 148200.0 86100.0 150150.0 ;
      RECT  92100.0 149550.0 90900.0 147750.0 ;
      RECT  92100.0 158850.0 90900.0 162450.0 ;
      RECT  89400.0 149550.0 88500.0 158850.0 ;
      RECT  92100.0 158850.0 90900.0 160050.0 ;
      RECT  89700.0 158850.0 88500.0 160050.0 ;
      RECT  89700.0 158850.0 88500.0 160050.0 ;
      RECT  92100.0 158850.0 90900.0 160050.0 ;
      RECT  92100.0 149550.0 90900.0 150750.0 ;
      RECT  89700.0 149550.0 88500.0 150750.0 ;
      RECT  89700.0 149550.0 88500.0 150750.0 ;
      RECT  92100.0 149550.0 90900.0 150750.0 ;
      RECT  87300.0 159450.0 86100.0 160650.0 ;
      RECT  87300.0 149550.0 86100.0 150750.0 ;
      RECT  91500.0 154200.0 90300.0 155400.0 ;
      RECT  91500.0 154200.0 90300.0 155400.0 ;
      RECT  88950.0 154350.0 88050.0 155250.0 ;
      RECT  93900.0 161550.0 84300.0 162450.0 ;
      RECT  93900.0 147750.0 84300.0 148650.0 ;
      RECT  87300.0 163950.0 86100.0 162000.0 ;
      RECT  87300.0 175800.0 86100.0 173850.0 ;
      RECT  92100.0 174450.0 90900.0 176250.0 ;
      RECT  92100.0 165150.0 90900.0 161550.0 ;
      RECT  89400.0 174450.0 88500.0 165150.0 ;
      RECT  92100.0 165150.0 90900.0 163950.0 ;
      RECT  89700.0 165150.0 88500.0 163950.0 ;
      RECT  89700.0 165150.0 88500.0 163950.0 ;
      RECT  92100.0 165150.0 90900.0 163950.0 ;
      RECT  92100.0 174450.0 90900.0 173250.0 ;
      RECT  89700.0 174450.0 88500.0 173250.0 ;
      RECT  89700.0 174450.0 88500.0 173250.0 ;
      RECT  92100.0 174450.0 90900.0 173250.0 ;
      RECT  87300.0 164550.0 86100.0 163350.0 ;
      RECT  87300.0 174450.0 86100.0 173250.0 ;
      RECT  91500.0 169800.0 90300.0 168600.0 ;
      RECT  91500.0 169800.0 90300.0 168600.0 ;
      RECT  88950.0 169650.0 88050.0 168750.0 ;
      RECT  93900.0 162450.0 84300.0 161550.0 ;
      RECT  93900.0 176250.0 84300.0 175350.0 ;
      RECT  87300.0 187650.0 86100.0 189600.0 ;
      RECT  87300.0 175800.0 86100.0 177750.0 ;
      RECT  92100.0 177150.0 90900.0 175350.0 ;
      RECT  92100.0 186450.0 90900.0 190050.0 ;
      RECT  89400.0 177150.0 88500.0 186450.0 ;
      RECT  92100.0 186450.0 90900.0 187650.0 ;
      RECT  89700.0 186450.0 88500.0 187650.0 ;
      RECT  89700.0 186450.0 88500.0 187650.0 ;
      RECT  92100.0 186450.0 90900.0 187650.0 ;
      RECT  92100.0 177150.0 90900.0 178350.0 ;
      RECT  89700.0 177150.0 88500.0 178350.0 ;
      RECT  89700.0 177150.0 88500.0 178350.0 ;
      RECT  92100.0 177150.0 90900.0 178350.0 ;
      RECT  87300.0 187050.0 86100.0 188250.0 ;
      RECT  87300.0 177150.0 86100.0 178350.0 ;
      RECT  91500.0 181800.0 90300.0 183000.0 ;
      RECT  91500.0 181800.0 90300.0 183000.0 ;
      RECT  88950.0 181950.0 88050.0 182850.0 ;
      RECT  93900.0 189150.0 84300.0 190050.0 ;
      RECT  93900.0 175350.0 84300.0 176250.0 ;
      RECT  87300.0 191550.0 86100.0 189600.0 ;
      RECT  87300.0 203400.0 86100.0 201450.0 ;
      RECT  92100.0 202050.0 90900.0 203850.0 ;
      RECT  92100.0 192750.0 90900.0 189150.0 ;
      RECT  89400.0 202050.0 88500.0 192750.0 ;
      RECT  92100.0 192750.0 90900.0 191550.0 ;
      RECT  89700.0 192750.0 88500.0 191550.0 ;
      RECT  89700.0 192750.0 88500.0 191550.0 ;
      RECT  92100.0 192750.0 90900.0 191550.0 ;
      RECT  92100.0 202050.0 90900.0 200850.0 ;
      RECT  89700.0 202050.0 88500.0 200850.0 ;
      RECT  89700.0 202050.0 88500.0 200850.0 ;
      RECT  92100.0 202050.0 90900.0 200850.0 ;
      RECT  87300.0 192150.0 86100.0 190950.0 ;
      RECT  87300.0 202050.0 86100.0 200850.0 ;
      RECT  91500.0 197400.0 90300.0 196200.0 ;
      RECT  91500.0 197400.0 90300.0 196200.0 ;
      RECT  88950.0 197250.0 88050.0 196350.0 ;
      RECT  93900.0 190050.0 84300.0 189150.0 ;
      RECT  93900.0 203850.0 84300.0 202950.0 ;
      RECT  106500.0 150150.0 105300.0 147750.0 ;
      RECT  106500.0 158850.0 105300.0 162450.0 ;
      RECT  101700.0 158850.0 100500.0 162450.0 ;
      RECT  99300.0 160050.0 98100.0 162000.0 ;
      RECT  99300.0 148200.0 98100.0 150150.0 ;
      RECT  106500.0 158850.0 105300.0 160050.0 ;
      RECT  104100.0 158850.0 102900.0 160050.0 ;
      RECT  104100.0 158850.0 102900.0 160050.0 ;
      RECT  106500.0 158850.0 105300.0 160050.0 ;
      RECT  104100.0 158850.0 102900.0 160050.0 ;
      RECT  101700.0 158850.0 100500.0 160050.0 ;
      RECT  101700.0 158850.0 100500.0 160050.0 ;
      RECT  104100.0 158850.0 102900.0 160050.0 ;
      RECT  106500.0 150150.0 105300.0 151350.0 ;
      RECT  104100.0 150150.0 102900.0 151350.0 ;
      RECT  104100.0 150150.0 102900.0 151350.0 ;
      RECT  106500.0 150150.0 105300.0 151350.0 ;
      RECT  104100.0 150150.0 102900.0 151350.0 ;
      RECT  101700.0 150150.0 100500.0 151350.0 ;
      RECT  101700.0 150150.0 100500.0 151350.0 ;
      RECT  104100.0 150150.0 102900.0 151350.0 ;
      RECT  99300.0 159450.0 98100.0 160650.0 ;
      RECT  99300.0 149550.0 98100.0 150750.0 ;
      RECT  101700.0 152700.0 102900.0 153900.0 ;
      RECT  104700.0 155400.0 105900.0 156600.0 ;
      RECT  104100.0 158850.0 102900.0 160050.0 ;
      RECT  101700.0 150150.0 100500.0 151350.0 ;
      RECT  100500.0 155400.0 101700.0 156600.0 ;
      RECT  105900.0 155400.0 104700.0 156600.0 ;
      RECT  102900.0 152700.0 101700.0 153900.0 ;
      RECT  101700.0 155400.0 100500.0 156600.0 ;
      RECT  108300.0 161550.0 93900.0 162450.0 ;
      RECT  108300.0 147750.0 93900.0 148650.0 ;
      RECT  106500.0 173850.0 105300.0 176250.0 ;
      RECT  106500.0 165150.0 105300.0 161550.0 ;
      RECT  101700.0 165150.0 100500.0 161550.0 ;
      RECT  99300.0 163950.0 98100.0 162000.0 ;
      RECT  99300.0 175800.0 98100.0 173850.0 ;
      RECT  106500.0 165150.0 105300.0 163950.0 ;
      RECT  104100.0 165150.0 102900.0 163950.0 ;
      RECT  104100.0 165150.0 102900.0 163950.0 ;
      RECT  106500.0 165150.0 105300.0 163950.0 ;
      RECT  104100.0 165150.0 102900.0 163950.0 ;
      RECT  101700.0 165150.0 100500.0 163950.0 ;
      RECT  101700.0 165150.0 100500.0 163950.0 ;
      RECT  104100.0 165150.0 102900.0 163950.0 ;
      RECT  106500.0 173850.0 105300.0 172650.0 ;
      RECT  104100.0 173850.0 102900.0 172650.0 ;
      RECT  104100.0 173850.0 102900.0 172650.0 ;
      RECT  106500.0 173850.0 105300.0 172650.0 ;
      RECT  104100.0 173850.0 102900.0 172650.0 ;
      RECT  101700.0 173850.0 100500.0 172650.0 ;
      RECT  101700.0 173850.0 100500.0 172650.0 ;
      RECT  104100.0 173850.0 102900.0 172650.0 ;
      RECT  99300.0 164550.0 98100.0 163350.0 ;
      RECT  99300.0 174450.0 98100.0 173250.0 ;
      RECT  101700.0 171300.0 102900.0 170100.0 ;
      RECT  104700.0 168600.0 105900.0 167400.0 ;
      RECT  104100.0 165150.0 102900.0 163950.0 ;
      RECT  101700.0 173850.0 100500.0 172650.0 ;
      RECT  100500.0 168600.0 101700.0 167400.0 ;
      RECT  105900.0 168600.0 104700.0 167400.0 ;
      RECT  102900.0 171300.0 101700.0 170100.0 ;
      RECT  101700.0 168600.0 100500.0 167400.0 ;
      RECT  108300.0 162450.0 93900.0 161550.0 ;
      RECT  108300.0 176250.0 93900.0 175350.0 ;
      RECT  106500.0 177750.0 105300.0 175350.0 ;
      RECT  106500.0 186450.0 105300.0 190050.0 ;
      RECT  101700.0 186450.0 100500.0 190050.0 ;
      RECT  99300.0 187650.0 98100.0 189600.0 ;
      RECT  99300.0 175800.0 98100.0 177750.0 ;
      RECT  106500.0 186450.0 105300.0 187650.0 ;
      RECT  104100.0 186450.0 102900.0 187650.0 ;
      RECT  104100.0 186450.0 102900.0 187650.0 ;
      RECT  106500.0 186450.0 105300.0 187650.0 ;
      RECT  104100.0 186450.0 102900.0 187650.0 ;
      RECT  101700.0 186450.0 100500.0 187650.0 ;
      RECT  101700.0 186450.0 100500.0 187650.0 ;
      RECT  104100.0 186450.0 102900.0 187650.0 ;
      RECT  106500.0 177750.0 105300.0 178950.0 ;
      RECT  104100.0 177750.0 102900.0 178950.0 ;
      RECT  104100.0 177750.0 102900.0 178950.0 ;
      RECT  106500.0 177750.0 105300.0 178950.0 ;
      RECT  104100.0 177750.0 102900.0 178950.0 ;
      RECT  101700.0 177750.0 100500.0 178950.0 ;
      RECT  101700.0 177750.0 100500.0 178950.0 ;
      RECT  104100.0 177750.0 102900.0 178950.0 ;
      RECT  99300.0 187050.0 98100.0 188250.0 ;
      RECT  99300.0 177150.0 98100.0 178350.0 ;
      RECT  101700.0 180300.0 102900.0 181500.0 ;
      RECT  104700.0 183000.0 105900.0 184200.0 ;
      RECT  104100.0 186450.0 102900.0 187650.0 ;
      RECT  101700.0 177750.0 100500.0 178950.0 ;
      RECT  100500.0 183000.0 101700.0 184200.0 ;
      RECT  105900.0 183000.0 104700.0 184200.0 ;
      RECT  102900.0 180300.0 101700.0 181500.0 ;
      RECT  101700.0 183000.0 100500.0 184200.0 ;
      RECT  108300.0 189150.0 93900.0 190050.0 ;
      RECT  108300.0 175350.0 93900.0 176250.0 ;
      RECT  106500.0 201450.0 105300.0 203850.0 ;
      RECT  106500.0 192750.0 105300.0 189150.0 ;
      RECT  101700.0 192750.0 100500.0 189150.0 ;
      RECT  99300.0 191550.0 98100.0 189600.0 ;
      RECT  99300.0 203400.0 98100.0 201450.0 ;
      RECT  106500.0 192750.0 105300.0 191550.0 ;
      RECT  104100.0 192750.0 102900.0 191550.0 ;
      RECT  104100.0 192750.0 102900.0 191550.0 ;
      RECT  106500.0 192750.0 105300.0 191550.0 ;
      RECT  104100.0 192750.0 102900.0 191550.0 ;
      RECT  101700.0 192750.0 100500.0 191550.0 ;
      RECT  101700.0 192750.0 100500.0 191550.0 ;
      RECT  104100.0 192750.0 102900.0 191550.0 ;
      RECT  106500.0 201450.0 105300.0 200250.0 ;
      RECT  104100.0 201450.0 102900.0 200250.0 ;
      RECT  104100.0 201450.0 102900.0 200250.0 ;
      RECT  106500.0 201450.0 105300.0 200250.0 ;
      RECT  104100.0 201450.0 102900.0 200250.0 ;
      RECT  101700.0 201450.0 100500.0 200250.0 ;
      RECT  101700.0 201450.0 100500.0 200250.0 ;
      RECT  104100.0 201450.0 102900.0 200250.0 ;
      RECT  99300.0 192150.0 98100.0 190950.0 ;
      RECT  99300.0 202050.0 98100.0 200850.0 ;
      RECT  101700.0 198900.0 102900.0 197700.0 ;
      RECT  104700.0 196200.0 105900.0 195000.0 ;
      RECT  104100.0 192750.0 102900.0 191550.0 ;
      RECT  101700.0 201450.0 100500.0 200250.0 ;
      RECT  100500.0 196200.0 101700.0 195000.0 ;
      RECT  105900.0 196200.0 104700.0 195000.0 ;
      RECT  102900.0 198900.0 101700.0 197700.0 ;
      RECT  101700.0 196200.0 100500.0 195000.0 ;
      RECT  108300.0 190050.0 93900.0 189150.0 ;
      RECT  108300.0 203850.0 93900.0 202950.0 ;
      RECT  119250.0 158700.0 120450.0 159900.0 ;
      RECT  137850.0 154200.0 139050.0 155400.0 ;
      RECT  116250.0 172500.0 117450.0 173700.0 ;
      RECT  134850.0 168600.0 136050.0 169800.0 ;
      RECT  137850.0 177300.0 139050.0 178500.0 ;
      RECT  113250.0 177300.0 114450.0 178500.0 ;
      RECT  134850.0 191100.0 136050.0 192300.0 ;
      RECT  110250.0 191100.0 111450.0 192300.0 ;
      RECT  119250.0 155400.0 120450.0 156600.0 ;
      RECT  116250.0 152700.0 117450.0 153900.0 ;
      RECT  113250.0 167400.0 114450.0 168600.0 ;
      RECT  116250.0 170100.0 117450.0 171300.0 ;
      RECT  119250.0 183000.0 120450.0 184200.0 ;
      RECT  110250.0 180300.0 111450.0 181500.0 ;
      RECT  113250.0 195000.0 114450.0 196200.0 ;
      RECT  110250.0 197700.0 111450.0 198900.0 ;
      RECT  88050.0 154350.0 84300.0 155250.0 ;
      RECT  88050.0 168750.0 84300.0 169650.0 ;
      RECT  88050.0 181950.0 84300.0 182850.0 ;
      RECT  88050.0 196350.0 84300.0 197250.0 ;
      RECT  138900.0 161550.0 84300.0 162450.0 ;
      RECT  138900.0 189150.0 84300.0 190050.0 ;
      RECT  138900.0 147750.0 84300.0 148650.0 ;
      RECT  138900.0 175350.0 84300.0 176250.0 ;
      RECT  138900.0 202950.0 84300.0 203850.0 ;
      RECT  122850.0 209550.0 121950.0 210450.0 ;
      RECT  122850.0 214050.0 121950.0 214950.0 ;
      RECT  127050.0 209550.0 122400.0 210450.0 ;
      RECT  122850.0 210000.0 121950.0 214500.0 ;
      RECT  122400.0 214050.0 119850.0 214950.0 ;
      RECT  138450.0 209550.0 130500.0 210450.0 ;
      RECT  122850.0 223950.0 121950.0 224850.0 ;
      RECT  122850.0 227850.0 121950.0 228750.0 ;
      RECT  127050.0 223950.0 122400.0 224850.0 ;
      RECT  122850.0 224400.0 121950.0 228300.0 ;
      RECT  122400.0 227850.0 116850.0 228750.0 ;
      RECT  135450.0 223950.0 130500.0 224850.0 ;
      RECT  138450.0 232650.0 113850.0 233550.0 ;
      RECT  135450.0 246450.0 110850.0 247350.0 ;
      RECT  119850.0 210750.0 105900.0 211650.0 ;
      RECT  116850.0 208050.0 102900.0 208950.0 ;
      RECT  113850.0 222750.0 105900.0 223650.0 ;
      RECT  116850.0 225450.0 102900.0 226350.0 ;
      RECT  119850.0 238350.0 105900.0 239250.0 ;
      RECT  110850.0 235650.0 102900.0 236550.0 ;
      RECT  113850.0 250350.0 105900.0 251250.0 ;
      RECT  110850.0 253050.0 102900.0 253950.0 ;
      RECT  96450.0 210750.0 95550.0 211650.0 ;
      RECT  96450.0 209550.0 95550.0 210450.0 ;
      RECT  100500.0 210750.0 96000.0 211650.0 ;
      RECT  96450.0 210000.0 95550.0 211200.0 ;
      RECT  96000.0 209550.0 91500.0 210450.0 ;
      RECT  96450.0 222750.0 95550.0 223650.0 ;
      RECT  96450.0 223950.0 95550.0 224850.0 ;
      RECT  100500.0 222750.0 96000.0 223650.0 ;
      RECT  96450.0 223200.0 95550.0 224400.0 ;
      RECT  96000.0 223950.0 91500.0 224850.0 ;
      RECT  96450.0 238350.0 95550.0 239250.0 ;
      RECT  96450.0 237150.0 95550.0 238050.0 ;
      RECT  100500.0 238350.0 96000.0 239250.0 ;
      RECT  96450.0 237600.0 95550.0 238800.0 ;
      RECT  96000.0 237150.0 91500.0 238050.0 ;
      RECT  96450.0 250350.0 95550.0 251250.0 ;
      RECT  96450.0 251550.0 95550.0 252450.0 ;
      RECT  100500.0 250350.0 96000.0 251250.0 ;
      RECT  96450.0 250800.0 95550.0 252000.0 ;
      RECT  96000.0 251550.0 91500.0 252450.0 ;
      RECT  126300.0 215250.0 125100.0 217200.0 ;
      RECT  126300.0 203400.0 125100.0 205350.0 ;
      RECT  131100.0 204750.0 129900.0 202950.0 ;
      RECT  131100.0 214050.0 129900.0 217650.0 ;
      RECT  128400.0 204750.0 127500.0 214050.0 ;
      RECT  131100.0 214050.0 129900.0 215250.0 ;
      RECT  128700.0 214050.0 127500.0 215250.0 ;
      RECT  128700.0 214050.0 127500.0 215250.0 ;
      RECT  131100.0 214050.0 129900.0 215250.0 ;
      RECT  131100.0 204750.0 129900.0 205950.0 ;
      RECT  128700.0 204750.0 127500.0 205950.0 ;
      RECT  128700.0 204750.0 127500.0 205950.0 ;
      RECT  131100.0 204750.0 129900.0 205950.0 ;
      RECT  126300.0 214650.0 125100.0 215850.0 ;
      RECT  126300.0 204750.0 125100.0 205950.0 ;
      RECT  130500.0 209400.0 129300.0 210600.0 ;
      RECT  130500.0 209400.0 129300.0 210600.0 ;
      RECT  127950.0 209550.0 127050.0 210450.0 ;
      RECT  132900.0 216750.0 123300.0 217650.0 ;
      RECT  132900.0 202950.0 123300.0 203850.0 ;
      RECT  126300.0 219150.0 125100.0 217200.0 ;
      RECT  126300.0 231000.0 125100.0 229050.0 ;
      RECT  131100.0 229650.0 129900.0 231450.0 ;
      RECT  131100.0 220350.0 129900.0 216750.0 ;
      RECT  128400.0 229650.0 127500.0 220350.0 ;
      RECT  131100.0 220350.0 129900.0 219150.0 ;
      RECT  128700.0 220350.0 127500.0 219150.0 ;
      RECT  128700.0 220350.0 127500.0 219150.0 ;
      RECT  131100.0 220350.0 129900.0 219150.0 ;
      RECT  131100.0 229650.0 129900.0 228450.0 ;
      RECT  128700.0 229650.0 127500.0 228450.0 ;
      RECT  128700.0 229650.0 127500.0 228450.0 ;
      RECT  131100.0 229650.0 129900.0 228450.0 ;
      RECT  126300.0 219750.0 125100.0 218550.0 ;
      RECT  126300.0 229650.0 125100.0 228450.0 ;
      RECT  130500.0 225000.0 129300.0 223800.0 ;
      RECT  130500.0 225000.0 129300.0 223800.0 ;
      RECT  127950.0 224850.0 127050.0 223950.0 ;
      RECT  132900.0 217650.0 123300.0 216750.0 ;
      RECT  132900.0 231450.0 123300.0 230550.0 ;
      RECT  87300.0 215250.0 86100.0 217200.0 ;
      RECT  87300.0 203400.0 86100.0 205350.0 ;
      RECT  92100.0 204750.0 90900.0 202950.0 ;
      RECT  92100.0 214050.0 90900.0 217650.0 ;
      RECT  89400.0 204750.0 88500.0 214050.0 ;
      RECT  92100.0 214050.0 90900.0 215250.0 ;
      RECT  89700.0 214050.0 88500.0 215250.0 ;
      RECT  89700.0 214050.0 88500.0 215250.0 ;
      RECT  92100.0 214050.0 90900.0 215250.0 ;
      RECT  92100.0 204750.0 90900.0 205950.0 ;
      RECT  89700.0 204750.0 88500.0 205950.0 ;
      RECT  89700.0 204750.0 88500.0 205950.0 ;
      RECT  92100.0 204750.0 90900.0 205950.0 ;
      RECT  87300.0 214650.0 86100.0 215850.0 ;
      RECT  87300.0 204750.0 86100.0 205950.0 ;
      RECT  91500.0 209400.0 90300.0 210600.0 ;
      RECT  91500.0 209400.0 90300.0 210600.0 ;
      RECT  88950.0 209550.0 88050.0 210450.0 ;
      RECT  93900.0 216750.0 84300.0 217650.0 ;
      RECT  93900.0 202950.0 84300.0 203850.0 ;
      RECT  87300.0 219150.0 86100.0 217200.0 ;
      RECT  87300.0 231000.0 86100.0 229050.0 ;
      RECT  92100.0 229650.0 90900.0 231450.0 ;
      RECT  92100.0 220350.0 90900.0 216750.0 ;
      RECT  89400.0 229650.0 88500.0 220350.0 ;
      RECT  92100.0 220350.0 90900.0 219150.0 ;
      RECT  89700.0 220350.0 88500.0 219150.0 ;
      RECT  89700.0 220350.0 88500.0 219150.0 ;
      RECT  92100.0 220350.0 90900.0 219150.0 ;
      RECT  92100.0 229650.0 90900.0 228450.0 ;
      RECT  89700.0 229650.0 88500.0 228450.0 ;
      RECT  89700.0 229650.0 88500.0 228450.0 ;
      RECT  92100.0 229650.0 90900.0 228450.0 ;
      RECT  87300.0 219750.0 86100.0 218550.0 ;
      RECT  87300.0 229650.0 86100.0 228450.0 ;
      RECT  91500.0 225000.0 90300.0 223800.0 ;
      RECT  91500.0 225000.0 90300.0 223800.0 ;
      RECT  88950.0 224850.0 88050.0 223950.0 ;
      RECT  93900.0 217650.0 84300.0 216750.0 ;
      RECT  93900.0 231450.0 84300.0 230550.0 ;
      RECT  87300.0 242850.0 86100.0 244800.0 ;
      RECT  87300.0 231000.0 86100.0 232950.0 ;
      RECT  92100.0 232350.0 90900.0 230550.0 ;
      RECT  92100.0 241650.0 90900.0 245250.0 ;
      RECT  89400.0 232350.0 88500.0 241650.0 ;
      RECT  92100.0 241650.0 90900.0 242850.0 ;
      RECT  89700.0 241650.0 88500.0 242850.0 ;
      RECT  89700.0 241650.0 88500.0 242850.0 ;
      RECT  92100.0 241650.0 90900.0 242850.0 ;
      RECT  92100.0 232350.0 90900.0 233550.0 ;
      RECT  89700.0 232350.0 88500.0 233550.0 ;
      RECT  89700.0 232350.0 88500.0 233550.0 ;
      RECT  92100.0 232350.0 90900.0 233550.0 ;
      RECT  87300.0 242250.0 86100.0 243450.0 ;
      RECT  87300.0 232350.0 86100.0 233550.0 ;
      RECT  91500.0 237000.0 90300.0 238200.0 ;
      RECT  91500.0 237000.0 90300.0 238200.0 ;
      RECT  88950.0 237150.0 88050.0 238050.0 ;
      RECT  93900.0 244350.0 84300.0 245250.0 ;
      RECT  93900.0 230550.0 84300.0 231450.0 ;
      RECT  87300.0 246750.0 86100.0 244800.0 ;
      RECT  87300.0 258600.0 86100.0 256650.0 ;
      RECT  92100.0 257250.0 90900.0 259050.0 ;
      RECT  92100.0 247950.0 90900.0 244350.0 ;
      RECT  89400.0 257250.0 88500.0 247950.0 ;
      RECT  92100.0 247950.0 90900.0 246750.0 ;
      RECT  89700.0 247950.0 88500.0 246750.0 ;
      RECT  89700.0 247950.0 88500.0 246750.0 ;
      RECT  92100.0 247950.0 90900.0 246750.0 ;
      RECT  92100.0 257250.0 90900.0 256050.0 ;
      RECT  89700.0 257250.0 88500.0 256050.0 ;
      RECT  89700.0 257250.0 88500.0 256050.0 ;
      RECT  92100.0 257250.0 90900.0 256050.0 ;
      RECT  87300.0 247350.0 86100.0 246150.0 ;
      RECT  87300.0 257250.0 86100.0 256050.0 ;
      RECT  91500.0 252600.0 90300.0 251400.0 ;
      RECT  91500.0 252600.0 90300.0 251400.0 ;
      RECT  88950.0 252450.0 88050.0 251550.0 ;
      RECT  93900.0 245250.0 84300.0 244350.0 ;
      RECT  93900.0 259050.0 84300.0 258150.0 ;
      RECT  106500.0 205350.0 105300.0 202950.0 ;
      RECT  106500.0 214050.0 105300.0 217650.0 ;
      RECT  101700.0 214050.0 100500.0 217650.0 ;
      RECT  99300.0 215250.0 98100.0 217200.0 ;
      RECT  99300.0 203400.0 98100.0 205350.0 ;
      RECT  106500.0 214050.0 105300.0 215250.0 ;
      RECT  104100.0 214050.0 102900.0 215250.0 ;
      RECT  104100.0 214050.0 102900.0 215250.0 ;
      RECT  106500.0 214050.0 105300.0 215250.0 ;
      RECT  104100.0 214050.0 102900.0 215250.0 ;
      RECT  101700.0 214050.0 100500.0 215250.0 ;
      RECT  101700.0 214050.0 100500.0 215250.0 ;
      RECT  104100.0 214050.0 102900.0 215250.0 ;
      RECT  106500.0 205350.0 105300.0 206550.0 ;
      RECT  104100.0 205350.0 102900.0 206550.0 ;
      RECT  104100.0 205350.0 102900.0 206550.0 ;
      RECT  106500.0 205350.0 105300.0 206550.0 ;
      RECT  104100.0 205350.0 102900.0 206550.0 ;
      RECT  101700.0 205350.0 100500.0 206550.0 ;
      RECT  101700.0 205350.0 100500.0 206550.0 ;
      RECT  104100.0 205350.0 102900.0 206550.0 ;
      RECT  99300.0 214650.0 98100.0 215850.0 ;
      RECT  99300.0 204750.0 98100.0 205950.0 ;
      RECT  101700.0 207900.0 102900.0 209100.0 ;
      RECT  104700.0 210600.0 105900.0 211800.0 ;
      RECT  104100.0 214050.0 102900.0 215250.0 ;
      RECT  101700.0 205350.0 100500.0 206550.0 ;
      RECT  100500.0 210600.0 101700.0 211800.0 ;
      RECT  105900.0 210600.0 104700.0 211800.0 ;
      RECT  102900.0 207900.0 101700.0 209100.0 ;
      RECT  101700.0 210600.0 100500.0 211800.0 ;
      RECT  108300.0 216750.0 93900.0 217650.0 ;
      RECT  108300.0 202950.0 93900.0 203850.0 ;
      RECT  106500.0 229050.0 105300.0 231450.0 ;
      RECT  106500.0 220350.0 105300.0 216750.0 ;
      RECT  101700.0 220350.0 100500.0 216750.0 ;
      RECT  99300.0 219150.0 98100.0 217200.0 ;
      RECT  99300.0 231000.0 98100.0 229050.0 ;
      RECT  106500.0 220350.0 105300.0 219150.0 ;
      RECT  104100.0 220350.0 102900.0 219150.0 ;
      RECT  104100.0 220350.0 102900.0 219150.0 ;
      RECT  106500.0 220350.0 105300.0 219150.0 ;
      RECT  104100.0 220350.0 102900.0 219150.0 ;
      RECT  101700.0 220350.0 100500.0 219150.0 ;
      RECT  101700.0 220350.0 100500.0 219150.0 ;
      RECT  104100.0 220350.0 102900.0 219150.0 ;
      RECT  106500.0 229050.0 105300.0 227850.0 ;
      RECT  104100.0 229050.0 102900.0 227850.0 ;
      RECT  104100.0 229050.0 102900.0 227850.0 ;
      RECT  106500.0 229050.0 105300.0 227850.0 ;
      RECT  104100.0 229050.0 102900.0 227850.0 ;
      RECT  101700.0 229050.0 100500.0 227850.0 ;
      RECT  101700.0 229050.0 100500.0 227850.0 ;
      RECT  104100.0 229050.0 102900.0 227850.0 ;
      RECT  99300.0 219750.0 98100.0 218550.0 ;
      RECT  99300.0 229650.0 98100.0 228450.0 ;
      RECT  101700.0 226500.0 102900.0 225300.0 ;
      RECT  104700.0 223800.0 105900.0 222600.0 ;
      RECT  104100.0 220350.0 102900.0 219150.0 ;
      RECT  101700.0 229050.0 100500.0 227850.0 ;
      RECT  100500.0 223800.0 101700.0 222600.0 ;
      RECT  105900.0 223800.0 104700.0 222600.0 ;
      RECT  102900.0 226500.0 101700.0 225300.0 ;
      RECT  101700.0 223800.0 100500.0 222600.0 ;
      RECT  108300.0 217650.0 93900.0 216750.0 ;
      RECT  108300.0 231450.0 93900.0 230550.0 ;
      RECT  106500.0 232950.0 105300.0 230550.0 ;
      RECT  106500.0 241650.0 105300.0 245250.0 ;
      RECT  101700.0 241650.0 100500.0 245250.0 ;
      RECT  99300.0 242850.0 98100.0 244800.0 ;
      RECT  99300.0 231000.0 98100.0 232950.0 ;
      RECT  106500.0 241650.0 105300.0 242850.0 ;
      RECT  104100.0 241650.0 102900.0 242850.0 ;
      RECT  104100.0 241650.0 102900.0 242850.0 ;
      RECT  106500.0 241650.0 105300.0 242850.0 ;
      RECT  104100.0 241650.0 102900.0 242850.0 ;
      RECT  101700.0 241650.0 100500.0 242850.0 ;
      RECT  101700.0 241650.0 100500.0 242850.0 ;
      RECT  104100.0 241650.0 102900.0 242850.0 ;
      RECT  106500.0 232950.0 105300.0 234150.0 ;
      RECT  104100.0 232950.0 102900.0 234150.0 ;
      RECT  104100.0 232950.0 102900.0 234150.0 ;
      RECT  106500.0 232950.0 105300.0 234150.0 ;
      RECT  104100.0 232950.0 102900.0 234150.0 ;
      RECT  101700.0 232950.0 100500.0 234150.0 ;
      RECT  101700.0 232950.0 100500.0 234150.0 ;
      RECT  104100.0 232950.0 102900.0 234150.0 ;
      RECT  99300.0 242250.0 98100.0 243450.0 ;
      RECT  99300.0 232350.0 98100.0 233550.0 ;
      RECT  101700.0 235500.0 102900.0 236700.0 ;
      RECT  104700.0 238200.0 105900.0 239400.0 ;
      RECT  104100.0 241650.0 102900.0 242850.0 ;
      RECT  101700.0 232950.0 100500.0 234150.0 ;
      RECT  100500.0 238200.0 101700.0 239400.0 ;
      RECT  105900.0 238200.0 104700.0 239400.0 ;
      RECT  102900.0 235500.0 101700.0 236700.0 ;
      RECT  101700.0 238200.0 100500.0 239400.0 ;
      RECT  108300.0 244350.0 93900.0 245250.0 ;
      RECT  108300.0 230550.0 93900.0 231450.0 ;
      RECT  106500.0 256650.0 105300.0 259050.0 ;
      RECT  106500.0 247950.0 105300.0 244350.0 ;
      RECT  101700.0 247950.0 100500.0 244350.0 ;
      RECT  99300.0 246750.0 98100.0 244800.0 ;
      RECT  99300.0 258600.0 98100.0 256650.0 ;
      RECT  106500.0 247950.0 105300.0 246750.0 ;
      RECT  104100.0 247950.0 102900.0 246750.0 ;
      RECT  104100.0 247950.0 102900.0 246750.0 ;
      RECT  106500.0 247950.0 105300.0 246750.0 ;
      RECT  104100.0 247950.0 102900.0 246750.0 ;
      RECT  101700.0 247950.0 100500.0 246750.0 ;
      RECT  101700.0 247950.0 100500.0 246750.0 ;
      RECT  104100.0 247950.0 102900.0 246750.0 ;
      RECT  106500.0 256650.0 105300.0 255450.0 ;
      RECT  104100.0 256650.0 102900.0 255450.0 ;
      RECT  104100.0 256650.0 102900.0 255450.0 ;
      RECT  106500.0 256650.0 105300.0 255450.0 ;
      RECT  104100.0 256650.0 102900.0 255450.0 ;
      RECT  101700.0 256650.0 100500.0 255450.0 ;
      RECT  101700.0 256650.0 100500.0 255450.0 ;
      RECT  104100.0 256650.0 102900.0 255450.0 ;
      RECT  99300.0 247350.0 98100.0 246150.0 ;
      RECT  99300.0 257250.0 98100.0 256050.0 ;
      RECT  101700.0 254100.0 102900.0 252900.0 ;
      RECT  104700.0 251400.0 105900.0 250200.0 ;
      RECT  104100.0 247950.0 102900.0 246750.0 ;
      RECT  101700.0 256650.0 100500.0 255450.0 ;
      RECT  100500.0 251400.0 101700.0 250200.0 ;
      RECT  105900.0 251400.0 104700.0 250200.0 ;
      RECT  102900.0 254100.0 101700.0 252900.0 ;
      RECT  101700.0 251400.0 100500.0 250200.0 ;
      RECT  108300.0 245250.0 93900.0 244350.0 ;
      RECT  108300.0 259050.0 93900.0 258150.0 ;
      RECT  119250.0 213900.0 120450.0 215100.0 ;
      RECT  137850.0 209400.0 139050.0 210600.0 ;
      RECT  116250.0 227700.0 117450.0 228900.0 ;
      RECT  134850.0 223800.0 136050.0 225000.0 ;
      RECT  137850.0 232500.0 139050.0 233700.0 ;
      RECT  113250.0 232500.0 114450.0 233700.0 ;
      RECT  134850.0 246300.0 136050.0 247500.0 ;
      RECT  110250.0 246300.0 111450.0 247500.0 ;
      RECT  119250.0 210600.0 120450.0 211800.0 ;
      RECT  116250.0 207900.0 117450.0 209100.0 ;
      RECT  113250.0 222600.0 114450.0 223800.0 ;
      RECT  116250.0 225300.0 117450.0 226500.0 ;
      RECT  119250.0 238200.0 120450.0 239400.0 ;
      RECT  110250.0 235500.0 111450.0 236700.0 ;
      RECT  113250.0 250200.0 114450.0 251400.0 ;
      RECT  110250.0 252900.0 111450.0 254100.0 ;
      RECT  88050.0 209550.0 84300.0 210450.0 ;
      RECT  88050.0 223950.0 84300.0 224850.0 ;
      RECT  88050.0 237150.0 84300.0 238050.0 ;
      RECT  88050.0 251550.0 84300.0 252450.0 ;
      RECT  138900.0 216750.0 84300.0 217650.0 ;
      RECT  138900.0 244350.0 84300.0 245250.0 ;
      RECT  138900.0 202950.0 84300.0 203850.0 ;
      RECT  138900.0 230550.0 84300.0 231450.0 ;
      RECT  138900.0 258150.0 84300.0 259050.0 ;
      RECT  122850.0 264750.0 121950.0 265650.0 ;
      RECT  122850.0 269250.0 121950.0 270150.0 ;
      RECT  127050.0 264750.0 122400.0 265650.0 ;
      RECT  122850.0 265200.0 121950.0 269700.0 ;
      RECT  122400.0 269250.0 119850.0 270150.0 ;
      RECT  138450.0 264750.0 130500.0 265650.0 ;
      RECT  122850.0 279150.0 121950.0 280050.0 ;
      RECT  122850.0 283050.0 121950.0 283950.0 ;
      RECT  127050.0 279150.0 122400.0 280050.0 ;
      RECT  122850.0 279600.0 121950.0 283500.0 ;
      RECT  122400.0 283050.0 116850.0 283950.0 ;
      RECT  135450.0 279150.0 130500.0 280050.0 ;
      RECT  138450.0 287850.0 113850.0 288750.0 ;
      RECT  135450.0 301650.0 110850.0 302550.0 ;
      RECT  119850.0 265950.0 105900.0 266850.0 ;
      RECT  116850.0 263250.0 102900.0 264150.0 ;
      RECT  113850.0 277950.0 105900.0 278850.0 ;
      RECT  116850.0 280650.0 102900.0 281550.0 ;
      RECT  119850.0 293550.0 105900.0 294450.0 ;
      RECT  110850.0 290850.0 102900.0 291750.0 ;
      RECT  113850.0 305550.0 105900.0 306450.0 ;
      RECT  110850.0 308250.0 102900.0 309150.0 ;
      RECT  96450.0 265950.0 95550.0 266850.0 ;
      RECT  96450.0 264750.0 95550.0 265650.0 ;
      RECT  100500.0 265950.0 96000.0 266850.0 ;
      RECT  96450.0 265200.0 95550.0 266400.0 ;
      RECT  96000.0 264750.0 91500.0 265650.0 ;
      RECT  96450.0 277950.0 95550.0 278850.0 ;
      RECT  96450.0 279150.0 95550.0 280050.0 ;
      RECT  100500.0 277950.0 96000.0 278850.0 ;
      RECT  96450.0 278400.0 95550.0 279600.0 ;
      RECT  96000.0 279150.0 91500.0 280050.0 ;
      RECT  96450.0 293550.0 95550.0 294450.0 ;
      RECT  96450.0 292350.0 95550.0 293250.0 ;
      RECT  100500.0 293550.0 96000.0 294450.0 ;
      RECT  96450.0 292800.0 95550.0 294000.0 ;
      RECT  96000.0 292350.0 91500.0 293250.0 ;
      RECT  96450.0 305550.0 95550.0 306450.0 ;
      RECT  96450.0 306750.0 95550.0 307650.0 ;
      RECT  100500.0 305550.0 96000.0 306450.0 ;
      RECT  96450.0 306000.0 95550.0 307200.0 ;
      RECT  96000.0 306750.0 91500.0 307650.0 ;
      RECT  126300.0 270450.0 125100.0 272400.0 ;
      RECT  126300.0 258600.0 125100.0 260550.0 ;
      RECT  131100.0 259950.0 129900.0 258150.0 ;
      RECT  131100.0 269250.0 129900.0 272850.0 ;
      RECT  128400.0 259950.0 127500.0 269250.0 ;
      RECT  131100.0 269250.0 129900.0 270450.0 ;
      RECT  128700.0 269250.0 127500.0 270450.0 ;
      RECT  128700.0 269250.0 127500.0 270450.0 ;
      RECT  131100.0 269250.0 129900.0 270450.0 ;
      RECT  131100.0 259950.0 129900.0 261150.0 ;
      RECT  128700.0 259950.0 127500.0 261150.0 ;
      RECT  128700.0 259950.0 127500.0 261150.0 ;
      RECT  131100.0 259950.0 129900.0 261150.0 ;
      RECT  126300.0 269850.0 125100.0 271050.0 ;
      RECT  126300.0 259950.0 125100.0 261150.0 ;
      RECT  130500.0 264600.0 129300.0 265800.0 ;
      RECT  130500.0 264600.0 129300.0 265800.0 ;
      RECT  127950.0 264750.0 127050.0 265650.0 ;
      RECT  132900.0 271950.0 123300.0 272850.0 ;
      RECT  132900.0 258150.0 123300.0 259050.0 ;
      RECT  126300.0 274350.0 125100.0 272400.0 ;
      RECT  126300.0 286200.0 125100.0 284250.0 ;
      RECT  131100.0 284850.0 129900.0 286650.0 ;
      RECT  131100.0 275550.0 129900.0 271950.0 ;
      RECT  128400.0 284850.0 127500.0 275550.0 ;
      RECT  131100.0 275550.0 129900.0 274350.0 ;
      RECT  128700.0 275550.0 127500.0 274350.0 ;
      RECT  128700.0 275550.0 127500.0 274350.0 ;
      RECT  131100.0 275550.0 129900.0 274350.0 ;
      RECT  131100.0 284850.0 129900.0 283650.0 ;
      RECT  128700.0 284850.0 127500.0 283650.0 ;
      RECT  128700.0 284850.0 127500.0 283650.0 ;
      RECT  131100.0 284850.0 129900.0 283650.0 ;
      RECT  126300.0 274950.0 125100.0 273750.0 ;
      RECT  126300.0 284850.0 125100.0 283650.0 ;
      RECT  130500.0 280200.0 129300.0 279000.0 ;
      RECT  130500.0 280200.0 129300.0 279000.0 ;
      RECT  127950.0 280050.0 127050.0 279150.0 ;
      RECT  132900.0 272850.0 123300.0 271950.0 ;
      RECT  132900.0 286650.0 123300.0 285750.0 ;
      RECT  87300.0 270450.0 86100.0 272400.0 ;
      RECT  87300.0 258600.0 86100.0 260550.0 ;
      RECT  92100.0 259950.0 90900.0 258150.0 ;
      RECT  92100.0 269250.0 90900.0 272850.0 ;
      RECT  89400.0 259950.0 88500.0 269250.0 ;
      RECT  92100.0 269250.0 90900.0 270450.0 ;
      RECT  89700.0 269250.0 88500.0 270450.0 ;
      RECT  89700.0 269250.0 88500.0 270450.0 ;
      RECT  92100.0 269250.0 90900.0 270450.0 ;
      RECT  92100.0 259950.0 90900.0 261150.0 ;
      RECT  89700.0 259950.0 88500.0 261150.0 ;
      RECT  89700.0 259950.0 88500.0 261150.0 ;
      RECT  92100.0 259950.0 90900.0 261150.0 ;
      RECT  87300.0 269850.0 86100.0 271050.0 ;
      RECT  87300.0 259950.0 86100.0 261150.0 ;
      RECT  91500.0 264600.0 90300.0 265800.0 ;
      RECT  91500.0 264600.0 90300.0 265800.0 ;
      RECT  88950.0 264750.0 88050.0 265650.0 ;
      RECT  93900.0 271950.0 84300.0 272850.0 ;
      RECT  93900.0 258150.0 84300.0 259050.0 ;
      RECT  87300.0 274350.0 86100.0 272400.0 ;
      RECT  87300.0 286200.0 86100.0 284250.0 ;
      RECT  92100.0 284850.0 90900.0 286650.0 ;
      RECT  92100.0 275550.0 90900.0 271950.0 ;
      RECT  89400.0 284850.0 88500.0 275550.0 ;
      RECT  92100.0 275550.0 90900.0 274350.0 ;
      RECT  89700.0 275550.0 88500.0 274350.0 ;
      RECT  89700.0 275550.0 88500.0 274350.0 ;
      RECT  92100.0 275550.0 90900.0 274350.0 ;
      RECT  92100.0 284850.0 90900.0 283650.0 ;
      RECT  89700.0 284850.0 88500.0 283650.0 ;
      RECT  89700.0 284850.0 88500.0 283650.0 ;
      RECT  92100.0 284850.0 90900.0 283650.0 ;
      RECT  87300.0 274950.0 86100.0 273750.0 ;
      RECT  87300.0 284850.0 86100.0 283650.0 ;
      RECT  91500.0 280200.0 90300.0 279000.0 ;
      RECT  91500.0 280200.0 90300.0 279000.0 ;
      RECT  88950.0 280050.0 88050.0 279150.0 ;
      RECT  93900.0 272850.0 84300.0 271950.0 ;
      RECT  93900.0 286650.0 84300.0 285750.0 ;
      RECT  87300.0 298050.0 86100.0 300000.0 ;
      RECT  87300.0 286200.0 86100.0 288150.0 ;
      RECT  92100.0 287550.0 90900.0 285750.0 ;
      RECT  92100.0 296850.0 90900.0 300450.0 ;
      RECT  89400.0 287550.0 88500.0 296850.0 ;
      RECT  92100.0 296850.0 90900.0 298050.0 ;
      RECT  89700.0 296850.0 88500.0 298050.0 ;
      RECT  89700.0 296850.0 88500.0 298050.0 ;
      RECT  92100.0 296850.0 90900.0 298050.0 ;
      RECT  92100.0 287550.0 90900.0 288750.0 ;
      RECT  89700.0 287550.0 88500.0 288750.0 ;
      RECT  89700.0 287550.0 88500.0 288750.0 ;
      RECT  92100.0 287550.0 90900.0 288750.0 ;
      RECT  87300.0 297450.0 86100.0 298650.0 ;
      RECT  87300.0 287550.0 86100.0 288750.0 ;
      RECT  91500.0 292200.0 90300.0 293400.0 ;
      RECT  91500.0 292200.0 90300.0 293400.0 ;
      RECT  88950.0 292350.0 88050.0 293250.0 ;
      RECT  93900.0 299550.0 84300.0 300450.0 ;
      RECT  93900.0 285750.0 84300.0 286650.0 ;
      RECT  87300.0 301950.0 86100.0 300000.0 ;
      RECT  87300.0 313800.0 86100.0 311850.0 ;
      RECT  92100.0 312450.0 90900.0 314250.0 ;
      RECT  92100.0 303150.0 90900.0 299550.0 ;
      RECT  89400.0 312450.0 88500.0 303150.0 ;
      RECT  92100.0 303150.0 90900.0 301950.0 ;
      RECT  89700.0 303150.0 88500.0 301950.0 ;
      RECT  89700.0 303150.0 88500.0 301950.0 ;
      RECT  92100.0 303150.0 90900.0 301950.0 ;
      RECT  92100.0 312450.0 90900.0 311250.0 ;
      RECT  89700.0 312450.0 88500.0 311250.0 ;
      RECT  89700.0 312450.0 88500.0 311250.0 ;
      RECT  92100.0 312450.0 90900.0 311250.0 ;
      RECT  87300.0 302550.0 86100.0 301350.0 ;
      RECT  87300.0 312450.0 86100.0 311250.0 ;
      RECT  91500.0 307800.0 90300.0 306600.0 ;
      RECT  91500.0 307800.0 90300.0 306600.0 ;
      RECT  88950.0 307650.0 88050.0 306750.0 ;
      RECT  93900.0 300450.0 84300.0 299550.0 ;
      RECT  93900.0 314250.0 84300.0 313350.0 ;
      RECT  106500.0 260550.0 105300.0 258150.0 ;
      RECT  106500.0 269250.0 105300.0 272850.0 ;
      RECT  101700.0 269250.0 100500.0 272850.0 ;
      RECT  99300.0 270450.0 98100.0 272400.0 ;
      RECT  99300.0 258600.0 98100.0 260550.0 ;
      RECT  106500.0 269250.0 105300.0 270450.0 ;
      RECT  104100.0 269250.0 102900.0 270450.0 ;
      RECT  104100.0 269250.0 102900.0 270450.0 ;
      RECT  106500.0 269250.0 105300.0 270450.0 ;
      RECT  104100.0 269250.0 102900.0 270450.0 ;
      RECT  101700.0 269250.0 100500.0 270450.0 ;
      RECT  101700.0 269250.0 100500.0 270450.0 ;
      RECT  104100.0 269250.0 102900.0 270450.0 ;
      RECT  106500.0 260550.0 105300.0 261750.0 ;
      RECT  104100.0 260550.0 102900.0 261750.0 ;
      RECT  104100.0 260550.0 102900.0 261750.0 ;
      RECT  106500.0 260550.0 105300.0 261750.0 ;
      RECT  104100.0 260550.0 102900.0 261750.0 ;
      RECT  101700.0 260550.0 100500.0 261750.0 ;
      RECT  101700.0 260550.0 100500.0 261750.0 ;
      RECT  104100.0 260550.0 102900.0 261750.0 ;
      RECT  99300.0 269850.0 98100.0 271050.0 ;
      RECT  99300.0 259950.0 98100.0 261150.0 ;
      RECT  101700.0 263100.0 102900.0 264300.0 ;
      RECT  104700.0 265800.0 105900.0 267000.0 ;
      RECT  104100.0 269250.0 102900.0 270450.0 ;
      RECT  101700.0 260550.0 100500.0 261750.0 ;
      RECT  100500.0 265800.0 101700.0 267000.0 ;
      RECT  105900.0 265800.0 104700.0 267000.0 ;
      RECT  102900.0 263100.0 101700.0 264300.0 ;
      RECT  101700.0 265800.0 100500.0 267000.0 ;
      RECT  108300.0 271950.0 93900.0 272850.0 ;
      RECT  108300.0 258150.0 93900.0 259050.0 ;
      RECT  106500.0 284250.0 105300.0 286650.0 ;
      RECT  106500.0 275550.0 105300.0 271950.0 ;
      RECT  101700.0 275550.0 100500.0 271950.0 ;
      RECT  99300.0 274350.0 98100.0 272400.0 ;
      RECT  99300.0 286200.0 98100.0 284250.0 ;
      RECT  106500.0 275550.0 105300.0 274350.0 ;
      RECT  104100.0 275550.0 102900.0 274350.0 ;
      RECT  104100.0 275550.0 102900.0 274350.0 ;
      RECT  106500.0 275550.0 105300.0 274350.0 ;
      RECT  104100.0 275550.0 102900.0 274350.0 ;
      RECT  101700.0 275550.0 100500.0 274350.0 ;
      RECT  101700.0 275550.0 100500.0 274350.0 ;
      RECT  104100.0 275550.0 102900.0 274350.0 ;
      RECT  106500.0 284250.0 105300.0 283050.0 ;
      RECT  104100.0 284250.0 102900.0 283050.0 ;
      RECT  104100.0 284250.0 102900.0 283050.0 ;
      RECT  106500.0 284250.0 105300.0 283050.0 ;
      RECT  104100.0 284250.0 102900.0 283050.0 ;
      RECT  101700.0 284250.0 100500.0 283050.0 ;
      RECT  101700.0 284250.0 100500.0 283050.0 ;
      RECT  104100.0 284250.0 102900.0 283050.0 ;
      RECT  99300.0 274950.0 98100.0 273750.0 ;
      RECT  99300.0 284850.0 98100.0 283650.0 ;
      RECT  101700.0 281700.0 102900.0 280500.0 ;
      RECT  104700.0 279000.0 105900.0 277800.0 ;
      RECT  104100.0 275550.0 102900.0 274350.0 ;
      RECT  101700.0 284250.0 100500.0 283050.0 ;
      RECT  100500.0 279000.0 101700.0 277800.0 ;
      RECT  105900.0 279000.0 104700.0 277800.0 ;
      RECT  102900.0 281700.0 101700.0 280500.0 ;
      RECT  101700.0 279000.0 100500.0 277800.0 ;
      RECT  108300.0 272850.0 93900.0 271950.0 ;
      RECT  108300.0 286650.0 93900.0 285750.0 ;
      RECT  106500.0 288150.0 105300.0 285750.0 ;
      RECT  106500.0 296850.0 105300.0 300450.0 ;
      RECT  101700.0 296850.0 100500.0 300450.0 ;
      RECT  99300.0 298050.0 98100.0 300000.0 ;
      RECT  99300.0 286200.0 98100.0 288150.0 ;
      RECT  106500.0 296850.0 105300.0 298050.0 ;
      RECT  104100.0 296850.0 102900.0 298050.0 ;
      RECT  104100.0 296850.0 102900.0 298050.0 ;
      RECT  106500.0 296850.0 105300.0 298050.0 ;
      RECT  104100.0 296850.0 102900.0 298050.0 ;
      RECT  101700.0 296850.0 100500.0 298050.0 ;
      RECT  101700.0 296850.0 100500.0 298050.0 ;
      RECT  104100.0 296850.0 102900.0 298050.0 ;
      RECT  106500.0 288150.0 105300.0 289350.0 ;
      RECT  104100.0 288150.0 102900.0 289350.0 ;
      RECT  104100.0 288150.0 102900.0 289350.0 ;
      RECT  106500.0 288150.0 105300.0 289350.0 ;
      RECT  104100.0 288150.0 102900.0 289350.0 ;
      RECT  101700.0 288150.0 100500.0 289350.0 ;
      RECT  101700.0 288150.0 100500.0 289350.0 ;
      RECT  104100.0 288150.0 102900.0 289350.0 ;
      RECT  99300.0 297450.0 98100.0 298650.0 ;
      RECT  99300.0 287550.0 98100.0 288750.0 ;
      RECT  101700.0 290700.0 102900.0 291900.0 ;
      RECT  104700.0 293400.0 105900.0 294600.0 ;
      RECT  104100.0 296850.0 102900.0 298050.0 ;
      RECT  101700.0 288150.0 100500.0 289350.0 ;
      RECT  100500.0 293400.0 101700.0 294600.0 ;
      RECT  105900.0 293400.0 104700.0 294600.0 ;
      RECT  102900.0 290700.0 101700.0 291900.0 ;
      RECT  101700.0 293400.0 100500.0 294600.0 ;
      RECT  108300.0 299550.0 93900.0 300450.0 ;
      RECT  108300.0 285750.0 93900.0 286650.0 ;
      RECT  106500.0 311850.0 105300.0 314250.0 ;
      RECT  106500.0 303150.0 105300.0 299550.0 ;
      RECT  101700.0 303150.0 100500.0 299550.0 ;
      RECT  99300.0 301950.0 98100.0 300000.0 ;
      RECT  99300.0 313800.0 98100.0 311850.0 ;
      RECT  106500.0 303150.0 105300.0 301950.0 ;
      RECT  104100.0 303150.0 102900.0 301950.0 ;
      RECT  104100.0 303150.0 102900.0 301950.0 ;
      RECT  106500.0 303150.0 105300.0 301950.0 ;
      RECT  104100.0 303150.0 102900.0 301950.0 ;
      RECT  101700.0 303150.0 100500.0 301950.0 ;
      RECT  101700.0 303150.0 100500.0 301950.0 ;
      RECT  104100.0 303150.0 102900.0 301950.0 ;
      RECT  106500.0 311850.0 105300.0 310650.0 ;
      RECT  104100.0 311850.0 102900.0 310650.0 ;
      RECT  104100.0 311850.0 102900.0 310650.0 ;
      RECT  106500.0 311850.0 105300.0 310650.0 ;
      RECT  104100.0 311850.0 102900.0 310650.0 ;
      RECT  101700.0 311850.0 100500.0 310650.0 ;
      RECT  101700.0 311850.0 100500.0 310650.0 ;
      RECT  104100.0 311850.0 102900.0 310650.0 ;
      RECT  99300.0 302550.0 98100.0 301350.0 ;
      RECT  99300.0 312450.0 98100.0 311250.0 ;
      RECT  101700.0 309300.0 102900.0 308100.0 ;
      RECT  104700.0 306600.0 105900.0 305400.0 ;
      RECT  104100.0 303150.0 102900.0 301950.0 ;
      RECT  101700.0 311850.0 100500.0 310650.0 ;
      RECT  100500.0 306600.0 101700.0 305400.0 ;
      RECT  105900.0 306600.0 104700.0 305400.0 ;
      RECT  102900.0 309300.0 101700.0 308100.0 ;
      RECT  101700.0 306600.0 100500.0 305400.0 ;
      RECT  108300.0 300450.0 93900.0 299550.0 ;
      RECT  108300.0 314250.0 93900.0 313350.0 ;
      RECT  119250.0 269100.0 120450.0 270300.0 ;
      RECT  137850.0 264600.0 139050.0 265800.0 ;
      RECT  116250.0 282900.0 117450.0 284100.0 ;
      RECT  134850.0 279000.0 136050.0 280200.0 ;
      RECT  137850.0 287700.0 139050.0 288900.0 ;
      RECT  113250.0 287700.0 114450.0 288900.0 ;
      RECT  134850.0 301500.0 136050.0 302700.0 ;
      RECT  110250.0 301500.0 111450.0 302700.0 ;
      RECT  119250.0 265800.0 120450.0 267000.0 ;
      RECT  116250.0 263100.0 117450.0 264300.0 ;
      RECT  113250.0 277800.0 114450.0 279000.0 ;
      RECT  116250.0 280500.0 117450.0 281700.0 ;
      RECT  119250.0 293400.0 120450.0 294600.0 ;
      RECT  110250.0 290700.0 111450.0 291900.0 ;
      RECT  113250.0 305400.0 114450.0 306600.0 ;
      RECT  110250.0 308100.0 111450.0 309300.0 ;
      RECT  88050.0 264750.0 84300.0 265650.0 ;
      RECT  88050.0 279150.0 84300.0 280050.0 ;
      RECT  88050.0 292350.0 84300.0 293250.0 ;
      RECT  88050.0 306750.0 84300.0 307650.0 ;
      RECT  138900.0 271950.0 84300.0 272850.0 ;
      RECT  138900.0 299550.0 84300.0 300450.0 ;
      RECT  138900.0 258150.0 84300.0 259050.0 ;
      RECT  138900.0 285750.0 84300.0 286650.0 ;
      RECT  138900.0 313350.0 84300.0 314250.0 ;
      RECT  86100.0 315750.0 87300.0 313350.0 ;
      RECT  86100.0 324450.0 87300.0 328050.0 ;
      RECT  90900.0 324450.0 92100.0 328050.0 ;
      RECT  95700.0 325650.0 96900.0 327600.0 ;
      RECT  95700.0 313800.0 96900.0 315750.0 ;
      RECT  86100.0 324450.0 87300.0 325650.0 ;
      RECT  88500.0 324450.0 89700.0 325650.0 ;
      RECT  88500.0 324450.0 89700.0 325650.0 ;
      RECT  86100.0 324450.0 87300.0 325650.0 ;
      RECT  88500.0 324450.0 89700.0 325650.0 ;
      RECT  90900.0 324450.0 92100.0 325650.0 ;
      RECT  90900.0 324450.0 92100.0 325650.0 ;
      RECT  88500.0 324450.0 89700.0 325650.0 ;
      RECT  90900.0 324450.0 92100.0 325650.0 ;
      RECT  93300.0 324450.0 94500.0 325650.0 ;
      RECT  93300.0 324450.0 94500.0 325650.0 ;
      RECT  90900.0 324450.0 92100.0 325650.0 ;
      RECT  86100.0 315750.0 87300.0 316950.0 ;
      RECT  88500.0 315750.0 89700.0 316950.0 ;
      RECT  88500.0 315750.0 89700.0 316950.0 ;
      RECT  86100.0 315750.0 87300.0 316950.0 ;
      RECT  88500.0 315750.0 89700.0 316950.0 ;
      RECT  90900.0 315750.0 92100.0 316950.0 ;
      RECT  90900.0 315750.0 92100.0 316950.0 ;
      RECT  88500.0 315750.0 89700.0 316950.0 ;
      RECT  90900.0 315750.0 92100.0 316950.0 ;
      RECT  93300.0 315750.0 94500.0 316950.0 ;
      RECT  93300.0 315750.0 94500.0 316950.0 ;
      RECT  90900.0 315750.0 92100.0 316950.0 ;
      RECT  95700.0 325050.0 96900.0 326250.0 ;
      RECT  95700.0 315150.0 96900.0 316350.0 ;
      RECT  93300.0 317850.0 92100.0 319050.0 ;
      RECT  90900.0 319800.0 89700.0 321000.0 ;
      RECT  88500.0 321750.0 87300.0 322950.0 ;
      RECT  88500.0 324450.0 89700.0 325650.0 ;
      RECT  93300.0 324450.0 94500.0 325650.0 ;
      RECT  93300.0 315750.0 94500.0 316950.0 ;
      RECT  93300.0 321750.0 94500.0 322950.0 ;
      RECT  87300.0 321750.0 88500.0 322950.0 ;
      RECT  89700.0 319800.0 90900.0 321000.0 ;
      RECT  92100.0 317850.0 93300.0 319050.0 ;
      RECT  93300.0 321750.0 94500.0 322950.0 ;
      RECT  84300.0 327150.0 99900.0 328050.0 ;
      RECT  84300.0 313350.0 99900.0 314250.0 ;
      RECT  86100.0 339450.0 87300.0 341850.0 ;
      RECT  86100.0 330750.0 87300.0 327150.0 ;
      RECT  90900.0 330750.0 92100.0 327150.0 ;
      RECT  95700.0 329550.0 96900.0 327600.0 ;
      RECT  95700.0 341400.0 96900.0 339450.0 ;
      RECT  86100.0 330750.0 87300.0 329550.0 ;
      RECT  88500.0 330750.0 89700.0 329550.0 ;
      RECT  88500.0 330750.0 89700.0 329550.0 ;
      RECT  86100.0 330750.0 87300.0 329550.0 ;
      RECT  88500.0 330750.0 89700.0 329550.0 ;
      RECT  90900.0 330750.0 92100.0 329550.0 ;
      RECT  90900.0 330750.0 92100.0 329550.0 ;
      RECT  88500.0 330750.0 89700.0 329550.0 ;
      RECT  90900.0 330750.0 92100.0 329550.0 ;
      RECT  93300.0 330750.0 94500.0 329550.0 ;
      RECT  93300.0 330750.0 94500.0 329550.0 ;
      RECT  90900.0 330750.0 92100.0 329550.0 ;
      RECT  86100.0 339450.0 87300.0 338250.0 ;
      RECT  88500.0 339450.0 89700.0 338250.0 ;
      RECT  88500.0 339450.0 89700.0 338250.0 ;
      RECT  86100.0 339450.0 87300.0 338250.0 ;
      RECT  88500.0 339450.0 89700.0 338250.0 ;
      RECT  90900.0 339450.0 92100.0 338250.0 ;
      RECT  90900.0 339450.0 92100.0 338250.0 ;
      RECT  88500.0 339450.0 89700.0 338250.0 ;
      RECT  90900.0 339450.0 92100.0 338250.0 ;
      RECT  93300.0 339450.0 94500.0 338250.0 ;
      RECT  93300.0 339450.0 94500.0 338250.0 ;
      RECT  90900.0 339450.0 92100.0 338250.0 ;
      RECT  95700.0 330150.0 96900.0 328950.0 ;
      RECT  95700.0 340050.0 96900.0 338850.0 ;
      RECT  93300.0 337350.0 92100.0 336150.0 ;
      RECT  90900.0 335400.0 89700.0 334200.0 ;
      RECT  88500.0 333450.0 87300.0 332250.0 ;
      RECT  88500.0 330750.0 89700.0 329550.0 ;
      RECT  93300.0 330750.0 94500.0 329550.0 ;
      RECT  93300.0 339450.0 94500.0 338250.0 ;
      RECT  93300.0 333450.0 94500.0 332250.0 ;
      RECT  87300.0 333450.0 88500.0 332250.0 ;
      RECT  89700.0 335400.0 90900.0 334200.0 ;
      RECT  92100.0 337350.0 93300.0 336150.0 ;
      RECT  93300.0 333450.0 94500.0 332250.0 ;
      RECT  84300.0 328050.0 99900.0 327150.0 ;
      RECT  84300.0 341850.0 99900.0 340950.0 ;
      RECT  86100.0 343350.0 87300.0 340950.0 ;
      RECT  86100.0 352050.0 87300.0 355650.0 ;
      RECT  90900.0 352050.0 92100.0 355650.0 ;
      RECT  95700.0 353250.0 96900.0 355200.0 ;
      RECT  95700.0 341400.0 96900.0 343350.0 ;
      RECT  86100.0 352050.0 87300.0 353250.0 ;
      RECT  88500.0 352050.0 89700.0 353250.0 ;
      RECT  88500.0 352050.0 89700.0 353250.0 ;
      RECT  86100.0 352050.0 87300.0 353250.0 ;
      RECT  88500.0 352050.0 89700.0 353250.0 ;
      RECT  90900.0 352050.0 92100.0 353250.0 ;
      RECT  90900.0 352050.0 92100.0 353250.0 ;
      RECT  88500.0 352050.0 89700.0 353250.0 ;
      RECT  90900.0 352050.0 92100.0 353250.0 ;
      RECT  93300.0 352050.0 94500.0 353250.0 ;
      RECT  93300.0 352050.0 94500.0 353250.0 ;
      RECT  90900.0 352050.0 92100.0 353250.0 ;
      RECT  86100.0 343350.0 87300.0 344550.0 ;
      RECT  88500.0 343350.0 89700.0 344550.0 ;
      RECT  88500.0 343350.0 89700.0 344550.0 ;
      RECT  86100.0 343350.0 87300.0 344550.0 ;
      RECT  88500.0 343350.0 89700.0 344550.0 ;
      RECT  90900.0 343350.0 92100.0 344550.0 ;
      RECT  90900.0 343350.0 92100.0 344550.0 ;
      RECT  88500.0 343350.0 89700.0 344550.0 ;
      RECT  90900.0 343350.0 92100.0 344550.0 ;
      RECT  93300.0 343350.0 94500.0 344550.0 ;
      RECT  93300.0 343350.0 94500.0 344550.0 ;
      RECT  90900.0 343350.0 92100.0 344550.0 ;
      RECT  95700.0 352650.0 96900.0 353850.0 ;
      RECT  95700.0 342750.0 96900.0 343950.0 ;
      RECT  93300.0 345450.0 92100.0 346650.0 ;
      RECT  90900.0 347400.0 89700.0 348600.0 ;
      RECT  88500.0 349350.0 87300.0 350550.0 ;
      RECT  88500.0 352050.0 89700.0 353250.0 ;
      RECT  93300.0 352050.0 94500.0 353250.0 ;
      RECT  93300.0 343350.0 94500.0 344550.0 ;
      RECT  93300.0 349350.0 94500.0 350550.0 ;
      RECT  87300.0 349350.0 88500.0 350550.0 ;
      RECT  89700.0 347400.0 90900.0 348600.0 ;
      RECT  92100.0 345450.0 93300.0 346650.0 ;
      RECT  93300.0 349350.0 94500.0 350550.0 ;
      RECT  84300.0 354750.0 99900.0 355650.0 ;
      RECT  84300.0 340950.0 99900.0 341850.0 ;
      RECT  86100.0 367050.0 87300.0 369450.0 ;
      RECT  86100.0 358350.0 87300.0 354750.0 ;
      RECT  90900.0 358350.0 92100.0 354750.0 ;
      RECT  95700.0 357150.0 96900.0 355200.0 ;
      RECT  95700.0 369000.0 96900.0 367050.0 ;
      RECT  86100.0 358350.0 87300.0 357150.0 ;
      RECT  88500.0 358350.0 89700.0 357150.0 ;
      RECT  88500.0 358350.0 89700.0 357150.0 ;
      RECT  86100.0 358350.0 87300.0 357150.0 ;
      RECT  88500.0 358350.0 89700.0 357150.0 ;
      RECT  90900.0 358350.0 92100.0 357150.0 ;
      RECT  90900.0 358350.0 92100.0 357150.0 ;
      RECT  88500.0 358350.0 89700.0 357150.0 ;
      RECT  90900.0 358350.0 92100.0 357150.0 ;
      RECT  93300.0 358350.0 94500.0 357150.0 ;
      RECT  93300.0 358350.0 94500.0 357150.0 ;
      RECT  90900.0 358350.0 92100.0 357150.0 ;
      RECT  86100.0 367050.0 87300.0 365850.0 ;
      RECT  88500.0 367050.0 89700.0 365850.0 ;
      RECT  88500.0 367050.0 89700.0 365850.0 ;
      RECT  86100.0 367050.0 87300.0 365850.0 ;
      RECT  88500.0 367050.0 89700.0 365850.0 ;
      RECT  90900.0 367050.0 92100.0 365850.0 ;
      RECT  90900.0 367050.0 92100.0 365850.0 ;
      RECT  88500.0 367050.0 89700.0 365850.0 ;
      RECT  90900.0 367050.0 92100.0 365850.0 ;
      RECT  93300.0 367050.0 94500.0 365850.0 ;
      RECT  93300.0 367050.0 94500.0 365850.0 ;
      RECT  90900.0 367050.0 92100.0 365850.0 ;
      RECT  95700.0 357750.0 96900.0 356550.0 ;
      RECT  95700.0 367650.0 96900.0 366450.0 ;
      RECT  93300.0 364950.0 92100.0 363750.0 ;
      RECT  90900.0 363000.0 89700.0 361800.0 ;
      RECT  88500.0 361050.0 87300.0 359850.0 ;
      RECT  88500.0 358350.0 89700.0 357150.0 ;
      RECT  93300.0 358350.0 94500.0 357150.0 ;
      RECT  93300.0 367050.0 94500.0 365850.0 ;
      RECT  93300.0 361050.0 94500.0 359850.0 ;
      RECT  87300.0 361050.0 88500.0 359850.0 ;
      RECT  89700.0 363000.0 90900.0 361800.0 ;
      RECT  92100.0 364950.0 93300.0 363750.0 ;
      RECT  93300.0 361050.0 94500.0 359850.0 ;
      RECT  84300.0 355650.0 99900.0 354750.0 ;
      RECT  84300.0 369450.0 99900.0 368550.0 ;
      RECT  86100.0 370950.0 87300.0 368550.0 ;
      RECT  86100.0 379650.0 87300.0 383250.0 ;
      RECT  90900.0 379650.0 92100.0 383250.0 ;
      RECT  95700.0 380850.0 96900.0 382800.0 ;
      RECT  95700.0 369000.0 96900.0 370950.0 ;
      RECT  86100.0 379650.0 87300.0 380850.0 ;
      RECT  88500.0 379650.0 89700.0 380850.0 ;
      RECT  88500.0 379650.0 89700.0 380850.0 ;
      RECT  86100.0 379650.0 87300.0 380850.0 ;
      RECT  88500.0 379650.0 89700.0 380850.0 ;
      RECT  90900.0 379650.0 92100.0 380850.0 ;
      RECT  90900.0 379650.0 92100.0 380850.0 ;
      RECT  88500.0 379650.0 89700.0 380850.0 ;
      RECT  90900.0 379650.0 92100.0 380850.0 ;
      RECT  93300.0 379650.0 94500.0 380850.0 ;
      RECT  93300.0 379650.0 94500.0 380850.0 ;
      RECT  90900.0 379650.0 92100.0 380850.0 ;
      RECT  86100.0 370950.0 87300.0 372150.0 ;
      RECT  88500.0 370950.0 89700.0 372150.0 ;
      RECT  88500.0 370950.0 89700.0 372150.0 ;
      RECT  86100.0 370950.0 87300.0 372150.0 ;
      RECT  88500.0 370950.0 89700.0 372150.0 ;
      RECT  90900.0 370950.0 92100.0 372150.0 ;
      RECT  90900.0 370950.0 92100.0 372150.0 ;
      RECT  88500.0 370950.0 89700.0 372150.0 ;
      RECT  90900.0 370950.0 92100.0 372150.0 ;
      RECT  93300.0 370950.0 94500.0 372150.0 ;
      RECT  93300.0 370950.0 94500.0 372150.0 ;
      RECT  90900.0 370950.0 92100.0 372150.0 ;
      RECT  95700.0 380250.0 96900.0 381450.0 ;
      RECT  95700.0 370350.0 96900.0 371550.0 ;
      RECT  93300.0 373050.0 92100.0 374250.0 ;
      RECT  90900.0 375000.0 89700.0 376200.0 ;
      RECT  88500.0 376950.0 87300.0 378150.0 ;
      RECT  88500.0 379650.0 89700.0 380850.0 ;
      RECT  93300.0 379650.0 94500.0 380850.0 ;
      RECT  93300.0 370950.0 94500.0 372150.0 ;
      RECT  93300.0 376950.0 94500.0 378150.0 ;
      RECT  87300.0 376950.0 88500.0 378150.0 ;
      RECT  89700.0 375000.0 90900.0 376200.0 ;
      RECT  92100.0 373050.0 93300.0 374250.0 ;
      RECT  93300.0 376950.0 94500.0 378150.0 ;
      RECT  84300.0 382350.0 99900.0 383250.0 ;
      RECT  84300.0 368550.0 99900.0 369450.0 ;
      RECT  86100.0 394650.0 87300.0 397050.0 ;
      RECT  86100.0 385950.0 87300.0 382350.0 ;
      RECT  90900.0 385950.0 92100.0 382350.0 ;
      RECT  95700.0 384750.0 96900.0 382800.0 ;
      RECT  95700.0 396600.0 96900.0 394650.0 ;
      RECT  86100.0 385950.0 87300.0 384750.0 ;
      RECT  88500.0 385950.0 89700.0 384750.0 ;
      RECT  88500.0 385950.0 89700.0 384750.0 ;
      RECT  86100.0 385950.0 87300.0 384750.0 ;
      RECT  88500.0 385950.0 89700.0 384750.0 ;
      RECT  90900.0 385950.0 92100.0 384750.0 ;
      RECT  90900.0 385950.0 92100.0 384750.0 ;
      RECT  88500.0 385950.0 89700.0 384750.0 ;
      RECT  90900.0 385950.0 92100.0 384750.0 ;
      RECT  93300.0 385950.0 94500.0 384750.0 ;
      RECT  93300.0 385950.0 94500.0 384750.0 ;
      RECT  90900.0 385950.0 92100.0 384750.0 ;
      RECT  86100.0 394650.0 87300.0 393450.0 ;
      RECT  88500.0 394650.0 89700.0 393450.0 ;
      RECT  88500.0 394650.0 89700.0 393450.0 ;
      RECT  86100.0 394650.0 87300.0 393450.0 ;
      RECT  88500.0 394650.0 89700.0 393450.0 ;
      RECT  90900.0 394650.0 92100.0 393450.0 ;
      RECT  90900.0 394650.0 92100.0 393450.0 ;
      RECT  88500.0 394650.0 89700.0 393450.0 ;
      RECT  90900.0 394650.0 92100.0 393450.0 ;
      RECT  93300.0 394650.0 94500.0 393450.0 ;
      RECT  93300.0 394650.0 94500.0 393450.0 ;
      RECT  90900.0 394650.0 92100.0 393450.0 ;
      RECT  95700.0 385350.0 96900.0 384150.0 ;
      RECT  95700.0 395250.0 96900.0 394050.0 ;
      RECT  93300.0 392550.0 92100.0 391350.0 ;
      RECT  90900.0 390600.0 89700.0 389400.0 ;
      RECT  88500.0 388650.0 87300.0 387450.0 ;
      RECT  88500.0 385950.0 89700.0 384750.0 ;
      RECT  93300.0 385950.0 94500.0 384750.0 ;
      RECT  93300.0 394650.0 94500.0 393450.0 ;
      RECT  93300.0 388650.0 94500.0 387450.0 ;
      RECT  87300.0 388650.0 88500.0 387450.0 ;
      RECT  89700.0 390600.0 90900.0 389400.0 ;
      RECT  92100.0 392550.0 93300.0 391350.0 ;
      RECT  93300.0 388650.0 94500.0 387450.0 ;
      RECT  84300.0 383250.0 99900.0 382350.0 ;
      RECT  84300.0 397050.0 99900.0 396150.0 ;
      RECT  86100.0 398550.0 87300.0 396150.0 ;
      RECT  86100.0 407250.0 87300.0 410850.0 ;
      RECT  90900.0 407250.0 92100.0 410850.0 ;
      RECT  95700.0 408450.0 96900.0 410400.0 ;
      RECT  95700.0 396600.0 96900.0 398550.0 ;
      RECT  86100.0 407250.0 87300.0 408450.0 ;
      RECT  88500.0 407250.0 89700.0 408450.0 ;
      RECT  88500.0 407250.0 89700.0 408450.0 ;
      RECT  86100.0 407250.0 87300.0 408450.0 ;
      RECT  88500.0 407250.0 89700.0 408450.0 ;
      RECT  90900.0 407250.0 92100.0 408450.0 ;
      RECT  90900.0 407250.0 92100.0 408450.0 ;
      RECT  88500.0 407250.0 89700.0 408450.0 ;
      RECT  90900.0 407250.0 92100.0 408450.0 ;
      RECT  93300.0 407250.0 94500.0 408450.0 ;
      RECT  93300.0 407250.0 94500.0 408450.0 ;
      RECT  90900.0 407250.0 92100.0 408450.0 ;
      RECT  86100.0 398550.0 87300.0 399750.0 ;
      RECT  88500.0 398550.0 89700.0 399750.0 ;
      RECT  88500.0 398550.0 89700.0 399750.0 ;
      RECT  86100.0 398550.0 87300.0 399750.0 ;
      RECT  88500.0 398550.0 89700.0 399750.0 ;
      RECT  90900.0 398550.0 92100.0 399750.0 ;
      RECT  90900.0 398550.0 92100.0 399750.0 ;
      RECT  88500.0 398550.0 89700.0 399750.0 ;
      RECT  90900.0 398550.0 92100.0 399750.0 ;
      RECT  93300.0 398550.0 94500.0 399750.0 ;
      RECT  93300.0 398550.0 94500.0 399750.0 ;
      RECT  90900.0 398550.0 92100.0 399750.0 ;
      RECT  95700.0 407850.0 96900.0 409050.0 ;
      RECT  95700.0 397950.0 96900.0 399150.0 ;
      RECT  93300.0 400650.0 92100.0 401850.0 ;
      RECT  90900.0 402600.0 89700.0 403800.0 ;
      RECT  88500.0 404550.0 87300.0 405750.0 ;
      RECT  88500.0 407250.0 89700.0 408450.0 ;
      RECT  93300.0 407250.0 94500.0 408450.0 ;
      RECT  93300.0 398550.0 94500.0 399750.0 ;
      RECT  93300.0 404550.0 94500.0 405750.0 ;
      RECT  87300.0 404550.0 88500.0 405750.0 ;
      RECT  89700.0 402600.0 90900.0 403800.0 ;
      RECT  92100.0 400650.0 93300.0 401850.0 ;
      RECT  93300.0 404550.0 94500.0 405750.0 ;
      RECT  84300.0 409950.0 99900.0 410850.0 ;
      RECT  84300.0 396150.0 99900.0 397050.0 ;
      RECT  86100.0 422250.0 87300.0 424650.0 ;
      RECT  86100.0 413550.0 87300.0 409950.0 ;
      RECT  90900.0 413550.0 92100.0 409950.0 ;
      RECT  95700.0 412350.0 96900.0 410400.0 ;
      RECT  95700.0 424200.0 96900.0 422250.0 ;
      RECT  86100.0 413550.0 87300.0 412350.0 ;
      RECT  88500.0 413550.0 89700.0 412350.0 ;
      RECT  88500.0 413550.0 89700.0 412350.0 ;
      RECT  86100.0 413550.0 87300.0 412350.0 ;
      RECT  88500.0 413550.0 89700.0 412350.0 ;
      RECT  90900.0 413550.0 92100.0 412350.0 ;
      RECT  90900.0 413550.0 92100.0 412350.0 ;
      RECT  88500.0 413550.0 89700.0 412350.0 ;
      RECT  90900.0 413550.0 92100.0 412350.0 ;
      RECT  93300.0 413550.0 94500.0 412350.0 ;
      RECT  93300.0 413550.0 94500.0 412350.0 ;
      RECT  90900.0 413550.0 92100.0 412350.0 ;
      RECT  86100.0 422250.0 87300.0 421050.0 ;
      RECT  88500.0 422250.0 89700.0 421050.0 ;
      RECT  88500.0 422250.0 89700.0 421050.0 ;
      RECT  86100.0 422250.0 87300.0 421050.0 ;
      RECT  88500.0 422250.0 89700.0 421050.0 ;
      RECT  90900.0 422250.0 92100.0 421050.0 ;
      RECT  90900.0 422250.0 92100.0 421050.0 ;
      RECT  88500.0 422250.0 89700.0 421050.0 ;
      RECT  90900.0 422250.0 92100.0 421050.0 ;
      RECT  93300.0 422250.0 94500.0 421050.0 ;
      RECT  93300.0 422250.0 94500.0 421050.0 ;
      RECT  90900.0 422250.0 92100.0 421050.0 ;
      RECT  95700.0 412950.0 96900.0 411750.0 ;
      RECT  95700.0 422850.0 96900.0 421650.0 ;
      RECT  93300.0 420150.0 92100.0 418950.0 ;
      RECT  90900.0 418200.0 89700.0 417000.0 ;
      RECT  88500.0 416250.0 87300.0 415050.0 ;
      RECT  88500.0 413550.0 89700.0 412350.0 ;
      RECT  93300.0 413550.0 94500.0 412350.0 ;
      RECT  93300.0 422250.0 94500.0 421050.0 ;
      RECT  93300.0 416250.0 94500.0 415050.0 ;
      RECT  87300.0 416250.0 88500.0 415050.0 ;
      RECT  89700.0 418200.0 90900.0 417000.0 ;
      RECT  92100.0 420150.0 93300.0 418950.0 ;
      RECT  93300.0 416250.0 94500.0 415050.0 ;
      RECT  84300.0 410850.0 99900.0 409950.0 ;
      RECT  84300.0 424650.0 99900.0 423750.0 ;
      RECT  86100.0 426150.0 87300.0 423750.0 ;
      RECT  86100.0 434850.0 87300.0 438450.0 ;
      RECT  90900.0 434850.0 92100.0 438450.0 ;
      RECT  95700.0 436050.0 96900.0 438000.0 ;
      RECT  95700.0 424200.0 96900.0 426150.0 ;
      RECT  86100.0 434850.0 87300.0 436050.0 ;
      RECT  88500.0 434850.0 89700.0 436050.0 ;
      RECT  88500.0 434850.0 89700.0 436050.0 ;
      RECT  86100.0 434850.0 87300.0 436050.0 ;
      RECT  88500.0 434850.0 89700.0 436050.0 ;
      RECT  90900.0 434850.0 92100.0 436050.0 ;
      RECT  90900.0 434850.0 92100.0 436050.0 ;
      RECT  88500.0 434850.0 89700.0 436050.0 ;
      RECT  90900.0 434850.0 92100.0 436050.0 ;
      RECT  93300.0 434850.0 94500.0 436050.0 ;
      RECT  93300.0 434850.0 94500.0 436050.0 ;
      RECT  90900.0 434850.0 92100.0 436050.0 ;
      RECT  86100.0 426150.0 87300.0 427350.0 ;
      RECT  88500.0 426150.0 89700.0 427350.0 ;
      RECT  88500.0 426150.0 89700.0 427350.0 ;
      RECT  86100.0 426150.0 87300.0 427350.0 ;
      RECT  88500.0 426150.0 89700.0 427350.0 ;
      RECT  90900.0 426150.0 92100.0 427350.0 ;
      RECT  90900.0 426150.0 92100.0 427350.0 ;
      RECT  88500.0 426150.0 89700.0 427350.0 ;
      RECT  90900.0 426150.0 92100.0 427350.0 ;
      RECT  93300.0 426150.0 94500.0 427350.0 ;
      RECT  93300.0 426150.0 94500.0 427350.0 ;
      RECT  90900.0 426150.0 92100.0 427350.0 ;
      RECT  95700.0 435450.0 96900.0 436650.0 ;
      RECT  95700.0 425550.0 96900.0 426750.0 ;
      RECT  93300.0 428250.0 92100.0 429450.0 ;
      RECT  90900.0 430200.0 89700.0 431400.0 ;
      RECT  88500.0 432150.0 87300.0 433350.0 ;
      RECT  88500.0 434850.0 89700.0 436050.0 ;
      RECT  93300.0 434850.0 94500.0 436050.0 ;
      RECT  93300.0 426150.0 94500.0 427350.0 ;
      RECT  93300.0 432150.0 94500.0 433350.0 ;
      RECT  87300.0 432150.0 88500.0 433350.0 ;
      RECT  89700.0 430200.0 90900.0 431400.0 ;
      RECT  92100.0 428250.0 93300.0 429450.0 ;
      RECT  93300.0 432150.0 94500.0 433350.0 ;
      RECT  84300.0 437550.0 99900.0 438450.0 ;
      RECT  84300.0 423750.0 99900.0 424650.0 ;
      RECT  86100.0 449850.0 87300.0 452250.0 ;
      RECT  86100.0 441150.0 87300.0 437550.0 ;
      RECT  90900.0 441150.0 92100.0 437550.0 ;
      RECT  95700.0 439950.0 96900.0 438000.0 ;
      RECT  95700.0 451800.0 96900.0 449850.0 ;
      RECT  86100.0 441150.0 87300.0 439950.0 ;
      RECT  88500.0 441150.0 89700.0 439950.0 ;
      RECT  88500.0 441150.0 89700.0 439950.0 ;
      RECT  86100.0 441150.0 87300.0 439950.0 ;
      RECT  88500.0 441150.0 89700.0 439950.0 ;
      RECT  90900.0 441150.0 92100.0 439950.0 ;
      RECT  90900.0 441150.0 92100.0 439950.0 ;
      RECT  88500.0 441150.0 89700.0 439950.0 ;
      RECT  90900.0 441150.0 92100.0 439950.0 ;
      RECT  93300.0 441150.0 94500.0 439950.0 ;
      RECT  93300.0 441150.0 94500.0 439950.0 ;
      RECT  90900.0 441150.0 92100.0 439950.0 ;
      RECT  86100.0 449850.0 87300.0 448650.0 ;
      RECT  88500.0 449850.0 89700.0 448650.0 ;
      RECT  88500.0 449850.0 89700.0 448650.0 ;
      RECT  86100.0 449850.0 87300.0 448650.0 ;
      RECT  88500.0 449850.0 89700.0 448650.0 ;
      RECT  90900.0 449850.0 92100.0 448650.0 ;
      RECT  90900.0 449850.0 92100.0 448650.0 ;
      RECT  88500.0 449850.0 89700.0 448650.0 ;
      RECT  90900.0 449850.0 92100.0 448650.0 ;
      RECT  93300.0 449850.0 94500.0 448650.0 ;
      RECT  93300.0 449850.0 94500.0 448650.0 ;
      RECT  90900.0 449850.0 92100.0 448650.0 ;
      RECT  95700.0 440550.0 96900.0 439350.0 ;
      RECT  95700.0 450450.0 96900.0 449250.0 ;
      RECT  93300.0 447750.0 92100.0 446550.0 ;
      RECT  90900.0 445800.0 89700.0 444600.0 ;
      RECT  88500.0 443850.0 87300.0 442650.0 ;
      RECT  88500.0 441150.0 89700.0 439950.0 ;
      RECT  93300.0 441150.0 94500.0 439950.0 ;
      RECT  93300.0 449850.0 94500.0 448650.0 ;
      RECT  93300.0 443850.0 94500.0 442650.0 ;
      RECT  87300.0 443850.0 88500.0 442650.0 ;
      RECT  89700.0 445800.0 90900.0 444600.0 ;
      RECT  92100.0 447750.0 93300.0 446550.0 ;
      RECT  93300.0 443850.0 94500.0 442650.0 ;
      RECT  84300.0 438450.0 99900.0 437550.0 ;
      RECT  84300.0 452250.0 99900.0 451350.0 ;
      RECT  86100.0 453750.0 87300.0 451350.0 ;
      RECT  86100.0 462450.0 87300.0 466050.0 ;
      RECT  90900.0 462450.0 92100.0 466050.0 ;
      RECT  95700.0 463650.0 96900.0 465600.0 ;
      RECT  95700.0 451800.0 96900.0 453750.0 ;
      RECT  86100.0 462450.0 87300.0 463650.0 ;
      RECT  88500.0 462450.0 89700.0 463650.0 ;
      RECT  88500.0 462450.0 89700.0 463650.0 ;
      RECT  86100.0 462450.0 87300.0 463650.0 ;
      RECT  88500.0 462450.0 89700.0 463650.0 ;
      RECT  90900.0 462450.0 92100.0 463650.0 ;
      RECT  90900.0 462450.0 92100.0 463650.0 ;
      RECT  88500.0 462450.0 89700.0 463650.0 ;
      RECT  90900.0 462450.0 92100.0 463650.0 ;
      RECT  93300.0 462450.0 94500.0 463650.0 ;
      RECT  93300.0 462450.0 94500.0 463650.0 ;
      RECT  90900.0 462450.0 92100.0 463650.0 ;
      RECT  86100.0 453750.0 87300.0 454950.0 ;
      RECT  88500.0 453750.0 89700.0 454950.0 ;
      RECT  88500.0 453750.0 89700.0 454950.0 ;
      RECT  86100.0 453750.0 87300.0 454950.0 ;
      RECT  88500.0 453750.0 89700.0 454950.0 ;
      RECT  90900.0 453750.0 92100.0 454950.0 ;
      RECT  90900.0 453750.0 92100.0 454950.0 ;
      RECT  88500.0 453750.0 89700.0 454950.0 ;
      RECT  90900.0 453750.0 92100.0 454950.0 ;
      RECT  93300.0 453750.0 94500.0 454950.0 ;
      RECT  93300.0 453750.0 94500.0 454950.0 ;
      RECT  90900.0 453750.0 92100.0 454950.0 ;
      RECT  95700.0 463050.0 96900.0 464250.0 ;
      RECT  95700.0 453150.0 96900.0 454350.0 ;
      RECT  93300.0 455850.0 92100.0 457050.0 ;
      RECT  90900.0 457800.0 89700.0 459000.0 ;
      RECT  88500.0 459750.0 87300.0 460950.0 ;
      RECT  88500.0 462450.0 89700.0 463650.0 ;
      RECT  93300.0 462450.0 94500.0 463650.0 ;
      RECT  93300.0 453750.0 94500.0 454950.0 ;
      RECT  93300.0 459750.0 94500.0 460950.0 ;
      RECT  87300.0 459750.0 88500.0 460950.0 ;
      RECT  89700.0 457800.0 90900.0 459000.0 ;
      RECT  92100.0 455850.0 93300.0 457050.0 ;
      RECT  93300.0 459750.0 94500.0 460950.0 ;
      RECT  84300.0 465150.0 99900.0 466050.0 ;
      RECT  84300.0 451350.0 99900.0 452250.0 ;
      RECT  86100.0 477450.0 87300.0 479850.0 ;
      RECT  86100.0 468750.0 87300.0 465150.0 ;
      RECT  90900.0 468750.0 92100.0 465150.0 ;
      RECT  95700.0 467550.0 96900.0 465600.0 ;
      RECT  95700.0 479400.0 96900.0 477450.0 ;
      RECT  86100.0 468750.0 87300.0 467550.0 ;
      RECT  88500.0 468750.0 89700.0 467550.0 ;
      RECT  88500.0 468750.0 89700.0 467550.0 ;
      RECT  86100.0 468750.0 87300.0 467550.0 ;
      RECT  88500.0 468750.0 89700.0 467550.0 ;
      RECT  90900.0 468750.0 92100.0 467550.0 ;
      RECT  90900.0 468750.0 92100.0 467550.0 ;
      RECT  88500.0 468750.0 89700.0 467550.0 ;
      RECT  90900.0 468750.0 92100.0 467550.0 ;
      RECT  93300.0 468750.0 94500.0 467550.0 ;
      RECT  93300.0 468750.0 94500.0 467550.0 ;
      RECT  90900.0 468750.0 92100.0 467550.0 ;
      RECT  86100.0 477450.0 87300.0 476250.0 ;
      RECT  88500.0 477450.0 89700.0 476250.0 ;
      RECT  88500.0 477450.0 89700.0 476250.0 ;
      RECT  86100.0 477450.0 87300.0 476250.0 ;
      RECT  88500.0 477450.0 89700.0 476250.0 ;
      RECT  90900.0 477450.0 92100.0 476250.0 ;
      RECT  90900.0 477450.0 92100.0 476250.0 ;
      RECT  88500.0 477450.0 89700.0 476250.0 ;
      RECT  90900.0 477450.0 92100.0 476250.0 ;
      RECT  93300.0 477450.0 94500.0 476250.0 ;
      RECT  93300.0 477450.0 94500.0 476250.0 ;
      RECT  90900.0 477450.0 92100.0 476250.0 ;
      RECT  95700.0 468150.0 96900.0 466950.0 ;
      RECT  95700.0 478050.0 96900.0 476850.0 ;
      RECT  93300.0 475350.0 92100.0 474150.0 ;
      RECT  90900.0 473400.0 89700.0 472200.0 ;
      RECT  88500.0 471450.0 87300.0 470250.0 ;
      RECT  88500.0 468750.0 89700.0 467550.0 ;
      RECT  93300.0 468750.0 94500.0 467550.0 ;
      RECT  93300.0 477450.0 94500.0 476250.0 ;
      RECT  93300.0 471450.0 94500.0 470250.0 ;
      RECT  87300.0 471450.0 88500.0 470250.0 ;
      RECT  89700.0 473400.0 90900.0 472200.0 ;
      RECT  92100.0 475350.0 93300.0 474150.0 ;
      RECT  93300.0 471450.0 94500.0 470250.0 ;
      RECT  84300.0 466050.0 99900.0 465150.0 ;
      RECT  84300.0 479850.0 99900.0 478950.0 ;
      RECT  86100.0 481350.0 87300.0 478950.0 ;
      RECT  86100.0 490050.0 87300.0 493650.0 ;
      RECT  90900.0 490050.0 92100.0 493650.0 ;
      RECT  95700.0 491250.0 96900.0 493200.0 ;
      RECT  95700.0 479400.0 96900.0 481350.0 ;
      RECT  86100.0 490050.0 87300.0 491250.0 ;
      RECT  88500.0 490050.0 89700.0 491250.0 ;
      RECT  88500.0 490050.0 89700.0 491250.0 ;
      RECT  86100.0 490050.0 87300.0 491250.0 ;
      RECT  88500.0 490050.0 89700.0 491250.0 ;
      RECT  90900.0 490050.0 92100.0 491250.0 ;
      RECT  90900.0 490050.0 92100.0 491250.0 ;
      RECT  88500.0 490050.0 89700.0 491250.0 ;
      RECT  90900.0 490050.0 92100.0 491250.0 ;
      RECT  93300.0 490050.0 94500.0 491250.0 ;
      RECT  93300.0 490050.0 94500.0 491250.0 ;
      RECT  90900.0 490050.0 92100.0 491250.0 ;
      RECT  86100.0 481350.0 87300.0 482550.0 ;
      RECT  88500.0 481350.0 89700.0 482550.0 ;
      RECT  88500.0 481350.0 89700.0 482550.0 ;
      RECT  86100.0 481350.0 87300.0 482550.0 ;
      RECT  88500.0 481350.0 89700.0 482550.0 ;
      RECT  90900.0 481350.0 92100.0 482550.0 ;
      RECT  90900.0 481350.0 92100.0 482550.0 ;
      RECT  88500.0 481350.0 89700.0 482550.0 ;
      RECT  90900.0 481350.0 92100.0 482550.0 ;
      RECT  93300.0 481350.0 94500.0 482550.0 ;
      RECT  93300.0 481350.0 94500.0 482550.0 ;
      RECT  90900.0 481350.0 92100.0 482550.0 ;
      RECT  95700.0 490650.0 96900.0 491850.0 ;
      RECT  95700.0 480750.0 96900.0 481950.0 ;
      RECT  93300.0 483450.0 92100.0 484650.0 ;
      RECT  90900.0 485400.0 89700.0 486600.0 ;
      RECT  88500.0 487350.0 87300.0 488550.0 ;
      RECT  88500.0 490050.0 89700.0 491250.0 ;
      RECT  93300.0 490050.0 94500.0 491250.0 ;
      RECT  93300.0 481350.0 94500.0 482550.0 ;
      RECT  93300.0 487350.0 94500.0 488550.0 ;
      RECT  87300.0 487350.0 88500.0 488550.0 ;
      RECT  89700.0 485400.0 90900.0 486600.0 ;
      RECT  92100.0 483450.0 93300.0 484650.0 ;
      RECT  93300.0 487350.0 94500.0 488550.0 ;
      RECT  84300.0 492750.0 99900.0 493650.0 ;
      RECT  84300.0 478950.0 99900.0 479850.0 ;
      RECT  86100.0 505050.0 87300.0 507450.0 ;
      RECT  86100.0 496350.0 87300.0 492750.0 ;
      RECT  90900.0 496350.0 92100.0 492750.0 ;
      RECT  95700.0 495150.0 96900.0 493200.0 ;
      RECT  95700.0 507000.0 96900.0 505050.0 ;
      RECT  86100.0 496350.0 87300.0 495150.0 ;
      RECT  88500.0 496350.0 89700.0 495150.0 ;
      RECT  88500.0 496350.0 89700.0 495150.0 ;
      RECT  86100.0 496350.0 87300.0 495150.0 ;
      RECT  88500.0 496350.0 89700.0 495150.0 ;
      RECT  90900.0 496350.0 92100.0 495150.0 ;
      RECT  90900.0 496350.0 92100.0 495150.0 ;
      RECT  88500.0 496350.0 89700.0 495150.0 ;
      RECT  90900.0 496350.0 92100.0 495150.0 ;
      RECT  93300.0 496350.0 94500.0 495150.0 ;
      RECT  93300.0 496350.0 94500.0 495150.0 ;
      RECT  90900.0 496350.0 92100.0 495150.0 ;
      RECT  86100.0 505050.0 87300.0 503850.0 ;
      RECT  88500.0 505050.0 89700.0 503850.0 ;
      RECT  88500.0 505050.0 89700.0 503850.0 ;
      RECT  86100.0 505050.0 87300.0 503850.0 ;
      RECT  88500.0 505050.0 89700.0 503850.0 ;
      RECT  90900.0 505050.0 92100.0 503850.0 ;
      RECT  90900.0 505050.0 92100.0 503850.0 ;
      RECT  88500.0 505050.0 89700.0 503850.0 ;
      RECT  90900.0 505050.0 92100.0 503850.0 ;
      RECT  93300.0 505050.0 94500.0 503850.0 ;
      RECT  93300.0 505050.0 94500.0 503850.0 ;
      RECT  90900.0 505050.0 92100.0 503850.0 ;
      RECT  95700.0 495750.0 96900.0 494550.0 ;
      RECT  95700.0 505650.0 96900.0 504450.0 ;
      RECT  93300.0 502950.0 92100.0 501750.0 ;
      RECT  90900.0 501000.0 89700.0 499800.0 ;
      RECT  88500.0 499050.0 87300.0 497850.0 ;
      RECT  88500.0 496350.0 89700.0 495150.0 ;
      RECT  93300.0 496350.0 94500.0 495150.0 ;
      RECT  93300.0 505050.0 94500.0 503850.0 ;
      RECT  93300.0 499050.0 94500.0 497850.0 ;
      RECT  87300.0 499050.0 88500.0 497850.0 ;
      RECT  89700.0 501000.0 90900.0 499800.0 ;
      RECT  92100.0 502950.0 93300.0 501750.0 ;
      RECT  93300.0 499050.0 94500.0 497850.0 ;
      RECT  84300.0 493650.0 99900.0 492750.0 ;
      RECT  84300.0 507450.0 99900.0 506550.0 ;
      RECT  86100.0 508950.0 87300.0 506550.0 ;
      RECT  86100.0 517650.0 87300.0 521250.0 ;
      RECT  90900.0 517650.0 92100.0 521250.0 ;
      RECT  95700.0 518850.0 96900.0 520800.0 ;
      RECT  95700.0 507000.0 96900.0 508950.0 ;
      RECT  86100.0 517650.0 87300.0 518850.0 ;
      RECT  88500.0 517650.0 89700.0 518850.0 ;
      RECT  88500.0 517650.0 89700.0 518850.0 ;
      RECT  86100.0 517650.0 87300.0 518850.0 ;
      RECT  88500.0 517650.0 89700.0 518850.0 ;
      RECT  90900.0 517650.0 92100.0 518850.0 ;
      RECT  90900.0 517650.0 92100.0 518850.0 ;
      RECT  88500.0 517650.0 89700.0 518850.0 ;
      RECT  90900.0 517650.0 92100.0 518850.0 ;
      RECT  93300.0 517650.0 94500.0 518850.0 ;
      RECT  93300.0 517650.0 94500.0 518850.0 ;
      RECT  90900.0 517650.0 92100.0 518850.0 ;
      RECT  86100.0 508950.0 87300.0 510150.0 ;
      RECT  88500.0 508950.0 89700.0 510150.0 ;
      RECT  88500.0 508950.0 89700.0 510150.0 ;
      RECT  86100.0 508950.0 87300.0 510150.0 ;
      RECT  88500.0 508950.0 89700.0 510150.0 ;
      RECT  90900.0 508950.0 92100.0 510150.0 ;
      RECT  90900.0 508950.0 92100.0 510150.0 ;
      RECT  88500.0 508950.0 89700.0 510150.0 ;
      RECT  90900.0 508950.0 92100.0 510150.0 ;
      RECT  93300.0 508950.0 94500.0 510150.0 ;
      RECT  93300.0 508950.0 94500.0 510150.0 ;
      RECT  90900.0 508950.0 92100.0 510150.0 ;
      RECT  95700.0 518250.0 96900.0 519450.0 ;
      RECT  95700.0 508350.0 96900.0 509550.0 ;
      RECT  93300.0 511050.0 92100.0 512250.0 ;
      RECT  90900.0 513000.0 89700.0 514200.0 ;
      RECT  88500.0 514950.0 87300.0 516150.0 ;
      RECT  88500.0 517650.0 89700.0 518850.0 ;
      RECT  93300.0 517650.0 94500.0 518850.0 ;
      RECT  93300.0 508950.0 94500.0 510150.0 ;
      RECT  93300.0 514950.0 94500.0 516150.0 ;
      RECT  87300.0 514950.0 88500.0 516150.0 ;
      RECT  89700.0 513000.0 90900.0 514200.0 ;
      RECT  92100.0 511050.0 93300.0 512250.0 ;
      RECT  93300.0 514950.0 94500.0 516150.0 ;
      RECT  84300.0 520350.0 99900.0 521250.0 ;
      RECT  84300.0 506550.0 99900.0 507450.0 ;
      RECT  86100.0 532650.0 87300.0 535050.0 ;
      RECT  86100.0 523950.0 87300.0 520350.0 ;
      RECT  90900.0 523950.0 92100.0 520350.0 ;
      RECT  95700.0 522750.0 96900.0 520800.0 ;
      RECT  95700.0 534600.0 96900.0 532650.0 ;
      RECT  86100.0 523950.0 87300.0 522750.0 ;
      RECT  88500.0 523950.0 89700.0 522750.0 ;
      RECT  88500.0 523950.0 89700.0 522750.0 ;
      RECT  86100.0 523950.0 87300.0 522750.0 ;
      RECT  88500.0 523950.0 89700.0 522750.0 ;
      RECT  90900.0 523950.0 92100.0 522750.0 ;
      RECT  90900.0 523950.0 92100.0 522750.0 ;
      RECT  88500.0 523950.0 89700.0 522750.0 ;
      RECT  90900.0 523950.0 92100.0 522750.0 ;
      RECT  93300.0 523950.0 94500.0 522750.0 ;
      RECT  93300.0 523950.0 94500.0 522750.0 ;
      RECT  90900.0 523950.0 92100.0 522750.0 ;
      RECT  86100.0 532650.0 87300.0 531450.0 ;
      RECT  88500.0 532650.0 89700.0 531450.0 ;
      RECT  88500.0 532650.0 89700.0 531450.0 ;
      RECT  86100.0 532650.0 87300.0 531450.0 ;
      RECT  88500.0 532650.0 89700.0 531450.0 ;
      RECT  90900.0 532650.0 92100.0 531450.0 ;
      RECT  90900.0 532650.0 92100.0 531450.0 ;
      RECT  88500.0 532650.0 89700.0 531450.0 ;
      RECT  90900.0 532650.0 92100.0 531450.0 ;
      RECT  93300.0 532650.0 94500.0 531450.0 ;
      RECT  93300.0 532650.0 94500.0 531450.0 ;
      RECT  90900.0 532650.0 92100.0 531450.0 ;
      RECT  95700.0 523350.0 96900.0 522150.0 ;
      RECT  95700.0 533250.0 96900.0 532050.0 ;
      RECT  93300.0 530550.0 92100.0 529350.0 ;
      RECT  90900.0 528600.0 89700.0 527400.0 ;
      RECT  88500.0 526650.0 87300.0 525450.0 ;
      RECT  88500.0 523950.0 89700.0 522750.0 ;
      RECT  93300.0 523950.0 94500.0 522750.0 ;
      RECT  93300.0 532650.0 94500.0 531450.0 ;
      RECT  93300.0 526650.0 94500.0 525450.0 ;
      RECT  87300.0 526650.0 88500.0 525450.0 ;
      RECT  89700.0 528600.0 90900.0 527400.0 ;
      RECT  92100.0 530550.0 93300.0 529350.0 ;
      RECT  93300.0 526650.0 94500.0 525450.0 ;
      RECT  84300.0 521250.0 99900.0 520350.0 ;
      RECT  84300.0 535050.0 99900.0 534150.0 ;
      RECT  86100.0 536550.0 87300.0 534150.0 ;
      RECT  86100.0 545250.0 87300.0 548850.0 ;
      RECT  90900.0 545250.0 92100.0 548850.0 ;
      RECT  95700.0 546450.0 96900.0 548400.0 ;
      RECT  95700.0 534600.0 96900.0 536550.0 ;
      RECT  86100.0 545250.0 87300.0 546450.0 ;
      RECT  88500.0 545250.0 89700.0 546450.0 ;
      RECT  88500.0 545250.0 89700.0 546450.0 ;
      RECT  86100.0 545250.0 87300.0 546450.0 ;
      RECT  88500.0 545250.0 89700.0 546450.0 ;
      RECT  90900.0 545250.0 92100.0 546450.0 ;
      RECT  90900.0 545250.0 92100.0 546450.0 ;
      RECT  88500.0 545250.0 89700.0 546450.0 ;
      RECT  90900.0 545250.0 92100.0 546450.0 ;
      RECT  93300.0 545250.0 94500.0 546450.0 ;
      RECT  93300.0 545250.0 94500.0 546450.0 ;
      RECT  90900.0 545250.0 92100.0 546450.0 ;
      RECT  86100.0 536550.0 87300.0 537750.0 ;
      RECT  88500.0 536550.0 89700.0 537750.0 ;
      RECT  88500.0 536550.0 89700.0 537750.0 ;
      RECT  86100.0 536550.0 87300.0 537750.0 ;
      RECT  88500.0 536550.0 89700.0 537750.0 ;
      RECT  90900.0 536550.0 92100.0 537750.0 ;
      RECT  90900.0 536550.0 92100.0 537750.0 ;
      RECT  88500.0 536550.0 89700.0 537750.0 ;
      RECT  90900.0 536550.0 92100.0 537750.0 ;
      RECT  93300.0 536550.0 94500.0 537750.0 ;
      RECT  93300.0 536550.0 94500.0 537750.0 ;
      RECT  90900.0 536550.0 92100.0 537750.0 ;
      RECT  95700.0 545850.0 96900.0 547050.0 ;
      RECT  95700.0 535950.0 96900.0 537150.0 ;
      RECT  93300.0 538650.0 92100.0 539850.0 ;
      RECT  90900.0 540600.0 89700.0 541800.0 ;
      RECT  88500.0 542550.0 87300.0 543750.0 ;
      RECT  88500.0 545250.0 89700.0 546450.0 ;
      RECT  93300.0 545250.0 94500.0 546450.0 ;
      RECT  93300.0 536550.0 94500.0 537750.0 ;
      RECT  93300.0 542550.0 94500.0 543750.0 ;
      RECT  87300.0 542550.0 88500.0 543750.0 ;
      RECT  89700.0 540600.0 90900.0 541800.0 ;
      RECT  92100.0 538650.0 93300.0 539850.0 ;
      RECT  93300.0 542550.0 94500.0 543750.0 ;
      RECT  84300.0 547950.0 99900.0 548850.0 ;
      RECT  84300.0 534150.0 99900.0 535050.0 ;
      RECT  86100.0 560250.0 87300.0 562650.0 ;
      RECT  86100.0 551550.0 87300.0 547950.0 ;
      RECT  90900.0 551550.0 92100.0 547950.0 ;
      RECT  95700.0 550350.0 96900.0 548400.0 ;
      RECT  95700.0 562200.0 96900.0 560250.0 ;
      RECT  86100.0 551550.0 87300.0 550350.0 ;
      RECT  88500.0 551550.0 89700.0 550350.0 ;
      RECT  88500.0 551550.0 89700.0 550350.0 ;
      RECT  86100.0 551550.0 87300.0 550350.0 ;
      RECT  88500.0 551550.0 89700.0 550350.0 ;
      RECT  90900.0 551550.0 92100.0 550350.0 ;
      RECT  90900.0 551550.0 92100.0 550350.0 ;
      RECT  88500.0 551550.0 89700.0 550350.0 ;
      RECT  90900.0 551550.0 92100.0 550350.0 ;
      RECT  93300.0 551550.0 94500.0 550350.0 ;
      RECT  93300.0 551550.0 94500.0 550350.0 ;
      RECT  90900.0 551550.0 92100.0 550350.0 ;
      RECT  86100.0 560250.0 87300.0 559050.0 ;
      RECT  88500.0 560250.0 89700.0 559050.0 ;
      RECT  88500.0 560250.0 89700.0 559050.0 ;
      RECT  86100.0 560250.0 87300.0 559050.0 ;
      RECT  88500.0 560250.0 89700.0 559050.0 ;
      RECT  90900.0 560250.0 92100.0 559050.0 ;
      RECT  90900.0 560250.0 92100.0 559050.0 ;
      RECT  88500.0 560250.0 89700.0 559050.0 ;
      RECT  90900.0 560250.0 92100.0 559050.0 ;
      RECT  93300.0 560250.0 94500.0 559050.0 ;
      RECT  93300.0 560250.0 94500.0 559050.0 ;
      RECT  90900.0 560250.0 92100.0 559050.0 ;
      RECT  95700.0 550950.0 96900.0 549750.0 ;
      RECT  95700.0 560850.0 96900.0 559650.0 ;
      RECT  93300.0 558150.0 92100.0 556950.0 ;
      RECT  90900.0 556200.0 89700.0 555000.0 ;
      RECT  88500.0 554250.0 87300.0 553050.0 ;
      RECT  88500.0 551550.0 89700.0 550350.0 ;
      RECT  93300.0 551550.0 94500.0 550350.0 ;
      RECT  93300.0 560250.0 94500.0 559050.0 ;
      RECT  93300.0 554250.0 94500.0 553050.0 ;
      RECT  87300.0 554250.0 88500.0 553050.0 ;
      RECT  89700.0 556200.0 90900.0 555000.0 ;
      RECT  92100.0 558150.0 93300.0 556950.0 ;
      RECT  93300.0 554250.0 94500.0 553050.0 ;
      RECT  84300.0 548850.0 99900.0 547950.0 ;
      RECT  84300.0 562650.0 99900.0 561750.0 ;
      RECT  86100.0 564150.0 87300.0 561750.0 ;
      RECT  86100.0 572850.0 87300.0 576450.0 ;
      RECT  90900.0 572850.0 92100.0 576450.0 ;
      RECT  95700.0 574050.0 96900.0 576000.0 ;
      RECT  95700.0 562200.0 96900.0 564150.0 ;
      RECT  86100.0 572850.0 87300.0 574050.0 ;
      RECT  88500.0 572850.0 89700.0 574050.0 ;
      RECT  88500.0 572850.0 89700.0 574050.0 ;
      RECT  86100.0 572850.0 87300.0 574050.0 ;
      RECT  88500.0 572850.0 89700.0 574050.0 ;
      RECT  90900.0 572850.0 92100.0 574050.0 ;
      RECT  90900.0 572850.0 92100.0 574050.0 ;
      RECT  88500.0 572850.0 89700.0 574050.0 ;
      RECT  90900.0 572850.0 92100.0 574050.0 ;
      RECT  93300.0 572850.0 94500.0 574050.0 ;
      RECT  93300.0 572850.0 94500.0 574050.0 ;
      RECT  90900.0 572850.0 92100.0 574050.0 ;
      RECT  86100.0 564150.0 87300.0 565350.0 ;
      RECT  88500.0 564150.0 89700.0 565350.0 ;
      RECT  88500.0 564150.0 89700.0 565350.0 ;
      RECT  86100.0 564150.0 87300.0 565350.0 ;
      RECT  88500.0 564150.0 89700.0 565350.0 ;
      RECT  90900.0 564150.0 92100.0 565350.0 ;
      RECT  90900.0 564150.0 92100.0 565350.0 ;
      RECT  88500.0 564150.0 89700.0 565350.0 ;
      RECT  90900.0 564150.0 92100.0 565350.0 ;
      RECT  93300.0 564150.0 94500.0 565350.0 ;
      RECT  93300.0 564150.0 94500.0 565350.0 ;
      RECT  90900.0 564150.0 92100.0 565350.0 ;
      RECT  95700.0 573450.0 96900.0 574650.0 ;
      RECT  95700.0 563550.0 96900.0 564750.0 ;
      RECT  93300.0 566250.0 92100.0 567450.0 ;
      RECT  90900.0 568200.0 89700.0 569400.0 ;
      RECT  88500.0 570150.0 87300.0 571350.0 ;
      RECT  88500.0 572850.0 89700.0 574050.0 ;
      RECT  93300.0 572850.0 94500.0 574050.0 ;
      RECT  93300.0 564150.0 94500.0 565350.0 ;
      RECT  93300.0 570150.0 94500.0 571350.0 ;
      RECT  87300.0 570150.0 88500.0 571350.0 ;
      RECT  89700.0 568200.0 90900.0 569400.0 ;
      RECT  92100.0 566250.0 93300.0 567450.0 ;
      RECT  93300.0 570150.0 94500.0 571350.0 ;
      RECT  84300.0 575550.0 99900.0 576450.0 ;
      RECT  84300.0 561750.0 99900.0 562650.0 ;
      RECT  86100.0 587850.0 87300.0 590250.0 ;
      RECT  86100.0 579150.0 87300.0 575550.0 ;
      RECT  90900.0 579150.0 92100.0 575550.0 ;
      RECT  95700.0 577950.0 96900.0 576000.0 ;
      RECT  95700.0 589800.0 96900.0 587850.0 ;
      RECT  86100.0 579150.0 87300.0 577950.0 ;
      RECT  88500.0 579150.0 89700.0 577950.0 ;
      RECT  88500.0 579150.0 89700.0 577950.0 ;
      RECT  86100.0 579150.0 87300.0 577950.0 ;
      RECT  88500.0 579150.0 89700.0 577950.0 ;
      RECT  90900.0 579150.0 92100.0 577950.0 ;
      RECT  90900.0 579150.0 92100.0 577950.0 ;
      RECT  88500.0 579150.0 89700.0 577950.0 ;
      RECT  90900.0 579150.0 92100.0 577950.0 ;
      RECT  93300.0 579150.0 94500.0 577950.0 ;
      RECT  93300.0 579150.0 94500.0 577950.0 ;
      RECT  90900.0 579150.0 92100.0 577950.0 ;
      RECT  86100.0 587850.0 87300.0 586650.0 ;
      RECT  88500.0 587850.0 89700.0 586650.0 ;
      RECT  88500.0 587850.0 89700.0 586650.0 ;
      RECT  86100.0 587850.0 87300.0 586650.0 ;
      RECT  88500.0 587850.0 89700.0 586650.0 ;
      RECT  90900.0 587850.0 92100.0 586650.0 ;
      RECT  90900.0 587850.0 92100.0 586650.0 ;
      RECT  88500.0 587850.0 89700.0 586650.0 ;
      RECT  90900.0 587850.0 92100.0 586650.0 ;
      RECT  93300.0 587850.0 94500.0 586650.0 ;
      RECT  93300.0 587850.0 94500.0 586650.0 ;
      RECT  90900.0 587850.0 92100.0 586650.0 ;
      RECT  95700.0 578550.0 96900.0 577350.0 ;
      RECT  95700.0 588450.0 96900.0 587250.0 ;
      RECT  93300.0 585750.0 92100.0 584550.0 ;
      RECT  90900.0 583800.0 89700.0 582600.0 ;
      RECT  88500.0 581850.0 87300.0 580650.0 ;
      RECT  88500.0 579150.0 89700.0 577950.0 ;
      RECT  93300.0 579150.0 94500.0 577950.0 ;
      RECT  93300.0 587850.0 94500.0 586650.0 ;
      RECT  93300.0 581850.0 94500.0 580650.0 ;
      RECT  87300.0 581850.0 88500.0 580650.0 ;
      RECT  89700.0 583800.0 90900.0 582600.0 ;
      RECT  92100.0 585750.0 93300.0 584550.0 ;
      RECT  93300.0 581850.0 94500.0 580650.0 ;
      RECT  84300.0 576450.0 99900.0 575550.0 ;
      RECT  84300.0 590250.0 99900.0 589350.0 ;
      RECT  86100.0 591750.0 87300.0 589350.0 ;
      RECT  86100.0 600450.0 87300.0 604050.0 ;
      RECT  90900.0 600450.0 92100.0 604050.0 ;
      RECT  95700.0 601650.0 96900.0 603600.0 ;
      RECT  95700.0 589800.0 96900.0 591750.0 ;
      RECT  86100.0 600450.0 87300.0 601650.0 ;
      RECT  88500.0 600450.0 89700.0 601650.0 ;
      RECT  88500.0 600450.0 89700.0 601650.0 ;
      RECT  86100.0 600450.0 87300.0 601650.0 ;
      RECT  88500.0 600450.0 89700.0 601650.0 ;
      RECT  90900.0 600450.0 92100.0 601650.0 ;
      RECT  90900.0 600450.0 92100.0 601650.0 ;
      RECT  88500.0 600450.0 89700.0 601650.0 ;
      RECT  90900.0 600450.0 92100.0 601650.0 ;
      RECT  93300.0 600450.0 94500.0 601650.0 ;
      RECT  93300.0 600450.0 94500.0 601650.0 ;
      RECT  90900.0 600450.0 92100.0 601650.0 ;
      RECT  86100.0 591750.0 87300.0 592950.0 ;
      RECT  88500.0 591750.0 89700.0 592950.0 ;
      RECT  88500.0 591750.0 89700.0 592950.0 ;
      RECT  86100.0 591750.0 87300.0 592950.0 ;
      RECT  88500.0 591750.0 89700.0 592950.0 ;
      RECT  90900.0 591750.0 92100.0 592950.0 ;
      RECT  90900.0 591750.0 92100.0 592950.0 ;
      RECT  88500.0 591750.0 89700.0 592950.0 ;
      RECT  90900.0 591750.0 92100.0 592950.0 ;
      RECT  93300.0 591750.0 94500.0 592950.0 ;
      RECT  93300.0 591750.0 94500.0 592950.0 ;
      RECT  90900.0 591750.0 92100.0 592950.0 ;
      RECT  95700.0 601050.0 96900.0 602250.0 ;
      RECT  95700.0 591150.0 96900.0 592350.0 ;
      RECT  93300.0 593850.0 92100.0 595050.0 ;
      RECT  90900.0 595800.0 89700.0 597000.0 ;
      RECT  88500.0 597750.0 87300.0 598950.0 ;
      RECT  88500.0 600450.0 89700.0 601650.0 ;
      RECT  93300.0 600450.0 94500.0 601650.0 ;
      RECT  93300.0 591750.0 94500.0 592950.0 ;
      RECT  93300.0 597750.0 94500.0 598950.0 ;
      RECT  87300.0 597750.0 88500.0 598950.0 ;
      RECT  89700.0 595800.0 90900.0 597000.0 ;
      RECT  92100.0 593850.0 93300.0 595050.0 ;
      RECT  93300.0 597750.0 94500.0 598950.0 ;
      RECT  84300.0 603150.0 99900.0 604050.0 ;
      RECT  84300.0 589350.0 99900.0 590250.0 ;
      RECT  86100.0 615450.0 87300.0 617850.0 ;
      RECT  86100.0 606750.0 87300.0 603150.0 ;
      RECT  90900.0 606750.0 92100.0 603150.0 ;
      RECT  95700.0 605550.0 96900.0 603600.0 ;
      RECT  95700.0 617400.0 96900.0 615450.0 ;
      RECT  86100.0 606750.0 87300.0 605550.0 ;
      RECT  88500.0 606750.0 89700.0 605550.0 ;
      RECT  88500.0 606750.0 89700.0 605550.0 ;
      RECT  86100.0 606750.0 87300.0 605550.0 ;
      RECT  88500.0 606750.0 89700.0 605550.0 ;
      RECT  90900.0 606750.0 92100.0 605550.0 ;
      RECT  90900.0 606750.0 92100.0 605550.0 ;
      RECT  88500.0 606750.0 89700.0 605550.0 ;
      RECT  90900.0 606750.0 92100.0 605550.0 ;
      RECT  93300.0 606750.0 94500.0 605550.0 ;
      RECT  93300.0 606750.0 94500.0 605550.0 ;
      RECT  90900.0 606750.0 92100.0 605550.0 ;
      RECT  86100.0 615450.0 87300.0 614250.0 ;
      RECT  88500.0 615450.0 89700.0 614250.0 ;
      RECT  88500.0 615450.0 89700.0 614250.0 ;
      RECT  86100.0 615450.0 87300.0 614250.0 ;
      RECT  88500.0 615450.0 89700.0 614250.0 ;
      RECT  90900.0 615450.0 92100.0 614250.0 ;
      RECT  90900.0 615450.0 92100.0 614250.0 ;
      RECT  88500.0 615450.0 89700.0 614250.0 ;
      RECT  90900.0 615450.0 92100.0 614250.0 ;
      RECT  93300.0 615450.0 94500.0 614250.0 ;
      RECT  93300.0 615450.0 94500.0 614250.0 ;
      RECT  90900.0 615450.0 92100.0 614250.0 ;
      RECT  95700.0 606150.0 96900.0 604950.0 ;
      RECT  95700.0 616050.0 96900.0 614850.0 ;
      RECT  93300.0 613350.0 92100.0 612150.0 ;
      RECT  90900.0 611400.0 89700.0 610200.0 ;
      RECT  88500.0 609450.0 87300.0 608250.0 ;
      RECT  88500.0 606750.0 89700.0 605550.0 ;
      RECT  93300.0 606750.0 94500.0 605550.0 ;
      RECT  93300.0 615450.0 94500.0 614250.0 ;
      RECT  93300.0 609450.0 94500.0 608250.0 ;
      RECT  87300.0 609450.0 88500.0 608250.0 ;
      RECT  89700.0 611400.0 90900.0 610200.0 ;
      RECT  92100.0 613350.0 93300.0 612150.0 ;
      RECT  93300.0 609450.0 94500.0 608250.0 ;
      RECT  84300.0 604050.0 99900.0 603150.0 ;
      RECT  84300.0 617850.0 99900.0 616950.0 ;
      RECT  86100.0 619350.0 87300.0 616950.0 ;
      RECT  86100.0 628050.0 87300.0 631650.0 ;
      RECT  90900.0 628050.0 92100.0 631650.0 ;
      RECT  95700.0 629250.0 96900.0 631200.0 ;
      RECT  95700.0 617400.0 96900.0 619350.0 ;
      RECT  86100.0 628050.0 87300.0 629250.0 ;
      RECT  88500.0 628050.0 89700.0 629250.0 ;
      RECT  88500.0 628050.0 89700.0 629250.0 ;
      RECT  86100.0 628050.0 87300.0 629250.0 ;
      RECT  88500.0 628050.0 89700.0 629250.0 ;
      RECT  90900.0 628050.0 92100.0 629250.0 ;
      RECT  90900.0 628050.0 92100.0 629250.0 ;
      RECT  88500.0 628050.0 89700.0 629250.0 ;
      RECT  90900.0 628050.0 92100.0 629250.0 ;
      RECT  93300.0 628050.0 94500.0 629250.0 ;
      RECT  93300.0 628050.0 94500.0 629250.0 ;
      RECT  90900.0 628050.0 92100.0 629250.0 ;
      RECT  86100.0 619350.0 87300.0 620550.0 ;
      RECT  88500.0 619350.0 89700.0 620550.0 ;
      RECT  88500.0 619350.0 89700.0 620550.0 ;
      RECT  86100.0 619350.0 87300.0 620550.0 ;
      RECT  88500.0 619350.0 89700.0 620550.0 ;
      RECT  90900.0 619350.0 92100.0 620550.0 ;
      RECT  90900.0 619350.0 92100.0 620550.0 ;
      RECT  88500.0 619350.0 89700.0 620550.0 ;
      RECT  90900.0 619350.0 92100.0 620550.0 ;
      RECT  93300.0 619350.0 94500.0 620550.0 ;
      RECT  93300.0 619350.0 94500.0 620550.0 ;
      RECT  90900.0 619350.0 92100.0 620550.0 ;
      RECT  95700.0 628650.0 96900.0 629850.0 ;
      RECT  95700.0 618750.0 96900.0 619950.0 ;
      RECT  93300.0 621450.0 92100.0 622650.0 ;
      RECT  90900.0 623400.0 89700.0 624600.0 ;
      RECT  88500.0 625350.0 87300.0 626550.0 ;
      RECT  88500.0 628050.0 89700.0 629250.0 ;
      RECT  93300.0 628050.0 94500.0 629250.0 ;
      RECT  93300.0 619350.0 94500.0 620550.0 ;
      RECT  93300.0 625350.0 94500.0 626550.0 ;
      RECT  87300.0 625350.0 88500.0 626550.0 ;
      RECT  89700.0 623400.0 90900.0 624600.0 ;
      RECT  92100.0 621450.0 93300.0 622650.0 ;
      RECT  93300.0 625350.0 94500.0 626550.0 ;
      RECT  84300.0 630750.0 99900.0 631650.0 ;
      RECT  84300.0 616950.0 99900.0 617850.0 ;
      RECT  86100.0 643050.0 87300.0 645450.0 ;
      RECT  86100.0 634350.0 87300.0 630750.0 ;
      RECT  90900.0 634350.0 92100.0 630750.0 ;
      RECT  95700.0 633150.0 96900.0 631200.0 ;
      RECT  95700.0 645000.0 96900.0 643050.0 ;
      RECT  86100.0 634350.0 87300.0 633150.0 ;
      RECT  88500.0 634350.0 89700.0 633150.0 ;
      RECT  88500.0 634350.0 89700.0 633150.0 ;
      RECT  86100.0 634350.0 87300.0 633150.0 ;
      RECT  88500.0 634350.0 89700.0 633150.0 ;
      RECT  90900.0 634350.0 92100.0 633150.0 ;
      RECT  90900.0 634350.0 92100.0 633150.0 ;
      RECT  88500.0 634350.0 89700.0 633150.0 ;
      RECT  90900.0 634350.0 92100.0 633150.0 ;
      RECT  93300.0 634350.0 94500.0 633150.0 ;
      RECT  93300.0 634350.0 94500.0 633150.0 ;
      RECT  90900.0 634350.0 92100.0 633150.0 ;
      RECT  86100.0 643050.0 87300.0 641850.0 ;
      RECT  88500.0 643050.0 89700.0 641850.0 ;
      RECT  88500.0 643050.0 89700.0 641850.0 ;
      RECT  86100.0 643050.0 87300.0 641850.0 ;
      RECT  88500.0 643050.0 89700.0 641850.0 ;
      RECT  90900.0 643050.0 92100.0 641850.0 ;
      RECT  90900.0 643050.0 92100.0 641850.0 ;
      RECT  88500.0 643050.0 89700.0 641850.0 ;
      RECT  90900.0 643050.0 92100.0 641850.0 ;
      RECT  93300.0 643050.0 94500.0 641850.0 ;
      RECT  93300.0 643050.0 94500.0 641850.0 ;
      RECT  90900.0 643050.0 92100.0 641850.0 ;
      RECT  95700.0 633750.0 96900.0 632550.0 ;
      RECT  95700.0 643650.0 96900.0 642450.0 ;
      RECT  93300.0 640950.0 92100.0 639750.0 ;
      RECT  90900.0 639000.0 89700.0 637800.0 ;
      RECT  88500.0 637050.0 87300.0 635850.0 ;
      RECT  88500.0 634350.0 89700.0 633150.0 ;
      RECT  93300.0 634350.0 94500.0 633150.0 ;
      RECT  93300.0 643050.0 94500.0 641850.0 ;
      RECT  93300.0 637050.0 94500.0 635850.0 ;
      RECT  87300.0 637050.0 88500.0 635850.0 ;
      RECT  89700.0 639000.0 90900.0 637800.0 ;
      RECT  92100.0 640950.0 93300.0 639750.0 ;
      RECT  93300.0 637050.0 94500.0 635850.0 ;
      RECT  84300.0 631650.0 99900.0 630750.0 ;
      RECT  84300.0 645450.0 99900.0 644550.0 ;
      RECT  86100.0 646950.0 87300.0 644550.0 ;
      RECT  86100.0 655650.0 87300.0 659250.0 ;
      RECT  90900.0 655650.0 92100.0 659250.0 ;
      RECT  95700.0 656850.0 96900.0 658800.0 ;
      RECT  95700.0 645000.0 96900.0 646950.0 ;
      RECT  86100.0 655650.0 87300.0 656850.0 ;
      RECT  88500.0 655650.0 89700.0 656850.0 ;
      RECT  88500.0 655650.0 89700.0 656850.0 ;
      RECT  86100.0 655650.0 87300.0 656850.0 ;
      RECT  88500.0 655650.0 89700.0 656850.0 ;
      RECT  90900.0 655650.0 92100.0 656850.0 ;
      RECT  90900.0 655650.0 92100.0 656850.0 ;
      RECT  88500.0 655650.0 89700.0 656850.0 ;
      RECT  90900.0 655650.0 92100.0 656850.0 ;
      RECT  93300.0 655650.0 94500.0 656850.0 ;
      RECT  93300.0 655650.0 94500.0 656850.0 ;
      RECT  90900.0 655650.0 92100.0 656850.0 ;
      RECT  86100.0 646950.0 87300.0 648150.0 ;
      RECT  88500.0 646950.0 89700.0 648150.0 ;
      RECT  88500.0 646950.0 89700.0 648150.0 ;
      RECT  86100.0 646950.0 87300.0 648150.0 ;
      RECT  88500.0 646950.0 89700.0 648150.0 ;
      RECT  90900.0 646950.0 92100.0 648150.0 ;
      RECT  90900.0 646950.0 92100.0 648150.0 ;
      RECT  88500.0 646950.0 89700.0 648150.0 ;
      RECT  90900.0 646950.0 92100.0 648150.0 ;
      RECT  93300.0 646950.0 94500.0 648150.0 ;
      RECT  93300.0 646950.0 94500.0 648150.0 ;
      RECT  90900.0 646950.0 92100.0 648150.0 ;
      RECT  95700.0 656250.0 96900.0 657450.0 ;
      RECT  95700.0 646350.0 96900.0 647550.0 ;
      RECT  93300.0 649050.0 92100.0 650250.0 ;
      RECT  90900.0 651000.0 89700.0 652200.0 ;
      RECT  88500.0 652950.0 87300.0 654150.0 ;
      RECT  88500.0 655650.0 89700.0 656850.0 ;
      RECT  93300.0 655650.0 94500.0 656850.0 ;
      RECT  93300.0 646950.0 94500.0 648150.0 ;
      RECT  93300.0 652950.0 94500.0 654150.0 ;
      RECT  87300.0 652950.0 88500.0 654150.0 ;
      RECT  89700.0 651000.0 90900.0 652200.0 ;
      RECT  92100.0 649050.0 93300.0 650250.0 ;
      RECT  93300.0 652950.0 94500.0 654150.0 ;
      RECT  84300.0 658350.0 99900.0 659250.0 ;
      RECT  84300.0 644550.0 99900.0 645450.0 ;
      RECT  86100.0 670650.0 87300.0 673050.0 ;
      RECT  86100.0 661950.0 87300.0 658350.0 ;
      RECT  90900.0 661950.0 92100.0 658350.0 ;
      RECT  95700.0 660750.0 96900.0 658800.0 ;
      RECT  95700.0 672600.0 96900.0 670650.0 ;
      RECT  86100.0 661950.0 87300.0 660750.0 ;
      RECT  88500.0 661950.0 89700.0 660750.0 ;
      RECT  88500.0 661950.0 89700.0 660750.0 ;
      RECT  86100.0 661950.0 87300.0 660750.0 ;
      RECT  88500.0 661950.0 89700.0 660750.0 ;
      RECT  90900.0 661950.0 92100.0 660750.0 ;
      RECT  90900.0 661950.0 92100.0 660750.0 ;
      RECT  88500.0 661950.0 89700.0 660750.0 ;
      RECT  90900.0 661950.0 92100.0 660750.0 ;
      RECT  93300.0 661950.0 94500.0 660750.0 ;
      RECT  93300.0 661950.0 94500.0 660750.0 ;
      RECT  90900.0 661950.0 92100.0 660750.0 ;
      RECT  86100.0 670650.0 87300.0 669450.0 ;
      RECT  88500.0 670650.0 89700.0 669450.0 ;
      RECT  88500.0 670650.0 89700.0 669450.0 ;
      RECT  86100.0 670650.0 87300.0 669450.0 ;
      RECT  88500.0 670650.0 89700.0 669450.0 ;
      RECT  90900.0 670650.0 92100.0 669450.0 ;
      RECT  90900.0 670650.0 92100.0 669450.0 ;
      RECT  88500.0 670650.0 89700.0 669450.0 ;
      RECT  90900.0 670650.0 92100.0 669450.0 ;
      RECT  93300.0 670650.0 94500.0 669450.0 ;
      RECT  93300.0 670650.0 94500.0 669450.0 ;
      RECT  90900.0 670650.0 92100.0 669450.0 ;
      RECT  95700.0 661350.0 96900.0 660150.0 ;
      RECT  95700.0 671250.0 96900.0 670050.0 ;
      RECT  93300.0 668550.0 92100.0 667350.0 ;
      RECT  90900.0 666600.0 89700.0 665400.0 ;
      RECT  88500.0 664650.0 87300.0 663450.0 ;
      RECT  88500.0 661950.0 89700.0 660750.0 ;
      RECT  93300.0 661950.0 94500.0 660750.0 ;
      RECT  93300.0 670650.0 94500.0 669450.0 ;
      RECT  93300.0 664650.0 94500.0 663450.0 ;
      RECT  87300.0 664650.0 88500.0 663450.0 ;
      RECT  89700.0 666600.0 90900.0 665400.0 ;
      RECT  92100.0 668550.0 93300.0 667350.0 ;
      RECT  93300.0 664650.0 94500.0 663450.0 ;
      RECT  84300.0 659250.0 99900.0 658350.0 ;
      RECT  84300.0 673050.0 99900.0 672150.0 ;
      RECT  86100.0 674550.0 87300.0 672150.0 ;
      RECT  86100.0 683250.0 87300.0 686850.0 ;
      RECT  90900.0 683250.0 92100.0 686850.0 ;
      RECT  95700.0 684450.0 96900.0 686400.0 ;
      RECT  95700.0 672600.0 96900.0 674550.0 ;
      RECT  86100.0 683250.0 87300.0 684450.0 ;
      RECT  88500.0 683250.0 89700.0 684450.0 ;
      RECT  88500.0 683250.0 89700.0 684450.0 ;
      RECT  86100.0 683250.0 87300.0 684450.0 ;
      RECT  88500.0 683250.0 89700.0 684450.0 ;
      RECT  90900.0 683250.0 92100.0 684450.0 ;
      RECT  90900.0 683250.0 92100.0 684450.0 ;
      RECT  88500.0 683250.0 89700.0 684450.0 ;
      RECT  90900.0 683250.0 92100.0 684450.0 ;
      RECT  93300.0 683250.0 94500.0 684450.0 ;
      RECT  93300.0 683250.0 94500.0 684450.0 ;
      RECT  90900.0 683250.0 92100.0 684450.0 ;
      RECT  86100.0 674550.0 87300.0 675750.0 ;
      RECT  88500.0 674550.0 89700.0 675750.0 ;
      RECT  88500.0 674550.0 89700.0 675750.0 ;
      RECT  86100.0 674550.0 87300.0 675750.0 ;
      RECT  88500.0 674550.0 89700.0 675750.0 ;
      RECT  90900.0 674550.0 92100.0 675750.0 ;
      RECT  90900.0 674550.0 92100.0 675750.0 ;
      RECT  88500.0 674550.0 89700.0 675750.0 ;
      RECT  90900.0 674550.0 92100.0 675750.0 ;
      RECT  93300.0 674550.0 94500.0 675750.0 ;
      RECT  93300.0 674550.0 94500.0 675750.0 ;
      RECT  90900.0 674550.0 92100.0 675750.0 ;
      RECT  95700.0 683850.0 96900.0 685050.0 ;
      RECT  95700.0 673950.0 96900.0 675150.0 ;
      RECT  93300.0 676650.0 92100.0 677850.0 ;
      RECT  90900.0 678600.0 89700.0 679800.0 ;
      RECT  88500.0 680550.0 87300.0 681750.0 ;
      RECT  88500.0 683250.0 89700.0 684450.0 ;
      RECT  93300.0 683250.0 94500.0 684450.0 ;
      RECT  93300.0 674550.0 94500.0 675750.0 ;
      RECT  93300.0 680550.0 94500.0 681750.0 ;
      RECT  87300.0 680550.0 88500.0 681750.0 ;
      RECT  89700.0 678600.0 90900.0 679800.0 ;
      RECT  92100.0 676650.0 93300.0 677850.0 ;
      RECT  93300.0 680550.0 94500.0 681750.0 ;
      RECT  84300.0 685950.0 99900.0 686850.0 ;
      RECT  84300.0 672150.0 99900.0 673050.0 ;
      RECT  86100.0 698250.0 87300.0 700650.0 ;
      RECT  86100.0 689550.0 87300.0 685950.0 ;
      RECT  90900.0 689550.0 92100.0 685950.0 ;
      RECT  95700.0 688350.0 96900.0 686400.0 ;
      RECT  95700.0 700200.0 96900.0 698250.0 ;
      RECT  86100.0 689550.0 87300.0 688350.0 ;
      RECT  88500.0 689550.0 89700.0 688350.0 ;
      RECT  88500.0 689550.0 89700.0 688350.0 ;
      RECT  86100.0 689550.0 87300.0 688350.0 ;
      RECT  88500.0 689550.0 89700.0 688350.0 ;
      RECT  90900.0 689550.0 92100.0 688350.0 ;
      RECT  90900.0 689550.0 92100.0 688350.0 ;
      RECT  88500.0 689550.0 89700.0 688350.0 ;
      RECT  90900.0 689550.0 92100.0 688350.0 ;
      RECT  93300.0 689550.0 94500.0 688350.0 ;
      RECT  93300.0 689550.0 94500.0 688350.0 ;
      RECT  90900.0 689550.0 92100.0 688350.0 ;
      RECT  86100.0 698250.0 87300.0 697050.0 ;
      RECT  88500.0 698250.0 89700.0 697050.0 ;
      RECT  88500.0 698250.0 89700.0 697050.0 ;
      RECT  86100.0 698250.0 87300.0 697050.0 ;
      RECT  88500.0 698250.0 89700.0 697050.0 ;
      RECT  90900.0 698250.0 92100.0 697050.0 ;
      RECT  90900.0 698250.0 92100.0 697050.0 ;
      RECT  88500.0 698250.0 89700.0 697050.0 ;
      RECT  90900.0 698250.0 92100.0 697050.0 ;
      RECT  93300.0 698250.0 94500.0 697050.0 ;
      RECT  93300.0 698250.0 94500.0 697050.0 ;
      RECT  90900.0 698250.0 92100.0 697050.0 ;
      RECT  95700.0 688950.0 96900.0 687750.0 ;
      RECT  95700.0 698850.0 96900.0 697650.0 ;
      RECT  93300.0 696150.0 92100.0 694950.0 ;
      RECT  90900.0 694200.0 89700.0 693000.0 ;
      RECT  88500.0 692250.0 87300.0 691050.0 ;
      RECT  88500.0 689550.0 89700.0 688350.0 ;
      RECT  93300.0 689550.0 94500.0 688350.0 ;
      RECT  93300.0 698250.0 94500.0 697050.0 ;
      RECT  93300.0 692250.0 94500.0 691050.0 ;
      RECT  87300.0 692250.0 88500.0 691050.0 ;
      RECT  89700.0 694200.0 90900.0 693000.0 ;
      RECT  92100.0 696150.0 93300.0 694950.0 ;
      RECT  93300.0 692250.0 94500.0 691050.0 ;
      RECT  84300.0 686850.0 99900.0 685950.0 ;
      RECT  84300.0 700650.0 99900.0 699750.0 ;
      RECT  86100.0 702150.0 87300.0 699750.0 ;
      RECT  86100.0 710850.0 87300.0 714450.0 ;
      RECT  90900.0 710850.0 92100.0 714450.0 ;
      RECT  95700.0 712050.0 96900.0 714000.0 ;
      RECT  95700.0 700200.0 96900.0 702150.0 ;
      RECT  86100.0 710850.0 87300.0 712050.0 ;
      RECT  88500.0 710850.0 89700.0 712050.0 ;
      RECT  88500.0 710850.0 89700.0 712050.0 ;
      RECT  86100.0 710850.0 87300.0 712050.0 ;
      RECT  88500.0 710850.0 89700.0 712050.0 ;
      RECT  90900.0 710850.0 92100.0 712050.0 ;
      RECT  90900.0 710850.0 92100.0 712050.0 ;
      RECT  88500.0 710850.0 89700.0 712050.0 ;
      RECT  90900.0 710850.0 92100.0 712050.0 ;
      RECT  93300.0 710850.0 94500.0 712050.0 ;
      RECT  93300.0 710850.0 94500.0 712050.0 ;
      RECT  90900.0 710850.0 92100.0 712050.0 ;
      RECT  86100.0 702150.0 87300.0 703350.0 ;
      RECT  88500.0 702150.0 89700.0 703350.0 ;
      RECT  88500.0 702150.0 89700.0 703350.0 ;
      RECT  86100.0 702150.0 87300.0 703350.0 ;
      RECT  88500.0 702150.0 89700.0 703350.0 ;
      RECT  90900.0 702150.0 92100.0 703350.0 ;
      RECT  90900.0 702150.0 92100.0 703350.0 ;
      RECT  88500.0 702150.0 89700.0 703350.0 ;
      RECT  90900.0 702150.0 92100.0 703350.0 ;
      RECT  93300.0 702150.0 94500.0 703350.0 ;
      RECT  93300.0 702150.0 94500.0 703350.0 ;
      RECT  90900.0 702150.0 92100.0 703350.0 ;
      RECT  95700.0 711450.0 96900.0 712650.0 ;
      RECT  95700.0 701550.0 96900.0 702750.0 ;
      RECT  93300.0 704250.0 92100.0 705450.0 ;
      RECT  90900.0 706200.0 89700.0 707400.0 ;
      RECT  88500.0 708150.0 87300.0 709350.0 ;
      RECT  88500.0 710850.0 89700.0 712050.0 ;
      RECT  93300.0 710850.0 94500.0 712050.0 ;
      RECT  93300.0 702150.0 94500.0 703350.0 ;
      RECT  93300.0 708150.0 94500.0 709350.0 ;
      RECT  87300.0 708150.0 88500.0 709350.0 ;
      RECT  89700.0 706200.0 90900.0 707400.0 ;
      RECT  92100.0 704250.0 93300.0 705450.0 ;
      RECT  93300.0 708150.0 94500.0 709350.0 ;
      RECT  84300.0 713550.0 99900.0 714450.0 ;
      RECT  84300.0 699750.0 99900.0 700650.0 ;
      RECT  86100.0 725850.0 87300.0 728250.0 ;
      RECT  86100.0 717150.0 87300.0 713550.0 ;
      RECT  90900.0 717150.0 92100.0 713550.0 ;
      RECT  95700.0 715950.0 96900.0 714000.0 ;
      RECT  95700.0 727800.0 96900.0 725850.0 ;
      RECT  86100.0 717150.0 87300.0 715950.0 ;
      RECT  88500.0 717150.0 89700.0 715950.0 ;
      RECT  88500.0 717150.0 89700.0 715950.0 ;
      RECT  86100.0 717150.0 87300.0 715950.0 ;
      RECT  88500.0 717150.0 89700.0 715950.0 ;
      RECT  90900.0 717150.0 92100.0 715950.0 ;
      RECT  90900.0 717150.0 92100.0 715950.0 ;
      RECT  88500.0 717150.0 89700.0 715950.0 ;
      RECT  90900.0 717150.0 92100.0 715950.0 ;
      RECT  93300.0 717150.0 94500.0 715950.0 ;
      RECT  93300.0 717150.0 94500.0 715950.0 ;
      RECT  90900.0 717150.0 92100.0 715950.0 ;
      RECT  86100.0 725850.0 87300.0 724650.0 ;
      RECT  88500.0 725850.0 89700.0 724650.0 ;
      RECT  88500.0 725850.0 89700.0 724650.0 ;
      RECT  86100.0 725850.0 87300.0 724650.0 ;
      RECT  88500.0 725850.0 89700.0 724650.0 ;
      RECT  90900.0 725850.0 92100.0 724650.0 ;
      RECT  90900.0 725850.0 92100.0 724650.0 ;
      RECT  88500.0 725850.0 89700.0 724650.0 ;
      RECT  90900.0 725850.0 92100.0 724650.0 ;
      RECT  93300.0 725850.0 94500.0 724650.0 ;
      RECT  93300.0 725850.0 94500.0 724650.0 ;
      RECT  90900.0 725850.0 92100.0 724650.0 ;
      RECT  95700.0 716550.0 96900.0 715350.0 ;
      RECT  95700.0 726450.0 96900.0 725250.0 ;
      RECT  93300.0 723750.0 92100.0 722550.0 ;
      RECT  90900.0 721800.0 89700.0 720600.0 ;
      RECT  88500.0 719850.0 87300.0 718650.0 ;
      RECT  88500.0 717150.0 89700.0 715950.0 ;
      RECT  93300.0 717150.0 94500.0 715950.0 ;
      RECT  93300.0 725850.0 94500.0 724650.0 ;
      RECT  93300.0 719850.0 94500.0 718650.0 ;
      RECT  87300.0 719850.0 88500.0 718650.0 ;
      RECT  89700.0 721800.0 90900.0 720600.0 ;
      RECT  92100.0 723750.0 93300.0 722550.0 ;
      RECT  93300.0 719850.0 94500.0 718650.0 ;
      RECT  84300.0 714450.0 99900.0 713550.0 ;
      RECT  84300.0 728250.0 99900.0 727350.0 ;
      RECT  86100.0 729750.0 87300.0 727350.0 ;
      RECT  86100.0 738450.0 87300.0 742050.0 ;
      RECT  90900.0 738450.0 92100.0 742050.0 ;
      RECT  95700.0 739650.0 96900.0 741600.0 ;
      RECT  95700.0 727800.0 96900.0 729750.0 ;
      RECT  86100.0 738450.0 87300.0 739650.0 ;
      RECT  88500.0 738450.0 89700.0 739650.0 ;
      RECT  88500.0 738450.0 89700.0 739650.0 ;
      RECT  86100.0 738450.0 87300.0 739650.0 ;
      RECT  88500.0 738450.0 89700.0 739650.0 ;
      RECT  90900.0 738450.0 92100.0 739650.0 ;
      RECT  90900.0 738450.0 92100.0 739650.0 ;
      RECT  88500.0 738450.0 89700.0 739650.0 ;
      RECT  90900.0 738450.0 92100.0 739650.0 ;
      RECT  93300.0 738450.0 94500.0 739650.0 ;
      RECT  93300.0 738450.0 94500.0 739650.0 ;
      RECT  90900.0 738450.0 92100.0 739650.0 ;
      RECT  86100.0 729750.0 87300.0 730950.0 ;
      RECT  88500.0 729750.0 89700.0 730950.0 ;
      RECT  88500.0 729750.0 89700.0 730950.0 ;
      RECT  86100.0 729750.0 87300.0 730950.0 ;
      RECT  88500.0 729750.0 89700.0 730950.0 ;
      RECT  90900.0 729750.0 92100.0 730950.0 ;
      RECT  90900.0 729750.0 92100.0 730950.0 ;
      RECT  88500.0 729750.0 89700.0 730950.0 ;
      RECT  90900.0 729750.0 92100.0 730950.0 ;
      RECT  93300.0 729750.0 94500.0 730950.0 ;
      RECT  93300.0 729750.0 94500.0 730950.0 ;
      RECT  90900.0 729750.0 92100.0 730950.0 ;
      RECT  95700.0 739050.0 96900.0 740250.0 ;
      RECT  95700.0 729150.0 96900.0 730350.0 ;
      RECT  93300.0 731850.0 92100.0 733050.0 ;
      RECT  90900.0 733800.0 89700.0 735000.0 ;
      RECT  88500.0 735750.0 87300.0 736950.0 ;
      RECT  88500.0 738450.0 89700.0 739650.0 ;
      RECT  93300.0 738450.0 94500.0 739650.0 ;
      RECT  93300.0 729750.0 94500.0 730950.0 ;
      RECT  93300.0 735750.0 94500.0 736950.0 ;
      RECT  87300.0 735750.0 88500.0 736950.0 ;
      RECT  89700.0 733800.0 90900.0 735000.0 ;
      RECT  92100.0 731850.0 93300.0 733050.0 ;
      RECT  93300.0 735750.0 94500.0 736950.0 ;
      RECT  84300.0 741150.0 99900.0 742050.0 ;
      RECT  84300.0 727350.0 99900.0 728250.0 ;
      RECT  86100.0 753450.0 87300.0 755850.0 ;
      RECT  86100.0 744750.0 87300.0 741150.0 ;
      RECT  90900.0 744750.0 92100.0 741150.0 ;
      RECT  95700.0 743550.0 96900.0 741600.0 ;
      RECT  95700.0 755400.0 96900.0 753450.0 ;
      RECT  86100.0 744750.0 87300.0 743550.0 ;
      RECT  88500.0 744750.0 89700.0 743550.0 ;
      RECT  88500.0 744750.0 89700.0 743550.0 ;
      RECT  86100.0 744750.0 87300.0 743550.0 ;
      RECT  88500.0 744750.0 89700.0 743550.0 ;
      RECT  90900.0 744750.0 92100.0 743550.0 ;
      RECT  90900.0 744750.0 92100.0 743550.0 ;
      RECT  88500.0 744750.0 89700.0 743550.0 ;
      RECT  90900.0 744750.0 92100.0 743550.0 ;
      RECT  93300.0 744750.0 94500.0 743550.0 ;
      RECT  93300.0 744750.0 94500.0 743550.0 ;
      RECT  90900.0 744750.0 92100.0 743550.0 ;
      RECT  86100.0 753450.0 87300.0 752250.0 ;
      RECT  88500.0 753450.0 89700.0 752250.0 ;
      RECT  88500.0 753450.0 89700.0 752250.0 ;
      RECT  86100.0 753450.0 87300.0 752250.0 ;
      RECT  88500.0 753450.0 89700.0 752250.0 ;
      RECT  90900.0 753450.0 92100.0 752250.0 ;
      RECT  90900.0 753450.0 92100.0 752250.0 ;
      RECT  88500.0 753450.0 89700.0 752250.0 ;
      RECT  90900.0 753450.0 92100.0 752250.0 ;
      RECT  93300.0 753450.0 94500.0 752250.0 ;
      RECT  93300.0 753450.0 94500.0 752250.0 ;
      RECT  90900.0 753450.0 92100.0 752250.0 ;
      RECT  95700.0 744150.0 96900.0 742950.0 ;
      RECT  95700.0 754050.0 96900.0 752850.0 ;
      RECT  93300.0 751350.0 92100.0 750150.0 ;
      RECT  90900.0 749400.0 89700.0 748200.0 ;
      RECT  88500.0 747450.0 87300.0 746250.0 ;
      RECT  88500.0 744750.0 89700.0 743550.0 ;
      RECT  93300.0 744750.0 94500.0 743550.0 ;
      RECT  93300.0 753450.0 94500.0 752250.0 ;
      RECT  93300.0 747450.0 94500.0 746250.0 ;
      RECT  87300.0 747450.0 88500.0 746250.0 ;
      RECT  89700.0 749400.0 90900.0 748200.0 ;
      RECT  92100.0 751350.0 93300.0 750150.0 ;
      RECT  93300.0 747450.0 94500.0 746250.0 ;
      RECT  84300.0 742050.0 99900.0 741150.0 ;
      RECT  84300.0 755850.0 99900.0 754950.0 ;
      RECT  86100.0 757350.0 87300.0 754950.0 ;
      RECT  86100.0 766050.0 87300.0 769650.0 ;
      RECT  90900.0 766050.0 92100.0 769650.0 ;
      RECT  95700.0 767250.0 96900.0 769200.0 ;
      RECT  95700.0 755400.0 96900.0 757350.0 ;
      RECT  86100.0 766050.0 87300.0 767250.0 ;
      RECT  88500.0 766050.0 89700.0 767250.0 ;
      RECT  88500.0 766050.0 89700.0 767250.0 ;
      RECT  86100.0 766050.0 87300.0 767250.0 ;
      RECT  88500.0 766050.0 89700.0 767250.0 ;
      RECT  90900.0 766050.0 92100.0 767250.0 ;
      RECT  90900.0 766050.0 92100.0 767250.0 ;
      RECT  88500.0 766050.0 89700.0 767250.0 ;
      RECT  90900.0 766050.0 92100.0 767250.0 ;
      RECT  93300.0 766050.0 94500.0 767250.0 ;
      RECT  93300.0 766050.0 94500.0 767250.0 ;
      RECT  90900.0 766050.0 92100.0 767250.0 ;
      RECT  86100.0 757350.0 87300.0 758550.0 ;
      RECT  88500.0 757350.0 89700.0 758550.0 ;
      RECT  88500.0 757350.0 89700.0 758550.0 ;
      RECT  86100.0 757350.0 87300.0 758550.0 ;
      RECT  88500.0 757350.0 89700.0 758550.0 ;
      RECT  90900.0 757350.0 92100.0 758550.0 ;
      RECT  90900.0 757350.0 92100.0 758550.0 ;
      RECT  88500.0 757350.0 89700.0 758550.0 ;
      RECT  90900.0 757350.0 92100.0 758550.0 ;
      RECT  93300.0 757350.0 94500.0 758550.0 ;
      RECT  93300.0 757350.0 94500.0 758550.0 ;
      RECT  90900.0 757350.0 92100.0 758550.0 ;
      RECT  95700.0 766650.0 96900.0 767850.0 ;
      RECT  95700.0 756750.0 96900.0 757950.0 ;
      RECT  93300.0 759450.0 92100.0 760650.0 ;
      RECT  90900.0 761400.0 89700.0 762600.0 ;
      RECT  88500.0 763350.0 87300.0 764550.0 ;
      RECT  88500.0 766050.0 89700.0 767250.0 ;
      RECT  93300.0 766050.0 94500.0 767250.0 ;
      RECT  93300.0 757350.0 94500.0 758550.0 ;
      RECT  93300.0 763350.0 94500.0 764550.0 ;
      RECT  87300.0 763350.0 88500.0 764550.0 ;
      RECT  89700.0 761400.0 90900.0 762600.0 ;
      RECT  92100.0 759450.0 93300.0 760650.0 ;
      RECT  93300.0 763350.0 94500.0 764550.0 ;
      RECT  84300.0 768750.0 99900.0 769650.0 ;
      RECT  84300.0 754950.0 99900.0 755850.0 ;
      RECT  86100.0 781050.0 87300.0 783450.0 ;
      RECT  86100.0 772350.0 87300.0 768750.0 ;
      RECT  90900.0 772350.0 92100.0 768750.0 ;
      RECT  95700.0 771150.0 96900.0 769200.0 ;
      RECT  95700.0 783000.0 96900.0 781050.0 ;
      RECT  86100.0 772350.0 87300.0 771150.0 ;
      RECT  88500.0 772350.0 89700.0 771150.0 ;
      RECT  88500.0 772350.0 89700.0 771150.0 ;
      RECT  86100.0 772350.0 87300.0 771150.0 ;
      RECT  88500.0 772350.0 89700.0 771150.0 ;
      RECT  90900.0 772350.0 92100.0 771150.0 ;
      RECT  90900.0 772350.0 92100.0 771150.0 ;
      RECT  88500.0 772350.0 89700.0 771150.0 ;
      RECT  90900.0 772350.0 92100.0 771150.0 ;
      RECT  93300.0 772350.0 94500.0 771150.0 ;
      RECT  93300.0 772350.0 94500.0 771150.0 ;
      RECT  90900.0 772350.0 92100.0 771150.0 ;
      RECT  86100.0 781050.0 87300.0 779850.0 ;
      RECT  88500.0 781050.0 89700.0 779850.0 ;
      RECT  88500.0 781050.0 89700.0 779850.0 ;
      RECT  86100.0 781050.0 87300.0 779850.0 ;
      RECT  88500.0 781050.0 89700.0 779850.0 ;
      RECT  90900.0 781050.0 92100.0 779850.0 ;
      RECT  90900.0 781050.0 92100.0 779850.0 ;
      RECT  88500.0 781050.0 89700.0 779850.0 ;
      RECT  90900.0 781050.0 92100.0 779850.0 ;
      RECT  93300.0 781050.0 94500.0 779850.0 ;
      RECT  93300.0 781050.0 94500.0 779850.0 ;
      RECT  90900.0 781050.0 92100.0 779850.0 ;
      RECT  95700.0 771750.0 96900.0 770550.0 ;
      RECT  95700.0 781650.0 96900.0 780450.0 ;
      RECT  93300.0 778950.0 92100.0 777750.0 ;
      RECT  90900.0 777000.0 89700.0 775800.0 ;
      RECT  88500.0 775050.0 87300.0 773850.0 ;
      RECT  88500.0 772350.0 89700.0 771150.0 ;
      RECT  93300.0 772350.0 94500.0 771150.0 ;
      RECT  93300.0 781050.0 94500.0 779850.0 ;
      RECT  93300.0 775050.0 94500.0 773850.0 ;
      RECT  87300.0 775050.0 88500.0 773850.0 ;
      RECT  89700.0 777000.0 90900.0 775800.0 ;
      RECT  92100.0 778950.0 93300.0 777750.0 ;
      RECT  93300.0 775050.0 94500.0 773850.0 ;
      RECT  84300.0 769650.0 99900.0 768750.0 ;
      RECT  84300.0 783450.0 99900.0 782550.0 ;
      RECT  86100.0 784950.0 87300.0 782550.0 ;
      RECT  86100.0 793650.0 87300.0 797250.0 ;
      RECT  90900.0 793650.0 92100.0 797250.0 ;
      RECT  95700.0 794850.0 96900.0 796800.0 ;
      RECT  95700.0 783000.0 96900.0 784950.0 ;
      RECT  86100.0 793650.0 87300.0 794850.0 ;
      RECT  88500.0 793650.0 89700.0 794850.0 ;
      RECT  88500.0 793650.0 89700.0 794850.0 ;
      RECT  86100.0 793650.0 87300.0 794850.0 ;
      RECT  88500.0 793650.0 89700.0 794850.0 ;
      RECT  90900.0 793650.0 92100.0 794850.0 ;
      RECT  90900.0 793650.0 92100.0 794850.0 ;
      RECT  88500.0 793650.0 89700.0 794850.0 ;
      RECT  90900.0 793650.0 92100.0 794850.0 ;
      RECT  93300.0 793650.0 94500.0 794850.0 ;
      RECT  93300.0 793650.0 94500.0 794850.0 ;
      RECT  90900.0 793650.0 92100.0 794850.0 ;
      RECT  86100.0 784950.0 87300.0 786150.0 ;
      RECT  88500.0 784950.0 89700.0 786150.0 ;
      RECT  88500.0 784950.0 89700.0 786150.0 ;
      RECT  86100.0 784950.0 87300.0 786150.0 ;
      RECT  88500.0 784950.0 89700.0 786150.0 ;
      RECT  90900.0 784950.0 92100.0 786150.0 ;
      RECT  90900.0 784950.0 92100.0 786150.0 ;
      RECT  88500.0 784950.0 89700.0 786150.0 ;
      RECT  90900.0 784950.0 92100.0 786150.0 ;
      RECT  93300.0 784950.0 94500.0 786150.0 ;
      RECT  93300.0 784950.0 94500.0 786150.0 ;
      RECT  90900.0 784950.0 92100.0 786150.0 ;
      RECT  95700.0 794250.0 96900.0 795450.0 ;
      RECT  95700.0 784350.0 96900.0 785550.0 ;
      RECT  93300.0 787050.0 92100.0 788250.0 ;
      RECT  90900.0 789000.0 89700.0 790200.0 ;
      RECT  88500.0 790950.0 87300.0 792150.0 ;
      RECT  88500.0 793650.0 89700.0 794850.0 ;
      RECT  93300.0 793650.0 94500.0 794850.0 ;
      RECT  93300.0 784950.0 94500.0 786150.0 ;
      RECT  93300.0 790950.0 94500.0 792150.0 ;
      RECT  87300.0 790950.0 88500.0 792150.0 ;
      RECT  89700.0 789000.0 90900.0 790200.0 ;
      RECT  92100.0 787050.0 93300.0 788250.0 ;
      RECT  93300.0 790950.0 94500.0 792150.0 ;
      RECT  84300.0 796350.0 99900.0 797250.0 ;
      RECT  84300.0 782550.0 99900.0 783450.0 ;
      RECT  86100.0 808650.0 87300.0 811050.0 ;
      RECT  86100.0 799950.0 87300.0 796350.0 ;
      RECT  90900.0 799950.0 92100.0 796350.0 ;
      RECT  95700.0 798750.0 96900.0 796800.0 ;
      RECT  95700.0 810600.0 96900.0 808650.0 ;
      RECT  86100.0 799950.0 87300.0 798750.0 ;
      RECT  88500.0 799950.0 89700.0 798750.0 ;
      RECT  88500.0 799950.0 89700.0 798750.0 ;
      RECT  86100.0 799950.0 87300.0 798750.0 ;
      RECT  88500.0 799950.0 89700.0 798750.0 ;
      RECT  90900.0 799950.0 92100.0 798750.0 ;
      RECT  90900.0 799950.0 92100.0 798750.0 ;
      RECT  88500.0 799950.0 89700.0 798750.0 ;
      RECT  90900.0 799950.0 92100.0 798750.0 ;
      RECT  93300.0 799950.0 94500.0 798750.0 ;
      RECT  93300.0 799950.0 94500.0 798750.0 ;
      RECT  90900.0 799950.0 92100.0 798750.0 ;
      RECT  86100.0 808650.0 87300.0 807450.0 ;
      RECT  88500.0 808650.0 89700.0 807450.0 ;
      RECT  88500.0 808650.0 89700.0 807450.0 ;
      RECT  86100.0 808650.0 87300.0 807450.0 ;
      RECT  88500.0 808650.0 89700.0 807450.0 ;
      RECT  90900.0 808650.0 92100.0 807450.0 ;
      RECT  90900.0 808650.0 92100.0 807450.0 ;
      RECT  88500.0 808650.0 89700.0 807450.0 ;
      RECT  90900.0 808650.0 92100.0 807450.0 ;
      RECT  93300.0 808650.0 94500.0 807450.0 ;
      RECT  93300.0 808650.0 94500.0 807450.0 ;
      RECT  90900.0 808650.0 92100.0 807450.0 ;
      RECT  95700.0 799350.0 96900.0 798150.0 ;
      RECT  95700.0 809250.0 96900.0 808050.0 ;
      RECT  93300.0 806550.0 92100.0 805350.0 ;
      RECT  90900.0 804600.0 89700.0 803400.0 ;
      RECT  88500.0 802650.0 87300.0 801450.0 ;
      RECT  88500.0 799950.0 89700.0 798750.0 ;
      RECT  93300.0 799950.0 94500.0 798750.0 ;
      RECT  93300.0 808650.0 94500.0 807450.0 ;
      RECT  93300.0 802650.0 94500.0 801450.0 ;
      RECT  87300.0 802650.0 88500.0 801450.0 ;
      RECT  89700.0 804600.0 90900.0 803400.0 ;
      RECT  92100.0 806550.0 93300.0 805350.0 ;
      RECT  93300.0 802650.0 94500.0 801450.0 ;
      RECT  84300.0 797250.0 99900.0 796350.0 ;
      RECT  84300.0 811050.0 99900.0 810150.0 ;
      RECT  86100.0 812550.0 87300.0 810150.0 ;
      RECT  86100.0 821250.0 87300.0 824850.0 ;
      RECT  90900.0 821250.0 92100.0 824850.0 ;
      RECT  95700.0 822450.0 96900.0 824400.0 ;
      RECT  95700.0 810600.0 96900.0 812550.0 ;
      RECT  86100.0 821250.0 87300.0 822450.0 ;
      RECT  88500.0 821250.0 89700.0 822450.0 ;
      RECT  88500.0 821250.0 89700.0 822450.0 ;
      RECT  86100.0 821250.0 87300.0 822450.0 ;
      RECT  88500.0 821250.0 89700.0 822450.0 ;
      RECT  90900.0 821250.0 92100.0 822450.0 ;
      RECT  90900.0 821250.0 92100.0 822450.0 ;
      RECT  88500.0 821250.0 89700.0 822450.0 ;
      RECT  90900.0 821250.0 92100.0 822450.0 ;
      RECT  93300.0 821250.0 94500.0 822450.0 ;
      RECT  93300.0 821250.0 94500.0 822450.0 ;
      RECT  90900.0 821250.0 92100.0 822450.0 ;
      RECT  86100.0 812550.0 87300.0 813750.0 ;
      RECT  88500.0 812550.0 89700.0 813750.0 ;
      RECT  88500.0 812550.0 89700.0 813750.0 ;
      RECT  86100.0 812550.0 87300.0 813750.0 ;
      RECT  88500.0 812550.0 89700.0 813750.0 ;
      RECT  90900.0 812550.0 92100.0 813750.0 ;
      RECT  90900.0 812550.0 92100.0 813750.0 ;
      RECT  88500.0 812550.0 89700.0 813750.0 ;
      RECT  90900.0 812550.0 92100.0 813750.0 ;
      RECT  93300.0 812550.0 94500.0 813750.0 ;
      RECT  93300.0 812550.0 94500.0 813750.0 ;
      RECT  90900.0 812550.0 92100.0 813750.0 ;
      RECT  95700.0 821850.0 96900.0 823050.0 ;
      RECT  95700.0 811950.0 96900.0 813150.0 ;
      RECT  93300.0 814650.0 92100.0 815850.0 ;
      RECT  90900.0 816600.0 89700.0 817800.0 ;
      RECT  88500.0 818550.0 87300.0 819750.0 ;
      RECT  88500.0 821250.0 89700.0 822450.0 ;
      RECT  93300.0 821250.0 94500.0 822450.0 ;
      RECT  93300.0 812550.0 94500.0 813750.0 ;
      RECT  93300.0 818550.0 94500.0 819750.0 ;
      RECT  87300.0 818550.0 88500.0 819750.0 ;
      RECT  89700.0 816600.0 90900.0 817800.0 ;
      RECT  92100.0 814650.0 93300.0 815850.0 ;
      RECT  93300.0 818550.0 94500.0 819750.0 ;
      RECT  84300.0 823950.0 99900.0 824850.0 ;
      RECT  84300.0 810150.0 99900.0 811050.0 ;
      RECT  86100.0 836250.0 87300.0 838650.0 ;
      RECT  86100.0 827550.0 87300.0 823950.0 ;
      RECT  90900.0 827550.0 92100.0 823950.0 ;
      RECT  95700.0 826350.0 96900.0 824400.0 ;
      RECT  95700.0 838200.0 96900.0 836250.0 ;
      RECT  86100.0 827550.0 87300.0 826350.0 ;
      RECT  88500.0 827550.0 89700.0 826350.0 ;
      RECT  88500.0 827550.0 89700.0 826350.0 ;
      RECT  86100.0 827550.0 87300.0 826350.0 ;
      RECT  88500.0 827550.0 89700.0 826350.0 ;
      RECT  90900.0 827550.0 92100.0 826350.0 ;
      RECT  90900.0 827550.0 92100.0 826350.0 ;
      RECT  88500.0 827550.0 89700.0 826350.0 ;
      RECT  90900.0 827550.0 92100.0 826350.0 ;
      RECT  93300.0 827550.0 94500.0 826350.0 ;
      RECT  93300.0 827550.0 94500.0 826350.0 ;
      RECT  90900.0 827550.0 92100.0 826350.0 ;
      RECT  86100.0 836250.0 87300.0 835050.0 ;
      RECT  88500.0 836250.0 89700.0 835050.0 ;
      RECT  88500.0 836250.0 89700.0 835050.0 ;
      RECT  86100.0 836250.0 87300.0 835050.0 ;
      RECT  88500.0 836250.0 89700.0 835050.0 ;
      RECT  90900.0 836250.0 92100.0 835050.0 ;
      RECT  90900.0 836250.0 92100.0 835050.0 ;
      RECT  88500.0 836250.0 89700.0 835050.0 ;
      RECT  90900.0 836250.0 92100.0 835050.0 ;
      RECT  93300.0 836250.0 94500.0 835050.0 ;
      RECT  93300.0 836250.0 94500.0 835050.0 ;
      RECT  90900.0 836250.0 92100.0 835050.0 ;
      RECT  95700.0 826950.0 96900.0 825750.0 ;
      RECT  95700.0 836850.0 96900.0 835650.0 ;
      RECT  93300.0 834150.0 92100.0 832950.0 ;
      RECT  90900.0 832200.0 89700.0 831000.0 ;
      RECT  88500.0 830250.0 87300.0 829050.0 ;
      RECT  88500.0 827550.0 89700.0 826350.0 ;
      RECT  93300.0 827550.0 94500.0 826350.0 ;
      RECT  93300.0 836250.0 94500.0 835050.0 ;
      RECT  93300.0 830250.0 94500.0 829050.0 ;
      RECT  87300.0 830250.0 88500.0 829050.0 ;
      RECT  89700.0 832200.0 90900.0 831000.0 ;
      RECT  92100.0 834150.0 93300.0 832950.0 ;
      RECT  93300.0 830250.0 94500.0 829050.0 ;
      RECT  84300.0 824850.0 99900.0 823950.0 ;
      RECT  84300.0 838650.0 99900.0 837750.0 ;
      RECT  86100.0 840150.0 87300.0 837750.0 ;
      RECT  86100.0 848850.0 87300.0 852450.0 ;
      RECT  90900.0 848850.0 92100.0 852450.0 ;
      RECT  95700.0 850050.0 96900.0 852000.0 ;
      RECT  95700.0 838200.0 96900.0 840150.0 ;
      RECT  86100.0 848850.0 87300.0 850050.0 ;
      RECT  88500.0 848850.0 89700.0 850050.0 ;
      RECT  88500.0 848850.0 89700.0 850050.0 ;
      RECT  86100.0 848850.0 87300.0 850050.0 ;
      RECT  88500.0 848850.0 89700.0 850050.0 ;
      RECT  90900.0 848850.0 92100.0 850050.0 ;
      RECT  90900.0 848850.0 92100.0 850050.0 ;
      RECT  88500.0 848850.0 89700.0 850050.0 ;
      RECT  90900.0 848850.0 92100.0 850050.0 ;
      RECT  93300.0 848850.0 94500.0 850050.0 ;
      RECT  93300.0 848850.0 94500.0 850050.0 ;
      RECT  90900.0 848850.0 92100.0 850050.0 ;
      RECT  86100.0 840150.0 87300.0 841350.0 ;
      RECT  88500.0 840150.0 89700.0 841350.0 ;
      RECT  88500.0 840150.0 89700.0 841350.0 ;
      RECT  86100.0 840150.0 87300.0 841350.0 ;
      RECT  88500.0 840150.0 89700.0 841350.0 ;
      RECT  90900.0 840150.0 92100.0 841350.0 ;
      RECT  90900.0 840150.0 92100.0 841350.0 ;
      RECT  88500.0 840150.0 89700.0 841350.0 ;
      RECT  90900.0 840150.0 92100.0 841350.0 ;
      RECT  93300.0 840150.0 94500.0 841350.0 ;
      RECT  93300.0 840150.0 94500.0 841350.0 ;
      RECT  90900.0 840150.0 92100.0 841350.0 ;
      RECT  95700.0 849450.0 96900.0 850650.0 ;
      RECT  95700.0 839550.0 96900.0 840750.0 ;
      RECT  93300.0 842250.0 92100.0 843450.0 ;
      RECT  90900.0 844200.0 89700.0 845400.0 ;
      RECT  88500.0 846150.0 87300.0 847350.0 ;
      RECT  88500.0 848850.0 89700.0 850050.0 ;
      RECT  93300.0 848850.0 94500.0 850050.0 ;
      RECT  93300.0 840150.0 94500.0 841350.0 ;
      RECT  93300.0 846150.0 94500.0 847350.0 ;
      RECT  87300.0 846150.0 88500.0 847350.0 ;
      RECT  89700.0 844200.0 90900.0 845400.0 ;
      RECT  92100.0 842250.0 93300.0 843450.0 ;
      RECT  93300.0 846150.0 94500.0 847350.0 ;
      RECT  84300.0 851550.0 99900.0 852450.0 ;
      RECT  84300.0 837750.0 99900.0 838650.0 ;
      RECT  86100.0 863850.0 87300.0 866250.0 ;
      RECT  86100.0 855150.0 87300.0 851550.0 ;
      RECT  90900.0 855150.0 92100.0 851550.0 ;
      RECT  95700.0 853950.0 96900.0 852000.0 ;
      RECT  95700.0 865800.0 96900.0 863850.0 ;
      RECT  86100.0 855150.0 87300.0 853950.0 ;
      RECT  88500.0 855150.0 89700.0 853950.0 ;
      RECT  88500.0 855150.0 89700.0 853950.0 ;
      RECT  86100.0 855150.0 87300.0 853950.0 ;
      RECT  88500.0 855150.0 89700.0 853950.0 ;
      RECT  90900.0 855150.0 92100.0 853950.0 ;
      RECT  90900.0 855150.0 92100.0 853950.0 ;
      RECT  88500.0 855150.0 89700.0 853950.0 ;
      RECT  90900.0 855150.0 92100.0 853950.0 ;
      RECT  93300.0 855150.0 94500.0 853950.0 ;
      RECT  93300.0 855150.0 94500.0 853950.0 ;
      RECT  90900.0 855150.0 92100.0 853950.0 ;
      RECT  86100.0 863850.0 87300.0 862650.0 ;
      RECT  88500.0 863850.0 89700.0 862650.0 ;
      RECT  88500.0 863850.0 89700.0 862650.0 ;
      RECT  86100.0 863850.0 87300.0 862650.0 ;
      RECT  88500.0 863850.0 89700.0 862650.0 ;
      RECT  90900.0 863850.0 92100.0 862650.0 ;
      RECT  90900.0 863850.0 92100.0 862650.0 ;
      RECT  88500.0 863850.0 89700.0 862650.0 ;
      RECT  90900.0 863850.0 92100.0 862650.0 ;
      RECT  93300.0 863850.0 94500.0 862650.0 ;
      RECT  93300.0 863850.0 94500.0 862650.0 ;
      RECT  90900.0 863850.0 92100.0 862650.0 ;
      RECT  95700.0 854550.0 96900.0 853350.0 ;
      RECT  95700.0 864450.0 96900.0 863250.0 ;
      RECT  93300.0 861750.0 92100.0 860550.0 ;
      RECT  90900.0 859800.0 89700.0 858600.0 ;
      RECT  88500.0 857850.0 87300.0 856650.0 ;
      RECT  88500.0 855150.0 89700.0 853950.0 ;
      RECT  93300.0 855150.0 94500.0 853950.0 ;
      RECT  93300.0 863850.0 94500.0 862650.0 ;
      RECT  93300.0 857850.0 94500.0 856650.0 ;
      RECT  87300.0 857850.0 88500.0 856650.0 ;
      RECT  89700.0 859800.0 90900.0 858600.0 ;
      RECT  92100.0 861750.0 93300.0 860550.0 ;
      RECT  93300.0 857850.0 94500.0 856650.0 ;
      RECT  84300.0 852450.0 99900.0 851550.0 ;
      RECT  84300.0 866250.0 99900.0 865350.0 ;
      RECT  86100.0 867750.0 87300.0 865350.0 ;
      RECT  86100.0 876450.0 87300.0 880050.0 ;
      RECT  90900.0 876450.0 92100.0 880050.0 ;
      RECT  95700.0 877650.0 96900.0 879600.0 ;
      RECT  95700.0 865800.0 96900.0 867750.0 ;
      RECT  86100.0 876450.0 87300.0 877650.0 ;
      RECT  88500.0 876450.0 89700.0 877650.0 ;
      RECT  88500.0 876450.0 89700.0 877650.0 ;
      RECT  86100.0 876450.0 87300.0 877650.0 ;
      RECT  88500.0 876450.0 89700.0 877650.0 ;
      RECT  90900.0 876450.0 92100.0 877650.0 ;
      RECT  90900.0 876450.0 92100.0 877650.0 ;
      RECT  88500.0 876450.0 89700.0 877650.0 ;
      RECT  90900.0 876450.0 92100.0 877650.0 ;
      RECT  93300.0 876450.0 94500.0 877650.0 ;
      RECT  93300.0 876450.0 94500.0 877650.0 ;
      RECT  90900.0 876450.0 92100.0 877650.0 ;
      RECT  86100.0 867750.0 87300.0 868950.0 ;
      RECT  88500.0 867750.0 89700.0 868950.0 ;
      RECT  88500.0 867750.0 89700.0 868950.0 ;
      RECT  86100.0 867750.0 87300.0 868950.0 ;
      RECT  88500.0 867750.0 89700.0 868950.0 ;
      RECT  90900.0 867750.0 92100.0 868950.0 ;
      RECT  90900.0 867750.0 92100.0 868950.0 ;
      RECT  88500.0 867750.0 89700.0 868950.0 ;
      RECT  90900.0 867750.0 92100.0 868950.0 ;
      RECT  93300.0 867750.0 94500.0 868950.0 ;
      RECT  93300.0 867750.0 94500.0 868950.0 ;
      RECT  90900.0 867750.0 92100.0 868950.0 ;
      RECT  95700.0 877050.0 96900.0 878250.0 ;
      RECT  95700.0 867150.0 96900.0 868350.0 ;
      RECT  93300.0 869850.0 92100.0 871050.0 ;
      RECT  90900.0 871800.0 89700.0 873000.0 ;
      RECT  88500.0 873750.0 87300.0 874950.0 ;
      RECT  88500.0 876450.0 89700.0 877650.0 ;
      RECT  93300.0 876450.0 94500.0 877650.0 ;
      RECT  93300.0 867750.0 94500.0 868950.0 ;
      RECT  93300.0 873750.0 94500.0 874950.0 ;
      RECT  87300.0 873750.0 88500.0 874950.0 ;
      RECT  89700.0 871800.0 90900.0 873000.0 ;
      RECT  92100.0 869850.0 93300.0 871050.0 ;
      RECT  93300.0 873750.0 94500.0 874950.0 ;
      RECT  84300.0 879150.0 99900.0 880050.0 ;
      RECT  84300.0 865350.0 99900.0 866250.0 ;
      RECT  86100.0 891450.0 87300.0 893850.0 ;
      RECT  86100.0 882750.0 87300.0 879150.0 ;
      RECT  90900.0 882750.0 92100.0 879150.0 ;
      RECT  95700.0 881550.0 96900.0 879600.0 ;
      RECT  95700.0 893400.0 96900.0 891450.0 ;
      RECT  86100.0 882750.0 87300.0 881550.0 ;
      RECT  88500.0 882750.0 89700.0 881550.0 ;
      RECT  88500.0 882750.0 89700.0 881550.0 ;
      RECT  86100.0 882750.0 87300.0 881550.0 ;
      RECT  88500.0 882750.0 89700.0 881550.0 ;
      RECT  90900.0 882750.0 92100.0 881550.0 ;
      RECT  90900.0 882750.0 92100.0 881550.0 ;
      RECT  88500.0 882750.0 89700.0 881550.0 ;
      RECT  90900.0 882750.0 92100.0 881550.0 ;
      RECT  93300.0 882750.0 94500.0 881550.0 ;
      RECT  93300.0 882750.0 94500.0 881550.0 ;
      RECT  90900.0 882750.0 92100.0 881550.0 ;
      RECT  86100.0 891450.0 87300.0 890250.0 ;
      RECT  88500.0 891450.0 89700.0 890250.0 ;
      RECT  88500.0 891450.0 89700.0 890250.0 ;
      RECT  86100.0 891450.0 87300.0 890250.0 ;
      RECT  88500.0 891450.0 89700.0 890250.0 ;
      RECT  90900.0 891450.0 92100.0 890250.0 ;
      RECT  90900.0 891450.0 92100.0 890250.0 ;
      RECT  88500.0 891450.0 89700.0 890250.0 ;
      RECT  90900.0 891450.0 92100.0 890250.0 ;
      RECT  93300.0 891450.0 94500.0 890250.0 ;
      RECT  93300.0 891450.0 94500.0 890250.0 ;
      RECT  90900.0 891450.0 92100.0 890250.0 ;
      RECT  95700.0 882150.0 96900.0 880950.0 ;
      RECT  95700.0 892050.0 96900.0 890850.0 ;
      RECT  93300.0 889350.0 92100.0 888150.0 ;
      RECT  90900.0 887400.0 89700.0 886200.0 ;
      RECT  88500.0 885450.0 87300.0 884250.0 ;
      RECT  88500.0 882750.0 89700.0 881550.0 ;
      RECT  93300.0 882750.0 94500.0 881550.0 ;
      RECT  93300.0 891450.0 94500.0 890250.0 ;
      RECT  93300.0 885450.0 94500.0 884250.0 ;
      RECT  87300.0 885450.0 88500.0 884250.0 ;
      RECT  89700.0 887400.0 90900.0 886200.0 ;
      RECT  92100.0 889350.0 93300.0 888150.0 ;
      RECT  93300.0 885450.0 94500.0 884250.0 ;
      RECT  84300.0 880050.0 99900.0 879150.0 ;
      RECT  84300.0 893850.0 99900.0 892950.0 ;
      RECT  86100.0 895350.0 87300.0 892950.0 ;
      RECT  86100.0 904050.0 87300.0 907650.0 ;
      RECT  90900.0 904050.0 92100.0 907650.0 ;
      RECT  95700.0 905250.0 96900.0 907200.0 ;
      RECT  95700.0 893400.0 96900.0 895350.0 ;
      RECT  86100.0 904050.0 87300.0 905250.0 ;
      RECT  88500.0 904050.0 89700.0 905250.0 ;
      RECT  88500.0 904050.0 89700.0 905250.0 ;
      RECT  86100.0 904050.0 87300.0 905250.0 ;
      RECT  88500.0 904050.0 89700.0 905250.0 ;
      RECT  90900.0 904050.0 92100.0 905250.0 ;
      RECT  90900.0 904050.0 92100.0 905250.0 ;
      RECT  88500.0 904050.0 89700.0 905250.0 ;
      RECT  90900.0 904050.0 92100.0 905250.0 ;
      RECT  93300.0 904050.0 94500.0 905250.0 ;
      RECT  93300.0 904050.0 94500.0 905250.0 ;
      RECT  90900.0 904050.0 92100.0 905250.0 ;
      RECT  86100.0 895350.0 87300.0 896550.0 ;
      RECT  88500.0 895350.0 89700.0 896550.0 ;
      RECT  88500.0 895350.0 89700.0 896550.0 ;
      RECT  86100.0 895350.0 87300.0 896550.0 ;
      RECT  88500.0 895350.0 89700.0 896550.0 ;
      RECT  90900.0 895350.0 92100.0 896550.0 ;
      RECT  90900.0 895350.0 92100.0 896550.0 ;
      RECT  88500.0 895350.0 89700.0 896550.0 ;
      RECT  90900.0 895350.0 92100.0 896550.0 ;
      RECT  93300.0 895350.0 94500.0 896550.0 ;
      RECT  93300.0 895350.0 94500.0 896550.0 ;
      RECT  90900.0 895350.0 92100.0 896550.0 ;
      RECT  95700.0 904650.0 96900.0 905850.0 ;
      RECT  95700.0 894750.0 96900.0 895950.0 ;
      RECT  93300.0 897450.0 92100.0 898650.0 ;
      RECT  90900.0 899400.0 89700.0 900600.0 ;
      RECT  88500.0 901350.0 87300.0 902550.0 ;
      RECT  88500.0 904050.0 89700.0 905250.0 ;
      RECT  93300.0 904050.0 94500.0 905250.0 ;
      RECT  93300.0 895350.0 94500.0 896550.0 ;
      RECT  93300.0 901350.0 94500.0 902550.0 ;
      RECT  87300.0 901350.0 88500.0 902550.0 ;
      RECT  89700.0 899400.0 90900.0 900600.0 ;
      RECT  92100.0 897450.0 93300.0 898650.0 ;
      RECT  93300.0 901350.0 94500.0 902550.0 ;
      RECT  84300.0 906750.0 99900.0 907650.0 ;
      RECT  84300.0 892950.0 99900.0 893850.0 ;
      RECT  86100.0 919050.0 87300.0 921450.0 ;
      RECT  86100.0 910350.0 87300.0 906750.0 ;
      RECT  90900.0 910350.0 92100.0 906750.0 ;
      RECT  95700.0 909150.0 96900.0 907200.0 ;
      RECT  95700.0 921000.0 96900.0 919050.0 ;
      RECT  86100.0 910350.0 87300.0 909150.0 ;
      RECT  88500.0 910350.0 89700.0 909150.0 ;
      RECT  88500.0 910350.0 89700.0 909150.0 ;
      RECT  86100.0 910350.0 87300.0 909150.0 ;
      RECT  88500.0 910350.0 89700.0 909150.0 ;
      RECT  90900.0 910350.0 92100.0 909150.0 ;
      RECT  90900.0 910350.0 92100.0 909150.0 ;
      RECT  88500.0 910350.0 89700.0 909150.0 ;
      RECT  90900.0 910350.0 92100.0 909150.0 ;
      RECT  93300.0 910350.0 94500.0 909150.0 ;
      RECT  93300.0 910350.0 94500.0 909150.0 ;
      RECT  90900.0 910350.0 92100.0 909150.0 ;
      RECT  86100.0 919050.0 87300.0 917850.0 ;
      RECT  88500.0 919050.0 89700.0 917850.0 ;
      RECT  88500.0 919050.0 89700.0 917850.0 ;
      RECT  86100.0 919050.0 87300.0 917850.0 ;
      RECT  88500.0 919050.0 89700.0 917850.0 ;
      RECT  90900.0 919050.0 92100.0 917850.0 ;
      RECT  90900.0 919050.0 92100.0 917850.0 ;
      RECT  88500.0 919050.0 89700.0 917850.0 ;
      RECT  90900.0 919050.0 92100.0 917850.0 ;
      RECT  93300.0 919050.0 94500.0 917850.0 ;
      RECT  93300.0 919050.0 94500.0 917850.0 ;
      RECT  90900.0 919050.0 92100.0 917850.0 ;
      RECT  95700.0 909750.0 96900.0 908550.0 ;
      RECT  95700.0 919650.0 96900.0 918450.0 ;
      RECT  93300.0 916950.0 92100.0 915750.0 ;
      RECT  90900.0 915000.0 89700.0 913800.0 ;
      RECT  88500.0 913050.0 87300.0 911850.0 ;
      RECT  88500.0 910350.0 89700.0 909150.0 ;
      RECT  93300.0 910350.0 94500.0 909150.0 ;
      RECT  93300.0 919050.0 94500.0 917850.0 ;
      RECT  93300.0 913050.0 94500.0 911850.0 ;
      RECT  87300.0 913050.0 88500.0 911850.0 ;
      RECT  89700.0 915000.0 90900.0 913800.0 ;
      RECT  92100.0 916950.0 93300.0 915750.0 ;
      RECT  93300.0 913050.0 94500.0 911850.0 ;
      RECT  84300.0 907650.0 99900.0 906750.0 ;
      RECT  84300.0 921450.0 99900.0 920550.0 ;
      RECT  86100.0 922950.0 87300.0 920550.0 ;
      RECT  86100.0 931650.0 87300.0 935250.0 ;
      RECT  90900.0 931650.0 92100.0 935250.0 ;
      RECT  95700.0 932850.0 96900.0 934800.0 ;
      RECT  95700.0 921000.0 96900.0 922950.0 ;
      RECT  86100.0 931650.0 87300.0 932850.0 ;
      RECT  88500.0 931650.0 89700.0 932850.0 ;
      RECT  88500.0 931650.0 89700.0 932850.0 ;
      RECT  86100.0 931650.0 87300.0 932850.0 ;
      RECT  88500.0 931650.0 89700.0 932850.0 ;
      RECT  90900.0 931650.0 92100.0 932850.0 ;
      RECT  90900.0 931650.0 92100.0 932850.0 ;
      RECT  88500.0 931650.0 89700.0 932850.0 ;
      RECT  90900.0 931650.0 92100.0 932850.0 ;
      RECT  93300.0 931650.0 94500.0 932850.0 ;
      RECT  93300.0 931650.0 94500.0 932850.0 ;
      RECT  90900.0 931650.0 92100.0 932850.0 ;
      RECT  86100.0 922950.0 87300.0 924150.0 ;
      RECT  88500.0 922950.0 89700.0 924150.0 ;
      RECT  88500.0 922950.0 89700.0 924150.0 ;
      RECT  86100.0 922950.0 87300.0 924150.0 ;
      RECT  88500.0 922950.0 89700.0 924150.0 ;
      RECT  90900.0 922950.0 92100.0 924150.0 ;
      RECT  90900.0 922950.0 92100.0 924150.0 ;
      RECT  88500.0 922950.0 89700.0 924150.0 ;
      RECT  90900.0 922950.0 92100.0 924150.0 ;
      RECT  93300.0 922950.0 94500.0 924150.0 ;
      RECT  93300.0 922950.0 94500.0 924150.0 ;
      RECT  90900.0 922950.0 92100.0 924150.0 ;
      RECT  95700.0 932250.0 96900.0 933450.0 ;
      RECT  95700.0 922350.0 96900.0 923550.0 ;
      RECT  93300.0 925050.0 92100.0 926250.0 ;
      RECT  90900.0 927000.0 89700.0 928200.0 ;
      RECT  88500.0 928950.0 87300.0 930150.0 ;
      RECT  88500.0 931650.0 89700.0 932850.0 ;
      RECT  93300.0 931650.0 94500.0 932850.0 ;
      RECT  93300.0 922950.0 94500.0 924150.0 ;
      RECT  93300.0 928950.0 94500.0 930150.0 ;
      RECT  87300.0 928950.0 88500.0 930150.0 ;
      RECT  89700.0 927000.0 90900.0 928200.0 ;
      RECT  92100.0 925050.0 93300.0 926250.0 ;
      RECT  93300.0 928950.0 94500.0 930150.0 ;
      RECT  84300.0 934350.0 99900.0 935250.0 ;
      RECT  84300.0 920550.0 99900.0 921450.0 ;
      RECT  86100.0 946650.0 87300.0 949050.0 ;
      RECT  86100.0 937950.0 87300.0 934350.0 ;
      RECT  90900.0 937950.0 92100.0 934350.0 ;
      RECT  95700.0 936750.0 96900.0 934800.0 ;
      RECT  95700.0 948600.0 96900.0 946650.0 ;
      RECT  86100.0 937950.0 87300.0 936750.0 ;
      RECT  88500.0 937950.0 89700.0 936750.0 ;
      RECT  88500.0 937950.0 89700.0 936750.0 ;
      RECT  86100.0 937950.0 87300.0 936750.0 ;
      RECT  88500.0 937950.0 89700.0 936750.0 ;
      RECT  90900.0 937950.0 92100.0 936750.0 ;
      RECT  90900.0 937950.0 92100.0 936750.0 ;
      RECT  88500.0 937950.0 89700.0 936750.0 ;
      RECT  90900.0 937950.0 92100.0 936750.0 ;
      RECT  93300.0 937950.0 94500.0 936750.0 ;
      RECT  93300.0 937950.0 94500.0 936750.0 ;
      RECT  90900.0 937950.0 92100.0 936750.0 ;
      RECT  86100.0 946650.0 87300.0 945450.0 ;
      RECT  88500.0 946650.0 89700.0 945450.0 ;
      RECT  88500.0 946650.0 89700.0 945450.0 ;
      RECT  86100.0 946650.0 87300.0 945450.0 ;
      RECT  88500.0 946650.0 89700.0 945450.0 ;
      RECT  90900.0 946650.0 92100.0 945450.0 ;
      RECT  90900.0 946650.0 92100.0 945450.0 ;
      RECT  88500.0 946650.0 89700.0 945450.0 ;
      RECT  90900.0 946650.0 92100.0 945450.0 ;
      RECT  93300.0 946650.0 94500.0 945450.0 ;
      RECT  93300.0 946650.0 94500.0 945450.0 ;
      RECT  90900.0 946650.0 92100.0 945450.0 ;
      RECT  95700.0 937350.0 96900.0 936150.0 ;
      RECT  95700.0 947250.0 96900.0 946050.0 ;
      RECT  93300.0 944550.0 92100.0 943350.0 ;
      RECT  90900.0 942600.0 89700.0 941400.0 ;
      RECT  88500.0 940650.0 87300.0 939450.0 ;
      RECT  88500.0 937950.0 89700.0 936750.0 ;
      RECT  93300.0 937950.0 94500.0 936750.0 ;
      RECT  93300.0 946650.0 94500.0 945450.0 ;
      RECT  93300.0 940650.0 94500.0 939450.0 ;
      RECT  87300.0 940650.0 88500.0 939450.0 ;
      RECT  89700.0 942600.0 90900.0 941400.0 ;
      RECT  92100.0 944550.0 93300.0 943350.0 ;
      RECT  93300.0 940650.0 94500.0 939450.0 ;
      RECT  84300.0 935250.0 99900.0 934350.0 ;
      RECT  84300.0 949050.0 99900.0 948150.0 ;
      RECT  86100.0 950550.0 87300.0 948150.0 ;
      RECT  86100.0 959250.0 87300.0 962850.0 ;
      RECT  90900.0 959250.0 92100.0 962850.0 ;
      RECT  95700.0 960450.0 96900.0 962400.0 ;
      RECT  95700.0 948600.0 96900.0 950550.0 ;
      RECT  86100.0 959250.0 87300.0 960450.0 ;
      RECT  88500.0 959250.0 89700.0 960450.0 ;
      RECT  88500.0 959250.0 89700.0 960450.0 ;
      RECT  86100.0 959250.0 87300.0 960450.0 ;
      RECT  88500.0 959250.0 89700.0 960450.0 ;
      RECT  90900.0 959250.0 92100.0 960450.0 ;
      RECT  90900.0 959250.0 92100.0 960450.0 ;
      RECT  88500.0 959250.0 89700.0 960450.0 ;
      RECT  90900.0 959250.0 92100.0 960450.0 ;
      RECT  93300.0 959250.0 94500.0 960450.0 ;
      RECT  93300.0 959250.0 94500.0 960450.0 ;
      RECT  90900.0 959250.0 92100.0 960450.0 ;
      RECT  86100.0 950550.0 87300.0 951750.0 ;
      RECT  88500.0 950550.0 89700.0 951750.0 ;
      RECT  88500.0 950550.0 89700.0 951750.0 ;
      RECT  86100.0 950550.0 87300.0 951750.0 ;
      RECT  88500.0 950550.0 89700.0 951750.0 ;
      RECT  90900.0 950550.0 92100.0 951750.0 ;
      RECT  90900.0 950550.0 92100.0 951750.0 ;
      RECT  88500.0 950550.0 89700.0 951750.0 ;
      RECT  90900.0 950550.0 92100.0 951750.0 ;
      RECT  93300.0 950550.0 94500.0 951750.0 ;
      RECT  93300.0 950550.0 94500.0 951750.0 ;
      RECT  90900.0 950550.0 92100.0 951750.0 ;
      RECT  95700.0 959850.0 96900.0 961050.0 ;
      RECT  95700.0 949950.0 96900.0 951150.0 ;
      RECT  93300.0 952650.0 92100.0 953850.0 ;
      RECT  90900.0 954600.0 89700.0 955800.0 ;
      RECT  88500.0 956550.0 87300.0 957750.0 ;
      RECT  88500.0 959250.0 89700.0 960450.0 ;
      RECT  93300.0 959250.0 94500.0 960450.0 ;
      RECT  93300.0 950550.0 94500.0 951750.0 ;
      RECT  93300.0 956550.0 94500.0 957750.0 ;
      RECT  87300.0 956550.0 88500.0 957750.0 ;
      RECT  89700.0 954600.0 90900.0 955800.0 ;
      RECT  92100.0 952650.0 93300.0 953850.0 ;
      RECT  93300.0 956550.0 94500.0 957750.0 ;
      RECT  84300.0 961950.0 99900.0 962850.0 ;
      RECT  84300.0 948150.0 99900.0 949050.0 ;
      RECT  86100.0 974250.0 87300.0 976650.0 ;
      RECT  86100.0 965550.0 87300.0 961950.0 ;
      RECT  90900.0 965550.0 92100.0 961950.0 ;
      RECT  95700.0 964350.0 96900.0 962400.0 ;
      RECT  95700.0 976200.0 96900.0 974250.0 ;
      RECT  86100.0 965550.0 87300.0 964350.0 ;
      RECT  88500.0 965550.0 89700.0 964350.0 ;
      RECT  88500.0 965550.0 89700.0 964350.0 ;
      RECT  86100.0 965550.0 87300.0 964350.0 ;
      RECT  88500.0 965550.0 89700.0 964350.0 ;
      RECT  90900.0 965550.0 92100.0 964350.0 ;
      RECT  90900.0 965550.0 92100.0 964350.0 ;
      RECT  88500.0 965550.0 89700.0 964350.0 ;
      RECT  90900.0 965550.0 92100.0 964350.0 ;
      RECT  93300.0 965550.0 94500.0 964350.0 ;
      RECT  93300.0 965550.0 94500.0 964350.0 ;
      RECT  90900.0 965550.0 92100.0 964350.0 ;
      RECT  86100.0 974250.0 87300.0 973050.0 ;
      RECT  88500.0 974250.0 89700.0 973050.0 ;
      RECT  88500.0 974250.0 89700.0 973050.0 ;
      RECT  86100.0 974250.0 87300.0 973050.0 ;
      RECT  88500.0 974250.0 89700.0 973050.0 ;
      RECT  90900.0 974250.0 92100.0 973050.0 ;
      RECT  90900.0 974250.0 92100.0 973050.0 ;
      RECT  88500.0 974250.0 89700.0 973050.0 ;
      RECT  90900.0 974250.0 92100.0 973050.0 ;
      RECT  93300.0 974250.0 94500.0 973050.0 ;
      RECT  93300.0 974250.0 94500.0 973050.0 ;
      RECT  90900.0 974250.0 92100.0 973050.0 ;
      RECT  95700.0 964950.0 96900.0 963750.0 ;
      RECT  95700.0 974850.0 96900.0 973650.0 ;
      RECT  93300.0 972150.0 92100.0 970950.0 ;
      RECT  90900.0 970200.0 89700.0 969000.0 ;
      RECT  88500.0 968250.0 87300.0 967050.0 ;
      RECT  88500.0 965550.0 89700.0 964350.0 ;
      RECT  93300.0 965550.0 94500.0 964350.0 ;
      RECT  93300.0 974250.0 94500.0 973050.0 ;
      RECT  93300.0 968250.0 94500.0 967050.0 ;
      RECT  87300.0 968250.0 88500.0 967050.0 ;
      RECT  89700.0 970200.0 90900.0 969000.0 ;
      RECT  92100.0 972150.0 93300.0 970950.0 ;
      RECT  93300.0 968250.0 94500.0 967050.0 ;
      RECT  84300.0 962850.0 99900.0 961950.0 ;
      RECT  84300.0 976650.0 99900.0 975750.0 ;
      RECT  86100.0 978150.0 87300.0 975750.0 ;
      RECT  86100.0 986850.0 87300.0 990450.0 ;
      RECT  90900.0 986850.0 92100.0 990450.0 ;
      RECT  95700.0 988050.0 96900.0 990000.0 ;
      RECT  95700.0 976200.0 96900.0 978150.0 ;
      RECT  86100.0 986850.0 87300.0 988050.0 ;
      RECT  88500.0 986850.0 89700.0 988050.0 ;
      RECT  88500.0 986850.0 89700.0 988050.0 ;
      RECT  86100.0 986850.0 87300.0 988050.0 ;
      RECT  88500.0 986850.0 89700.0 988050.0 ;
      RECT  90900.0 986850.0 92100.0 988050.0 ;
      RECT  90900.0 986850.0 92100.0 988050.0 ;
      RECT  88500.0 986850.0 89700.0 988050.0 ;
      RECT  90900.0 986850.0 92100.0 988050.0 ;
      RECT  93300.0 986850.0 94500.0 988050.0 ;
      RECT  93300.0 986850.0 94500.0 988050.0 ;
      RECT  90900.0 986850.0 92100.0 988050.0 ;
      RECT  86100.0 978150.0 87300.0 979350.0 ;
      RECT  88500.0 978150.0 89700.0 979350.0 ;
      RECT  88500.0 978150.0 89700.0 979350.0 ;
      RECT  86100.0 978150.0 87300.0 979350.0 ;
      RECT  88500.0 978150.0 89700.0 979350.0 ;
      RECT  90900.0 978150.0 92100.0 979350.0 ;
      RECT  90900.0 978150.0 92100.0 979350.0 ;
      RECT  88500.0 978150.0 89700.0 979350.0 ;
      RECT  90900.0 978150.0 92100.0 979350.0 ;
      RECT  93300.0 978150.0 94500.0 979350.0 ;
      RECT  93300.0 978150.0 94500.0 979350.0 ;
      RECT  90900.0 978150.0 92100.0 979350.0 ;
      RECT  95700.0 987450.0 96900.0 988650.0 ;
      RECT  95700.0 977550.0 96900.0 978750.0 ;
      RECT  93300.0 980250.0 92100.0 981450.0 ;
      RECT  90900.0 982200.0 89700.0 983400.0 ;
      RECT  88500.0 984150.0 87300.0 985350.0 ;
      RECT  88500.0 986850.0 89700.0 988050.0 ;
      RECT  93300.0 986850.0 94500.0 988050.0 ;
      RECT  93300.0 978150.0 94500.0 979350.0 ;
      RECT  93300.0 984150.0 94500.0 985350.0 ;
      RECT  87300.0 984150.0 88500.0 985350.0 ;
      RECT  89700.0 982200.0 90900.0 983400.0 ;
      RECT  92100.0 980250.0 93300.0 981450.0 ;
      RECT  93300.0 984150.0 94500.0 985350.0 ;
      RECT  84300.0 989550.0 99900.0 990450.0 ;
      RECT  84300.0 975750.0 99900.0 976650.0 ;
      RECT  86100.0 1001850.0 87300.0 1004250.0 ;
      RECT  86100.0 993150.0 87300.0 989550.0 ;
      RECT  90900.0 993150.0 92100.0 989550.0 ;
      RECT  95700.0 991950.0 96900.0 990000.0 ;
      RECT  95700.0 1003800.0 96900.0 1001850.0 ;
      RECT  86100.0 993150.0 87300.0 991950.0 ;
      RECT  88500.0 993150.0 89700.0 991950.0 ;
      RECT  88500.0 993150.0 89700.0 991950.0 ;
      RECT  86100.0 993150.0 87300.0 991950.0 ;
      RECT  88500.0 993150.0 89700.0 991950.0 ;
      RECT  90900.0 993150.0 92100.0 991950.0 ;
      RECT  90900.0 993150.0 92100.0 991950.0 ;
      RECT  88500.0 993150.0 89700.0 991950.0 ;
      RECT  90900.0 993150.0 92100.0 991950.0 ;
      RECT  93300.0 993150.0 94500.0 991950.0 ;
      RECT  93300.0 993150.0 94500.0 991950.0 ;
      RECT  90900.0 993150.0 92100.0 991950.0 ;
      RECT  86100.0 1001850.0 87300.0 1000650.0 ;
      RECT  88500.0 1001850.0 89700.0 1000650.0 ;
      RECT  88500.0 1001850.0 89700.0 1000650.0 ;
      RECT  86100.0 1001850.0 87300.0 1000650.0 ;
      RECT  88500.0 1001850.0 89700.0 1000650.0 ;
      RECT  90900.0 1001850.0 92100.0 1000650.0 ;
      RECT  90900.0 1001850.0 92100.0 1000650.0 ;
      RECT  88500.0 1001850.0 89700.0 1000650.0 ;
      RECT  90900.0 1001850.0 92100.0 1000650.0 ;
      RECT  93300.0 1001850.0 94500.0 1000650.0 ;
      RECT  93300.0 1001850.0 94500.0 1000650.0 ;
      RECT  90900.0 1001850.0 92100.0 1000650.0 ;
      RECT  95700.0 992550.0 96900.0 991350.0 ;
      RECT  95700.0 1002450.0 96900.0 1001250.0 ;
      RECT  93300.0 999750.0 92100.0 998550.0 ;
      RECT  90900.0 997800.0 89700.0 996600.0 ;
      RECT  88500.0 995850.0 87300.0 994650.0 ;
      RECT  88500.0 993150.0 89700.0 991950.0 ;
      RECT  93300.0 993150.0 94500.0 991950.0 ;
      RECT  93300.0 1001850.0 94500.0 1000650.0 ;
      RECT  93300.0 995850.0 94500.0 994650.0 ;
      RECT  87300.0 995850.0 88500.0 994650.0 ;
      RECT  89700.0 997800.0 90900.0 996600.0 ;
      RECT  92100.0 999750.0 93300.0 998550.0 ;
      RECT  93300.0 995850.0 94500.0 994650.0 ;
      RECT  84300.0 990450.0 99900.0 989550.0 ;
      RECT  84300.0 1004250.0 99900.0 1003350.0 ;
      RECT  86100.0 1005750.0 87300.0 1003350.0 ;
      RECT  86100.0 1014450.0 87300.0 1018050.0 ;
      RECT  90900.0 1014450.0 92100.0 1018050.0 ;
      RECT  95700.0 1015650.0 96900.0 1017600.0 ;
      RECT  95700.0 1003800.0 96900.0 1005750.0 ;
      RECT  86100.0 1014450.0 87300.0 1015650.0 ;
      RECT  88500.0 1014450.0 89700.0 1015650.0 ;
      RECT  88500.0 1014450.0 89700.0 1015650.0 ;
      RECT  86100.0 1014450.0 87300.0 1015650.0 ;
      RECT  88500.0 1014450.0 89700.0 1015650.0 ;
      RECT  90900.0 1014450.0 92100.0 1015650.0 ;
      RECT  90900.0 1014450.0 92100.0 1015650.0 ;
      RECT  88500.0 1014450.0 89700.0 1015650.0 ;
      RECT  90900.0 1014450.0 92100.0 1015650.0 ;
      RECT  93300.0 1014450.0 94500.0 1015650.0 ;
      RECT  93300.0 1014450.0 94500.0 1015650.0 ;
      RECT  90900.0 1014450.0 92100.0 1015650.0 ;
      RECT  86100.0 1005750.0 87300.0 1006950.0 ;
      RECT  88500.0 1005750.0 89700.0 1006950.0 ;
      RECT  88500.0 1005750.0 89700.0 1006950.0 ;
      RECT  86100.0 1005750.0 87300.0 1006950.0 ;
      RECT  88500.0 1005750.0 89700.0 1006950.0 ;
      RECT  90900.0 1005750.0 92100.0 1006950.0 ;
      RECT  90900.0 1005750.0 92100.0 1006950.0 ;
      RECT  88500.0 1005750.0 89700.0 1006950.0 ;
      RECT  90900.0 1005750.0 92100.0 1006950.0 ;
      RECT  93300.0 1005750.0 94500.0 1006950.0 ;
      RECT  93300.0 1005750.0 94500.0 1006950.0 ;
      RECT  90900.0 1005750.0 92100.0 1006950.0 ;
      RECT  95700.0 1015050.0 96900.0 1016250.0 ;
      RECT  95700.0 1005150.0 96900.0 1006350.0 ;
      RECT  93300.0 1007850.0 92100.0 1009050.0 ;
      RECT  90900.0 1009800.0 89700.0 1011000.0 ;
      RECT  88500.0 1011750.0 87300.0 1012950.0 ;
      RECT  88500.0 1014450.0 89700.0 1015650.0 ;
      RECT  93300.0 1014450.0 94500.0 1015650.0 ;
      RECT  93300.0 1005750.0 94500.0 1006950.0 ;
      RECT  93300.0 1011750.0 94500.0 1012950.0 ;
      RECT  87300.0 1011750.0 88500.0 1012950.0 ;
      RECT  89700.0 1009800.0 90900.0 1011000.0 ;
      RECT  92100.0 1007850.0 93300.0 1009050.0 ;
      RECT  93300.0 1011750.0 94500.0 1012950.0 ;
      RECT  84300.0 1017150.0 99900.0 1018050.0 ;
      RECT  84300.0 1003350.0 99900.0 1004250.0 ;
      RECT  86100.0 1029450.0 87300.0 1031850.0 ;
      RECT  86100.0 1020750.0 87300.0 1017150.0 ;
      RECT  90900.0 1020750.0 92100.0 1017150.0 ;
      RECT  95700.0 1019550.0 96900.0 1017600.0 ;
      RECT  95700.0 1031400.0 96900.0 1029450.0 ;
      RECT  86100.0 1020750.0 87300.0 1019550.0 ;
      RECT  88500.0 1020750.0 89700.0 1019550.0 ;
      RECT  88500.0 1020750.0 89700.0 1019550.0 ;
      RECT  86100.0 1020750.0 87300.0 1019550.0 ;
      RECT  88500.0 1020750.0 89700.0 1019550.0 ;
      RECT  90900.0 1020750.0 92100.0 1019550.0 ;
      RECT  90900.0 1020750.0 92100.0 1019550.0 ;
      RECT  88500.0 1020750.0 89700.0 1019550.0 ;
      RECT  90900.0 1020750.0 92100.0 1019550.0 ;
      RECT  93300.0 1020750.0 94500.0 1019550.0 ;
      RECT  93300.0 1020750.0 94500.0 1019550.0 ;
      RECT  90900.0 1020750.0 92100.0 1019550.0 ;
      RECT  86100.0 1029450.0 87300.0 1028250.0 ;
      RECT  88500.0 1029450.0 89700.0 1028250.0 ;
      RECT  88500.0 1029450.0 89700.0 1028250.0 ;
      RECT  86100.0 1029450.0 87300.0 1028250.0 ;
      RECT  88500.0 1029450.0 89700.0 1028250.0 ;
      RECT  90900.0 1029450.0 92100.0 1028250.0 ;
      RECT  90900.0 1029450.0 92100.0 1028250.0 ;
      RECT  88500.0 1029450.0 89700.0 1028250.0 ;
      RECT  90900.0 1029450.0 92100.0 1028250.0 ;
      RECT  93300.0 1029450.0 94500.0 1028250.0 ;
      RECT  93300.0 1029450.0 94500.0 1028250.0 ;
      RECT  90900.0 1029450.0 92100.0 1028250.0 ;
      RECT  95700.0 1020150.0 96900.0 1018950.0 ;
      RECT  95700.0 1030050.0 96900.0 1028850.0 ;
      RECT  93300.0 1027350.0 92100.0 1026150.0 ;
      RECT  90900.0 1025400.0 89700.0 1024200.0 ;
      RECT  88500.0 1023450.0 87300.0 1022250.0 ;
      RECT  88500.0 1020750.0 89700.0 1019550.0 ;
      RECT  93300.0 1020750.0 94500.0 1019550.0 ;
      RECT  93300.0 1029450.0 94500.0 1028250.0 ;
      RECT  93300.0 1023450.0 94500.0 1022250.0 ;
      RECT  87300.0 1023450.0 88500.0 1022250.0 ;
      RECT  89700.0 1025400.0 90900.0 1024200.0 ;
      RECT  92100.0 1027350.0 93300.0 1026150.0 ;
      RECT  93300.0 1023450.0 94500.0 1022250.0 ;
      RECT  84300.0 1018050.0 99900.0 1017150.0 ;
      RECT  84300.0 1031850.0 99900.0 1030950.0 ;
      RECT  86100.0 1033350.0 87300.0 1030950.0 ;
      RECT  86100.0 1042050.0 87300.0 1045650.0 ;
      RECT  90900.0 1042050.0 92100.0 1045650.0 ;
      RECT  95700.0 1043250.0 96900.0 1045200.0 ;
      RECT  95700.0 1031400.0 96900.0 1033350.0 ;
      RECT  86100.0 1042050.0 87300.0 1043250.0 ;
      RECT  88500.0 1042050.0 89700.0 1043250.0 ;
      RECT  88500.0 1042050.0 89700.0 1043250.0 ;
      RECT  86100.0 1042050.0 87300.0 1043250.0 ;
      RECT  88500.0 1042050.0 89700.0 1043250.0 ;
      RECT  90900.0 1042050.0 92100.0 1043250.0 ;
      RECT  90900.0 1042050.0 92100.0 1043250.0 ;
      RECT  88500.0 1042050.0 89700.0 1043250.0 ;
      RECT  90900.0 1042050.0 92100.0 1043250.0 ;
      RECT  93300.0 1042050.0 94500.0 1043250.0 ;
      RECT  93300.0 1042050.0 94500.0 1043250.0 ;
      RECT  90900.0 1042050.0 92100.0 1043250.0 ;
      RECT  86100.0 1033350.0 87300.0 1034550.0 ;
      RECT  88500.0 1033350.0 89700.0 1034550.0 ;
      RECT  88500.0 1033350.0 89700.0 1034550.0 ;
      RECT  86100.0 1033350.0 87300.0 1034550.0 ;
      RECT  88500.0 1033350.0 89700.0 1034550.0 ;
      RECT  90900.0 1033350.0 92100.0 1034550.0 ;
      RECT  90900.0 1033350.0 92100.0 1034550.0 ;
      RECT  88500.0 1033350.0 89700.0 1034550.0 ;
      RECT  90900.0 1033350.0 92100.0 1034550.0 ;
      RECT  93300.0 1033350.0 94500.0 1034550.0 ;
      RECT  93300.0 1033350.0 94500.0 1034550.0 ;
      RECT  90900.0 1033350.0 92100.0 1034550.0 ;
      RECT  95700.0 1042650.0 96900.0 1043850.0 ;
      RECT  95700.0 1032750.0 96900.0 1033950.0 ;
      RECT  93300.0 1035450.0 92100.0 1036650.0 ;
      RECT  90900.0 1037400.0 89700.0 1038600.0 ;
      RECT  88500.0 1039350.0 87300.0 1040550.0 ;
      RECT  88500.0 1042050.0 89700.0 1043250.0 ;
      RECT  93300.0 1042050.0 94500.0 1043250.0 ;
      RECT  93300.0 1033350.0 94500.0 1034550.0 ;
      RECT  93300.0 1039350.0 94500.0 1040550.0 ;
      RECT  87300.0 1039350.0 88500.0 1040550.0 ;
      RECT  89700.0 1037400.0 90900.0 1038600.0 ;
      RECT  92100.0 1035450.0 93300.0 1036650.0 ;
      RECT  93300.0 1039350.0 94500.0 1040550.0 ;
      RECT  84300.0 1044750.0 99900.0 1045650.0 ;
      RECT  84300.0 1030950.0 99900.0 1031850.0 ;
      RECT  86100.0 1057050.0 87300.0 1059450.0 ;
      RECT  86100.0 1048350.0 87300.0 1044750.0 ;
      RECT  90900.0 1048350.0 92100.0 1044750.0 ;
      RECT  95700.0 1047150.0 96900.0 1045200.0 ;
      RECT  95700.0 1059000.0 96900.0 1057050.0 ;
      RECT  86100.0 1048350.0 87300.0 1047150.0 ;
      RECT  88500.0 1048350.0 89700.0 1047150.0 ;
      RECT  88500.0 1048350.0 89700.0 1047150.0 ;
      RECT  86100.0 1048350.0 87300.0 1047150.0 ;
      RECT  88500.0 1048350.0 89700.0 1047150.0 ;
      RECT  90900.0 1048350.0 92100.0 1047150.0 ;
      RECT  90900.0 1048350.0 92100.0 1047150.0 ;
      RECT  88500.0 1048350.0 89700.0 1047150.0 ;
      RECT  90900.0 1048350.0 92100.0 1047150.0 ;
      RECT  93300.0 1048350.0 94500.0 1047150.0 ;
      RECT  93300.0 1048350.0 94500.0 1047150.0 ;
      RECT  90900.0 1048350.0 92100.0 1047150.0 ;
      RECT  86100.0 1057050.0 87300.0 1055850.0 ;
      RECT  88500.0 1057050.0 89700.0 1055850.0 ;
      RECT  88500.0 1057050.0 89700.0 1055850.0 ;
      RECT  86100.0 1057050.0 87300.0 1055850.0 ;
      RECT  88500.0 1057050.0 89700.0 1055850.0 ;
      RECT  90900.0 1057050.0 92100.0 1055850.0 ;
      RECT  90900.0 1057050.0 92100.0 1055850.0 ;
      RECT  88500.0 1057050.0 89700.0 1055850.0 ;
      RECT  90900.0 1057050.0 92100.0 1055850.0 ;
      RECT  93300.0 1057050.0 94500.0 1055850.0 ;
      RECT  93300.0 1057050.0 94500.0 1055850.0 ;
      RECT  90900.0 1057050.0 92100.0 1055850.0 ;
      RECT  95700.0 1047750.0 96900.0 1046550.0 ;
      RECT  95700.0 1057650.0 96900.0 1056450.0 ;
      RECT  93300.0 1054950.0 92100.0 1053750.0 ;
      RECT  90900.0 1053000.0 89700.0 1051800.0 ;
      RECT  88500.0 1051050.0 87300.0 1049850.0 ;
      RECT  88500.0 1048350.0 89700.0 1047150.0 ;
      RECT  93300.0 1048350.0 94500.0 1047150.0 ;
      RECT  93300.0 1057050.0 94500.0 1055850.0 ;
      RECT  93300.0 1051050.0 94500.0 1049850.0 ;
      RECT  87300.0 1051050.0 88500.0 1049850.0 ;
      RECT  89700.0 1053000.0 90900.0 1051800.0 ;
      RECT  92100.0 1054950.0 93300.0 1053750.0 ;
      RECT  93300.0 1051050.0 94500.0 1049850.0 ;
      RECT  84300.0 1045650.0 99900.0 1044750.0 ;
      RECT  84300.0 1059450.0 99900.0 1058550.0 ;
      RECT  86100.0 1060950.0 87300.0 1058550.0 ;
      RECT  86100.0 1069650.0 87300.0 1073250.0 ;
      RECT  90900.0 1069650.0 92100.0 1073250.0 ;
      RECT  95700.0 1070850.0 96900.0 1072800.0 ;
      RECT  95700.0 1059000.0 96900.0 1060950.0 ;
      RECT  86100.0 1069650.0 87300.0 1070850.0 ;
      RECT  88500.0 1069650.0 89700.0 1070850.0 ;
      RECT  88500.0 1069650.0 89700.0 1070850.0 ;
      RECT  86100.0 1069650.0 87300.0 1070850.0 ;
      RECT  88500.0 1069650.0 89700.0 1070850.0 ;
      RECT  90900.0 1069650.0 92100.0 1070850.0 ;
      RECT  90900.0 1069650.0 92100.0 1070850.0 ;
      RECT  88500.0 1069650.0 89700.0 1070850.0 ;
      RECT  90900.0 1069650.0 92100.0 1070850.0 ;
      RECT  93300.0 1069650.0 94500.0 1070850.0 ;
      RECT  93300.0 1069650.0 94500.0 1070850.0 ;
      RECT  90900.0 1069650.0 92100.0 1070850.0 ;
      RECT  86100.0 1060950.0 87300.0 1062150.0 ;
      RECT  88500.0 1060950.0 89700.0 1062150.0 ;
      RECT  88500.0 1060950.0 89700.0 1062150.0 ;
      RECT  86100.0 1060950.0 87300.0 1062150.0 ;
      RECT  88500.0 1060950.0 89700.0 1062150.0 ;
      RECT  90900.0 1060950.0 92100.0 1062150.0 ;
      RECT  90900.0 1060950.0 92100.0 1062150.0 ;
      RECT  88500.0 1060950.0 89700.0 1062150.0 ;
      RECT  90900.0 1060950.0 92100.0 1062150.0 ;
      RECT  93300.0 1060950.0 94500.0 1062150.0 ;
      RECT  93300.0 1060950.0 94500.0 1062150.0 ;
      RECT  90900.0 1060950.0 92100.0 1062150.0 ;
      RECT  95700.0 1070250.0 96900.0 1071450.0 ;
      RECT  95700.0 1060350.0 96900.0 1061550.0 ;
      RECT  93300.0 1063050.0 92100.0 1064250.0 ;
      RECT  90900.0 1065000.0 89700.0 1066200.0 ;
      RECT  88500.0 1066950.0 87300.0 1068150.0 ;
      RECT  88500.0 1069650.0 89700.0 1070850.0 ;
      RECT  93300.0 1069650.0 94500.0 1070850.0 ;
      RECT  93300.0 1060950.0 94500.0 1062150.0 ;
      RECT  93300.0 1066950.0 94500.0 1068150.0 ;
      RECT  87300.0 1066950.0 88500.0 1068150.0 ;
      RECT  89700.0 1065000.0 90900.0 1066200.0 ;
      RECT  92100.0 1063050.0 93300.0 1064250.0 ;
      RECT  93300.0 1066950.0 94500.0 1068150.0 ;
      RECT  84300.0 1072350.0 99900.0 1073250.0 ;
      RECT  84300.0 1058550.0 99900.0 1059450.0 ;
      RECT  86100.0 1084650.0 87300.0 1087050.0 ;
      RECT  86100.0 1075950.0 87300.0 1072350.0 ;
      RECT  90900.0 1075950.0 92100.0 1072350.0 ;
      RECT  95700.0 1074750.0 96900.0 1072800.0 ;
      RECT  95700.0 1086600.0 96900.0 1084650.0 ;
      RECT  86100.0 1075950.0 87300.0 1074750.0 ;
      RECT  88500.0 1075950.0 89700.0 1074750.0 ;
      RECT  88500.0 1075950.0 89700.0 1074750.0 ;
      RECT  86100.0 1075950.0 87300.0 1074750.0 ;
      RECT  88500.0 1075950.0 89700.0 1074750.0 ;
      RECT  90900.0 1075950.0 92100.0 1074750.0 ;
      RECT  90900.0 1075950.0 92100.0 1074750.0 ;
      RECT  88500.0 1075950.0 89700.0 1074750.0 ;
      RECT  90900.0 1075950.0 92100.0 1074750.0 ;
      RECT  93300.0 1075950.0 94500.0 1074750.0 ;
      RECT  93300.0 1075950.0 94500.0 1074750.0 ;
      RECT  90900.0 1075950.0 92100.0 1074750.0 ;
      RECT  86100.0 1084650.0 87300.0 1083450.0 ;
      RECT  88500.0 1084650.0 89700.0 1083450.0 ;
      RECT  88500.0 1084650.0 89700.0 1083450.0 ;
      RECT  86100.0 1084650.0 87300.0 1083450.0 ;
      RECT  88500.0 1084650.0 89700.0 1083450.0 ;
      RECT  90900.0 1084650.0 92100.0 1083450.0 ;
      RECT  90900.0 1084650.0 92100.0 1083450.0 ;
      RECT  88500.0 1084650.0 89700.0 1083450.0 ;
      RECT  90900.0 1084650.0 92100.0 1083450.0 ;
      RECT  93300.0 1084650.0 94500.0 1083450.0 ;
      RECT  93300.0 1084650.0 94500.0 1083450.0 ;
      RECT  90900.0 1084650.0 92100.0 1083450.0 ;
      RECT  95700.0 1075350.0 96900.0 1074150.0 ;
      RECT  95700.0 1085250.0 96900.0 1084050.0 ;
      RECT  93300.0 1082550.0 92100.0 1081350.0 ;
      RECT  90900.0 1080600.0 89700.0 1079400.0 ;
      RECT  88500.0 1078650.0 87300.0 1077450.0 ;
      RECT  88500.0 1075950.0 89700.0 1074750.0 ;
      RECT  93300.0 1075950.0 94500.0 1074750.0 ;
      RECT  93300.0 1084650.0 94500.0 1083450.0 ;
      RECT  93300.0 1078650.0 94500.0 1077450.0 ;
      RECT  87300.0 1078650.0 88500.0 1077450.0 ;
      RECT  89700.0 1080600.0 90900.0 1079400.0 ;
      RECT  92100.0 1082550.0 93300.0 1081350.0 ;
      RECT  93300.0 1078650.0 94500.0 1077450.0 ;
      RECT  84300.0 1073250.0 99900.0 1072350.0 ;
      RECT  84300.0 1087050.0 99900.0 1086150.0 ;
      RECT  86100.0 1088550.0 87300.0 1086150.0 ;
      RECT  86100.0 1097250.0 87300.0 1100850.0 ;
      RECT  90900.0 1097250.0 92100.0 1100850.0 ;
      RECT  95700.0 1098450.0 96900.0 1100400.0 ;
      RECT  95700.0 1086600.0 96900.0 1088550.0 ;
      RECT  86100.0 1097250.0 87300.0 1098450.0 ;
      RECT  88500.0 1097250.0 89700.0 1098450.0 ;
      RECT  88500.0 1097250.0 89700.0 1098450.0 ;
      RECT  86100.0 1097250.0 87300.0 1098450.0 ;
      RECT  88500.0 1097250.0 89700.0 1098450.0 ;
      RECT  90900.0 1097250.0 92100.0 1098450.0 ;
      RECT  90900.0 1097250.0 92100.0 1098450.0 ;
      RECT  88500.0 1097250.0 89700.0 1098450.0 ;
      RECT  90900.0 1097250.0 92100.0 1098450.0 ;
      RECT  93300.0 1097250.0 94500.0 1098450.0 ;
      RECT  93300.0 1097250.0 94500.0 1098450.0 ;
      RECT  90900.0 1097250.0 92100.0 1098450.0 ;
      RECT  86100.0 1088550.0 87300.0 1089750.0 ;
      RECT  88500.0 1088550.0 89700.0 1089750.0 ;
      RECT  88500.0 1088550.0 89700.0 1089750.0 ;
      RECT  86100.0 1088550.0 87300.0 1089750.0 ;
      RECT  88500.0 1088550.0 89700.0 1089750.0 ;
      RECT  90900.0 1088550.0 92100.0 1089750.0 ;
      RECT  90900.0 1088550.0 92100.0 1089750.0 ;
      RECT  88500.0 1088550.0 89700.0 1089750.0 ;
      RECT  90900.0 1088550.0 92100.0 1089750.0 ;
      RECT  93300.0 1088550.0 94500.0 1089750.0 ;
      RECT  93300.0 1088550.0 94500.0 1089750.0 ;
      RECT  90900.0 1088550.0 92100.0 1089750.0 ;
      RECT  95700.0 1097850.0 96900.0 1099050.0 ;
      RECT  95700.0 1087950.0 96900.0 1089150.0 ;
      RECT  93300.0 1090650.0 92100.0 1091850.0 ;
      RECT  90900.0 1092600.0 89700.0 1093800.0 ;
      RECT  88500.0 1094550.0 87300.0 1095750.0 ;
      RECT  88500.0 1097250.0 89700.0 1098450.0 ;
      RECT  93300.0 1097250.0 94500.0 1098450.0 ;
      RECT  93300.0 1088550.0 94500.0 1089750.0 ;
      RECT  93300.0 1094550.0 94500.0 1095750.0 ;
      RECT  87300.0 1094550.0 88500.0 1095750.0 ;
      RECT  89700.0 1092600.0 90900.0 1093800.0 ;
      RECT  92100.0 1090650.0 93300.0 1091850.0 ;
      RECT  93300.0 1094550.0 94500.0 1095750.0 ;
      RECT  84300.0 1099950.0 99900.0 1100850.0 ;
      RECT  84300.0 1086150.0 99900.0 1087050.0 ;
      RECT  86100.0 1112250.0 87300.0 1114650.0 ;
      RECT  86100.0 1103550.0 87300.0 1099950.0 ;
      RECT  90900.0 1103550.0 92100.0 1099950.0 ;
      RECT  95700.0 1102350.0 96900.0 1100400.0 ;
      RECT  95700.0 1114200.0 96900.0 1112250.0 ;
      RECT  86100.0 1103550.0 87300.0 1102350.0 ;
      RECT  88500.0 1103550.0 89700.0 1102350.0 ;
      RECT  88500.0 1103550.0 89700.0 1102350.0 ;
      RECT  86100.0 1103550.0 87300.0 1102350.0 ;
      RECT  88500.0 1103550.0 89700.0 1102350.0 ;
      RECT  90900.0 1103550.0 92100.0 1102350.0 ;
      RECT  90900.0 1103550.0 92100.0 1102350.0 ;
      RECT  88500.0 1103550.0 89700.0 1102350.0 ;
      RECT  90900.0 1103550.0 92100.0 1102350.0 ;
      RECT  93300.0 1103550.0 94500.0 1102350.0 ;
      RECT  93300.0 1103550.0 94500.0 1102350.0 ;
      RECT  90900.0 1103550.0 92100.0 1102350.0 ;
      RECT  86100.0 1112250.0 87300.0 1111050.0 ;
      RECT  88500.0 1112250.0 89700.0 1111050.0 ;
      RECT  88500.0 1112250.0 89700.0 1111050.0 ;
      RECT  86100.0 1112250.0 87300.0 1111050.0 ;
      RECT  88500.0 1112250.0 89700.0 1111050.0 ;
      RECT  90900.0 1112250.0 92100.0 1111050.0 ;
      RECT  90900.0 1112250.0 92100.0 1111050.0 ;
      RECT  88500.0 1112250.0 89700.0 1111050.0 ;
      RECT  90900.0 1112250.0 92100.0 1111050.0 ;
      RECT  93300.0 1112250.0 94500.0 1111050.0 ;
      RECT  93300.0 1112250.0 94500.0 1111050.0 ;
      RECT  90900.0 1112250.0 92100.0 1111050.0 ;
      RECT  95700.0 1102950.0 96900.0 1101750.0 ;
      RECT  95700.0 1112850.0 96900.0 1111650.0 ;
      RECT  93300.0 1110150.0 92100.0 1108950.0 ;
      RECT  90900.0 1108200.0 89700.0 1107000.0 ;
      RECT  88500.0 1106250.0 87300.0 1105050.0 ;
      RECT  88500.0 1103550.0 89700.0 1102350.0 ;
      RECT  93300.0 1103550.0 94500.0 1102350.0 ;
      RECT  93300.0 1112250.0 94500.0 1111050.0 ;
      RECT  93300.0 1106250.0 94500.0 1105050.0 ;
      RECT  87300.0 1106250.0 88500.0 1105050.0 ;
      RECT  89700.0 1108200.0 90900.0 1107000.0 ;
      RECT  92100.0 1110150.0 93300.0 1108950.0 ;
      RECT  93300.0 1106250.0 94500.0 1105050.0 ;
      RECT  84300.0 1100850.0 99900.0 1099950.0 ;
      RECT  84300.0 1114650.0 99900.0 1113750.0 ;
      RECT  86100.0 1116150.0 87300.0 1113750.0 ;
      RECT  86100.0 1124850.0 87300.0 1128450.0 ;
      RECT  90900.0 1124850.0 92100.0 1128450.0 ;
      RECT  95700.0 1126050.0 96900.0 1128000.0 ;
      RECT  95700.0 1114200.0 96900.0 1116150.0 ;
      RECT  86100.0 1124850.0 87300.0 1126050.0 ;
      RECT  88500.0 1124850.0 89700.0 1126050.0 ;
      RECT  88500.0 1124850.0 89700.0 1126050.0 ;
      RECT  86100.0 1124850.0 87300.0 1126050.0 ;
      RECT  88500.0 1124850.0 89700.0 1126050.0 ;
      RECT  90900.0 1124850.0 92100.0 1126050.0 ;
      RECT  90900.0 1124850.0 92100.0 1126050.0 ;
      RECT  88500.0 1124850.0 89700.0 1126050.0 ;
      RECT  90900.0 1124850.0 92100.0 1126050.0 ;
      RECT  93300.0 1124850.0 94500.0 1126050.0 ;
      RECT  93300.0 1124850.0 94500.0 1126050.0 ;
      RECT  90900.0 1124850.0 92100.0 1126050.0 ;
      RECT  86100.0 1116150.0 87300.0 1117350.0 ;
      RECT  88500.0 1116150.0 89700.0 1117350.0 ;
      RECT  88500.0 1116150.0 89700.0 1117350.0 ;
      RECT  86100.0 1116150.0 87300.0 1117350.0 ;
      RECT  88500.0 1116150.0 89700.0 1117350.0 ;
      RECT  90900.0 1116150.0 92100.0 1117350.0 ;
      RECT  90900.0 1116150.0 92100.0 1117350.0 ;
      RECT  88500.0 1116150.0 89700.0 1117350.0 ;
      RECT  90900.0 1116150.0 92100.0 1117350.0 ;
      RECT  93300.0 1116150.0 94500.0 1117350.0 ;
      RECT  93300.0 1116150.0 94500.0 1117350.0 ;
      RECT  90900.0 1116150.0 92100.0 1117350.0 ;
      RECT  95700.0 1125450.0 96900.0 1126650.0 ;
      RECT  95700.0 1115550.0 96900.0 1116750.0 ;
      RECT  93300.0 1118250.0 92100.0 1119450.0 ;
      RECT  90900.0 1120200.0 89700.0 1121400.0 ;
      RECT  88500.0 1122150.0 87300.0 1123350.0 ;
      RECT  88500.0 1124850.0 89700.0 1126050.0 ;
      RECT  93300.0 1124850.0 94500.0 1126050.0 ;
      RECT  93300.0 1116150.0 94500.0 1117350.0 ;
      RECT  93300.0 1122150.0 94500.0 1123350.0 ;
      RECT  87300.0 1122150.0 88500.0 1123350.0 ;
      RECT  89700.0 1120200.0 90900.0 1121400.0 ;
      RECT  92100.0 1118250.0 93300.0 1119450.0 ;
      RECT  93300.0 1122150.0 94500.0 1123350.0 ;
      RECT  84300.0 1127550.0 99900.0 1128450.0 ;
      RECT  84300.0 1113750.0 99900.0 1114650.0 ;
      RECT  86100.0 1139850.0 87300.0 1142250.0 ;
      RECT  86100.0 1131150.0 87300.0 1127550.0 ;
      RECT  90900.0 1131150.0 92100.0 1127550.0 ;
      RECT  95700.0 1129950.0 96900.0 1128000.0 ;
      RECT  95700.0 1141800.0 96900.0 1139850.0 ;
      RECT  86100.0 1131150.0 87300.0 1129950.0 ;
      RECT  88500.0 1131150.0 89700.0 1129950.0 ;
      RECT  88500.0 1131150.0 89700.0 1129950.0 ;
      RECT  86100.0 1131150.0 87300.0 1129950.0 ;
      RECT  88500.0 1131150.0 89700.0 1129950.0 ;
      RECT  90900.0 1131150.0 92100.0 1129950.0 ;
      RECT  90900.0 1131150.0 92100.0 1129950.0 ;
      RECT  88500.0 1131150.0 89700.0 1129950.0 ;
      RECT  90900.0 1131150.0 92100.0 1129950.0 ;
      RECT  93300.0 1131150.0 94500.0 1129950.0 ;
      RECT  93300.0 1131150.0 94500.0 1129950.0 ;
      RECT  90900.0 1131150.0 92100.0 1129950.0 ;
      RECT  86100.0 1139850.0 87300.0 1138650.0 ;
      RECT  88500.0 1139850.0 89700.0 1138650.0 ;
      RECT  88500.0 1139850.0 89700.0 1138650.0 ;
      RECT  86100.0 1139850.0 87300.0 1138650.0 ;
      RECT  88500.0 1139850.0 89700.0 1138650.0 ;
      RECT  90900.0 1139850.0 92100.0 1138650.0 ;
      RECT  90900.0 1139850.0 92100.0 1138650.0 ;
      RECT  88500.0 1139850.0 89700.0 1138650.0 ;
      RECT  90900.0 1139850.0 92100.0 1138650.0 ;
      RECT  93300.0 1139850.0 94500.0 1138650.0 ;
      RECT  93300.0 1139850.0 94500.0 1138650.0 ;
      RECT  90900.0 1139850.0 92100.0 1138650.0 ;
      RECT  95700.0 1130550.0 96900.0 1129350.0 ;
      RECT  95700.0 1140450.0 96900.0 1139250.0 ;
      RECT  93300.0 1137750.0 92100.0 1136550.0 ;
      RECT  90900.0 1135800.0 89700.0 1134600.0 ;
      RECT  88500.0 1133850.0 87300.0 1132650.0 ;
      RECT  88500.0 1131150.0 89700.0 1129950.0 ;
      RECT  93300.0 1131150.0 94500.0 1129950.0 ;
      RECT  93300.0 1139850.0 94500.0 1138650.0 ;
      RECT  93300.0 1133850.0 94500.0 1132650.0 ;
      RECT  87300.0 1133850.0 88500.0 1132650.0 ;
      RECT  89700.0 1135800.0 90900.0 1134600.0 ;
      RECT  92100.0 1137750.0 93300.0 1136550.0 ;
      RECT  93300.0 1133850.0 94500.0 1132650.0 ;
      RECT  84300.0 1128450.0 99900.0 1127550.0 ;
      RECT  84300.0 1142250.0 99900.0 1141350.0 ;
      RECT  86100.0 1143750.0 87300.0 1141350.0 ;
      RECT  86100.0 1152450.0 87300.0 1156050.0 ;
      RECT  90900.0 1152450.0 92100.0 1156050.0 ;
      RECT  95700.0 1153650.0 96900.0 1155600.0 ;
      RECT  95700.0 1141800.0 96900.0 1143750.0 ;
      RECT  86100.0 1152450.0 87300.0 1153650.0 ;
      RECT  88500.0 1152450.0 89700.0 1153650.0 ;
      RECT  88500.0 1152450.0 89700.0 1153650.0 ;
      RECT  86100.0 1152450.0 87300.0 1153650.0 ;
      RECT  88500.0 1152450.0 89700.0 1153650.0 ;
      RECT  90900.0 1152450.0 92100.0 1153650.0 ;
      RECT  90900.0 1152450.0 92100.0 1153650.0 ;
      RECT  88500.0 1152450.0 89700.0 1153650.0 ;
      RECT  90900.0 1152450.0 92100.0 1153650.0 ;
      RECT  93300.0 1152450.0 94500.0 1153650.0 ;
      RECT  93300.0 1152450.0 94500.0 1153650.0 ;
      RECT  90900.0 1152450.0 92100.0 1153650.0 ;
      RECT  86100.0 1143750.0 87300.0 1144950.0 ;
      RECT  88500.0 1143750.0 89700.0 1144950.0 ;
      RECT  88500.0 1143750.0 89700.0 1144950.0 ;
      RECT  86100.0 1143750.0 87300.0 1144950.0 ;
      RECT  88500.0 1143750.0 89700.0 1144950.0 ;
      RECT  90900.0 1143750.0 92100.0 1144950.0 ;
      RECT  90900.0 1143750.0 92100.0 1144950.0 ;
      RECT  88500.0 1143750.0 89700.0 1144950.0 ;
      RECT  90900.0 1143750.0 92100.0 1144950.0 ;
      RECT  93300.0 1143750.0 94500.0 1144950.0 ;
      RECT  93300.0 1143750.0 94500.0 1144950.0 ;
      RECT  90900.0 1143750.0 92100.0 1144950.0 ;
      RECT  95700.0 1153050.0 96900.0 1154250.0 ;
      RECT  95700.0 1143150.0 96900.0 1144350.0 ;
      RECT  93300.0 1145850.0 92100.0 1147050.0 ;
      RECT  90900.0 1147800.0 89700.0 1149000.0 ;
      RECT  88500.0 1149750.0 87300.0 1150950.0 ;
      RECT  88500.0 1152450.0 89700.0 1153650.0 ;
      RECT  93300.0 1152450.0 94500.0 1153650.0 ;
      RECT  93300.0 1143750.0 94500.0 1144950.0 ;
      RECT  93300.0 1149750.0 94500.0 1150950.0 ;
      RECT  87300.0 1149750.0 88500.0 1150950.0 ;
      RECT  89700.0 1147800.0 90900.0 1149000.0 ;
      RECT  92100.0 1145850.0 93300.0 1147050.0 ;
      RECT  93300.0 1149750.0 94500.0 1150950.0 ;
      RECT  84300.0 1155150.0 99900.0 1156050.0 ;
      RECT  84300.0 1141350.0 99900.0 1142250.0 ;
      RECT  86100.0 1167450.0 87300.0 1169850.0 ;
      RECT  86100.0 1158750.0 87300.0 1155150.0 ;
      RECT  90900.0 1158750.0 92100.0 1155150.0 ;
      RECT  95700.0 1157550.0 96900.0 1155600.0 ;
      RECT  95700.0 1169400.0 96900.0 1167450.0 ;
      RECT  86100.0 1158750.0 87300.0 1157550.0 ;
      RECT  88500.0 1158750.0 89700.0 1157550.0 ;
      RECT  88500.0 1158750.0 89700.0 1157550.0 ;
      RECT  86100.0 1158750.0 87300.0 1157550.0 ;
      RECT  88500.0 1158750.0 89700.0 1157550.0 ;
      RECT  90900.0 1158750.0 92100.0 1157550.0 ;
      RECT  90900.0 1158750.0 92100.0 1157550.0 ;
      RECT  88500.0 1158750.0 89700.0 1157550.0 ;
      RECT  90900.0 1158750.0 92100.0 1157550.0 ;
      RECT  93300.0 1158750.0 94500.0 1157550.0 ;
      RECT  93300.0 1158750.0 94500.0 1157550.0 ;
      RECT  90900.0 1158750.0 92100.0 1157550.0 ;
      RECT  86100.0 1167450.0 87300.0 1166250.0 ;
      RECT  88500.0 1167450.0 89700.0 1166250.0 ;
      RECT  88500.0 1167450.0 89700.0 1166250.0 ;
      RECT  86100.0 1167450.0 87300.0 1166250.0 ;
      RECT  88500.0 1167450.0 89700.0 1166250.0 ;
      RECT  90900.0 1167450.0 92100.0 1166250.0 ;
      RECT  90900.0 1167450.0 92100.0 1166250.0 ;
      RECT  88500.0 1167450.0 89700.0 1166250.0 ;
      RECT  90900.0 1167450.0 92100.0 1166250.0 ;
      RECT  93300.0 1167450.0 94500.0 1166250.0 ;
      RECT  93300.0 1167450.0 94500.0 1166250.0 ;
      RECT  90900.0 1167450.0 92100.0 1166250.0 ;
      RECT  95700.0 1158150.0 96900.0 1156950.0 ;
      RECT  95700.0 1168050.0 96900.0 1166850.0 ;
      RECT  93300.0 1165350.0 92100.0 1164150.0 ;
      RECT  90900.0 1163400.0 89700.0 1162200.0 ;
      RECT  88500.0 1161450.0 87300.0 1160250.0 ;
      RECT  88500.0 1158750.0 89700.0 1157550.0 ;
      RECT  93300.0 1158750.0 94500.0 1157550.0 ;
      RECT  93300.0 1167450.0 94500.0 1166250.0 ;
      RECT  93300.0 1161450.0 94500.0 1160250.0 ;
      RECT  87300.0 1161450.0 88500.0 1160250.0 ;
      RECT  89700.0 1163400.0 90900.0 1162200.0 ;
      RECT  92100.0 1165350.0 93300.0 1164150.0 ;
      RECT  93300.0 1161450.0 94500.0 1160250.0 ;
      RECT  84300.0 1156050.0 99900.0 1155150.0 ;
      RECT  84300.0 1169850.0 99900.0 1168950.0 ;
      RECT  86100.0 1171350.0 87300.0 1168950.0 ;
      RECT  86100.0 1180050.0 87300.0 1183650.0 ;
      RECT  90900.0 1180050.0 92100.0 1183650.0 ;
      RECT  95700.0 1181250.0 96900.0 1183200.0 ;
      RECT  95700.0 1169400.0 96900.0 1171350.0 ;
      RECT  86100.0 1180050.0 87300.0 1181250.0 ;
      RECT  88500.0 1180050.0 89700.0 1181250.0 ;
      RECT  88500.0 1180050.0 89700.0 1181250.0 ;
      RECT  86100.0 1180050.0 87300.0 1181250.0 ;
      RECT  88500.0 1180050.0 89700.0 1181250.0 ;
      RECT  90900.0 1180050.0 92100.0 1181250.0 ;
      RECT  90900.0 1180050.0 92100.0 1181250.0 ;
      RECT  88500.0 1180050.0 89700.0 1181250.0 ;
      RECT  90900.0 1180050.0 92100.0 1181250.0 ;
      RECT  93300.0 1180050.0 94500.0 1181250.0 ;
      RECT  93300.0 1180050.0 94500.0 1181250.0 ;
      RECT  90900.0 1180050.0 92100.0 1181250.0 ;
      RECT  86100.0 1171350.0 87300.0 1172550.0 ;
      RECT  88500.0 1171350.0 89700.0 1172550.0 ;
      RECT  88500.0 1171350.0 89700.0 1172550.0 ;
      RECT  86100.0 1171350.0 87300.0 1172550.0 ;
      RECT  88500.0 1171350.0 89700.0 1172550.0 ;
      RECT  90900.0 1171350.0 92100.0 1172550.0 ;
      RECT  90900.0 1171350.0 92100.0 1172550.0 ;
      RECT  88500.0 1171350.0 89700.0 1172550.0 ;
      RECT  90900.0 1171350.0 92100.0 1172550.0 ;
      RECT  93300.0 1171350.0 94500.0 1172550.0 ;
      RECT  93300.0 1171350.0 94500.0 1172550.0 ;
      RECT  90900.0 1171350.0 92100.0 1172550.0 ;
      RECT  95700.0 1180650.0 96900.0 1181850.0 ;
      RECT  95700.0 1170750.0 96900.0 1171950.0 ;
      RECT  93300.0 1173450.0 92100.0 1174650.0 ;
      RECT  90900.0 1175400.0 89700.0 1176600.0 ;
      RECT  88500.0 1177350.0 87300.0 1178550.0 ;
      RECT  88500.0 1180050.0 89700.0 1181250.0 ;
      RECT  93300.0 1180050.0 94500.0 1181250.0 ;
      RECT  93300.0 1171350.0 94500.0 1172550.0 ;
      RECT  93300.0 1177350.0 94500.0 1178550.0 ;
      RECT  87300.0 1177350.0 88500.0 1178550.0 ;
      RECT  89700.0 1175400.0 90900.0 1176600.0 ;
      RECT  92100.0 1173450.0 93300.0 1174650.0 ;
      RECT  93300.0 1177350.0 94500.0 1178550.0 ;
      RECT  84300.0 1182750.0 99900.0 1183650.0 ;
      RECT  84300.0 1168950.0 99900.0 1169850.0 ;
      RECT  86100.0 1195050.0 87300.0 1197450.0 ;
      RECT  86100.0 1186350.0 87300.0 1182750.0 ;
      RECT  90900.0 1186350.0 92100.0 1182750.0 ;
      RECT  95700.0 1185150.0 96900.0 1183200.0 ;
      RECT  95700.0 1197000.0 96900.0 1195050.0 ;
      RECT  86100.0 1186350.0 87300.0 1185150.0 ;
      RECT  88500.0 1186350.0 89700.0 1185150.0 ;
      RECT  88500.0 1186350.0 89700.0 1185150.0 ;
      RECT  86100.0 1186350.0 87300.0 1185150.0 ;
      RECT  88500.0 1186350.0 89700.0 1185150.0 ;
      RECT  90900.0 1186350.0 92100.0 1185150.0 ;
      RECT  90900.0 1186350.0 92100.0 1185150.0 ;
      RECT  88500.0 1186350.0 89700.0 1185150.0 ;
      RECT  90900.0 1186350.0 92100.0 1185150.0 ;
      RECT  93300.0 1186350.0 94500.0 1185150.0 ;
      RECT  93300.0 1186350.0 94500.0 1185150.0 ;
      RECT  90900.0 1186350.0 92100.0 1185150.0 ;
      RECT  86100.0 1195050.0 87300.0 1193850.0 ;
      RECT  88500.0 1195050.0 89700.0 1193850.0 ;
      RECT  88500.0 1195050.0 89700.0 1193850.0 ;
      RECT  86100.0 1195050.0 87300.0 1193850.0 ;
      RECT  88500.0 1195050.0 89700.0 1193850.0 ;
      RECT  90900.0 1195050.0 92100.0 1193850.0 ;
      RECT  90900.0 1195050.0 92100.0 1193850.0 ;
      RECT  88500.0 1195050.0 89700.0 1193850.0 ;
      RECT  90900.0 1195050.0 92100.0 1193850.0 ;
      RECT  93300.0 1195050.0 94500.0 1193850.0 ;
      RECT  93300.0 1195050.0 94500.0 1193850.0 ;
      RECT  90900.0 1195050.0 92100.0 1193850.0 ;
      RECT  95700.0 1185750.0 96900.0 1184550.0 ;
      RECT  95700.0 1195650.0 96900.0 1194450.0 ;
      RECT  93300.0 1192950.0 92100.0 1191750.0 ;
      RECT  90900.0 1191000.0 89700.0 1189800.0 ;
      RECT  88500.0 1189050.0 87300.0 1187850.0 ;
      RECT  88500.0 1186350.0 89700.0 1185150.0 ;
      RECT  93300.0 1186350.0 94500.0 1185150.0 ;
      RECT  93300.0 1195050.0 94500.0 1193850.0 ;
      RECT  93300.0 1189050.0 94500.0 1187850.0 ;
      RECT  87300.0 1189050.0 88500.0 1187850.0 ;
      RECT  89700.0 1191000.0 90900.0 1189800.0 ;
      RECT  92100.0 1192950.0 93300.0 1191750.0 ;
      RECT  93300.0 1189050.0 94500.0 1187850.0 ;
      RECT  84300.0 1183650.0 99900.0 1182750.0 ;
      RECT  84300.0 1197450.0 99900.0 1196550.0 ;
      RECT  106500.0 325650.0 107700.0 327600.0 ;
      RECT  106500.0 313800.0 107700.0 315750.0 ;
      RECT  101700.0 315150.0 102900.0 313350.0 ;
      RECT  101700.0 324450.0 102900.0 328050.0 ;
      RECT  104400.0 315150.0 105300.0 324450.0 ;
      RECT  101700.0 324450.0 102900.0 325650.0 ;
      RECT  104100.0 324450.0 105300.0 325650.0 ;
      RECT  104100.0 324450.0 105300.0 325650.0 ;
      RECT  101700.0 324450.0 102900.0 325650.0 ;
      RECT  101700.0 315150.0 102900.0 316350.0 ;
      RECT  104100.0 315150.0 105300.0 316350.0 ;
      RECT  104100.0 315150.0 105300.0 316350.0 ;
      RECT  101700.0 315150.0 102900.0 316350.0 ;
      RECT  106500.0 325050.0 107700.0 326250.0 ;
      RECT  106500.0 315150.0 107700.0 316350.0 ;
      RECT  102300.0 319800.0 103500.0 321000.0 ;
      RECT  102300.0 319800.0 103500.0 321000.0 ;
      RECT  104850.0 319950.0 105750.0 320850.0 ;
      RECT  99900.0 327150.0 109500.0 328050.0 ;
      RECT  99900.0 313350.0 109500.0 314250.0 ;
      RECT  106500.0 329550.0 107700.0 327600.0 ;
      RECT  106500.0 341400.0 107700.0 339450.0 ;
      RECT  101700.0 340050.0 102900.0 341850.0 ;
      RECT  101700.0 330750.0 102900.0 327150.0 ;
      RECT  104400.0 340050.0 105300.0 330750.0 ;
      RECT  101700.0 330750.0 102900.0 329550.0 ;
      RECT  104100.0 330750.0 105300.0 329550.0 ;
      RECT  104100.0 330750.0 105300.0 329550.0 ;
      RECT  101700.0 330750.0 102900.0 329550.0 ;
      RECT  101700.0 340050.0 102900.0 338850.0 ;
      RECT  104100.0 340050.0 105300.0 338850.0 ;
      RECT  104100.0 340050.0 105300.0 338850.0 ;
      RECT  101700.0 340050.0 102900.0 338850.0 ;
      RECT  106500.0 330150.0 107700.0 328950.0 ;
      RECT  106500.0 340050.0 107700.0 338850.0 ;
      RECT  102300.0 335400.0 103500.0 334200.0 ;
      RECT  102300.0 335400.0 103500.0 334200.0 ;
      RECT  104850.0 335250.0 105750.0 334350.0 ;
      RECT  99900.0 328050.0 109500.0 327150.0 ;
      RECT  99900.0 341850.0 109500.0 340950.0 ;
      RECT  106500.0 353250.0 107700.0 355200.0 ;
      RECT  106500.0 341400.0 107700.0 343350.0 ;
      RECT  101700.0 342750.0 102900.0 340950.0 ;
      RECT  101700.0 352050.0 102900.0 355650.0 ;
      RECT  104400.0 342750.0 105300.0 352050.0 ;
      RECT  101700.0 352050.0 102900.0 353250.0 ;
      RECT  104100.0 352050.0 105300.0 353250.0 ;
      RECT  104100.0 352050.0 105300.0 353250.0 ;
      RECT  101700.0 352050.0 102900.0 353250.0 ;
      RECT  101700.0 342750.0 102900.0 343950.0 ;
      RECT  104100.0 342750.0 105300.0 343950.0 ;
      RECT  104100.0 342750.0 105300.0 343950.0 ;
      RECT  101700.0 342750.0 102900.0 343950.0 ;
      RECT  106500.0 352650.0 107700.0 353850.0 ;
      RECT  106500.0 342750.0 107700.0 343950.0 ;
      RECT  102300.0 347400.0 103500.0 348600.0 ;
      RECT  102300.0 347400.0 103500.0 348600.0 ;
      RECT  104850.0 347550.0 105750.0 348450.0 ;
      RECT  99900.0 354750.0 109500.0 355650.0 ;
      RECT  99900.0 340950.0 109500.0 341850.0 ;
      RECT  106500.0 357150.0 107700.0 355200.0 ;
      RECT  106500.0 369000.0 107700.0 367050.0 ;
      RECT  101700.0 367650.0 102900.0 369450.0 ;
      RECT  101700.0 358350.0 102900.0 354750.0 ;
      RECT  104400.0 367650.0 105300.0 358350.0 ;
      RECT  101700.0 358350.0 102900.0 357150.0 ;
      RECT  104100.0 358350.0 105300.0 357150.0 ;
      RECT  104100.0 358350.0 105300.0 357150.0 ;
      RECT  101700.0 358350.0 102900.0 357150.0 ;
      RECT  101700.0 367650.0 102900.0 366450.0 ;
      RECT  104100.0 367650.0 105300.0 366450.0 ;
      RECT  104100.0 367650.0 105300.0 366450.0 ;
      RECT  101700.0 367650.0 102900.0 366450.0 ;
      RECT  106500.0 357750.0 107700.0 356550.0 ;
      RECT  106500.0 367650.0 107700.0 366450.0 ;
      RECT  102300.0 363000.0 103500.0 361800.0 ;
      RECT  102300.0 363000.0 103500.0 361800.0 ;
      RECT  104850.0 362850.0 105750.0 361950.0 ;
      RECT  99900.0 355650.0 109500.0 354750.0 ;
      RECT  99900.0 369450.0 109500.0 368550.0 ;
      RECT  106500.0 380850.0 107700.0 382800.0 ;
      RECT  106500.0 369000.0 107700.0 370950.0 ;
      RECT  101700.0 370350.0 102900.0 368550.0 ;
      RECT  101700.0 379650.0 102900.0 383250.0 ;
      RECT  104400.0 370350.0 105300.0 379650.0 ;
      RECT  101700.0 379650.0 102900.0 380850.0 ;
      RECT  104100.0 379650.0 105300.0 380850.0 ;
      RECT  104100.0 379650.0 105300.0 380850.0 ;
      RECT  101700.0 379650.0 102900.0 380850.0 ;
      RECT  101700.0 370350.0 102900.0 371550.0 ;
      RECT  104100.0 370350.0 105300.0 371550.0 ;
      RECT  104100.0 370350.0 105300.0 371550.0 ;
      RECT  101700.0 370350.0 102900.0 371550.0 ;
      RECT  106500.0 380250.0 107700.0 381450.0 ;
      RECT  106500.0 370350.0 107700.0 371550.0 ;
      RECT  102300.0 375000.0 103500.0 376200.0 ;
      RECT  102300.0 375000.0 103500.0 376200.0 ;
      RECT  104850.0 375150.0 105750.0 376050.0 ;
      RECT  99900.0 382350.0 109500.0 383250.0 ;
      RECT  99900.0 368550.0 109500.0 369450.0 ;
      RECT  106500.0 384750.0 107700.0 382800.0 ;
      RECT  106500.0 396600.0 107700.0 394650.0 ;
      RECT  101700.0 395250.0 102900.0 397050.0 ;
      RECT  101700.0 385950.0 102900.0 382350.0 ;
      RECT  104400.0 395250.0 105300.0 385950.0 ;
      RECT  101700.0 385950.0 102900.0 384750.0 ;
      RECT  104100.0 385950.0 105300.0 384750.0 ;
      RECT  104100.0 385950.0 105300.0 384750.0 ;
      RECT  101700.0 385950.0 102900.0 384750.0 ;
      RECT  101700.0 395250.0 102900.0 394050.0 ;
      RECT  104100.0 395250.0 105300.0 394050.0 ;
      RECT  104100.0 395250.0 105300.0 394050.0 ;
      RECT  101700.0 395250.0 102900.0 394050.0 ;
      RECT  106500.0 385350.0 107700.0 384150.0 ;
      RECT  106500.0 395250.0 107700.0 394050.0 ;
      RECT  102300.0 390600.0 103500.0 389400.0 ;
      RECT  102300.0 390600.0 103500.0 389400.0 ;
      RECT  104850.0 390450.0 105750.0 389550.0 ;
      RECT  99900.0 383250.0 109500.0 382350.0 ;
      RECT  99900.0 397050.0 109500.0 396150.0 ;
      RECT  106500.0 408450.0 107700.0 410400.0 ;
      RECT  106500.0 396600.0 107700.0 398550.0 ;
      RECT  101700.0 397950.0 102900.0 396150.0 ;
      RECT  101700.0 407250.0 102900.0 410850.0 ;
      RECT  104400.0 397950.0 105300.0 407250.0 ;
      RECT  101700.0 407250.0 102900.0 408450.0 ;
      RECT  104100.0 407250.0 105300.0 408450.0 ;
      RECT  104100.0 407250.0 105300.0 408450.0 ;
      RECT  101700.0 407250.0 102900.0 408450.0 ;
      RECT  101700.0 397950.0 102900.0 399150.0 ;
      RECT  104100.0 397950.0 105300.0 399150.0 ;
      RECT  104100.0 397950.0 105300.0 399150.0 ;
      RECT  101700.0 397950.0 102900.0 399150.0 ;
      RECT  106500.0 407850.0 107700.0 409050.0 ;
      RECT  106500.0 397950.0 107700.0 399150.0 ;
      RECT  102300.0 402600.0 103500.0 403800.0 ;
      RECT  102300.0 402600.0 103500.0 403800.0 ;
      RECT  104850.0 402750.0 105750.0 403650.0 ;
      RECT  99900.0 409950.0 109500.0 410850.0 ;
      RECT  99900.0 396150.0 109500.0 397050.0 ;
      RECT  106500.0 412350.0 107700.0 410400.0 ;
      RECT  106500.0 424200.0 107700.0 422250.0 ;
      RECT  101700.0 422850.0 102900.0 424650.0 ;
      RECT  101700.0 413550.0 102900.0 409950.0 ;
      RECT  104400.0 422850.0 105300.0 413550.0 ;
      RECT  101700.0 413550.0 102900.0 412350.0 ;
      RECT  104100.0 413550.0 105300.0 412350.0 ;
      RECT  104100.0 413550.0 105300.0 412350.0 ;
      RECT  101700.0 413550.0 102900.0 412350.0 ;
      RECT  101700.0 422850.0 102900.0 421650.0 ;
      RECT  104100.0 422850.0 105300.0 421650.0 ;
      RECT  104100.0 422850.0 105300.0 421650.0 ;
      RECT  101700.0 422850.0 102900.0 421650.0 ;
      RECT  106500.0 412950.0 107700.0 411750.0 ;
      RECT  106500.0 422850.0 107700.0 421650.0 ;
      RECT  102300.0 418200.0 103500.0 417000.0 ;
      RECT  102300.0 418200.0 103500.0 417000.0 ;
      RECT  104850.0 418050.0 105750.0 417150.0 ;
      RECT  99900.0 410850.0 109500.0 409950.0 ;
      RECT  99900.0 424650.0 109500.0 423750.0 ;
      RECT  106500.0 436050.0 107700.0 438000.0 ;
      RECT  106500.0 424200.0 107700.0 426150.0 ;
      RECT  101700.0 425550.0 102900.0 423750.0 ;
      RECT  101700.0 434850.0 102900.0 438450.0 ;
      RECT  104400.0 425550.0 105300.0 434850.0 ;
      RECT  101700.0 434850.0 102900.0 436050.0 ;
      RECT  104100.0 434850.0 105300.0 436050.0 ;
      RECT  104100.0 434850.0 105300.0 436050.0 ;
      RECT  101700.0 434850.0 102900.0 436050.0 ;
      RECT  101700.0 425550.0 102900.0 426750.0 ;
      RECT  104100.0 425550.0 105300.0 426750.0 ;
      RECT  104100.0 425550.0 105300.0 426750.0 ;
      RECT  101700.0 425550.0 102900.0 426750.0 ;
      RECT  106500.0 435450.0 107700.0 436650.0 ;
      RECT  106500.0 425550.0 107700.0 426750.0 ;
      RECT  102300.0 430200.0 103500.0 431400.0 ;
      RECT  102300.0 430200.0 103500.0 431400.0 ;
      RECT  104850.0 430350.0 105750.0 431250.0 ;
      RECT  99900.0 437550.0 109500.0 438450.0 ;
      RECT  99900.0 423750.0 109500.0 424650.0 ;
      RECT  106500.0 439950.0 107700.0 438000.0 ;
      RECT  106500.0 451800.0 107700.0 449850.0 ;
      RECT  101700.0 450450.0 102900.0 452250.0 ;
      RECT  101700.0 441150.0 102900.0 437550.0 ;
      RECT  104400.0 450450.0 105300.0 441150.0 ;
      RECT  101700.0 441150.0 102900.0 439950.0 ;
      RECT  104100.0 441150.0 105300.0 439950.0 ;
      RECT  104100.0 441150.0 105300.0 439950.0 ;
      RECT  101700.0 441150.0 102900.0 439950.0 ;
      RECT  101700.0 450450.0 102900.0 449250.0 ;
      RECT  104100.0 450450.0 105300.0 449250.0 ;
      RECT  104100.0 450450.0 105300.0 449250.0 ;
      RECT  101700.0 450450.0 102900.0 449250.0 ;
      RECT  106500.0 440550.0 107700.0 439350.0 ;
      RECT  106500.0 450450.0 107700.0 449250.0 ;
      RECT  102300.0 445800.0 103500.0 444600.0 ;
      RECT  102300.0 445800.0 103500.0 444600.0 ;
      RECT  104850.0 445650.0 105750.0 444750.0 ;
      RECT  99900.0 438450.0 109500.0 437550.0 ;
      RECT  99900.0 452250.0 109500.0 451350.0 ;
      RECT  106500.0 463650.0 107700.0 465600.0 ;
      RECT  106500.0 451800.0 107700.0 453750.0 ;
      RECT  101700.0 453150.0 102900.0 451350.0 ;
      RECT  101700.0 462450.0 102900.0 466050.0 ;
      RECT  104400.0 453150.0 105300.0 462450.0 ;
      RECT  101700.0 462450.0 102900.0 463650.0 ;
      RECT  104100.0 462450.0 105300.0 463650.0 ;
      RECT  104100.0 462450.0 105300.0 463650.0 ;
      RECT  101700.0 462450.0 102900.0 463650.0 ;
      RECT  101700.0 453150.0 102900.0 454350.0 ;
      RECT  104100.0 453150.0 105300.0 454350.0 ;
      RECT  104100.0 453150.0 105300.0 454350.0 ;
      RECT  101700.0 453150.0 102900.0 454350.0 ;
      RECT  106500.0 463050.0 107700.0 464250.0 ;
      RECT  106500.0 453150.0 107700.0 454350.0 ;
      RECT  102300.0 457800.0 103500.0 459000.0 ;
      RECT  102300.0 457800.0 103500.0 459000.0 ;
      RECT  104850.0 457950.0 105750.0 458850.0 ;
      RECT  99900.0 465150.0 109500.0 466050.0 ;
      RECT  99900.0 451350.0 109500.0 452250.0 ;
      RECT  106500.0 467550.0 107700.0 465600.0 ;
      RECT  106500.0 479400.0 107700.0 477450.0 ;
      RECT  101700.0 478050.0 102900.0 479850.0 ;
      RECT  101700.0 468750.0 102900.0 465150.0 ;
      RECT  104400.0 478050.0 105300.0 468750.0 ;
      RECT  101700.0 468750.0 102900.0 467550.0 ;
      RECT  104100.0 468750.0 105300.0 467550.0 ;
      RECT  104100.0 468750.0 105300.0 467550.0 ;
      RECT  101700.0 468750.0 102900.0 467550.0 ;
      RECT  101700.0 478050.0 102900.0 476850.0 ;
      RECT  104100.0 478050.0 105300.0 476850.0 ;
      RECT  104100.0 478050.0 105300.0 476850.0 ;
      RECT  101700.0 478050.0 102900.0 476850.0 ;
      RECT  106500.0 468150.0 107700.0 466950.0 ;
      RECT  106500.0 478050.0 107700.0 476850.0 ;
      RECT  102300.0 473400.0 103500.0 472200.0 ;
      RECT  102300.0 473400.0 103500.0 472200.0 ;
      RECT  104850.0 473250.0 105750.0 472350.0 ;
      RECT  99900.0 466050.0 109500.0 465150.0 ;
      RECT  99900.0 479850.0 109500.0 478950.0 ;
      RECT  106500.0 491250.0 107700.0 493200.0 ;
      RECT  106500.0 479400.0 107700.0 481350.0 ;
      RECT  101700.0 480750.0 102900.0 478950.0 ;
      RECT  101700.0 490050.0 102900.0 493650.0 ;
      RECT  104400.0 480750.0 105300.0 490050.0 ;
      RECT  101700.0 490050.0 102900.0 491250.0 ;
      RECT  104100.0 490050.0 105300.0 491250.0 ;
      RECT  104100.0 490050.0 105300.0 491250.0 ;
      RECT  101700.0 490050.0 102900.0 491250.0 ;
      RECT  101700.0 480750.0 102900.0 481950.0 ;
      RECT  104100.0 480750.0 105300.0 481950.0 ;
      RECT  104100.0 480750.0 105300.0 481950.0 ;
      RECT  101700.0 480750.0 102900.0 481950.0 ;
      RECT  106500.0 490650.0 107700.0 491850.0 ;
      RECT  106500.0 480750.0 107700.0 481950.0 ;
      RECT  102300.0 485400.0 103500.0 486600.0 ;
      RECT  102300.0 485400.0 103500.0 486600.0 ;
      RECT  104850.0 485550.0 105750.0 486450.0 ;
      RECT  99900.0 492750.0 109500.0 493650.0 ;
      RECT  99900.0 478950.0 109500.0 479850.0 ;
      RECT  106500.0 495150.0 107700.0 493200.0 ;
      RECT  106500.0 507000.0 107700.0 505050.0 ;
      RECT  101700.0 505650.0 102900.0 507450.0 ;
      RECT  101700.0 496350.0 102900.0 492750.0 ;
      RECT  104400.0 505650.0 105300.0 496350.0 ;
      RECT  101700.0 496350.0 102900.0 495150.0 ;
      RECT  104100.0 496350.0 105300.0 495150.0 ;
      RECT  104100.0 496350.0 105300.0 495150.0 ;
      RECT  101700.0 496350.0 102900.0 495150.0 ;
      RECT  101700.0 505650.0 102900.0 504450.0 ;
      RECT  104100.0 505650.0 105300.0 504450.0 ;
      RECT  104100.0 505650.0 105300.0 504450.0 ;
      RECT  101700.0 505650.0 102900.0 504450.0 ;
      RECT  106500.0 495750.0 107700.0 494550.0 ;
      RECT  106500.0 505650.0 107700.0 504450.0 ;
      RECT  102300.0 501000.0 103500.0 499800.0 ;
      RECT  102300.0 501000.0 103500.0 499800.0 ;
      RECT  104850.0 500850.0 105750.0 499950.0 ;
      RECT  99900.0 493650.0 109500.0 492750.0 ;
      RECT  99900.0 507450.0 109500.0 506550.0 ;
      RECT  106500.0 518850.0 107700.0 520800.0 ;
      RECT  106500.0 507000.0 107700.0 508950.0 ;
      RECT  101700.0 508350.0 102900.0 506550.0 ;
      RECT  101700.0 517650.0 102900.0 521250.0 ;
      RECT  104400.0 508350.0 105300.0 517650.0 ;
      RECT  101700.0 517650.0 102900.0 518850.0 ;
      RECT  104100.0 517650.0 105300.0 518850.0 ;
      RECT  104100.0 517650.0 105300.0 518850.0 ;
      RECT  101700.0 517650.0 102900.0 518850.0 ;
      RECT  101700.0 508350.0 102900.0 509550.0 ;
      RECT  104100.0 508350.0 105300.0 509550.0 ;
      RECT  104100.0 508350.0 105300.0 509550.0 ;
      RECT  101700.0 508350.0 102900.0 509550.0 ;
      RECT  106500.0 518250.0 107700.0 519450.0 ;
      RECT  106500.0 508350.0 107700.0 509550.0 ;
      RECT  102300.0 513000.0 103500.0 514200.0 ;
      RECT  102300.0 513000.0 103500.0 514200.0 ;
      RECT  104850.0 513150.0 105750.0 514050.0 ;
      RECT  99900.0 520350.0 109500.0 521250.0 ;
      RECT  99900.0 506550.0 109500.0 507450.0 ;
      RECT  106500.0 522750.0 107700.0 520800.0 ;
      RECT  106500.0 534600.0 107700.0 532650.0 ;
      RECT  101700.0 533250.0 102900.0 535050.0 ;
      RECT  101700.0 523950.0 102900.0 520350.0 ;
      RECT  104400.0 533250.0 105300.0 523950.0 ;
      RECT  101700.0 523950.0 102900.0 522750.0 ;
      RECT  104100.0 523950.0 105300.0 522750.0 ;
      RECT  104100.0 523950.0 105300.0 522750.0 ;
      RECT  101700.0 523950.0 102900.0 522750.0 ;
      RECT  101700.0 533250.0 102900.0 532050.0 ;
      RECT  104100.0 533250.0 105300.0 532050.0 ;
      RECT  104100.0 533250.0 105300.0 532050.0 ;
      RECT  101700.0 533250.0 102900.0 532050.0 ;
      RECT  106500.0 523350.0 107700.0 522150.0 ;
      RECT  106500.0 533250.0 107700.0 532050.0 ;
      RECT  102300.0 528600.0 103500.0 527400.0 ;
      RECT  102300.0 528600.0 103500.0 527400.0 ;
      RECT  104850.0 528450.0 105750.0 527550.0 ;
      RECT  99900.0 521250.0 109500.0 520350.0 ;
      RECT  99900.0 535050.0 109500.0 534150.0 ;
      RECT  106500.0 546450.0 107700.0 548400.0 ;
      RECT  106500.0 534600.0 107700.0 536550.0 ;
      RECT  101700.0 535950.0 102900.0 534150.0 ;
      RECT  101700.0 545250.0 102900.0 548850.0 ;
      RECT  104400.0 535950.0 105300.0 545250.0 ;
      RECT  101700.0 545250.0 102900.0 546450.0 ;
      RECT  104100.0 545250.0 105300.0 546450.0 ;
      RECT  104100.0 545250.0 105300.0 546450.0 ;
      RECT  101700.0 545250.0 102900.0 546450.0 ;
      RECT  101700.0 535950.0 102900.0 537150.0 ;
      RECT  104100.0 535950.0 105300.0 537150.0 ;
      RECT  104100.0 535950.0 105300.0 537150.0 ;
      RECT  101700.0 535950.0 102900.0 537150.0 ;
      RECT  106500.0 545850.0 107700.0 547050.0 ;
      RECT  106500.0 535950.0 107700.0 537150.0 ;
      RECT  102300.0 540600.0 103500.0 541800.0 ;
      RECT  102300.0 540600.0 103500.0 541800.0 ;
      RECT  104850.0 540750.0 105750.0 541650.0 ;
      RECT  99900.0 547950.0 109500.0 548850.0 ;
      RECT  99900.0 534150.0 109500.0 535050.0 ;
      RECT  106500.0 550350.0 107700.0 548400.0 ;
      RECT  106500.0 562200.0 107700.0 560250.0 ;
      RECT  101700.0 560850.0 102900.0 562650.0 ;
      RECT  101700.0 551550.0 102900.0 547950.0 ;
      RECT  104400.0 560850.0 105300.0 551550.0 ;
      RECT  101700.0 551550.0 102900.0 550350.0 ;
      RECT  104100.0 551550.0 105300.0 550350.0 ;
      RECT  104100.0 551550.0 105300.0 550350.0 ;
      RECT  101700.0 551550.0 102900.0 550350.0 ;
      RECT  101700.0 560850.0 102900.0 559650.0 ;
      RECT  104100.0 560850.0 105300.0 559650.0 ;
      RECT  104100.0 560850.0 105300.0 559650.0 ;
      RECT  101700.0 560850.0 102900.0 559650.0 ;
      RECT  106500.0 550950.0 107700.0 549750.0 ;
      RECT  106500.0 560850.0 107700.0 559650.0 ;
      RECT  102300.0 556200.0 103500.0 555000.0 ;
      RECT  102300.0 556200.0 103500.0 555000.0 ;
      RECT  104850.0 556050.0 105750.0 555150.0 ;
      RECT  99900.0 548850.0 109500.0 547950.0 ;
      RECT  99900.0 562650.0 109500.0 561750.0 ;
      RECT  106500.0 574050.0 107700.0 576000.0 ;
      RECT  106500.0 562200.0 107700.0 564150.0 ;
      RECT  101700.0 563550.0 102900.0 561750.0 ;
      RECT  101700.0 572850.0 102900.0 576450.0 ;
      RECT  104400.0 563550.0 105300.0 572850.0 ;
      RECT  101700.0 572850.0 102900.0 574050.0 ;
      RECT  104100.0 572850.0 105300.0 574050.0 ;
      RECT  104100.0 572850.0 105300.0 574050.0 ;
      RECT  101700.0 572850.0 102900.0 574050.0 ;
      RECT  101700.0 563550.0 102900.0 564750.0 ;
      RECT  104100.0 563550.0 105300.0 564750.0 ;
      RECT  104100.0 563550.0 105300.0 564750.0 ;
      RECT  101700.0 563550.0 102900.0 564750.0 ;
      RECT  106500.0 573450.0 107700.0 574650.0 ;
      RECT  106500.0 563550.0 107700.0 564750.0 ;
      RECT  102300.0 568200.0 103500.0 569400.0 ;
      RECT  102300.0 568200.0 103500.0 569400.0 ;
      RECT  104850.0 568350.0 105750.0 569250.0 ;
      RECT  99900.0 575550.0 109500.0 576450.0 ;
      RECT  99900.0 561750.0 109500.0 562650.0 ;
      RECT  106500.0 577950.0 107700.0 576000.0 ;
      RECT  106500.0 589800.0 107700.0 587850.0 ;
      RECT  101700.0 588450.0 102900.0 590250.0 ;
      RECT  101700.0 579150.0 102900.0 575550.0 ;
      RECT  104400.0 588450.0 105300.0 579150.0 ;
      RECT  101700.0 579150.0 102900.0 577950.0 ;
      RECT  104100.0 579150.0 105300.0 577950.0 ;
      RECT  104100.0 579150.0 105300.0 577950.0 ;
      RECT  101700.0 579150.0 102900.0 577950.0 ;
      RECT  101700.0 588450.0 102900.0 587250.0 ;
      RECT  104100.0 588450.0 105300.0 587250.0 ;
      RECT  104100.0 588450.0 105300.0 587250.0 ;
      RECT  101700.0 588450.0 102900.0 587250.0 ;
      RECT  106500.0 578550.0 107700.0 577350.0 ;
      RECT  106500.0 588450.0 107700.0 587250.0 ;
      RECT  102300.0 583800.0 103500.0 582600.0 ;
      RECT  102300.0 583800.0 103500.0 582600.0 ;
      RECT  104850.0 583650.0 105750.0 582750.0 ;
      RECT  99900.0 576450.0 109500.0 575550.0 ;
      RECT  99900.0 590250.0 109500.0 589350.0 ;
      RECT  106500.0 601650.0 107700.0 603600.0 ;
      RECT  106500.0 589800.0 107700.0 591750.0 ;
      RECT  101700.0 591150.0 102900.0 589350.0 ;
      RECT  101700.0 600450.0 102900.0 604050.0 ;
      RECT  104400.0 591150.0 105300.0 600450.0 ;
      RECT  101700.0 600450.0 102900.0 601650.0 ;
      RECT  104100.0 600450.0 105300.0 601650.0 ;
      RECT  104100.0 600450.0 105300.0 601650.0 ;
      RECT  101700.0 600450.0 102900.0 601650.0 ;
      RECT  101700.0 591150.0 102900.0 592350.0 ;
      RECT  104100.0 591150.0 105300.0 592350.0 ;
      RECT  104100.0 591150.0 105300.0 592350.0 ;
      RECT  101700.0 591150.0 102900.0 592350.0 ;
      RECT  106500.0 601050.0 107700.0 602250.0 ;
      RECT  106500.0 591150.0 107700.0 592350.0 ;
      RECT  102300.0 595800.0 103500.0 597000.0 ;
      RECT  102300.0 595800.0 103500.0 597000.0 ;
      RECT  104850.0 595950.0 105750.0 596850.0 ;
      RECT  99900.0 603150.0 109500.0 604050.0 ;
      RECT  99900.0 589350.0 109500.0 590250.0 ;
      RECT  106500.0 605550.0 107700.0 603600.0 ;
      RECT  106500.0 617400.0 107700.0 615450.0 ;
      RECT  101700.0 616050.0 102900.0 617850.0 ;
      RECT  101700.0 606750.0 102900.0 603150.0 ;
      RECT  104400.0 616050.0 105300.0 606750.0 ;
      RECT  101700.0 606750.0 102900.0 605550.0 ;
      RECT  104100.0 606750.0 105300.0 605550.0 ;
      RECT  104100.0 606750.0 105300.0 605550.0 ;
      RECT  101700.0 606750.0 102900.0 605550.0 ;
      RECT  101700.0 616050.0 102900.0 614850.0 ;
      RECT  104100.0 616050.0 105300.0 614850.0 ;
      RECT  104100.0 616050.0 105300.0 614850.0 ;
      RECT  101700.0 616050.0 102900.0 614850.0 ;
      RECT  106500.0 606150.0 107700.0 604950.0 ;
      RECT  106500.0 616050.0 107700.0 614850.0 ;
      RECT  102300.0 611400.0 103500.0 610200.0 ;
      RECT  102300.0 611400.0 103500.0 610200.0 ;
      RECT  104850.0 611250.0 105750.0 610350.0 ;
      RECT  99900.0 604050.0 109500.0 603150.0 ;
      RECT  99900.0 617850.0 109500.0 616950.0 ;
      RECT  106500.0 629250.0 107700.0 631200.0 ;
      RECT  106500.0 617400.0 107700.0 619350.0 ;
      RECT  101700.0 618750.0 102900.0 616950.0 ;
      RECT  101700.0 628050.0 102900.0 631650.0 ;
      RECT  104400.0 618750.0 105300.0 628050.0 ;
      RECT  101700.0 628050.0 102900.0 629250.0 ;
      RECT  104100.0 628050.0 105300.0 629250.0 ;
      RECT  104100.0 628050.0 105300.0 629250.0 ;
      RECT  101700.0 628050.0 102900.0 629250.0 ;
      RECT  101700.0 618750.0 102900.0 619950.0 ;
      RECT  104100.0 618750.0 105300.0 619950.0 ;
      RECT  104100.0 618750.0 105300.0 619950.0 ;
      RECT  101700.0 618750.0 102900.0 619950.0 ;
      RECT  106500.0 628650.0 107700.0 629850.0 ;
      RECT  106500.0 618750.0 107700.0 619950.0 ;
      RECT  102300.0 623400.0 103500.0 624600.0 ;
      RECT  102300.0 623400.0 103500.0 624600.0 ;
      RECT  104850.0 623550.0 105750.0 624450.0 ;
      RECT  99900.0 630750.0 109500.0 631650.0 ;
      RECT  99900.0 616950.0 109500.0 617850.0 ;
      RECT  106500.0 633150.0 107700.0 631200.0 ;
      RECT  106500.0 645000.0 107700.0 643050.0 ;
      RECT  101700.0 643650.0 102900.0 645450.0 ;
      RECT  101700.0 634350.0 102900.0 630750.0 ;
      RECT  104400.0 643650.0 105300.0 634350.0 ;
      RECT  101700.0 634350.0 102900.0 633150.0 ;
      RECT  104100.0 634350.0 105300.0 633150.0 ;
      RECT  104100.0 634350.0 105300.0 633150.0 ;
      RECT  101700.0 634350.0 102900.0 633150.0 ;
      RECT  101700.0 643650.0 102900.0 642450.0 ;
      RECT  104100.0 643650.0 105300.0 642450.0 ;
      RECT  104100.0 643650.0 105300.0 642450.0 ;
      RECT  101700.0 643650.0 102900.0 642450.0 ;
      RECT  106500.0 633750.0 107700.0 632550.0 ;
      RECT  106500.0 643650.0 107700.0 642450.0 ;
      RECT  102300.0 639000.0 103500.0 637800.0 ;
      RECT  102300.0 639000.0 103500.0 637800.0 ;
      RECT  104850.0 638850.0 105750.0 637950.0 ;
      RECT  99900.0 631650.0 109500.0 630750.0 ;
      RECT  99900.0 645450.0 109500.0 644550.0 ;
      RECT  106500.0 656850.0 107700.0 658800.0 ;
      RECT  106500.0 645000.0 107700.0 646950.0 ;
      RECT  101700.0 646350.0 102900.0 644550.0 ;
      RECT  101700.0 655650.0 102900.0 659250.0 ;
      RECT  104400.0 646350.0 105300.0 655650.0 ;
      RECT  101700.0 655650.0 102900.0 656850.0 ;
      RECT  104100.0 655650.0 105300.0 656850.0 ;
      RECT  104100.0 655650.0 105300.0 656850.0 ;
      RECT  101700.0 655650.0 102900.0 656850.0 ;
      RECT  101700.0 646350.0 102900.0 647550.0 ;
      RECT  104100.0 646350.0 105300.0 647550.0 ;
      RECT  104100.0 646350.0 105300.0 647550.0 ;
      RECT  101700.0 646350.0 102900.0 647550.0 ;
      RECT  106500.0 656250.0 107700.0 657450.0 ;
      RECT  106500.0 646350.0 107700.0 647550.0 ;
      RECT  102300.0 651000.0 103500.0 652200.0 ;
      RECT  102300.0 651000.0 103500.0 652200.0 ;
      RECT  104850.0 651150.0 105750.0 652050.0 ;
      RECT  99900.0 658350.0 109500.0 659250.0 ;
      RECT  99900.0 644550.0 109500.0 645450.0 ;
      RECT  106500.0 660750.0 107700.0 658800.0 ;
      RECT  106500.0 672600.0 107700.0 670650.0 ;
      RECT  101700.0 671250.0 102900.0 673050.0 ;
      RECT  101700.0 661950.0 102900.0 658350.0 ;
      RECT  104400.0 671250.0 105300.0 661950.0 ;
      RECT  101700.0 661950.0 102900.0 660750.0 ;
      RECT  104100.0 661950.0 105300.0 660750.0 ;
      RECT  104100.0 661950.0 105300.0 660750.0 ;
      RECT  101700.0 661950.0 102900.0 660750.0 ;
      RECT  101700.0 671250.0 102900.0 670050.0 ;
      RECT  104100.0 671250.0 105300.0 670050.0 ;
      RECT  104100.0 671250.0 105300.0 670050.0 ;
      RECT  101700.0 671250.0 102900.0 670050.0 ;
      RECT  106500.0 661350.0 107700.0 660150.0 ;
      RECT  106500.0 671250.0 107700.0 670050.0 ;
      RECT  102300.0 666600.0 103500.0 665400.0 ;
      RECT  102300.0 666600.0 103500.0 665400.0 ;
      RECT  104850.0 666450.0 105750.0 665550.0 ;
      RECT  99900.0 659250.0 109500.0 658350.0 ;
      RECT  99900.0 673050.0 109500.0 672150.0 ;
      RECT  106500.0 684450.0 107700.0 686400.0 ;
      RECT  106500.0 672600.0 107700.0 674550.0 ;
      RECT  101700.0 673950.0 102900.0 672150.0 ;
      RECT  101700.0 683250.0 102900.0 686850.0 ;
      RECT  104400.0 673950.0 105300.0 683250.0 ;
      RECT  101700.0 683250.0 102900.0 684450.0 ;
      RECT  104100.0 683250.0 105300.0 684450.0 ;
      RECT  104100.0 683250.0 105300.0 684450.0 ;
      RECT  101700.0 683250.0 102900.0 684450.0 ;
      RECT  101700.0 673950.0 102900.0 675150.0 ;
      RECT  104100.0 673950.0 105300.0 675150.0 ;
      RECT  104100.0 673950.0 105300.0 675150.0 ;
      RECT  101700.0 673950.0 102900.0 675150.0 ;
      RECT  106500.0 683850.0 107700.0 685050.0 ;
      RECT  106500.0 673950.0 107700.0 675150.0 ;
      RECT  102300.0 678600.0 103500.0 679800.0 ;
      RECT  102300.0 678600.0 103500.0 679800.0 ;
      RECT  104850.0 678750.0 105750.0 679650.0 ;
      RECT  99900.0 685950.0 109500.0 686850.0 ;
      RECT  99900.0 672150.0 109500.0 673050.0 ;
      RECT  106500.0 688350.0 107700.0 686400.0 ;
      RECT  106500.0 700200.0 107700.0 698250.0 ;
      RECT  101700.0 698850.0 102900.0 700650.0 ;
      RECT  101700.0 689550.0 102900.0 685950.0 ;
      RECT  104400.0 698850.0 105300.0 689550.0 ;
      RECT  101700.0 689550.0 102900.0 688350.0 ;
      RECT  104100.0 689550.0 105300.0 688350.0 ;
      RECT  104100.0 689550.0 105300.0 688350.0 ;
      RECT  101700.0 689550.0 102900.0 688350.0 ;
      RECT  101700.0 698850.0 102900.0 697650.0 ;
      RECT  104100.0 698850.0 105300.0 697650.0 ;
      RECT  104100.0 698850.0 105300.0 697650.0 ;
      RECT  101700.0 698850.0 102900.0 697650.0 ;
      RECT  106500.0 688950.0 107700.0 687750.0 ;
      RECT  106500.0 698850.0 107700.0 697650.0 ;
      RECT  102300.0 694200.0 103500.0 693000.0 ;
      RECT  102300.0 694200.0 103500.0 693000.0 ;
      RECT  104850.0 694050.0 105750.0 693150.0 ;
      RECT  99900.0 686850.0 109500.0 685950.0 ;
      RECT  99900.0 700650.0 109500.0 699750.0 ;
      RECT  106500.0 712050.0 107700.0 714000.0 ;
      RECT  106500.0 700200.0 107700.0 702150.0 ;
      RECT  101700.0 701550.0 102900.0 699750.0 ;
      RECT  101700.0 710850.0 102900.0 714450.0 ;
      RECT  104400.0 701550.0 105300.0 710850.0 ;
      RECT  101700.0 710850.0 102900.0 712050.0 ;
      RECT  104100.0 710850.0 105300.0 712050.0 ;
      RECT  104100.0 710850.0 105300.0 712050.0 ;
      RECT  101700.0 710850.0 102900.0 712050.0 ;
      RECT  101700.0 701550.0 102900.0 702750.0 ;
      RECT  104100.0 701550.0 105300.0 702750.0 ;
      RECT  104100.0 701550.0 105300.0 702750.0 ;
      RECT  101700.0 701550.0 102900.0 702750.0 ;
      RECT  106500.0 711450.0 107700.0 712650.0 ;
      RECT  106500.0 701550.0 107700.0 702750.0 ;
      RECT  102300.0 706200.0 103500.0 707400.0 ;
      RECT  102300.0 706200.0 103500.0 707400.0 ;
      RECT  104850.0 706350.0 105750.0 707250.0 ;
      RECT  99900.0 713550.0 109500.0 714450.0 ;
      RECT  99900.0 699750.0 109500.0 700650.0 ;
      RECT  106500.0 715950.0 107700.0 714000.0 ;
      RECT  106500.0 727800.0 107700.0 725850.0 ;
      RECT  101700.0 726450.0 102900.0 728250.0 ;
      RECT  101700.0 717150.0 102900.0 713550.0 ;
      RECT  104400.0 726450.0 105300.0 717150.0 ;
      RECT  101700.0 717150.0 102900.0 715950.0 ;
      RECT  104100.0 717150.0 105300.0 715950.0 ;
      RECT  104100.0 717150.0 105300.0 715950.0 ;
      RECT  101700.0 717150.0 102900.0 715950.0 ;
      RECT  101700.0 726450.0 102900.0 725250.0 ;
      RECT  104100.0 726450.0 105300.0 725250.0 ;
      RECT  104100.0 726450.0 105300.0 725250.0 ;
      RECT  101700.0 726450.0 102900.0 725250.0 ;
      RECT  106500.0 716550.0 107700.0 715350.0 ;
      RECT  106500.0 726450.0 107700.0 725250.0 ;
      RECT  102300.0 721800.0 103500.0 720600.0 ;
      RECT  102300.0 721800.0 103500.0 720600.0 ;
      RECT  104850.0 721650.0 105750.0 720750.0 ;
      RECT  99900.0 714450.0 109500.0 713550.0 ;
      RECT  99900.0 728250.0 109500.0 727350.0 ;
      RECT  106500.0 739650.0 107700.0 741600.0 ;
      RECT  106500.0 727800.0 107700.0 729750.0 ;
      RECT  101700.0 729150.0 102900.0 727350.0 ;
      RECT  101700.0 738450.0 102900.0 742050.0 ;
      RECT  104400.0 729150.0 105300.0 738450.0 ;
      RECT  101700.0 738450.0 102900.0 739650.0 ;
      RECT  104100.0 738450.0 105300.0 739650.0 ;
      RECT  104100.0 738450.0 105300.0 739650.0 ;
      RECT  101700.0 738450.0 102900.0 739650.0 ;
      RECT  101700.0 729150.0 102900.0 730350.0 ;
      RECT  104100.0 729150.0 105300.0 730350.0 ;
      RECT  104100.0 729150.0 105300.0 730350.0 ;
      RECT  101700.0 729150.0 102900.0 730350.0 ;
      RECT  106500.0 739050.0 107700.0 740250.0 ;
      RECT  106500.0 729150.0 107700.0 730350.0 ;
      RECT  102300.0 733800.0 103500.0 735000.0 ;
      RECT  102300.0 733800.0 103500.0 735000.0 ;
      RECT  104850.0 733950.0 105750.0 734850.0 ;
      RECT  99900.0 741150.0 109500.0 742050.0 ;
      RECT  99900.0 727350.0 109500.0 728250.0 ;
      RECT  106500.0 743550.0 107700.0 741600.0 ;
      RECT  106500.0 755400.0 107700.0 753450.0 ;
      RECT  101700.0 754050.0 102900.0 755850.0 ;
      RECT  101700.0 744750.0 102900.0 741150.0 ;
      RECT  104400.0 754050.0 105300.0 744750.0 ;
      RECT  101700.0 744750.0 102900.0 743550.0 ;
      RECT  104100.0 744750.0 105300.0 743550.0 ;
      RECT  104100.0 744750.0 105300.0 743550.0 ;
      RECT  101700.0 744750.0 102900.0 743550.0 ;
      RECT  101700.0 754050.0 102900.0 752850.0 ;
      RECT  104100.0 754050.0 105300.0 752850.0 ;
      RECT  104100.0 754050.0 105300.0 752850.0 ;
      RECT  101700.0 754050.0 102900.0 752850.0 ;
      RECT  106500.0 744150.0 107700.0 742950.0 ;
      RECT  106500.0 754050.0 107700.0 752850.0 ;
      RECT  102300.0 749400.0 103500.0 748200.0 ;
      RECT  102300.0 749400.0 103500.0 748200.0 ;
      RECT  104850.0 749250.0 105750.0 748350.0 ;
      RECT  99900.0 742050.0 109500.0 741150.0 ;
      RECT  99900.0 755850.0 109500.0 754950.0 ;
      RECT  106500.0 767250.0 107700.0 769200.0 ;
      RECT  106500.0 755400.0 107700.0 757350.0 ;
      RECT  101700.0 756750.0 102900.0 754950.0 ;
      RECT  101700.0 766050.0 102900.0 769650.0 ;
      RECT  104400.0 756750.0 105300.0 766050.0 ;
      RECT  101700.0 766050.0 102900.0 767250.0 ;
      RECT  104100.0 766050.0 105300.0 767250.0 ;
      RECT  104100.0 766050.0 105300.0 767250.0 ;
      RECT  101700.0 766050.0 102900.0 767250.0 ;
      RECT  101700.0 756750.0 102900.0 757950.0 ;
      RECT  104100.0 756750.0 105300.0 757950.0 ;
      RECT  104100.0 756750.0 105300.0 757950.0 ;
      RECT  101700.0 756750.0 102900.0 757950.0 ;
      RECT  106500.0 766650.0 107700.0 767850.0 ;
      RECT  106500.0 756750.0 107700.0 757950.0 ;
      RECT  102300.0 761400.0 103500.0 762600.0 ;
      RECT  102300.0 761400.0 103500.0 762600.0 ;
      RECT  104850.0 761550.0 105750.0 762450.0 ;
      RECT  99900.0 768750.0 109500.0 769650.0 ;
      RECT  99900.0 754950.0 109500.0 755850.0 ;
      RECT  106500.0 771150.0 107700.0 769200.0 ;
      RECT  106500.0 783000.0 107700.0 781050.0 ;
      RECT  101700.0 781650.0 102900.0 783450.0 ;
      RECT  101700.0 772350.0 102900.0 768750.0 ;
      RECT  104400.0 781650.0 105300.0 772350.0 ;
      RECT  101700.0 772350.0 102900.0 771150.0 ;
      RECT  104100.0 772350.0 105300.0 771150.0 ;
      RECT  104100.0 772350.0 105300.0 771150.0 ;
      RECT  101700.0 772350.0 102900.0 771150.0 ;
      RECT  101700.0 781650.0 102900.0 780450.0 ;
      RECT  104100.0 781650.0 105300.0 780450.0 ;
      RECT  104100.0 781650.0 105300.0 780450.0 ;
      RECT  101700.0 781650.0 102900.0 780450.0 ;
      RECT  106500.0 771750.0 107700.0 770550.0 ;
      RECT  106500.0 781650.0 107700.0 780450.0 ;
      RECT  102300.0 777000.0 103500.0 775800.0 ;
      RECT  102300.0 777000.0 103500.0 775800.0 ;
      RECT  104850.0 776850.0 105750.0 775950.0 ;
      RECT  99900.0 769650.0 109500.0 768750.0 ;
      RECT  99900.0 783450.0 109500.0 782550.0 ;
      RECT  106500.0 794850.0 107700.0 796800.0 ;
      RECT  106500.0 783000.0 107700.0 784950.0 ;
      RECT  101700.0 784350.0 102900.0 782550.0 ;
      RECT  101700.0 793650.0 102900.0 797250.0 ;
      RECT  104400.0 784350.0 105300.0 793650.0 ;
      RECT  101700.0 793650.0 102900.0 794850.0 ;
      RECT  104100.0 793650.0 105300.0 794850.0 ;
      RECT  104100.0 793650.0 105300.0 794850.0 ;
      RECT  101700.0 793650.0 102900.0 794850.0 ;
      RECT  101700.0 784350.0 102900.0 785550.0 ;
      RECT  104100.0 784350.0 105300.0 785550.0 ;
      RECT  104100.0 784350.0 105300.0 785550.0 ;
      RECT  101700.0 784350.0 102900.0 785550.0 ;
      RECT  106500.0 794250.0 107700.0 795450.0 ;
      RECT  106500.0 784350.0 107700.0 785550.0 ;
      RECT  102300.0 789000.0 103500.0 790200.0 ;
      RECT  102300.0 789000.0 103500.0 790200.0 ;
      RECT  104850.0 789150.0 105750.0 790050.0 ;
      RECT  99900.0 796350.0 109500.0 797250.0 ;
      RECT  99900.0 782550.0 109500.0 783450.0 ;
      RECT  106500.0 798750.0 107700.0 796800.0 ;
      RECT  106500.0 810600.0 107700.0 808650.0 ;
      RECT  101700.0 809250.0 102900.0 811050.0 ;
      RECT  101700.0 799950.0 102900.0 796350.0 ;
      RECT  104400.0 809250.0 105300.0 799950.0 ;
      RECT  101700.0 799950.0 102900.0 798750.0 ;
      RECT  104100.0 799950.0 105300.0 798750.0 ;
      RECT  104100.0 799950.0 105300.0 798750.0 ;
      RECT  101700.0 799950.0 102900.0 798750.0 ;
      RECT  101700.0 809250.0 102900.0 808050.0 ;
      RECT  104100.0 809250.0 105300.0 808050.0 ;
      RECT  104100.0 809250.0 105300.0 808050.0 ;
      RECT  101700.0 809250.0 102900.0 808050.0 ;
      RECT  106500.0 799350.0 107700.0 798150.0 ;
      RECT  106500.0 809250.0 107700.0 808050.0 ;
      RECT  102300.0 804600.0 103500.0 803400.0 ;
      RECT  102300.0 804600.0 103500.0 803400.0 ;
      RECT  104850.0 804450.0 105750.0 803550.0 ;
      RECT  99900.0 797250.0 109500.0 796350.0 ;
      RECT  99900.0 811050.0 109500.0 810150.0 ;
      RECT  106500.0 822450.0 107700.0 824400.0 ;
      RECT  106500.0 810600.0 107700.0 812550.0 ;
      RECT  101700.0 811950.0 102900.0 810150.0 ;
      RECT  101700.0 821250.0 102900.0 824850.0 ;
      RECT  104400.0 811950.0 105300.0 821250.0 ;
      RECT  101700.0 821250.0 102900.0 822450.0 ;
      RECT  104100.0 821250.0 105300.0 822450.0 ;
      RECT  104100.0 821250.0 105300.0 822450.0 ;
      RECT  101700.0 821250.0 102900.0 822450.0 ;
      RECT  101700.0 811950.0 102900.0 813150.0 ;
      RECT  104100.0 811950.0 105300.0 813150.0 ;
      RECT  104100.0 811950.0 105300.0 813150.0 ;
      RECT  101700.0 811950.0 102900.0 813150.0 ;
      RECT  106500.0 821850.0 107700.0 823050.0 ;
      RECT  106500.0 811950.0 107700.0 813150.0 ;
      RECT  102300.0 816600.0 103500.0 817800.0 ;
      RECT  102300.0 816600.0 103500.0 817800.0 ;
      RECT  104850.0 816750.0 105750.0 817650.0 ;
      RECT  99900.0 823950.0 109500.0 824850.0 ;
      RECT  99900.0 810150.0 109500.0 811050.0 ;
      RECT  106500.0 826350.0 107700.0 824400.0 ;
      RECT  106500.0 838200.0 107700.0 836250.0 ;
      RECT  101700.0 836850.0 102900.0 838650.0 ;
      RECT  101700.0 827550.0 102900.0 823950.0 ;
      RECT  104400.0 836850.0 105300.0 827550.0 ;
      RECT  101700.0 827550.0 102900.0 826350.0 ;
      RECT  104100.0 827550.0 105300.0 826350.0 ;
      RECT  104100.0 827550.0 105300.0 826350.0 ;
      RECT  101700.0 827550.0 102900.0 826350.0 ;
      RECT  101700.0 836850.0 102900.0 835650.0 ;
      RECT  104100.0 836850.0 105300.0 835650.0 ;
      RECT  104100.0 836850.0 105300.0 835650.0 ;
      RECT  101700.0 836850.0 102900.0 835650.0 ;
      RECT  106500.0 826950.0 107700.0 825750.0 ;
      RECT  106500.0 836850.0 107700.0 835650.0 ;
      RECT  102300.0 832200.0 103500.0 831000.0 ;
      RECT  102300.0 832200.0 103500.0 831000.0 ;
      RECT  104850.0 832050.0 105750.0 831150.0 ;
      RECT  99900.0 824850.0 109500.0 823950.0 ;
      RECT  99900.0 838650.0 109500.0 837750.0 ;
      RECT  106500.0 850050.0 107700.0 852000.0 ;
      RECT  106500.0 838200.0 107700.0 840150.0 ;
      RECT  101700.0 839550.0 102900.0 837750.0 ;
      RECT  101700.0 848850.0 102900.0 852450.0 ;
      RECT  104400.0 839550.0 105300.0 848850.0 ;
      RECT  101700.0 848850.0 102900.0 850050.0 ;
      RECT  104100.0 848850.0 105300.0 850050.0 ;
      RECT  104100.0 848850.0 105300.0 850050.0 ;
      RECT  101700.0 848850.0 102900.0 850050.0 ;
      RECT  101700.0 839550.0 102900.0 840750.0 ;
      RECT  104100.0 839550.0 105300.0 840750.0 ;
      RECT  104100.0 839550.0 105300.0 840750.0 ;
      RECT  101700.0 839550.0 102900.0 840750.0 ;
      RECT  106500.0 849450.0 107700.0 850650.0 ;
      RECT  106500.0 839550.0 107700.0 840750.0 ;
      RECT  102300.0 844200.0 103500.0 845400.0 ;
      RECT  102300.0 844200.0 103500.0 845400.0 ;
      RECT  104850.0 844350.0 105750.0 845250.0 ;
      RECT  99900.0 851550.0 109500.0 852450.0 ;
      RECT  99900.0 837750.0 109500.0 838650.0 ;
      RECT  106500.0 853950.0 107700.0 852000.0 ;
      RECT  106500.0 865800.0 107700.0 863850.0 ;
      RECT  101700.0 864450.0 102900.0 866250.0 ;
      RECT  101700.0 855150.0 102900.0 851550.0 ;
      RECT  104400.0 864450.0 105300.0 855150.0 ;
      RECT  101700.0 855150.0 102900.0 853950.0 ;
      RECT  104100.0 855150.0 105300.0 853950.0 ;
      RECT  104100.0 855150.0 105300.0 853950.0 ;
      RECT  101700.0 855150.0 102900.0 853950.0 ;
      RECT  101700.0 864450.0 102900.0 863250.0 ;
      RECT  104100.0 864450.0 105300.0 863250.0 ;
      RECT  104100.0 864450.0 105300.0 863250.0 ;
      RECT  101700.0 864450.0 102900.0 863250.0 ;
      RECT  106500.0 854550.0 107700.0 853350.0 ;
      RECT  106500.0 864450.0 107700.0 863250.0 ;
      RECT  102300.0 859800.0 103500.0 858600.0 ;
      RECT  102300.0 859800.0 103500.0 858600.0 ;
      RECT  104850.0 859650.0 105750.0 858750.0 ;
      RECT  99900.0 852450.0 109500.0 851550.0 ;
      RECT  99900.0 866250.0 109500.0 865350.0 ;
      RECT  106500.0 877650.0 107700.0 879600.0 ;
      RECT  106500.0 865800.0 107700.0 867750.0 ;
      RECT  101700.0 867150.0 102900.0 865350.0 ;
      RECT  101700.0 876450.0 102900.0 880050.0 ;
      RECT  104400.0 867150.0 105300.0 876450.0 ;
      RECT  101700.0 876450.0 102900.0 877650.0 ;
      RECT  104100.0 876450.0 105300.0 877650.0 ;
      RECT  104100.0 876450.0 105300.0 877650.0 ;
      RECT  101700.0 876450.0 102900.0 877650.0 ;
      RECT  101700.0 867150.0 102900.0 868350.0 ;
      RECT  104100.0 867150.0 105300.0 868350.0 ;
      RECT  104100.0 867150.0 105300.0 868350.0 ;
      RECT  101700.0 867150.0 102900.0 868350.0 ;
      RECT  106500.0 877050.0 107700.0 878250.0 ;
      RECT  106500.0 867150.0 107700.0 868350.0 ;
      RECT  102300.0 871800.0 103500.0 873000.0 ;
      RECT  102300.0 871800.0 103500.0 873000.0 ;
      RECT  104850.0 871950.0 105750.0 872850.0 ;
      RECT  99900.0 879150.0 109500.0 880050.0 ;
      RECT  99900.0 865350.0 109500.0 866250.0 ;
      RECT  106500.0 881550.0 107700.0 879600.0 ;
      RECT  106500.0 893400.0 107700.0 891450.0 ;
      RECT  101700.0 892050.0 102900.0 893850.0 ;
      RECT  101700.0 882750.0 102900.0 879150.0 ;
      RECT  104400.0 892050.0 105300.0 882750.0 ;
      RECT  101700.0 882750.0 102900.0 881550.0 ;
      RECT  104100.0 882750.0 105300.0 881550.0 ;
      RECT  104100.0 882750.0 105300.0 881550.0 ;
      RECT  101700.0 882750.0 102900.0 881550.0 ;
      RECT  101700.0 892050.0 102900.0 890850.0 ;
      RECT  104100.0 892050.0 105300.0 890850.0 ;
      RECT  104100.0 892050.0 105300.0 890850.0 ;
      RECT  101700.0 892050.0 102900.0 890850.0 ;
      RECT  106500.0 882150.0 107700.0 880950.0 ;
      RECT  106500.0 892050.0 107700.0 890850.0 ;
      RECT  102300.0 887400.0 103500.0 886200.0 ;
      RECT  102300.0 887400.0 103500.0 886200.0 ;
      RECT  104850.0 887250.0 105750.0 886350.0 ;
      RECT  99900.0 880050.0 109500.0 879150.0 ;
      RECT  99900.0 893850.0 109500.0 892950.0 ;
      RECT  106500.0 905250.0 107700.0 907200.0 ;
      RECT  106500.0 893400.0 107700.0 895350.0 ;
      RECT  101700.0 894750.0 102900.0 892950.0 ;
      RECT  101700.0 904050.0 102900.0 907650.0 ;
      RECT  104400.0 894750.0 105300.0 904050.0 ;
      RECT  101700.0 904050.0 102900.0 905250.0 ;
      RECT  104100.0 904050.0 105300.0 905250.0 ;
      RECT  104100.0 904050.0 105300.0 905250.0 ;
      RECT  101700.0 904050.0 102900.0 905250.0 ;
      RECT  101700.0 894750.0 102900.0 895950.0 ;
      RECT  104100.0 894750.0 105300.0 895950.0 ;
      RECT  104100.0 894750.0 105300.0 895950.0 ;
      RECT  101700.0 894750.0 102900.0 895950.0 ;
      RECT  106500.0 904650.0 107700.0 905850.0 ;
      RECT  106500.0 894750.0 107700.0 895950.0 ;
      RECT  102300.0 899400.0 103500.0 900600.0 ;
      RECT  102300.0 899400.0 103500.0 900600.0 ;
      RECT  104850.0 899550.0 105750.0 900450.0 ;
      RECT  99900.0 906750.0 109500.0 907650.0 ;
      RECT  99900.0 892950.0 109500.0 893850.0 ;
      RECT  106500.0 909150.0 107700.0 907200.0 ;
      RECT  106500.0 921000.0 107700.0 919050.0 ;
      RECT  101700.0 919650.0 102900.0 921450.0 ;
      RECT  101700.0 910350.0 102900.0 906750.0 ;
      RECT  104400.0 919650.0 105300.0 910350.0 ;
      RECT  101700.0 910350.0 102900.0 909150.0 ;
      RECT  104100.0 910350.0 105300.0 909150.0 ;
      RECT  104100.0 910350.0 105300.0 909150.0 ;
      RECT  101700.0 910350.0 102900.0 909150.0 ;
      RECT  101700.0 919650.0 102900.0 918450.0 ;
      RECT  104100.0 919650.0 105300.0 918450.0 ;
      RECT  104100.0 919650.0 105300.0 918450.0 ;
      RECT  101700.0 919650.0 102900.0 918450.0 ;
      RECT  106500.0 909750.0 107700.0 908550.0 ;
      RECT  106500.0 919650.0 107700.0 918450.0 ;
      RECT  102300.0 915000.0 103500.0 913800.0 ;
      RECT  102300.0 915000.0 103500.0 913800.0 ;
      RECT  104850.0 914850.0 105750.0 913950.0 ;
      RECT  99900.0 907650.0 109500.0 906750.0 ;
      RECT  99900.0 921450.0 109500.0 920550.0 ;
      RECT  106500.0 932850.0 107700.0 934800.0 ;
      RECT  106500.0 921000.0 107700.0 922950.0 ;
      RECT  101700.0 922350.0 102900.0 920550.0 ;
      RECT  101700.0 931650.0 102900.0 935250.0 ;
      RECT  104400.0 922350.0 105300.0 931650.0 ;
      RECT  101700.0 931650.0 102900.0 932850.0 ;
      RECT  104100.0 931650.0 105300.0 932850.0 ;
      RECT  104100.0 931650.0 105300.0 932850.0 ;
      RECT  101700.0 931650.0 102900.0 932850.0 ;
      RECT  101700.0 922350.0 102900.0 923550.0 ;
      RECT  104100.0 922350.0 105300.0 923550.0 ;
      RECT  104100.0 922350.0 105300.0 923550.0 ;
      RECT  101700.0 922350.0 102900.0 923550.0 ;
      RECT  106500.0 932250.0 107700.0 933450.0 ;
      RECT  106500.0 922350.0 107700.0 923550.0 ;
      RECT  102300.0 927000.0 103500.0 928200.0 ;
      RECT  102300.0 927000.0 103500.0 928200.0 ;
      RECT  104850.0 927150.0 105750.0 928050.0 ;
      RECT  99900.0 934350.0 109500.0 935250.0 ;
      RECT  99900.0 920550.0 109500.0 921450.0 ;
      RECT  106500.0 936750.0 107700.0 934800.0 ;
      RECT  106500.0 948600.0 107700.0 946650.0 ;
      RECT  101700.0 947250.0 102900.0 949050.0 ;
      RECT  101700.0 937950.0 102900.0 934350.0 ;
      RECT  104400.0 947250.0 105300.0 937950.0 ;
      RECT  101700.0 937950.0 102900.0 936750.0 ;
      RECT  104100.0 937950.0 105300.0 936750.0 ;
      RECT  104100.0 937950.0 105300.0 936750.0 ;
      RECT  101700.0 937950.0 102900.0 936750.0 ;
      RECT  101700.0 947250.0 102900.0 946050.0 ;
      RECT  104100.0 947250.0 105300.0 946050.0 ;
      RECT  104100.0 947250.0 105300.0 946050.0 ;
      RECT  101700.0 947250.0 102900.0 946050.0 ;
      RECT  106500.0 937350.0 107700.0 936150.0 ;
      RECT  106500.0 947250.0 107700.0 946050.0 ;
      RECT  102300.0 942600.0 103500.0 941400.0 ;
      RECT  102300.0 942600.0 103500.0 941400.0 ;
      RECT  104850.0 942450.0 105750.0 941550.0 ;
      RECT  99900.0 935250.0 109500.0 934350.0 ;
      RECT  99900.0 949050.0 109500.0 948150.0 ;
      RECT  106500.0 960450.0 107700.0 962400.0 ;
      RECT  106500.0 948600.0 107700.0 950550.0 ;
      RECT  101700.0 949950.0 102900.0 948150.0 ;
      RECT  101700.0 959250.0 102900.0 962850.0 ;
      RECT  104400.0 949950.0 105300.0 959250.0 ;
      RECT  101700.0 959250.0 102900.0 960450.0 ;
      RECT  104100.0 959250.0 105300.0 960450.0 ;
      RECT  104100.0 959250.0 105300.0 960450.0 ;
      RECT  101700.0 959250.0 102900.0 960450.0 ;
      RECT  101700.0 949950.0 102900.0 951150.0 ;
      RECT  104100.0 949950.0 105300.0 951150.0 ;
      RECT  104100.0 949950.0 105300.0 951150.0 ;
      RECT  101700.0 949950.0 102900.0 951150.0 ;
      RECT  106500.0 959850.0 107700.0 961050.0 ;
      RECT  106500.0 949950.0 107700.0 951150.0 ;
      RECT  102300.0 954600.0 103500.0 955800.0 ;
      RECT  102300.0 954600.0 103500.0 955800.0 ;
      RECT  104850.0 954750.0 105750.0 955650.0 ;
      RECT  99900.0 961950.0 109500.0 962850.0 ;
      RECT  99900.0 948150.0 109500.0 949050.0 ;
      RECT  106500.0 964350.0 107700.0 962400.0 ;
      RECT  106500.0 976200.0 107700.0 974250.0 ;
      RECT  101700.0 974850.0 102900.0 976650.0 ;
      RECT  101700.0 965550.0 102900.0 961950.0 ;
      RECT  104400.0 974850.0 105300.0 965550.0 ;
      RECT  101700.0 965550.0 102900.0 964350.0 ;
      RECT  104100.0 965550.0 105300.0 964350.0 ;
      RECT  104100.0 965550.0 105300.0 964350.0 ;
      RECT  101700.0 965550.0 102900.0 964350.0 ;
      RECT  101700.0 974850.0 102900.0 973650.0 ;
      RECT  104100.0 974850.0 105300.0 973650.0 ;
      RECT  104100.0 974850.0 105300.0 973650.0 ;
      RECT  101700.0 974850.0 102900.0 973650.0 ;
      RECT  106500.0 964950.0 107700.0 963750.0 ;
      RECT  106500.0 974850.0 107700.0 973650.0 ;
      RECT  102300.0 970200.0 103500.0 969000.0 ;
      RECT  102300.0 970200.0 103500.0 969000.0 ;
      RECT  104850.0 970050.0 105750.0 969150.0 ;
      RECT  99900.0 962850.0 109500.0 961950.0 ;
      RECT  99900.0 976650.0 109500.0 975750.0 ;
      RECT  106500.0 988050.0 107700.0 990000.0 ;
      RECT  106500.0 976200.0 107700.0 978150.0 ;
      RECT  101700.0 977550.0 102900.0 975750.0 ;
      RECT  101700.0 986850.0 102900.0 990450.0 ;
      RECT  104400.0 977550.0 105300.0 986850.0 ;
      RECT  101700.0 986850.0 102900.0 988050.0 ;
      RECT  104100.0 986850.0 105300.0 988050.0 ;
      RECT  104100.0 986850.0 105300.0 988050.0 ;
      RECT  101700.0 986850.0 102900.0 988050.0 ;
      RECT  101700.0 977550.0 102900.0 978750.0 ;
      RECT  104100.0 977550.0 105300.0 978750.0 ;
      RECT  104100.0 977550.0 105300.0 978750.0 ;
      RECT  101700.0 977550.0 102900.0 978750.0 ;
      RECT  106500.0 987450.0 107700.0 988650.0 ;
      RECT  106500.0 977550.0 107700.0 978750.0 ;
      RECT  102300.0 982200.0 103500.0 983400.0 ;
      RECT  102300.0 982200.0 103500.0 983400.0 ;
      RECT  104850.0 982350.0 105750.0 983250.0 ;
      RECT  99900.0 989550.0 109500.0 990450.0 ;
      RECT  99900.0 975750.0 109500.0 976650.0 ;
      RECT  106500.0 991950.0 107700.0 990000.0 ;
      RECT  106500.0 1003800.0 107700.0 1001850.0 ;
      RECT  101700.0 1002450.0 102900.0 1004250.0 ;
      RECT  101700.0 993150.0 102900.0 989550.0 ;
      RECT  104400.0 1002450.0 105300.0 993150.0 ;
      RECT  101700.0 993150.0 102900.0 991950.0 ;
      RECT  104100.0 993150.0 105300.0 991950.0 ;
      RECT  104100.0 993150.0 105300.0 991950.0 ;
      RECT  101700.0 993150.0 102900.0 991950.0 ;
      RECT  101700.0 1002450.0 102900.0 1001250.0 ;
      RECT  104100.0 1002450.0 105300.0 1001250.0 ;
      RECT  104100.0 1002450.0 105300.0 1001250.0 ;
      RECT  101700.0 1002450.0 102900.0 1001250.0 ;
      RECT  106500.0 992550.0 107700.0 991350.0 ;
      RECT  106500.0 1002450.0 107700.0 1001250.0 ;
      RECT  102300.0 997800.0 103500.0 996600.0 ;
      RECT  102300.0 997800.0 103500.0 996600.0 ;
      RECT  104850.0 997650.0 105750.0 996750.0 ;
      RECT  99900.0 990450.0 109500.0 989550.0 ;
      RECT  99900.0 1004250.0 109500.0 1003350.0 ;
      RECT  106500.0 1015650.0 107700.0 1017600.0 ;
      RECT  106500.0 1003800.0 107700.0 1005750.0 ;
      RECT  101700.0 1005150.0 102900.0 1003350.0 ;
      RECT  101700.0 1014450.0 102900.0 1018050.0 ;
      RECT  104400.0 1005150.0 105300.0 1014450.0 ;
      RECT  101700.0 1014450.0 102900.0 1015650.0 ;
      RECT  104100.0 1014450.0 105300.0 1015650.0 ;
      RECT  104100.0 1014450.0 105300.0 1015650.0 ;
      RECT  101700.0 1014450.0 102900.0 1015650.0 ;
      RECT  101700.0 1005150.0 102900.0 1006350.0 ;
      RECT  104100.0 1005150.0 105300.0 1006350.0 ;
      RECT  104100.0 1005150.0 105300.0 1006350.0 ;
      RECT  101700.0 1005150.0 102900.0 1006350.0 ;
      RECT  106500.0 1015050.0 107700.0 1016250.0 ;
      RECT  106500.0 1005150.0 107700.0 1006350.0 ;
      RECT  102300.0 1009800.0 103500.0 1011000.0 ;
      RECT  102300.0 1009800.0 103500.0 1011000.0 ;
      RECT  104850.0 1009950.0 105750.0 1010850.0 ;
      RECT  99900.0 1017150.0 109500.0 1018050.0 ;
      RECT  99900.0 1003350.0 109500.0 1004250.0 ;
      RECT  106500.0 1019550.0 107700.0 1017600.0 ;
      RECT  106500.0 1031400.0 107700.0 1029450.0 ;
      RECT  101700.0 1030050.0 102900.0 1031850.0 ;
      RECT  101700.0 1020750.0 102900.0 1017150.0 ;
      RECT  104400.0 1030050.0 105300.0 1020750.0 ;
      RECT  101700.0 1020750.0 102900.0 1019550.0 ;
      RECT  104100.0 1020750.0 105300.0 1019550.0 ;
      RECT  104100.0 1020750.0 105300.0 1019550.0 ;
      RECT  101700.0 1020750.0 102900.0 1019550.0 ;
      RECT  101700.0 1030050.0 102900.0 1028850.0 ;
      RECT  104100.0 1030050.0 105300.0 1028850.0 ;
      RECT  104100.0 1030050.0 105300.0 1028850.0 ;
      RECT  101700.0 1030050.0 102900.0 1028850.0 ;
      RECT  106500.0 1020150.0 107700.0 1018950.0 ;
      RECT  106500.0 1030050.0 107700.0 1028850.0 ;
      RECT  102300.0 1025400.0 103500.0 1024200.0 ;
      RECT  102300.0 1025400.0 103500.0 1024200.0 ;
      RECT  104850.0 1025250.0 105750.0 1024350.0 ;
      RECT  99900.0 1018050.0 109500.0 1017150.0 ;
      RECT  99900.0 1031850.0 109500.0 1030950.0 ;
      RECT  106500.0 1043250.0 107700.0 1045200.0 ;
      RECT  106500.0 1031400.0 107700.0 1033350.0 ;
      RECT  101700.0 1032750.0 102900.0 1030950.0 ;
      RECT  101700.0 1042050.0 102900.0 1045650.0 ;
      RECT  104400.0 1032750.0 105300.0 1042050.0 ;
      RECT  101700.0 1042050.0 102900.0 1043250.0 ;
      RECT  104100.0 1042050.0 105300.0 1043250.0 ;
      RECT  104100.0 1042050.0 105300.0 1043250.0 ;
      RECT  101700.0 1042050.0 102900.0 1043250.0 ;
      RECT  101700.0 1032750.0 102900.0 1033950.0 ;
      RECT  104100.0 1032750.0 105300.0 1033950.0 ;
      RECT  104100.0 1032750.0 105300.0 1033950.0 ;
      RECT  101700.0 1032750.0 102900.0 1033950.0 ;
      RECT  106500.0 1042650.0 107700.0 1043850.0 ;
      RECT  106500.0 1032750.0 107700.0 1033950.0 ;
      RECT  102300.0 1037400.0 103500.0 1038600.0 ;
      RECT  102300.0 1037400.0 103500.0 1038600.0 ;
      RECT  104850.0 1037550.0 105750.0 1038450.0 ;
      RECT  99900.0 1044750.0 109500.0 1045650.0 ;
      RECT  99900.0 1030950.0 109500.0 1031850.0 ;
      RECT  106500.0 1047150.0 107700.0 1045200.0 ;
      RECT  106500.0 1059000.0 107700.0 1057050.0 ;
      RECT  101700.0 1057650.0 102900.0 1059450.0 ;
      RECT  101700.0 1048350.0 102900.0 1044750.0 ;
      RECT  104400.0 1057650.0 105300.0 1048350.0 ;
      RECT  101700.0 1048350.0 102900.0 1047150.0 ;
      RECT  104100.0 1048350.0 105300.0 1047150.0 ;
      RECT  104100.0 1048350.0 105300.0 1047150.0 ;
      RECT  101700.0 1048350.0 102900.0 1047150.0 ;
      RECT  101700.0 1057650.0 102900.0 1056450.0 ;
      RECT  104100.0 1057650.0 105300.0 1056450.0 ;
      RECT  104100.0 1057650.0 105300.0 1056450.0 ;
      RECT  101700.0 1057650.0 102900.0 1056450.0 ;
      RECT  106500.0 1047750.0 107700.0 1046550.0 ;
      RECT  106500.0 1057650.0 107700.0 1056450.0 ;
      RECT  102300.0 1053000.0 103500.0 1051800.0 ;
      RECT  102300.0 1053000.0 103500.0 1051800.0 ;
      RECT  104850.0 1052850.0 105750.0 1051950.0 ;
      RECT  99900.0 1045650.0 109500.0 1044750.0 ;
      RECT  99900.0 1059450.0 109500.0 1058550.0 ;
      RECT  106500.0 1070850.0 107700.0 1072800.0 ;
      RECT  106500.0 1059000.0 107700.0 1060950.0 ;
      RECT  101700.0 1060350.0 102900.0 1058550.0 ;
      RECT  101700.0 1069650.0 102900.0 1073250.0 ;
      RECT  104400.0 1060350.0 105300.0 1069650.0 ;
      RECT  101700.0 1069650.0 102900.0 1070850.0 ;
      RECT  104100.0 1069650.0 105300.0 1070850.0 ;
      RECT  104100.0 1069650.0 105300.0 1070850.0 ;
      RECT  101700.0 1069650.0 102900.0 1070850.0 ;
      RECT  101700.0 1060350.0 102900.0 1061550.0 ;
      RECT  104100.0 1060350.0 105300.0 1061550.0 ;
      RECT  104100.0 1060350.0 105300.0 1061550.0 ;
      RECT  101700.0 1060350.0 102900.0 1061550.0 ;
      RECT  106500.0 1070250.0 107700.0 1071450.0 ;
      RECT  106500.0 1060350.0 107700.0 1061550.0 ;
      RECT  102300.0 1065000.0 103500.0 1066200.0 ;
      RECT  102300.0 1065000.0 103500.0 1066200.0 ;
      RECT  104850.0 1065150.0 105750.0 1066050.0 ;
      RECT  99900.0 1072350.0 109500.0 1073250.0 ;
      RECT  99900.0 1058550.0 109500.0 1059450.0 ;
      RECT  106500.0 1074750.0 107700.0 1072800.0 ;
      RECT  106500.0 1086600.0 107700.0 1084650.0 ;
      RECT  101700.0 1085250.0 102900.0 1087050.0 ;
      RECT  101700.0 1075950.0 102900.0 1072350.0 ;
      RECT  104400.0 1085250.0 105300.0 1075950.0 ;
      RECT  101700.0 1075950.0 102900.0 1074750.0 ;
      RECT  104100.0 1075950.0 105300.0 1074750.0 ;
      RECT  104100.0 1075950.0 105300.0 1074750.0 ;
      RECT  101700.0 1075950.0 102900.0 1074750.0 ;
      RECT  101700.0 1085250.0 102900.0 1084050.0 ;
      RECT  104100.0 1085250.0 105300.0 1084050.0 ;
      RECT  104100.0 1085250.0 105300.0 1084050.0 ;
      RECT  101700.0 1085250.0 102900.0 1084050.0 ;
      RECT  106500.0 1075350.0 107700.0 1074150.0 ;
      RECT  106500.0 1085250.0 107700.0 1084050.0 ;
      RECT  102300.0 1080600.0 103500.0 1079400.0 ;
      RECT  102300.0 1080600.0 103500.0 1079400.0 ;
      RECT  104850.0 1080450.0 105750.0 1079550.0 ;
      RECT  99900.0 1073250.0 109500.0 1072350.0 ;
      RECT  99900.0 1087050.0 109500.0 1086150.0 ;
      RECT  106500.0 1098450.0 107700.0 1100400.0 ;
      RECT  106500.0 1086600.0 107700.0 1088550.0 ;
      RECT  101700.0 1087950.0 102900.0 1086150.0 ;
      RECT  101700.0 1097250.0 102900.0 1100850.0 ;
      RECT  104400.0 1087950.0 105300.0 1097250.0 ;
      RECT  101700.0 1097250.0 102900.0 1098450.0 ;
      RECT  104100.0 1097250.0 105300.0 1098450.0 ;
      RECT  104100.0 1097250.0 105300.0 1098450.0 ;
      RECT  101700.0 1097250.0 102900.0 1098450.0 ;
      RECT  101700.0 1087950.0 102900.0 1089150.0 ;
      RECT  104100.0 1087950.0 105300.0 1089150.0 ;
      RECT  104100.0 1087950.0 105300.0 1089150.0 ;
      RECT  101700.0 1087950.0 102900.0 1089150.0 ;
      RECT  106500.0 1097850.0 107700.0 1099050.0 ;
      RECT  106500.0 1087950.0 107700.0 1089150.0 ;
      RECT  102300.0 1092600.0 103500.0 1093800.0 ;
      RECT  102300.0 1092600.0 103500.0 1093800.0 ;
      RECT  104850.0 1092750.0 105750.0 1093650.0 ;
      RECT  99900.0 1099950.0 109500.0 1100850.0 ;
      RECT  99900.0 1086150.0 109500.0 1087050.0 ;
      RECT  106500.0 1102350.0 107700.0 1100400.0 ;
      RECT  106500.0 1114200.0 107700.0 1112250.0 ;
      RECT  101700.0 1112850.0 102900.0 1114650.0 ;
      RECT  101700.0 1103550.0 102900.0 1099950.0 ;
      RECT  104400.0 1112850.0 105300.0 1103550.0 ;
      RECT  101700.0 1103550.0 102900.0 1102350.0 ;
      RECT  104100.0 1103550.0 105300.0 1102350.0 ;
      RECT  104100.0 1103550.0 105300.0 1102350.0 ;
      RECT  101700.0 1103550.0 102900.0 1102350.0 ;
      RECT  101700.0 1112850.0 102900.0 1111650.0 ;
      RECT  104100.0 1112850.0 105300.0 1111650.0 ;
      RECT  104100.0 1112850.0 105300.0 1111650.0 ;
      RECT  101700.0 1112850.0 102900.0 1111650.0 ;
      RECT  106500.0 1102950.0 107700.0 1101750.0 ;
      RECT  106500.0 1112850.0 107700.0 1111650.0 ;
      RECT  102300.0 1108200.0 103500.0 1107000.0 ;
      RECT  102300.0 1108200.0 103500.0 1107000.0 ;
      RECT  104850.0 1108050.0 105750.0 1107150.0 ;
      RECT  99900.0 1100850.0 109500.0 1099950.0 ;
      RECT  99900.0 1114650.0 109500.0 1113750.0 ;
      RECT  106500.0 1126050.0 107700.0 1128000.0 ;
      RECT  106500.0 1114200.0 107700.0 1116150.0 ;
      RECT  101700.0 1115550.0 102900.0 1113750.0 ;
      RECT  101700.0 1124850.0 102900.0 1128450.0 ;
      RECT  104400.0 1115550.0 105300.0 1124850.0 ;
      RECT  101700.0 1124850.0 102900.0 1126050.0 ;
      RECT  104100.0 1124850.0 105300.0 1126050.0 ;
      RECT  104100.0 1124850.0 105300.0 1126050.0 ;
      RECT  101700.0 1124850.0 102900.0 1126050.0 ;
      RECT  101700.0 1115550.0 102900.0 1116750.0 ;
      RECT  104100.0 1115550.0 105300.0 1116750.0 ;
      RECT  104100.0 1115550.0 105300.0 1116750.0 ;
      RECT  101700.0 1115550.0 102900.0 1116750.0 ;
      RECT  106500.0 1125450.0 107700.0 1126650.0 ;
      RECT  106500.0 1115550.0 107700.0 1116750.0 ;
      RECT  102300.0 1120200.0 103500.0 1121400.0 ;
      RECT  102300.0 1120200.0 103500.0 1121400.0 ;
      RECT  104850.0 1120350.0 105750.0 1121250.0 ;
      RECT  99900.0 1127550.0 109500.0 1128450.0 ;
      RECT  99900.0 1113750.0 109500.0 1114650.0 ;
      RECT  106500.0 1129950.0 107700.0 1128000.0 ;
      RECT  106500.0 1141800.0 107700.0 1139850.0 ;
      RECT  101700.0 1140450.0 102900.0 1142250.0 ;
      RECT  101700.0 1131150.0 102900.0 1127550.0 ;
      RECT  104400.0 1140450.0 105300.0 1131150.0 ;
      RECT  101700.0 1131150.0 102900.0 1129950.0 ;
      RECT  104100.0 1131150.0 105300.0 1129950.0 ;
      RECT  104100.0 1131150.0 105300.0 1129950.0 ;
      RECT  101700.0 1131150.0 102900.0 1129950.0 ;
      RECT  101700.0 1140450.0 102900.0 1139250.0 ;
      RECT  104100.0 1140450.0 105300.0 1139250.0 ;
      RECT  104100.0 1140450.0 105300.0 1139250.0 ;
      RECT  101700.0 1140450.0 102900.0 1139250.0 ;
      RECT  106500.0 1130550.0 107700.0 1129350.0 ;
      RECT  106500.0 1140450.0 107700.0 1139250.0 ;
      RECT  102300.0 1135800.0 103500.0 1134600.0 ;
      RECT  102300.0 1135800.0 103500.0 1134600.0 ;
      RECT  104850.0 1135650.0 105750.0 1134750.0 ;
      RECT  99900.0 1128450.0 109500.0 1127550.0 ;
      RECT  99900.0 1142250.0 109500.0 1141350.0 ;
      RECT  106500.0 1153650.0 107700.0 1155600.0 ;
      RECT  106500.0 1141800.0 107700.0 1143750.0 ;
      RECT  101700.0 1143150.0 102900.0 1141350.0 ;
      RECT  101700.0 1152450.0 102900.0 1156050.0 ;
      RECT  104400.0 1143150.0 105300.0 1152450.0 ;
      RECT  101700.0 1152450.0 102900.0 1153650.0 ;
      RECT  104100.0 1152450.0 105300.0 1153650.0 ;
      RECT  104100.0 1152450.0 105300.0 1153650.0 ;
      RECT  101700.0 1152450.0 102900.0 1153650.0 ;
      RECT  101700.0 1143150.0 102900.0 1144350.0 ;
      RECT  104100.0 1143150.0 105300.0 1144350.0 ;
      RECT  104100.0 1143150.0 105300.0 1144350.0 ;
      RECT  101700.0 1143150.0 102900.0 1144350.0 ;
      RECT  106500.0 1153050.0 107700.0 1154250.0 ;
      RECT  106500.0 1143150.0 107700.0 1144350.0 ;
      RECT  102300.0 1147800.0 103500.0 1149000.0 ;
      RECT  102300.0 1147800.0 103500.0 1149000.0 ;
      RECT  104850.0 1147950.0 105750.0 1148850.0 ;
      RECT  99900.0 1155150.0 109500.0 1156050.0 ;
      RECT  99900.0 1141350.0 109500.0 1142250.0 ;
      RECT  106500.0 1157550.0 107700.0 1155600.0 ;
      RECT  106500.0 1169400.0 107700.0 1167450.0 ;
      RECT  101700.0 1168050.0 102900.0 1169850.0 ;
      RECT  101700.0 1158750.0 102900.0 1155150.0 ;
      RECT  104400.0 1168050.0 105300.0 1158750.0 ;
      RECT  101700.0 1158750.0 102900.0 1157550.0 ;
      RECT  104100.0 1158750.0 105300.0 1157550.0 ;
      RECT  104100.0 1158750.0 105300.0 1157550.0 ;
      RECT  101700.0 1158750.0 102900.0 1157550.0 ;
      RECT  101700.0 1168050.0 102900.0 1166850.0 ;
      RECT  104100.0 1168050.0 105300.0 1166850.0 ;
      RECT  104100.0 1168050.0 105300.0 1166850.0 ;
      RECT  101700.0 1168050.0 102900.0 1166850.0 ;
      RECT  106500.0 1158150.0 107700.0 1156950.0 ;
      RECT  106500.0 1168050.0 107700.0 1166850.0 ;
      RECT  102300.0 1163400.0 103500.0 1162200.0 ;
      RECT  102300.0 1163400.0 103500.0 1162200.0 ;
      RECT  104850.0 1163250.0 105750.0 1162350.0 ;
      RECT  99900.0 1156050.0 109500.0 1155150.0 ;
      RECT  99900.0 1169850.0 109500.0 1168950.0 ;
      RECT  106500.0 1181250.0 107700.0 1183200.0 ;
      RECT  106500.0 1169400.0 107700.0 1171350.0 ;
      RECT  101700.0 1170750.0 102900.0 1168950.0 ;
      RECT  101700.0 1180050.0 102900.0 1183650.0 ;
      RECT  104400.0 1170750.0 105300.0 1180050.0 ;
      RECT  101700.0 1180050.0 102900.0 1181250.0 ;
      RECT  104100.0 1180050.0 105300.0 1181250.0 ;
      RECT  104100.0 1180050.0 105300.0 1181250.0 ;
      RECT  101700.0 1180050.0 102900.0 1181250.0 ;
      RECT  101700.0 1170750.0 102900.0 1171950.0 ;
      RECT  104100.0 1170750.0 105300.0 1171950.0 ;
      RECT  104100.0 1170750.0 105300.0 1171950.0 ;
      RECT  101700.0 1170750.0 102900.0 1171950.0 ;
      RECT  106500.0 1180650.0 107700.0 1181850.0 ;
      RECT  106500.0 1170750.0 107700.0 1171950.0 ;
      RECT  102300.0 1175400.0 103500.0 1176600.0 ;
      RECT  102300.0 1175400.0 103500.0 1176600.0 ;
      RECT  104850.0 1175550.0 105750.0 1176450.0 ;
      RECT  99900.0 1182750.0 109500.0 1183650.0 ;
      RECT  99900.0 1168950.0 109500.0 1169850.0 ;
      RECT  106500.0 1185150.0 107700.0 1183200.0 ;
      RECT  106500.0 1197000.0 107700.0 1195050.0 ;
      RECT  101700.0 1195650.0 102900.0 1197450.0 ;
      RECT  101700.0 1186350.0 102900.0 1182750.0 ;
      RECT  104400.0 1195650.0 105300.0 1186350.0 ;
      RECT  101700.0 1186350.0 102900.0 1185150.0 ;
      RECT  104100.0 1186350.0 105300.0 1185150.0 ;
      RECT  104100.0 1186350.0 105300.0 1185150.0 ;
      RECT  101700.0 1186350.0 102900.0 1185150.0 ;
      RECT  101700.0 1195650.0 102900.0 1194450.0 ;
      RECT  104100.0 1195650.0 105300.0 1194450.0 ;
      RECT  104100.0 1195650.0 105300.0 1194450.0 ;
      RECT  101700.0 1195650.0 102900.0 1194450.0 ;
      RECT  106500.0 1185750.0 107700.0 1184550.0 ;
      RECT  106500.0 1195650.0 107700.0 1194450.0 ;
      RECT  102300.0 1191000.0 103500.0 1189800.0 ;
      RECT  102300.0 1191000.0 103500.0 1189800.0 ;
      RECT  104850.0 1190850.0 105750.0 1189950.0 ;
      RECT  99900.0 1183650.0 109500.0 1182750.0 ;
      RECT  99900.0 1197450.0 109500.0 1196550.0 ;
      RECT  60150.0 154200.0 58950.0 155400.0 ;
      RECT  62250.0 168600.0 61050.0 169800.0 ;
      RECT  64350.0 181800.0 63150.0 183000.0 ;
      RECT  66450.0 196200.0 65250.0 197400.0 ;
      RECT  68550.0 209400.0 67350.0 210600.0 ;
      RECT  70650.0 223800.0 69450.0 225000.0 ;
      RECT  72750.0 237000.0 71550.0 238200.0 ;
      RECT  74850.0 251400.0 73650.0 252600.0 ;
      RECT  76950.0 264600.0 75750.0 265800.0 ;
      RECT  79050.0 279000.0 77850.0 280200.0 ;
      RECT  81150.0 292200.0 79950.0 293400.0 ;
      RECT  83250.0 306600.0 82050.0 307800.0 ;
      RECT  60150.0 321750.0 58950.0 322950.0 ;
      RECT  68550.0 319800.0 67350.0 321000.0 ;
      RECT  76950.0 317850.0 75750.0 319050.0 ;
      RECT  60150.0 332250.0 58950.0 333450.0 ;
      RECT  68550.0 334200.0 67350.0 335400.0 ;
      RECT  79050.0 336150.0 77850.0 337350.0 ;
      RECT  60150.0 349350.0 58950.0 350550.0 ;
      RECT  68550.0 347400.0 67350.0 348600.0 ;
      RECT  81150.0 345450.0 79950.0 346650.0 ;
      RECT  60150.0 359850.0 58950.0 361050.0 ;
      RECT  68550.0 361800.0 67350.0 363000.0 ;
      RECT  83250.0 363750.0 82050.0 364950.0 ;
      RECT  60150.0 376950.0 58950.0 378150.0 ;
      RECT  70650.0 375000.0 69450.0 376200.0 ;
      RECT  76950.0 373050.0 75750.0 374250.0 ;
      RECT  60150.0 387450.0 58950.0 388650.0 ;
      RECT  70650.0 389400.0 69450.0 390600.0 ;
      RECT  79050.0 391350.0 77850.0 392550.0 ;
      RECT  60150.0 404550.0 58950.0 405750.0 ;
      RECT  70650.0 402600.0 69450.0 403800.0 ;
      RECT  81150.0 400650.0 79950.0 401850.0 ;
      RECT  60150.0 415050.0 58950.0 416250.0 ;
      RECT  70650.0 417000.0 69450.0 418200.0 ;
      RECT  83250.0 418950.0 82050.0 420150.0 ;
      RECT  60150.0 432150.0 58950.0 433350.0 ;
      RECT  72750.0 430200.0 71550.0 431400.0 ;
      RECT  76950.0 428250.0 75750.0 429450.0 ;
      RECT  60150.0 442650.0 58950.0 443850.0 ;
      RECT  72750.0 444600.0 71550.0 445800.0 ;
      RECT  79050.0 446550.0 77850.0 447750.0 ;
      RECT  60150.0 459750.0 58950.0 460950.0 ;
      RECT  72750.0 457800.0 71550.0 459000.0 ;
      RECT  81150.0 455850.0 79950.0 457050.0 ;
      RECT  60150.0 470250.0 58950.0 471450.0 ;
      RECT  72750.0 472200.0 71550.0 473400.0 ;
      RECT  83250.0 474150.0 82050.0 475350.0 ;
      RECT  60150.0 487350.0 58950.0 488550.0 ;
      RECT  74850.0 485400.0 73650.0 486600.0 ;
      RECT  76950.0 483450.0 75750.0 484650.0 ;
      RECT  60150.0 497850.0 58950.0 499050.0 ;
      RECT  74850.0 499800.0 73650.0 501000.0 ;
      RECT  79050.0 501750.0 77850.0 502950.0 ;
      RECT  60150.0 514950.0 58950.0 516150.0 ;
      RECT  74850.0 513000.0 73650.0 514200.0 ;
      RECT  81150.0 511050.0 79950.0 512250.0 ;
      RECT  60150.0 525450.0 58950.0 526650.0 ;
      RECT  74850.0 527400.0 73650.0 528600.0 ;
      RECT  83250.0 529350.0 82050.0 530550.0 ;
      RECT  62250.0 542550.0 61050.0 543750.0 ;
      RECT  68550.0 540600.0 67350.0 541800.0 ;
      RECT  76950.0 538650.0 75750.0 539850.0 ;
      RECT  62250.0 553050.0 61050.0 554250.0 ;
      RECT  68550.0 555000.0 67350.0 556200.0 ;
      RECT  79050.0 556950.0 77850.0 558150.0 ;
      RECT  62250.0 570150.0 61050.0 571350.0 ;
      RECT  68550.0 568200.0 67350.0 569400.0 ;
      RECT  81150.0 566250.0 79950.0 567450.0 ;
      RECT  62250.0 580650.0 61050.0 581850.0 ;
      RECT  68550.0 582600.0 67350.0 583800.0 ;
      RECT  83250.0 584550.0 82050.0 585750.0 ;
      RECT  62250.0 597750.0 61050.0 598950.0 ;
      RECT  70650.0 595800.0 69450.0 597000.0 ;
      RECT  76950.0 593850.0 75750.0 595050.0 ;
      RECT  62250.0 608250.0 61050.0 609450.0 ;
      RECT  70650.0 610200.0 69450.0 611400.0 ;
      RECT  79050.0 612150.0 77850.0 613350.0 ;
      RECT  62250.0 625350.0 61050.0 626550.0 ;
      RECT  70650.0 623400.0 69450.0 624600.0 ;
      RECT  81150.0 621450.0 79950.0 622650.0 ;
      RECT  62250.0 635850.0 61050.0 637050.0 ;
      RECT  70650.0 637800.0 69450.0 639000.0 ;
      RECT  83250.0 639750.0 82050.0 640950.0 ;
      RECT  62250.0 652950.0 61050.0 654150.0 ;
      RECT  72750.0 651000.0 71550.0 652200.0 ;
      RECT  76950.0 649050.0 75750.0 650250.0 ;
      RECT  62250.0 663450.0 61050.0 664650.0 ;
      RECT  72750.0 665400.0 71550.0 666600.0 ;
      RECT  79050.0 667350.0 77850.0 668550.0 ;
      RECT  62250.0 680550.0 61050.0 681750.0 ;
      RECT  72750.0 678600.0 71550.0 679800.0 ;
      RECT  81150.0 676650.0 79950.0 677850.0 ;
      RECT  62250.0 691050.0 61050.0 692250.0 ;
      RECT  72750.0 693000.0 71550.0 694200.0 ;
      RECT  83250.0 694950.0 82050.0 696150.0 ;
      RECT  62250.0 708150.0 61050.0 709350.0 ;
      RECT  74850.0 706200.0 73650.0 707400.0 ;
      RECT  76950.0 704250.0 75750.0 705450.0 ;
      RECT  62250.0 718650.0 61050.0 719850.0 ;
      RECT  74850.0 720600.0 73650.0 721800.0 ;
      RECT  79050.0 722550.0 77850.0 723750.0 ;
      RECT  62250.0 735750.0 61050.0 736950.0 ;
      RECT  74850.0 733800.0 73650.0 735000.0 ;
      RECT  81150.0 731850.0 79950.0 733050.0 ;
      RECT  62250.0 746250.0 61050.0 747450.0 ;
      RECT  74850.0 748200.0 73650.0 749400.0 ;
      RECT  83250.0 750150.0 82050.0 751350.0 ;
      RECT  64350.0 763350.0 63150.0 764550.0 ;
      RECT  68550.0 761400.0 67350.0 762600.0 ;
      RECT  76950.0 759450.0 75750.0 760650.0 ;
      RECT  64350.0 773850.0 63150.0 775050.0 ;
      RECT  68550.0 775800.0 67350.0 777000.0 ;
      RECT  79050.0 777750.0 77850.0 778950.0 ;
      RECT  64350.0 790950.0 63150.0 792150.0 ;
      RECT  68550.0 789000.0 67350.0 790200.0 ;
      RECT  81150.0 787050.0 79950.0 788250.0 ;
      RECT  64350.0 801450.0 63150.0 802650.0 ;
      RECT  68550.0 803400.0 67350.0 804600.0 ;
      RECT  83250.0 805350.0 82050.0 806550.0 ;
      RECT  64350.0 818550.0 63150.0 819750.0 ;
      RECT  70650.0 816600.0 69450.0 817800.0 ;
      RECT  76950.0 814650.0 75750.0 815850.0 ;
      RECT  64350.0 829050.0 63150.0 830250.0 ;
      RECT  70650.0 831000.0 69450.0 832200.0 ;
      RECT  79050.0 832950.0 77850.0 834150.0 ;
      RECT  64350.0 846150.0 63150.0 847350.0 ;
      RECT  70650.0 844200.0 69450.0 845400.0 ;
      RECT  81150.0 842250.0 79950.0 843450.0 ;
      RECT  64350.0 856650.0 63150.0 857850.0 ;
      RECT  70650.0 858600.0 69450.0 859800.0 ;
      RECT  83250.0 860550.0 82050.0 861750.0 ;
      RECT  64350.0 873750.0 63150.0 874950.0 ;
      RECT  72750.0 871800.0 71550.0 873000.0 ;
      RECT  76950.0 869850.0 75750.0 871050.0 ;
      RECT  64350.0 884250.0 63150.0 885450.0 ;
      RECT  72750.0 886200.0 71550.0 887400.0 ;
      RECT  79050.0 888150.0 77850.0 889350.0 ;
      RECT  64350.0 901350.0 63150.0 902550.0 ;
      RECT  72750.0 899400.0 71550.0 900600.0 ;
      RECT  81150.0 897450.0 79950.0 898650.0 ;
      RECT  64350.0 911850.0 63150.0 913050.0 ;
      RECT  72750.0 913800.0 71550.0 915000.0 ;
      RECT  83250.0 915750.0 82050.0 916950.0 ;
      RECT  64350.0 928950.0 63150.0 930150.0 ;
      RECT  74850.0 927000.0 73650.0 928200.0 ;
      RECT  76950.0 925050.0 75750.0 926250.0 ;
      RECT  64350.0 939450.0 63150.0 940650.0 ;
      RECT  74850.0 941400.0 73650.0 942600.0 ;
      RECT  79050.0 943350.0 77850.0 944550.0 ;
      RECT  64350.0 956550.0 63150.0 957750.0 ;
      RECT  74850.0 954600.0 73650.0 955800.0 ;
      RECT  81150.0 952650.0 79950.0 953850.0 ;
      RECT  64350.0 967050.0 63150.0 968250.0 ;
      RECT  74850.0 969000.0 73650.0 970200.0 ;
      RECT  83250.0 970950.0 82050.0 972150.0 ;
      RECT  66450.0 984150.0 65250.0 985350.0 ;
      RECT  68550.0 982200.0 67350.0 983400.0 ;
      RECT  76950.0 980250.0 75750.0 981450.0 ;
      RECT  66450.0 994650.0 65250.0 995850.0 ;
      RECT  68550.0 996600.0 67350.0 997800.0 ;
      RECT  79050.0 998550.0 77850.0 999750.0 ;
      RECT  66450.0 1011750.0 65250.0 1012950.0 ;
      RECT  68550.0 1009800.0 67350.0 1011000.0 ;
      RECT  81150.0 1007850.0 79950.0 1009050.0 ;
      RECT  66450.0 1022250.0 65250.0 1023450.0 ;
      RECT  68550.0 1024200.0 67350.0 1025400.0 ;
      RECT  83250.0 1026150.0 82050.0 1027350.0 ;
      RECT  66450.0 1039350.0 65250.0 1040550.0 ;
      RECT  70650.0 1037400.0 69450.0 1038600.0 ;
      RECT  76950.0 1035450.0 75750.0 1036650.0 ;
      RECT  66450.0 1049850.0 65250.0 1051050.0 ;
      RECT  70650.0 1051800.0 69450.0 1053000.0 ;
      RECT  79050.0 1053750.0 77850.0 1054950.0 ;
      RECT  66450.0 1066950.0 65250.0 1068150.0 ;
      RECT  70650.0 1065000.0 69450.0 1066200.0 ;
      RECT  81150.0 1063050.0 79950.0 1064250.0 ;
      RECT  66450.0 1077450.0 65250.0 1078650.0 ;
      RECT  70650.0 1079400.0 69450.0 1080600.0 ;
      RECT  83250.0 1081350.0 82050.0 1082550.0 ;
      RECT  66450.0 1094550.0 65250.0 1095750.0 ;
      RECT  72750.0 1092600.0 71550.0 1093800.0 ;
      RECT  76950.0 1090650.0 75750.0 1091850.0 ;
      RECT  66450.0 1105050.0 65250.0 1106250.0 ;
      RECT  72750.0 1107000.0 71550.0 1108200.0 ;
      RECT  79050.0 1108950.0 77850.0 1110150.0 ;
      RECT  66450.0 1122150.0 65250.0 1123350.0 ;
      RECT  72750.0 1120200.0 71550.0 1121400.0 ;
      RECT  81150.0 1118250.0 79950.0 1119450.0 ;
      RECT  66450.0 1132650.0 65250.0 1133850.0 ;
      RECT  72750.0 1134600.0 71550.0 1135800.0 ;
      RECT  83250.0 1136550.0 82050.0 1137750.0 ;
      RECT  66450.0 1149750.0 65250.0 1150950.0 ;
      RECT  74850.0 1147800.0 73650.0 1149000.0 ;
      RECT  76950.0 1145850.0 75750.0 1147050.0 ;
      RECT  66450.0 1160250.0 65250.0 1161450.0 ;
      RECT  74850.0 1162200.0 73650.0 1163400.0 ;
      RECT  79050.0 1164150.0 77850.0 1165350.0 ;
      RECT  66450.0 1177350.0 65250.0 1178550.0 ;
      RECT  74850.0 1175400.0 73650.0 1176600.0 ;
      RECT  81150.0 1173450.0 79950.0 1174650.0 ;
      RECT  66450.0 1187850.0 65250.0 1189050.0 ;
      RECT  74850.0 1189800.0 73650.0 1191000.0 ;
      RECT  83250.0 1191750.0 82050.0 1192950.0 ;
      RECT  104850.0 319950.0 105750.0 320850.0 ;
      RECT  104850.0 334350.0 105750.0 335250.0 ;
      RECT  104850.0 347550.0 105750.0 348450.0 ;
      RECT  104850.0 361950.0 105750.0 362850.0 ;
      RECT  104850.0 375150.0 105750.0 376050.0 ;
      RECT  104850.0 389550.0 105750.0 390450.0 ;
      RECT  104850.0 402750.0 105750.0 403650.0 ;
      RECT  104850.0 417150.0 105750.0 418050.0 ;
      RECT  104850.0 430350.0 105750.0 431250.0 ;
      RECT  104850.0 444750.0 105750.0 445650.0 ;
      RECT  104850.0 457950.0 105750.0 458850.0 ;
      RECT  104850.0 472350.0 105750.0 473250.0 ;
      RECT  104850.0 485550.0 105750.0 486450.0 ;
      RECT  104850.0 499950.0 105750.0 500850.0 ;
      RECT  104850.0 513150.0 105750.0 514050.0 ;
      RECT  104850.0 527550.0 105750.0 528450.0 ;
      RECT  104850.0 540750.0 105750.0 541650.0 ;
      RECT  104850.0 555150.0 105750.0 556050.0 ;
      RECT  104850.0 568350.0 105750.0 569250.0 ;
      RECT  104850.0 582750.0 105750.0 583650.0 ;
      RECT  104850.0 595950.0 105750.0 596850.0 ;
      RECT  104850.0 610350.0 105750.0 611250.0 ;
      RECT  104850.0 623550.0 105750.0 624450.0 ;
      RECT  104850.0 637950.0 105750.0 638850.0 ;
      RECT  104850.0 651150.0 105750.0 652050.0 ;
      RECT  104850.0 665550.0 105750.0 666450.0 ;
      RECT  104850.0 678750.0 105750.0 679650.0 ;
      RECT  104850.0 693150.0 105750.0 694050.0 ;
      RECT  104850.0 706350.0 105750.0 707250.0 ;
      RECT  104850.0 720750.0 105750.0 721650.0 ;
      RECT  104850.0 733950.0 105750.0 734850.0 ;
      RECT  104850.0 748350.0 105750.0 749250.0 ;
      RECT  104850.0 761550.0 105750.0 762450.0 ;
      RECT  104850.0 775950.0 105750.0 776850.0 ;
      RECT  104850.0 789150.0 105750.0 790050.0 ;
      RECT  104850.0 803550.0 105750.0 804450.0 ;
      RECT  104850.0 816750.0 105750.0 817650.0 ;
      RECT  104850.0 831150.0 105750.0 832050.0 ;
      RECT  104850.0 844350.0 105750.0 845250.0 ;
      RECT  104850.0 858750.0 105750.0 859650.0 ;
      RECT  104850.0 871950.0 105750.0 872850.0 ;
      RECT  104850.0 886350.0 105750.0 887250.0 ;
      RECT  104850.0 899550.0 105750.0 900450.0 ;
      RECT  104850.0 913950.0 105750.0 914850.0 ;
      RECT  104850.0 927150.0 105750.0 928050.0 ;
      RECT  104850.0 941550.0 105750.0 942450.0 ;
      RECT  104850.0 954750.0 105750.0 955650.0 ;
      RECT  104850.0 969150.0 105750.0 970050.0 ;
      RECT  104850.0 982350.0 105750.0 983250.0 ;
      RECT  104850.0 996750.0 105750.0 997650.0 ;
      RECT  104850.0 1009950.0 105750.0 1010850.0 ;
      RECT  104850.0 1024350.0 105750.0 1025250.0 ;
      RECT  104850.0 1037550.0 105750.0 1038450.0 ;
      RECT  104850.0 1051950.0 105750.0 1052850.0 ;
      RECT  104850.0 1065150.0 105750.0 1066050.0 ;
      RECT  104850.0 1079550.0 105750.0 1080450.0 ;
      RECT  104850.0 1092750.0 105750.0 1093650.0 ;
      RECT  104850.0 1107150.0 105750.0 1108050.0 ;
      RECT  104850.0 1120350.0 105750.0 1121250.0 ;
      RECT  104850.0 1134750.0 105750.0 1135650.0 ;
      RECT  104850.0 1147950.0 105750.0 1148850.0 ;
      RECT  104850.0 1162350.0 105750.0 1163250.0 ;
      RECT  104850.0 1175550.0 105750.0 1176450.0 ;
      RECT  104850.0 1189950.0 105750.0 1190850.0 ;
      RECT  59100.0 161550.0 138900.0 162450.0 ;
      RECT  59100.0 189150.0 138900.0 190050.0 ;
      RECT  59100.0 216750.0 138900.0 217650.0 ;
      RECT  59100.0 244350.0 138900.0 245250.0 ;
      RECT  59100.0 271950.0 138900.0 272850.0 ;
      RECT  59100.0 299550.0 138900.0 300450.0 ;
      RECT  59100.0 327150.0 138900.0 328050.0 ;
      RECT  59100.0 354750.0 138900.0 355650.0 ;
      RECT  59100.0 382350.0 138900.0 383250.0 ;
      RECT  59100.0 409950.0 138900.0 410850.0 ;
      RECT  59100.0 437550.0 138900.0 438450.0 ;
      RECT  59100.0 465150.0 138900.0 466050.0 ;
      RECT  59100.0 492750.0 138900.0 493650.0 ;
      RECT  59100.0 520350.0 138900.0 521250.0 ;
      RECT  59100.0 547950.0 138900.0 548850.0 ;
      RECT  59100.0 575550.0 138900.0 576450.0 ;
      RECT  59100.0 603150.0 138900.0 604050.0 ;
      RECT  59100.0 630750.0 138900.0 631650.0 ;
      RECT  59100.0 658350.0 138900.0 659250.0 ;
      RECT  59100.0 685950.0 138900.0 686850.0 ;
      RECT  59100.0 713550.0 138900.0 714450.0 ;
      RECT  59100.0 741150.0 138900.0 742050.0 ;
      RECT  59100.0 768750.0 138900.0 769650.0 ;
      RECT  59100.0 796350.0 138900.0 797250.0 ;
      RECT  59100.0 823950.0 138900.0 824850.0 ;
      RECT  59100.0 851550.0 138900.0 852450.0 ;
      RECT  59100.0 879150.0 138900.0 880050.0 ;
      RECT  59100.0 906750.0 138900.0 907650.0 ;
      RECT  59100.0 934350.0 138900.0 935250.0 ;
      RECT  59100.0 961950.0 138900.0 962850.0 ;
      RECT  59100.0 989550.0 138900.0 990450.0 ;
      RECT  59100.0 1017150.0 138900.0 1018050.0 ;
      RECT  59100.0 1044750.0 138900.0 1045650.0 ;
      RECT  59100.0 1072350.0 138900.0 1073250.0 ;
      RECT  59100.0 1099950.0 138900.0 1100850.0 ;
      RECT  59100.0 1127550.0 138900.0 1128450.0 ;
      RECT  59100.0 1155150.0 138900.0 1156050.0 ;
      RECT  59100.0 1182750.0 138900.0 1183650.0 ;
      RECT  59100.0 147750.0 138900.0 148650.0 ;
      RECT  59100.0 175350.0 138900.0 176250.0 ;
      RECT  59100.0 202950.0 138900.0 203850.0 ;
      RECT  59100.0 230550.0 138900.0 231450.0 ;
      RECT  59100.0 258150.0 138900.0 259050.0 ;
      RECT  59100.0 285750.0 138900.0 286650.0 ;
      RECT  59100.0 313350.0 138900.0 314250.0 ;
      RECT  59100.0 340950.0 138900.0 341850.0 ;
      RECT  59100.0 368550.0 138900.0 369450.0 ;
      RECT  59100.0 396150.0 138900.0 397050.0 ;
      RECT  59100.0 423750.0 138900.0 424650.0 ;
      RECT  59100.0 451350.0 138900.0 452250.0 ;
      RECT  59100.0 478950.0 138900.0 479850.0 ;
      RECT  59100.0 506550.0 138900.0 507450.0 ;
      RECT  59100.0 534150.0 138900.0 535050.0 ;
      RECT  59100.0 561750.0 138900.0 562650.0 ;
      RECT  59100.0 589350.0 138900.0 590250.0 ;
      RECT  59100.0 616950.0 138900.0 617850.0 ;
      RECT  59100.0 644550.0 138900.0 645450.0 ;
      RECT  59100.0 672150.0 138900.0 673050.0 ;
      RECT  59100.0 699750.0 138900.0 700650.0 ;
      RECT  59100.0 727350.0 138900.0 728250.0 ;
      RECT  59100.0 754950.0 138900.0 755850.0 ;
      RECT  59100.0 782550.0 138900.0 783450.0 ;
      RECT  59100.0 810150.0 138900.0 811050.0 ;
      RECT  59100.0 837750.0 138900.0 838650.0 ;
      RECT  59100.0 865350.0 138900.0 866250.0 ;
      RECT  59100.0 892950.0 138900.0 893850.0 ;
      RECT  59100.0 920550.0 138900.0 921450.0 ;
      RECT  59100.0 948150.0 138900.0 949050.0 ;
      RECT  59100.0 975750.0 138900.0 976650.0 ;
      RECT  59100.0 1003350.0 138900.0 1004250.0 ;
      RECT  59100.0 1030950.0 138900.0 1031850.0 ;
      RECT  59100.0 1058550.0 138900.0 1059450.0 ;
      RECT  59100.0 1086150.0 138900.0 1087050.0 ;
      RECT  59100.0 1113750.0 138900.0 1114650.0 ;
      RECT  59100.0 1141350.0 138900.0 1142250.0 ;
      RECT  59100.0 1168950.0 138900.0 1169850.0 ;
      RECT  59100.0 1196550.0 138900.0 1197450.0 ;
      RECT  112650.0 319950.0 118200.0 320850.0 ;
      RECT  120750.0 321150.0 121650.0 322050.0 ;
      RECT  120750.0 319950.0 121650.0 320850.0 ;
      RECT  120750.0 320850.0 121650.0 321600.0 ;
      RECT  121200.0 321150.0 127800.0 322050.0 ;
      RECT  127800.0 321150.0 129000.0 322050.0 ;
      RECT  137250.0 321150.0 138150.0 322050.0 ;
      RECT  137250.0 319950.0 138150.0 320850.0 ;
      RECT  133200.0 321150.0 137700.0 322050.0 ;
      RECT  137250.0 320400.0 138150.0 321600.0 ;
      RECT  137700.0 319950.0 142200.0 320850.0 ;
      RECT  112650.0 334350.0 118200.0 335250.0 ;
      RECT  120750.0 333150.0 121650.0 334050.0 ;
      RECT  120750.0 334350.0 121650.0 335250.0 ;
      RECT  120750.0 333600.0 121650.0 335250.0 ;
      RECT  121200.0 333150.0 127800.0 334050.0 ;
      RECT  127800.0 333150.0 129000.0 334050.0 ;
      RECT  137250.0 333150.0 138150.0 334050.0 ;
      RECT  137250.0 334350.0 138150.0 335250.0 ;
      RECT  133200.0 333150.0 137700.0 334050.0 ;
      RECT  137250.0 333600.0 138150.0 334800.0 ;
      RECT  137700.0 334350.0 142200.0 335250.0 ;
      RECT  112650.0 347550.0 118200.0 348450.0 ;
      RECT  120750.0 348750.0 121650.0 349650.0 ;
      RECT  120750.0 347550.0 121650.0 348450.0 ;
      RECT  120750.0 348450.0 121650.0 349200.0 ;
      RECT  121200.0 348750.0 127800.0 349650.0 ;
      RECT  127800.0 348750.0 129000.0 349650.0 ;
      RECT  137250.0 348750.0 138150.0 349650.0 ;
      RECT  137250.0 347550.0 138150.0 348450.0 ;
      RECT  133200.0 348750.0 137700.0 349650.0 ;
      RECT  137250.0 348000.0 138150.0 349200.0 ;
      RECT  137700.0 347550.0 142200.0 348450.0 ;
      RECT  112650.0 361950.0 118200.0 362850.0 ;
      RECT  120750.0 360750.0 121650.0 361650.0 ;
      RECT  120750.0 361950.0 121650.0 362850.0 ;
      RECT  120750.0 361200.0 121650.0 362850.0 ;
      RECT  121200.0 360750.0 127800.0 361650.0 ;
      RECT  127800.0 360750.0 129000.0 361650.0 ;
      RECT  137250.0 360750.0 138150.0 361650.0 ;
      RECT  137250.0 361950.0 138150.0 362850.0 ;
      RECT  133200.0 360750.0 137700.0 361650.0 ;
      RECT  137250.0 361200.0 138150.0 362400.0 ;
      RECT  137700.0 361950.0 142200.0 362850.0 ;
      RECT  112650.0 375150.0 118200.0 376050.0 ;
      RECT  120750.0 376350.0 121650.0 377250.0 ;
      RECT  120750.0 375150.0 121650.0 376050.0 ;
      RECT  120750.0 376050.0 121650.0 376800.0 ;
      RECT  121200.0 376350.0 127800.0 377250.0 ;
      RECT  127800.0 376350.0 129000.0 377250.0 ;
      RECT  137250.0 376350.0 138150.0 377250.0 ;
      RECT  137250.0 375150.0 138150.0 376050.0 ;
      RECT  133200.0 376350.0 137700.0 377250.0 ;
      RECT  137250.0 375600.0 138150.0 376800.0 ;
      RECT  137700.0 375150.0 142200.0 376050.0 ;
      RECT  112650.0 389550.0 118200.0 390450.0 ;
      RECT  120750.0 388350.0 121650.0 389250.0 ;
      RECT  120750.0 389550.0 121650.0 390450.0 ;
      RECT  120750.0 388800.0 121650.0 390450.0 ;
      RECT  121200.0 388350.0 127800.0 389250.0 ;
      RECT  127800.0 388350.0 129000.0 389250.0 ;
      RECT  137250.0 388350.0 138150.0 389250.0 ;
      RECT  137250.0 389550.0 138150.0 390450.0 ;
      RECT  133200.0 388350.0 137700.0 389250.0 ;
      RECT  137250.0 388800.0 138150.0 390000.0 ;
      RECT  137700.0 389550.0 142200.0 390450.0 ;
      RECT  112650.0 402750.0 118200.0 403650.0 ;
      RECT  120750.0 403950.0 121650.0 404850.0 ;
      RECT  120750.0 402750.0 121650.0 403650.0 ;
      RECT  120750.0 403650.0 121650.0 404400.0 ;
      RECT  121200.0 403950.0 127800.0 404850.0 ;
      RECT  127800.0 403950.0 129000.0 404850.0 ;
      RECT  137250.0 403950.0 138150.0 404850.0 ;
      RECT  137250.0 402750.0 138150.0 403650.0 ;
      RECT  133200.0 403950.0 137700.0 404850.0 ;
      RECT  137250.0 403200.0 138150.0 404400.0 ;
      RECT  137700.0 402750.0 142200.0 403650.0 ;
      RECT  112650.0 417150.0 118200.0 418050.0 ;
      RECT  120750.0 415950.0 121650.0 416850.0 ;
      RECT  120750.0 417150.0 121650.0 418050.0 ;
      RECT  120750.0 416400.0 121650.0 418050.0 ;
      RECT  121200.0 415950.0 127800.0 416850.0 ;
      RECT  127800.0 415950.0 129000.0 416850.0 ;
      RECT  137250.0 415950.0 138150.0 416850.0 ;
      RECT  137250.0 417150.0 138150.0 418050.0 ;
      RECT  133200.0 415950.0 137700.0 416850.0 ;
      RECT  137250.0 416400.0 138150.0 417600.0 ;
      RECT  137700.0 417150.0 142200.0 418050.0 ;
      RECT  112650.0 430350.0 118200.0 431250.0 ;
      RECT  120750.0 431550.0 121650.0 432450.0 ;
      RECT  120750.0 430350.0 121650.0 431250.0 ;
      RECT  120750.0 431250.0 121650.0 432000.0 ;
      RECT  121200.0 431550.0 127800.0 432450.0 ;
      RECT  127800.0 431550.0 129000.0 432450.0 ;
      RECT  137250.0 431550.0 138150.0 432450.0 ;
      RECT  137250.0 430350.0 138150.0 431250.0 ;
      RECT  133200.0 431550.0 137700.0 432450.0 ;
      RECT  137250.0 430800.0 138150.0 432000.0 ;
      RECT  137700.0 430350.0 142200.0 431250.0 ;
      RECT  112650.0 444750.0 118200.0 445650.0 ;
      RECT  120750.0 443550.0 121650.0 444450.0 ;
      RECT  120750.0 444750.0 121650.0 445650.0 ;
      RECT  120750.0 444000.0 121650.0 445650.0 ;
      RECT  121200.0 443550.0 127800.0 444450.0 ;
      RECT  127800.0 443550.0 129000.0 444450.0 ;
      RECT  137250.0 443550.0 138150.0 444450.0 ;
      RECT  137250.0 444750.0 138150.0 445650.0 ;
      RECT  133200.0 443550.0 137700.0 444450.0 ;
      RECT  137250.0 444000.0 138150.0 445200.0 ;
      RECT  137700.0 444750.0 142200.0 445650.0 ;
      RECT  112650.0 457950.0 118200.0 458850.0 ;
      RECT  120750.0 459150.0 121650.0 460050.0 ;
      RECT  120750.0 457950.0 121650.0 458850.0 ;
      RECT  120750.0 458850.0 121650.0 459600.0 ;
      RECT  121200.0 459150.0 127800.0 460050.0 ;
      RECT  127800.0 459150.0 129000.0 460050.0 ;
      RECT  137250.0 459150.0 138150.0 460050.0 ;
      RECT  137250.0 457950.0 138150.0 458850.0 ;
      RECT  133200.0 459150.0 137700.0 460050.0 ;
      RECT  137250.0 458400.0 138150.0 459600.0 ;
      RECT  137700.0 457950.0 142200.0 458850.0 ;
      RECT  112650.0 472350.0 118200.0 473250.0 ;
      RECT  120750.0 471150.0 121650.0 472050.0 ;
      RECT  120750.0 472350.0 121650.0 473250.0 ;
      RECT  120750.0 471600.0 121650.0 473250.0 ;
      RECT  121200.0 471150.0 127800.0 472050.0 ;
      RECT  127800.0 471150.0 129000.0 472050.0 ;
      RECT  137250.0 471150.0 138150.0 472050.0 ;
      RECT  137250.0 472350.0 138150.0 473250.0 ;
      RECT  133200.0 471150.0 137700.0 472050.0 ;
      RECT  137250.0 471600.0 138150.0 472800.0 ;
      RECT  137700.0 472350.0 142200.0 473250.0 ;
      RECT  112650.0 485550.0 118200.0 486450.0 ;
      RECT  120750.0 486750.0 121650.0 487650.0 ;
      RECT  120750.0 485550.0 121650.0 486450.0 ;
      RECT  120750.0 486450.0 121650.0 487200.0 ;
      RECT  121200.0 486750.0 127800.0 487650.0 ;
      RECT  127800.0 486750.0 129000.0 487650.0 ;
      RECT  137250.0 486750.0 138150.0 487650.0 ;
      RECT  137250.0 485550.0 138150.0 486450.0 ;
      RECT  133200.0 486750.0 137700.0 487650.0 ;
      RECT  137250.0 486000.0 138150.0 487200.0 ;
      RECT  137700.0 485550.0 142200.0 486450.0 ;
      RECT  112650.0 499950.0 118200.0 500850.0 ;
      RECT  120750.0 498750.0 121650.0 499650.0 ;
      RECT  120750.0 499950.0 121650.0 500850.0 ;
      RECT  120750.0 499200.0 121650.0 500850.0 ;
      RECT  121200.0 498750.0 127800.0 499650.0 ;
      RECT  127800.0 498750.0 129000.0 499650.0 ;
      RECT  137250.0 498750.0 138150.0 499650.0 ;
      RECT  137250.0 499950.0 138150.0 500850.0 ;
      RECT  133200.0 498750.0 137700.0 499650.0 ;
      RECT  137250.0 499200.0 138150.0 500400.0 ;
      RECT  137700.0 499950.0 142200.0 500850.0 ;
      RECT  112650.0 513150.0 118200.0 514050.0 ;
      RECT  120750.0 514350.0 121650.0 515250.0 ;
      RECT  120750.0 513150.0 121650.0 514050.0 ;
      RECT  120750.0 514050.0 121650.0 514800.0 ;
      RECT  121200.0 514350.0 127800.0 515250.0 ;
      RECT  127800.0 514350.0 129000.0 515250.0 ;
      RECT  137250.0 514350.0 138150.0 515250.0 ;
      RECT  137250.0 513150.0 138150.0 514050.0 ;
      RECT  133200.0 514350.0 137700.0 515250.0 ;
      RECT  137250.0 513600.0 138150.0 514800.0 ;
      RECT  137700.0 513150.0 142200.0 514050.0 ;
      RECT  112650.0 527550.0 118200.0 528450.0 ;
      RECT  120750.0 526350.0 121650.0 527250.0 ;
      RECT  120750.0 527550.0 121650.0 528450.0 ;
      RECT  120750.0 526800.0 121650.0 528450.0 ;
      RECT  121200.0 526350.0 127800.0 527250.0 ;
      RECT  127800.0 526350.0 129000.0 527250.0 ;
      RECT  137250.0 526350.0 138150.0 527250.0 ;
      RECT  137250.0 527550.0 138150.0 528450.0 ;
      RECT  133200.0 526350.0 137700.0 527250.0 ;
      RECT  137250.0 526800.0 138150.0 528000.0 ;
      RECT  137700.0 527550.0 142200.0 528450.0 ;
      RECT  112650.0 540750.0 118200.0 541650.0 ;
      RECT  120750.0 541950.0 121650.0 542850.0 ;
      RECT  120750.0 540750.0 121650.0 541650.0 ;
      RECT  120750.0 541650.0 121650.0 542400.0 ;
      RECT  121200.0 541950.0 127800.0 542850.0 ;
      RECT  127800.0 541950.0 129000.0 542850.0 ;
      RECT  137250.0 541950.0 138150.0 542850.0 ;
      RECT  137250.0 540750.0 138150.0 541650.0 ;
      RECT  133200.0 541950.0 137700.0 542850.0 ;
      RECT  137250.0 541200.0 138150.0 542400.0 ;
      RECT  137700.0 540750.0 142200.0 541650.0 ;
      RECT  112650.0 555150.0 118200.0 556050.0 ;
      RECT  120750.0 553950.0 121650.0 554850.0 ;
      RECT  120750.0 555150.0 121650.0 556050.0 ;
      RECT  120750.0 554400.0 121650.0 556050.0 ;
      RECT  121200.0 553950.0 127800.0 554850.0 ;
      RECT  127800.0 553950.0 129000.0 554850.0 ;
      RECT  137250.0 553950.0 138150.0 554850.0 ;
      RECT  137250.0 555150.0 138150.0 556050.0 ;
      RECT  133200.0 553950.0 137700.0 554850.0 ;
      RECT  137250.0 554400.0 138150.0 555600.0 ;
      RECT  137700.0 555150.0 142200.0 556050.0 ;
      RECT  112650.0 568350.0 118200.0 569250.0 ;
      RECT  120750.0 569550.0 121650.0 570450.0 ;
      RECT  120750.0 568350.0 121650.0 569250.0 ;
      RECT  120750.0 569250.0 121650.0 570000.0 ;
      RECT  121200.0 569550.0 127800.0 570450.0 ;
      RECT  127800.0 569550.0 129000.0 570450.0 ;
      RECT  137250.0 569550.0 138150.0 570450.0 ;
      RECT  137250.0 568350.0 138150.0 569250.0 ;
      RECT  133200.0 569550.0 137700.0 570450.0 ;
      RECT  137250.0 568800.0 138150.0 570000.0 ;
      RECT  137700.0 568350.0 142200.0 569250.0 ;
      RECT  112650.0 582750.0 118200.0 583650.0 ;
      RECT  120750.0 581550.0 121650.0 582450.0 ;
      RECT  120750.0 582750.0 121650.0 583650.0 ;
      RECT  120750.0 582000.0 121650.0 583650.0 ;
      RECT  121200.0 581550.0 127800.0 582450.0 ;
      RECT  127800.0 581550.0 129000.0 582450.0 ;
      RECT  137250.0 581550.0 138150.0 582450.0 ;
      RECT  137250.0 582750.0 138150.0 583650.0 ;
      RECT  133200.0 581550.0 137700.0 582450.0 ;
      RECT  137250.0 582000.0 138150.0 583200.0 ;
      RECT  137700.0 582750.0 142200.0 583650.0 ;
      RECT  112650.0 595950.0 118200.0 596850.0 ;
      RECT  120750.0 597150.0 121650.0 598050.0 ;
      RECT  120750.0 595950.0 121650.0 596850.0 ;
      RECT  120750.0 596850.0 121650.0 597600.0 ;
      RECT  121200.0 597150.0 127800.0 598050.0 ;
      RECT  127800.0 597150.0 129000.0 598050.0 ;
      RECT  137250.0 597150.0 138150.0 598050.0 ;
      RECT  137250.0 595950.0 138150.0 596850.0 ;
      RECT  133200.0 597150.0 137700.0 598050.0 ;
      RECT  137250.0 596400.0 138150.0 597600.0 ;
      RECT  137700.0 595950.0 142200.0 596850.0 ;
      RECT  112650.0 610350.0 118200.0 611250.0 ;
      RECT  120750.0 609150.0 121650.0 610050.0 ;
      RECT  120750.0 610350.0 121650.0 611250.0 ;
      RECT  120750.0 609600.0 121650.0 611250.0 ;
      RECT  121200.0 609150.0 127800.0 610050.0 ;
      RECT  127800.0 609150.0 129000.0 610050.0 ;
      RECT  137250.0 609150.0 138150.0 610050.0 ;
      RECT  137250.0 610350.0 138150.0 611250.0 ;
      RECT  133200.0 609150.0 137700.0 610050.0 ;
      RECT  137250.0 609600.0 138150.0 610800.0 ;
      RECT  137700.0 610350.0 142200.0 611250.0 ;
      RECT  112650.0 623550.0 118200.0 624450.0 ;
      RECT  120750.0 624750.0 121650.0 625650.0 ;
      RECT  120750.0 623550.0 121650.0 624450.0 ;
      RECT  120750.0 624450.0 121650.0 625200.0 ;
      RECT  121200.0 624750.0 127800.0 625650.0 ;
      RECT  127800.0 624750.0 129000.0 625650.0 ;
      RECT  137250.0 624750.0 138150.0 625650.0 ;
      RECT  137250.0 623550.0 138150.0 624450.0 ;
      RECT  133200.0 624750.0 137700.0 625650.0 ;
      RECT  137250.0 624000.0 138150.0 625200.0 ;
      RECT  137700.0 623550.0 142200.0 624450.0 ;
      RECT  112650.0 637950.0 118200.0 638850.0 ;
      RECT  120750.0 636750.0 121650.0 637650.0 ;
      RECT  120750.0 637950.0 121650.0 638850.0 ;
      RECT  120750.0 637200.0 121650.0 638850.0 ;
      RECT  121200.0 636750.0 127800.0 637650.0 ;
      RECT  127800.0 636750.0 129000.0 637650.0 ;
      RECT  137250.0 636750.0 138150.0 637650.0 ;
      RECT  137250.0 637950.0 138150.0 638850.0 ;
      RECT  133200.0 636750.0 137700.0 637650.0 ;
      RECT  137250.0 637200.0 138150.0 638400.0 ;
      RECT  137700.0 637950.0 142200.0 638850.0 ;
      RECT  112650.0 651150.0 118200.0 652050.0 ;
      RECT  120750.0 652350.0 121650.0 653250.0 ;
      RECT  120750.0 651150.0 121650.0 652050.0 ;
      RECT  120750.0 652050.0 121650.0 652800.0 ;
      RECT  121200.0 652350.0 127800.0 653250.0 ;
      RECT  127800.0 652350.0 129000.0 653250.0 ;
      RECT  137250.0 652350.0 138150.0 653250.0 ;
      RECT  137250.0 651150.0 138150.0 652050.0 ;
      RECT  133200.0 652350.0 137700.0 653250.0 ;
      RECT  137250.0 651600.0 138150.0 652800.0 ;
      RECT  137700.0 651150.0 142200.0 652050.0 ;
      RECT  112650.0 665550.0 118200.0 666450.0 ;
      RECT  120750.0 664350.0 121650.0 665250.0 ;
      RECT  120750.0 665550.0 121650.0 666450.0 ;
      RECT  120750.0 664800.0 121650.0 666450.0 ;
      RECT  121200.0 664350.0 127800.0 665250.0 ;
      RECT  127800.0 664350.0 129000.0 665250.0 ;
      RECT  137250.0 664350.0 138150.0 665250.0 ;
      RECT  137250.0 665550.0 138150.0 666450.0 ;
      RECT  133200.0 664350.0 137700.0 665250.0 ;
      RECT  137250.0 664800.0 138150.0 666000.0 ;
      RECT  137700.0 665550.0 142200.0 666450.0 ;
      RECT  112650.0 678750.0 118200.0 679650.0 ;
      RECT  120750.0 679950.0 121650.0 680850.0 ;
      RECT  120750.0 678750.0 121650.0 679650.0 ;
      RECT  120750.0 679650.0 121650.0 680400.0 ;
      RECT  121200.0 679950.0 127800.0 680850.0 ;
      RECT  127800.0 679950.0 129000.0 680850.0 ;
      RECT  137250.0 679950.0 138150.0 680850.0 ;
      RECT  137250.0 678750.0 138150.0 679650.0 ;
      RECT  133200.0 679950.0 137700.0 680850.0 ;
      RECT  137250.0 679200.0 138150.0 680400.0 ;
      RECT  137700.0 678750.0 142200.0 679650.0 ;
      RECT  112650.0 693150.0 118200.0 694050.0 ;
      RECT  120750.0 691950.0 121650.0 692850.0 ;
      RECT  120750.0 693150.0 121650.0 694050.0 ;
      RECT  120750.0 692400.0 121650.0 694050.0 ;
      RECT  121200.0 691950.0 127800.0 692850.0 ;
      RECT  127800.0 691950.0 129000.0 692850.0 ;
      RECT  137250.0 691950.0 138150.0 692850.0 ;
      RECT  137250.0 693150.0 138150.0 694050.0 ;
      RECT  133200.0 691950.0 137700.0 692850.0 ;
      RECT  137250.0 692400.0 138150.0 693600.0 ;
      RECT  137700.0 693150.0 142200.0 694050.0 ;
      RECT  112650.0 706350.0 118200.0 707250.0 ;
      RECT  120750.0 707550.0 121650.0 708450.0 ;
      RECT  120750.0 706350.0 121650.0 707250.0 ;
      RECT  120750.0 707250.0 121650.0 708000.0 ;
      RECT  121200.0 707550.0 127800.0 708450.0 ;
      RECT  127800.0 707550.0 129000.0 708450.0 ;
      RECT  137250.0 707550.0 138150.0 708450.0 ;
      RECT  137250.0 706350.0 138150.0 707250.0 ;
      RECT  133200.0 707550.0 137700.0 708450.0 ;
      RECT  137250.0 706800.0 138150.0 708000.0 ;
      RECT  137700.0 706350.0 142200.0 707250.0 ;
      RECT  112650.0 720750.0 118200.0 721650.0 ;
      RECT  120750.0 719550.0 121650.0 720450.0 ;
      RECT  120750.0 720750.0 121650.0 721650.0 ;
      RECT  120750.0 720000.0 121650.0 721650.0 ;
      RECT  121200.0 719550.0 127800.0 720450.0 ;
      RECT  127800.0 719550.0 129000.0 720450.0 ;
      RECT  137250.0 719550.0 138150.0 720450.0 ;
      RECT  137250.0 720750.0 138150.0 721650.0 ;
      RECT  133200.0 719550.0 137700.0 720450.0 ;
      RECT  137250.0 720000.0 138150.0 721200.0 ;
      RECT  137700.0 720750.0 142200.0 721650.0 ;
      RECT  112650.0 733950.0 118200.0 734850.0 ;
      RECT  120750.0 735150.0 121650.0 736050.0 ;
      RECT  120750.0 733950.0 121650.0 734850.0 ;
      RECT  120750.0 734850.0 121650.0 735600.0 ;
      RECT  121200.0 735150.0 127800.0 736050.0 ;
      RECT  127800.0 735150.0 129000.0 736050.0 ;
      RECT  137250.0 735150.0 138150.0 736050.0 ;
      RECT  137250.0 733950.0 138150.0 734850.0 ;
      RECT  133200.0 735150.0 137700.0 736050.0 ;
      RECT  137250.0 734400.0 138150.0 735600.0 ;
      RECT  137700.0 733950.0 142200.0 734850.0 ;
      RECT  112650.0 748350.0 118200.0 749250.0 ;
      RECT  120750.0 747150.0 121650.0 748050.0 ;
      RECT  120750.0 748350.0 121650.0 749250.0 ;
      RECT  120750.0 747600.0 121650.0 749250.0 ;
      RECT  121200.0 747150.0 127800.0 748050.0 ;
      RECT  127800.0 747150.0 129000.0 748050.0 ;
      RECT  137250.0 747150.0 138150.0 748050.0 ;
      RECT  137250.0 748350.0 138150.0 749250.0 ;
      RECT  133200.0 747150.0 137700.0 748050.0 ;
      RECT  137250.0 747600.0 138150.0 748800.0 ;
      RECT  137700.0 748350.0 142200.0 749250.0 ;
      RECT  112650.0 761550.0 118200.0 762450.0 ;
      RECT  120750.0 762750.0 121650.0 763650.0 ;
      RECT  120750.0 761550.0 121650.0 762450.0 ;
      RECT  120750.0 762450.0 121650.0 763200.0 ;
      RECT  121200.0 762750.0 127800.0 763650.0 ;
      RECT  127800.0 762750.0 129000.0 763650.0 ;
      RECT  137250.0 762750.0 138150.0 763650.0 ;
      RECT  137250.0 761550.0 138150.0 762450.0 ;
      RECT  133200.0 762750.0 137700.0 763650.0 ;
      RECT  137250.0 762000.0 138150.0 763200.0 ;
      RECT  137700.0 761550.0 142200.0 762450.0 ;
      RECT  112650.0 775950.0 118200.0 776850.0 ;
      RECT  120750.0 774750.0 121650.0 775650.0 ;
      RECT  120750.0 775950.0 121650.0 776850.0 ;
      RECT  120750.0 775200.0 121650.0 776850.0 ;
      RECT  121200.0 774750.0 127800.0 775650.0 ;
      RECT  127800.0 774750.0 129000.0 775650.0 ;
      RECT  137250.0 774750.0 138150.0 775650.0 ;
      RECT  137250.0 775950.0 138150.0 776850.0 ;
      RECT  133200.0 774750.0 137700.0 775650.0 ;
      RECT  137250.0 775200.0 138150.0 776400.0 ;
      RECT  137700.0 775950.0 142200.0 776850.0 ;
      RECT  112650.0 789150.0 118200.0 790050.0 ;
      RECT  120750.0 790350.0 121650.0 791250.0 ;
      RECT  120750.0 789150.0 121650.0 790050.0 ;
      RECT  120750.0 790050.0 121650.0 790800.0 ;
      RECT  121200.0 790350.0 127800.0 791250.0 ;
      RECT  127800.0 790350.0 129000.0 791250.0 ;
      RECT  137250.0 790350.0 138150.0 791250.0 ;
      RECT  137250.0 789150.0 138150.0 790050.0 ;
      RECT  133200.0 790350.0 137700.0 791250.0 ;
      RECT  137250.0 789600.0 138150.0 790800.0 ;
      RECT  137700.0 789150.0 142200.0 790050.0 ;
      RECT  112650.0 803550.0 118200.0 804450.0 ;
      RECT  120750.0 802350.0 121650.0 803250.0 ;
      RECT  120750.0 803550.0 121650.0 804450.0 ;
      RECT  120750.0 802800.0 121650.0 804450.0 ;
      RECT  121200.0 802350.0 127800.0 803250.0 ;
      RECT  127800.0 802350.0 129000.0 803250.0 ;
      RECT  137250.0 802350.0 138150.0 803250.0 ;
      RECT  137250.0 803550.0 138150.0 804450.0 ;
      RECT  133200.0 802350.0 137700.0 803250.0 ;
      RECT  137250.0 802800.0 138150.0 804000.0 ;
      RECT  137700.0 803550.0 142200.0 804450.0 ;
      RECT  112650.0 816750.0 118200.0 817650.0 ;
      RECT  120750.0 817950.0 121650.0 818850.0 ;
      RECT  120750.0 816750.0 121650.0 817650.0 ;
      RECT  120750.0 817650.0 121650.0 818400.0 ;
      RECT  121200.0 817950.0 127800.0 818850.0 ;
      RECT  127800.0 817950.0 129000.0 818850.0 ;
      RECT  137250.0 817950.0 138150.0 818850.0 ;
      RECT  137250.0 816750.0 138150.0 817650.0 ;
      RECT  133200.0 817950.0 137700.0 818850.0 ;
      RECT  137250.0 817200.0 138150.0 818400.0 ;
      RECT  137700.0 816750.0 142200.0 817650.0 ;
      RECT  112650.0 831150.0 118200.0 832050.0 ;
      RECT  120750.0 829950.0 121650.0 830850.0 ;
      RECT  120750.0 831150.0 121650.0 832050.0 ;
      RECT  120750.0 830400.0 121650.0 832050.0 ;
      RECT  121200.0 829950.0 127800.0 830850.0 ;
      RECT  127800.0 829950.0 129000.0 830850.0 ;
      RECT  137250.0 829950.0 138150.0 830850.0 ;
      RECT  137250.0 831150.0 138150.0 832050.0 ;
      RECT  133200.0 829950.0 137700.0 830850.0 ;
      RECT  137250.0 830400.0 138150.0 831600.0 ;
      RECT  137700.0 831150.0 142200.0 832050.0 ;
      RECT  112650.0 844350.0 118200.0 845250.0 ;
      RECT  120750.0 845550.0 121650.0 846450.0 ;
      RECT  120750.0 844350.0 121650.0 845250.0 ;
      RECT  120750.0 845250.0 121650.0 846000.0 ;
      RECT  121200.0 845550.0 127800.0 846450.0 ;
      RECT  127800.0 845550.0 129000.0 846450.0 ;
      RECT  137250.0 845550.0 138150.0 846450.0 ;
      RECT  137250.0 844350.0 138150.0 845250.0 ;
      RECT  133200.0 845550.0 137700.0 846450.0 ;
      RECT  137250.0 844800.0 138150.0 846000.0 ;
      RECT  137700.0 844350.0 142200.0 845250.0 ;
      RECT  112650.0 858750.0 118200.0 859650.0 ;
      RECT  120750.0 857550.0 121650.0 858450.0 ;
      RECT  120750.0 858750.0 121650.0 859650.0 ;
      RECT  120750.0 858000.0 121650.0 859650.0 ;
      RECT  121200.0 857550.0 127800.0 858450.0 ;
      RECT  127800.0 857550.0 129000.0 858450.0 ;
      RECT  137250.0 857550.0 138150.0 858450.0 ;
      RECT  137250.0 858750.0 138150.0 859650.0 ;
      RECT  133200.0 857550.0 137700.0 858450.0 ;
      RECT  137250.0 858000.0 138150.0 859200.0 ;
      RECT  137700.0 858750.0 142200.0 859650.0 ;
      RECT  112650.0 871950.0 118200.0 872850.0 ;
      RECT  120750.0 873150.0 121650.0 874050.0 ;
      RECT  120750.0 871950.0 121650.0 872850.0 ;
      RECT  120750.0 872850.0 121650.0 873600.0 ;
      RECT  121200.0 873150.0 127800.0 874050.0 ;
      RECT  127800.0 873150.0 129000.0 874050.0 ;
      RECT  137250.0 873150.0 138150.0 874050.0 ;
      RECT  137250.0 871950.0 138150.0 872850.0 ;
      RECT  133200.0 873150.0 137700.0 874050.0 ;
      RECT  137250.0 872400.0 138150.0 873600.0 ;
      RECT  137700.0 871950.0 142200.0 872850.0 ;
      RECT  112650.0 886350.0 118200.0 887250.0 ;
      RECT  120750.0 885150.0 121650.0 886050.0 ;
      RECT  120750.0 886350.0 121650.0 887250.0 ;
      RECT  120750.0 885600.0 121650.0 887250.0 ;
      RECT  121200.0 885150.0 127800.0 886050.0 ;
      RECT  127800.0 885150.0 129000.0 886050.0 ;
      RECT  137250.0 885150.0 138150.0 886050.0 ;
      RECT  137250.0 886350.0 138150.0 887250.0 ;
      RECT  133200.0 885150.0 137700.0 886050.0 ;
      RECT  137250.0 885600.0 138150.0 886800.0 ;
      RECT  137700.0 886350.0 142200.0 887250.0 ;
      RECT  112650.0 899550.0 118200.0 900450.0 ;
      RECT  120750.0 900750.0 121650.0 901650.0 ;
      RECT  120750.0 899550.0 121650.0 900450.0 ;
      RECT  120750.0 900450.0 121650.0 901200.0 ;
      RECT  121200.0 900750.0 127800.0 901650.0 ;
      RECT  127800.0 900750.0 129000.0 901650.0 ;
      RECT  137250.0 900750.0 138150.0 901650.0 ;
      RECT  137250.0 899550.0 138150.0 900450.0 ;
      RECT  133200.0 900750.0 137700.0 901650.0 ;
      RECT  137250.0 900000.0 138150.0 901200.0 ;
      RECT  137700.0 899550.0 142200.0 900450.0 ;
      RECT  112650.0 913950.0 118200.0 914850.0 ;
      RECT  120750.0 912750.0 121650.0 913650.0 ;
      RECT  120750.0 913950.0 121650.0 914850.0 ;
      RECT  120750.0 913200.0 121650.0 914850.0 ;
      RECT  121200.0 912750.0 127800.0 913650.0 ;
      RECT  127800.0 912750.0 129000.0 913650.0 ;
      RECT  137250.0 912750.0 138150.0 913650.0 ;
      RECT  137250.0 913950.0 138150.0 914850.0 ;
      RECT  133200.0 912750.0 137700.0 913650.0 ;
      RECT  137250.0 913200.0 138150.0 914400.0 ;
      RECT  137700.0 913950.0 142200.0 914850.0 ;
      RECT  112650.0 927150.0 118200.0 928050.0 ;
      RECT  120750.0 928350.0 121650.0 929250.0 ;
      RECT  120750.0 927150.0 121650.0 928050.0 ;
      RECT  120750.0 928050.0 121650.0 928800.0 ;
      RECT  121200.0 928350.0 127800.0 929250.0 ;
      RECT  127800.0 928350.0 129000.0 929250.0 ;
      RECT  137250.0 928350.0 138150.0 929250.0 ;
      RECT  137250.0 927150.0 138150.0 928050.0 ;
      RECT  133200.0 928350.0 137700.0 929250.0 ;
      RECT  137250.0 927600.0 138150.0 928800.0 ;
      RECT  137700.0 927150.0 142200.0 928050.0 ;
      RECT  112650.0 941550.0 118200.0 942450.0 ;
      RECT  120750.0 940350.0 121650.0 941250.0 ;
      RECT  120750.0 941550.0 121650.0 942450.0 ;
      RECT  120750.0 940800.0 121650.0 942450.0 ;
      RECT  121200.0 940350.0 127800.0 941250.0 ;
      RECT  127800.0 940350.0 129000.0 941250.0 ;
      RECT  137250.0 940350.0 138150.0 941250.0 ;
      RECT  137250.0 941550.0 138150.0 942450.0 ;
      RECT  133200.0 940350.0 137700.0 941250.0 ;
      RECT  137250.0 940800.0 138150.0 942000.0 ;
      RECT  137700.0 941550.0 142200.0 942450.0 ;
      RECT  112650.0 954750.0 118200.0 955650.0 ;
      RECT  120750.0 955950.0 121650.0 956850.0 ;
      RECT  120750.0 954750.0 121650.0 955650.0 ;
      RECT  120750.0 955650.0 121650.0 956400.0 ;
      RECT  121200.0 955950.0 127800.0 956850.0 ;
      RECT  127800.0 955950.0 129000.0 956850.0 ;
      RECT  137250.0 955950.0 138150.0 956850.0 ;
      RECT  137250.0 954750.0 138150.0 955650.0 ;
      RECT  133200.0 955950.0 137700.0 956850.0 ;
      RECT  137250.0 955200.0 138150.0 956400.0 ;
      RECT  137700.0 954750.0 142200.0 955650.0 ;
      RECT  112650.0 969150.0 118200.0 970050.0 ;
      RECT  120750.0 967950.0 121650.0 968850.0 ;
      RECT  120750.0 969150.0 121650.0 970050.0 ;
      RECT  120750.0 968400.0 121650.0 970050.0 ;
      RECT  121200.0 967950.0 127800.0 968850.0 ;
      RECT  127800.0 967950.0 129000.0 968850.0 ;
      RECT  137250.0 967950.0 138150.0 968850.0 ;
      RECT  137250.0 969150.0 138150.0 970050.0 ;
      RECT  133200.0 967950.0 137700.0 968850.0 ;
      RECT  137250.0 968400.0 138150.0 969600.0 ;
      RECT  137700.0 969150.0 142200.0 970050.0 ;
      RECT  112650.0 982350.0 118200.0 983250.0 ;
      RECT  120750.0 983550.0 121650.0 984450.0 ;
      RECT  120750.0 982350.0 121650.0 983250.0 ;
      RECT  120750.0 983250.0 121650.0 984000.0 ;
      RECT  121200.0 983550.0 127800.0 984450.0 ;
      RECT  127800.0 983550.0 129000.0 984450.0 ;
      RECT  137250.0 983550.0 138150.0 984450.0 ;
      RECT  137250.0 982350.0 138150.0 983250.0 ;
      RECT  133200.0 983550.0 137700.0 984450.0 ;
      RECT  137250.0 982800.0 138150.0 984000.0 ;
      RECT  137700.0 982350.0 142200.0 983250.0 ;
      RECT  112650.0 996750.0 118200.0 997650.0 ;
      RECT  120750.0 995550.0 121650.0 996450.0 ;
      RECT  120750.0 996750.0 121650.0 997650.0 ;
      RECT  120750.0 996000.0 121650.0 997650.0 ;
      RECT  121200.0 995550.0 127800.0 996450.0 ;
      RECT  127800.0 995550.0 129000.0 996450.0 ;
      RECT  137250.0 995550.0 138150.0 996450.0 ;
      RECT  137250.0 996750.0 138150.0 997650.0 ;
      RECT  133200.0 995550.0 137700.0 996450.0 ;
      RECT  137250.0 996000.0 138150.0 997200.0 ;
      RECT  137700.0 996750.0 142200.0 997650.0 ;
      RECT  112650.0 1009950.0 118200.0 1010850.0 ;
      RECT  120750.0 1011150.0 121650.0 1012050.0 ;
      RECT  120750.0 1009950.0 121650.0 1010850.0 ;
      RECT  120750.0 1010850.0 121650.0 1011600.0 ;
      RECT  121200.0 1011150.0 127800.0 1012050.0 ;
      RECT  127800.0 1011150.0 129000.0 1012050.0 ;
      RECT  137250.0 1011150.0 138150.0 1012050.0 ;
      RECT  137250.0 1009950.0 138150.0 1010850.0 ;
      RECT  133200.0 1011150.0 137700.0 1012050.0 ;
      RECT  137250.0 1010400.0 138150.0 1011600.0 ;
      RECT  137700.0 1009950.0 142200.0 1010850.0 ;
      RECT  112650.0 1024350.0 118200.0 1025250.0 ;
      RECT  120750.0 1023150.0 121650.0 1024050.0 ;
      RECT  120750.0 1024350.0 121650.0 1025250.0 ;
      RECT  120750.0 1023600.0 121650.0 1025250.0 ;
      RECT  121200.0 1023150.0 127800.0 1024050.0 ;
      RECT  127800.0 1023150.0 129000.0 1024050.0 ;
      RECT  137250.0 1023150.0 138150.0 1024050.0 ;
      RECT  137250.0 1024350.0 138150.0 1025250.0 ;
      RECT  133200.0 1023150.0 137700.0 1024050.0 ;
      RECT  137250.0 1023600.0 138150.0 1024800.0 ;
      RECT  137700.0 1024350.0 142200.0 1025250.0 ;
      RECT  112650.0 1037550.0 118200.0 1038450.0 ;
      RECT  120750.0 1038750.0 121650.0 1039650.0 ;
      RECT  120750.0 1037550.0 121650.0 1038450.0 ;
      RECT  120750.0 1038450.0 121650.0 1039200.0 ;
      RECT  121200.0 1038750.0 127800.0 1039650.0 ;
      RECT  127800.0 1038750.0 129000.0 1039650.0 ;
      RECT  137250.0 1038750.0 138150.0 1039650.0 ;
      RECT  137250.0 1037550.0 138150.0 1038450.0 ;
      RECT  133200.0 1038750.0 137700.0 1039650.0 ;
      RECT  137250.0 1038000.0 138150.0 1039200.0 ;
      RECT  137700.0 1037550.0 142200.0 1038450.0 ;
      RECT  112650.0 1051950.0 118200.0 1052850.0 ;
      RECT  120750.0 1050750.0 121650.0 1051650.0 ;
      RECT  120750.0 1051950.0 121650.0 1052850.0 ;
      RECT  120750.0 1051200.0 121650.0 1052850.0 ;
      RECT  121200.0 1050750.0 127800.0 1051650.0 ;
      RECT  127800.0 1050750.0 129000.0 1051650.0 ;
      RECT  137250.0 1050750.0 138150.0 1051650.0 ;
      RECT  137250.0 1051950.0 138150.0 1052850.0 ;
      RECT  133200.0 1050750.0 137700.0 1051650.0 ;
      RECT  137250.0 1051200.0 138150.0 1052400.0 ;
      RECT  137700.0 1051950.0 142200.0 1052850.0 ;
      RECT  112650.0 1065150.0 118200.0 1066050.0 ;
      RECT  120750.0 1066350.0 121650.0 1067250.0 ;
      RECT  120750.0 1065150.0 121650.0 1066050.0 ;
      RECT  120750.0 1066050.0 121650.0 1066800.0 ;
      RECT  121200.0 1066350.0 127800.0 1067250.0 ;
      RECT  127800.0 1066350.0 129000.0 1067250.0 ;
      RECT  137250.0 1066350.0 138150.0 1067250.0 ;
      RECT  137250.0 1065150.0 138150.0 1066050.0 ;
      RECT  133200.0 1066350.0 137700.0 1067250.0 ;
      RECT  137250.0 1065600.0 138150.0 1066800.0 ;
      RECT  137700.0 1065150.0 142200.0 1066050.0 ;
      RECT  112650.0 1079550.0 118200.0 1080450.0 ;
      RECT  120750.0 1078350.0 121650.0 1079250.0 ;
      RECT  120750.0 1079550.0 121650.0 1080450.0 ;
      RECT  120750.0 1078800.0 121650.0 1080450.0 ;
      RECT  121200.0 1078350.0 127800.0 1079250.0 ;
      RECT  127800.0 1078350.0 129000.0 1079250.0 ;
      RECT  137250.0 1078350.0 138150.0 1079250.0 ;
      RECT  137250.0 1079550.0 138150.0 1080450.0 ;
      RECT  133200.0 1078350.0 137700.0 1079250.0 ;
      RECT  137250.0 1078800.0 138150.0 1080000.0 ;
      RECT  137700.0 1079550.0 142200.0 1080450.0 ;
      RECT  112650.0 1092750.0 118200.0 1093650.0 ;
      RECT  120750.0 1093950.0 121650.0 1094850.0 ;
      RECT  120750.0 1092750.0 121650.0 1093650.0 ;
      RECT  120750.0 1093650.0 121650.0 1094400.0 ;
      RECT  121200.0 1093950.0 127800.0 1094850.0 ;
      RECT  127800.0 1093950.0 129000.0 1094850.0 ;
      RECT  137250.0 1093950.0 138150.0 1094850.0 ;
      RECT  137250.0 1092750.0 138150.0 1093650.0 ;
      RECT  133200.0 1093950.0 137700.0 1094850.0 ;
      RECT  137250.0 1093200.0 138150.0 1094400.0 ;
      RECT  137700.0 1092750.0 142200.0 1093650.0 ;
      RECT  112650.0 1107150.0 118200.0 1108050.0 ;
      RECT  120750.0 1105950.0 121650.0 1106850.0 ;
      RECT  120750.0 1107150.0 121650.0 1108050.0 ;
      RECT  120750.0 1106400.0 121650.0 1108050.0 ;
      RECT  121200.0 1105950.0 127800.0 1106850.0 ;
      RECT  127800.0 1105950.0 129000.0 1106850.0 ;
      RECT  137250.0 1105950.0 138150.0 1106850.0 ;
      RECT  137250.0 1107150.0 138150.0 1108050.0 ;
      RECT  133200.0 1105950.0 137700.0 1106850.0 ;
      RECT  137250.0 1106400.0 138150.0 1107600.0 ;
      RECT  137700.0 1107150.0 142200.0 1108050.0 ;
      RECT  112650.0 1120350.0 118200.0 1121250.0 ;
      RECT  120750.0 1121550.0 121650.0 1122450.0 ;
      RECT  120750.0 1120350.0 121650.0 1121250.0 ;
      RECT  120750.0 1121250.0 121650.0 1122000.0 ;
      RECT  121200.0 1121550.0 127800.0 1122450.0 ;
      RECT  127800.0 1121550.0 129000.0 1122450.0 ;
      RECT  137250.0 1121550.0 138150.0 1122450.0 ;
      RECT  137250.0 1120350.0 138150.0 1121250.0 ;
      RECT  133200.0 1121550.0 137700.0 1122450.0 ;
      RECT  137250.0 1120800.0 138150.0 1122000.0 ;
      RECT  137700.0 1120350.0 142200.0 1121250.0 ;
      RECT  112650.0 1134750.0 118200.0 1135650.0 ;
      RECT  120750.0 1133550.0 121650.0 1134450.0 ;
      RECT  120750.0 1134750.0 121650.0 1135650.0 ;
      RECT  120750.0 1134000.0 121650.0 1135650.0 ;
      RECT  121200.0 1133550.0 127800.0 1134450.0 ;
      RECT  127800.0 1133550.0 129000.0 1134450.0 ;
      RECT  137250.0 1133550.0 138150.0 1134450.0 ;
      RECT  137250.0 1134750.0 138150.0 1135650.0 ;
      RECT  133200.0 1133550.0 137700.0 1134450.0 ;
      RECT  137250.0 1134000.0 138150.0 1135200.0 ;
      RECT  137700.0 1134750.0 142200.0 1135650.0 ;
      RECT  112650.0 1147950.0 118200.0 1148850.0 ;
      RECT  120750.0 1149150.0 121650.0 1150050.0 ;
      RECT  120750.0 1147950.0 121650.0 1148850.0 ;
      RECT  120750.0 1148850.0 121650.0 1149600.0 ;
      RECT  121200.0 1149150.0 127800.0 1150050.0 ;
      RECT  127800.0 1149150.0 129000.0 1150050.0 ;
      RECT  137250.0 1149150.0 138150.0 1150050.0 ;
      RECT  137250.0 1147950.0 138150.0 1148850.0 ;
      RECT  133200.0 1149150.0 137700.0 1150050.0 ;
      RECT  137250.0 1148400.0 138150.0 1149600.0 ;
      RECT  137700.0 1147950.0 142200.0 1148850.0 ;
      RECT  112650.0 1162350.0 118200.0 1163250.0 ;
      RECT  120750.0 1161150.0 121650.0 1162050.0 ;
      RECT  120750.0 1162350.0 121650.0 1163250.0 ;
      RECT  120750.0 1161600.0 121650.0 1163250.0 ;
      RECT  121200.0 1161150.0 127800.0 1162050.0 ;
      RECT  127800.0 1161150.0 129000.0 1162050.0 ;
      RECT  137250.0 1161150.0 138150.0 1162050.0 ;
      RECT  137250.0 1162350.0 138150.0 1163250.0 ;
      RECT  133200.0 1161150.0 137700.0 1162050.0 ;
      RECT  137250.0 1161600.0 138150.0 1162800.0 ;
      RECT  137700.0 1162350.0 142200.0 1163250.0 ;
      RECT  112650.0 1175550.0 118200.0 1176450.0 ;
      RECT  120750.0 1176750.0 121650.0 1177650.0 ;
      RECT  120750.0 1175550.0 121650.0 1176450.0 ;
      RECT  120750.0 1176450.0 121650.0 1177200.0 ;
      RECT  121200.0 1176750.0 127800.0 1177650.0 ;
      RECT  127800.0 1176750.0 129000.0 1177650.0 ;
      RECT  137250.0 1176750.0 138150.0 1177650.0 ;
      RECT  137250.0 1175550.0 138150.0 1176450.0 ;
      RECT  133200.0 1176750.0 137700.0 1177650.0 ;
      RECT  137250.0 1176000.0 138150.0 1177200.0 ;
      RECT  137700.0 1175550.0 142200.0 1176450.0 ;
      RECT  112650.0 1189950.0 118200.0 1190850.0 ;
      RECT  120750.0 1188750.0 121650.0 1189650.0 ;
      RECT  120750.0 1189950.0 121650.0 1190850.0 ;
      RECT  120750.0 1189200.0 121650.0 1190850.0 ;
      RECT  121200.0 1188750.0 127800.0 1189650.0 ;
      RECT  127800.0 1188750.0 129000.0 1189650.0 ;
      RECT  137250.0 1188750.0 138150.0 1189650.0 ;
      RECT  137250.0 1189950.0 138150.0 1190850.0 ;
      RECT  133200.0 1188750.0 137700.0 1189650.0 ;
      RECT  137250.0 1189200.0 138150.0 1190400.0 ;
      RECT  137700.0 1189950.0 142200.0 1190850.0 ;
      RECT  122400.0 325650.0 123600.0 327600.0 ;
      RECT  122400.0 313800.0 123600.0 315750.0 ;
      RECT  117600.0 315150.0 118800.0 313350.0 ;
      RECT  117600.0 324450.0 118800.0 328050.0 ;
      RECT  120300.0 315150.0 121200.0 324450.0 ;
      RECT  117600.0 324450.0 118800.0 325650.0 ;
      RECT  120000.0 324450.0 121200.0 325650.0 ;
      RECT  120000.0 324450.0 121200.0 325650.0 ;
      RECT  117600.0 324450.0 118800.0 325650.0 ;
      RECT  117600.0 315150.0 118800.0 316350.0 ;
      RECT  120000.0 315150.0 121200.0 316350.0 ;
      RECT  120000.0 315150.0 121200.0 316350.0 ;
      RECT  117600.0 315150.0 118800.0 316350.0 ;
      RECT  122400.0 325050.0 123600.0 326250.0 ;
      RECT  122400.0 315150.0 123600.0 316350.0 ;
      RECT  118200.0 319800.0 119400.0 321000.0 ;
      RECT  118200.0 319800.0 119400.0 321000.0 ;
      RECT  120750.0 319950.0 121650.0 320850.0 ;
      RECT  115800.0 327150.0 125400.0 328050.0 ;
      RECT  115800.0 313350.0 125400.0 314250.0 ;
      RECT  127200.0 315750.0 128400.0 313350.0 ;
      RECT  127200.0 324450.0 128400.0 328050.0 ;
      RECT  132000.0 324450.0 133200.0 328050.0 ;
      RECT  134400.0 325650.0 135600.0 327600.0 ;
      RECT  134400.0 313800.0 135600.0 315750.0 ;
      RECT  127200.0 324450.0 128400.0 325650.0 ;
      RECT  129600.0 324450.0 130800.0 325650.0 ;
      RECT  129600.0 324450.0 130800.0 325650.0 ;
      RECT  127200.0 324450.0 128400.0 325650.0 ;
      RECT  129600.0 324450.0 130800.0 325650.0 ;
      RECT  132000.0 324450.0 133200.0 325650.0 ;
      RECT  132000.0 324450.0 133200.0 325650.0 ;
      RECT  129600.0 324450.0 130800.0 325650.0 ;
      RECT  127200.0 315750.0 128400.0 316950.0 ;
      RECT  129600.0 315750.0 130800.0 316950.0 ;
      RECT  129600.0 315750.0 130800.0 316950.0 ;
      RECT  127200.0 315750.0 128400.0 316950.0 ;
      RECT  129600.0 315750.0 130800.0 316950.0 ;
      RECT  132000.0 315750.0 133200.0 316950.0 ;
      RECT  132000.0 315750.0 133200.0 316950.0 ;
      RECT  129600.0 315750.0 130800.0 316950.0 ;
      RECT  134400.0 325050.0 135600.0 326250.0 ;
      RECT  134400.0 315150.0 135600.0 316350.0 ;
      RECT  132000.0 318300.0 130800.0 319500.0 ;
      RECT  129000.0 321000.0 127800.0 322200.0 ;
      RECT  129600.0 324450.0 130800.0 325650.0 ;
      RECT  132000.0 315750.0 133200.0 316950.0 ;
      RECT  133200.0 321000.0 132000.0 322200.0 ;
      RECT  127800.0 321000.0 129000.0 322200.0 ;
      RECT  130800.0 318300.0 132000.0 319500.0 ;
      RECT  132000.0 321000.0 133200.0 322200.0 ;
      RECT  125400.0 327150.0 139800.0 328050.0 ;
      RECT  125400.0 313350.0 139800.0 314250.0 ;
      RECT  146400.0 325650.0 147600.0 327600.0 ;
      RECT  146400.0 313800.0 147600.0 315750.0 ;
      RECT  141600.0 315150.0 142800.0 313350.0 ;
      RECT  141600.0 324450.0 142800.0 328050.0 ;
      RECT  144300.0 315150.0 145200.0 324450.0 ;
      RECT  141600.0 324450.0 142800.0 325650.0 ;
      RECT  144000.0 324450.0 145200.0 325650.0 ;
      RECT  144000.0 324450.0 145200.0 325650.0 ;
      RECT  141600.0 324450.0 142800.0 325650.0 ;
      RECT  141600.0 315150.0 142800.0 316350.0 ;
      RECT  144000.0 315150.0 145200.0 316350.0 ;
      RECT  144000.0 315150.0 145200.0 316350.0 ;
      RECT  141600.0 315150.0 142800.0 316350.0 ;
      RECT  146400.0 325050.0 147600.0 326250.0 ;
      RECT  146400.0 315150.0 147600.0 316350.0 ;
      RECT  142200.0 319800.0 143400.0 321000.0 ;
      RECT  142200.0 319800.0 143400.0 321000.0 ;
      RECT  144750.0 319950.0 145650.0 320850.0 ;
      RECT  139800.0 327150.0 149400.0 328050.0 ;
      RECT  139800.0 313350.0 149400.0 314250.0 ;
      RECT  112050.0 319800.0 113250.0 321000.0 ;
      RECT  114000.0 317400.0 115200.0 318600.0 ;
      RECT  130800.0 318300.0 129600.0 319500.0 ;
      RECT  122400.0 329550.0 123600.0 327600.0 ;
      RECT  122400.0 341400.0 123600.0 339450.0 ;
      RECT  117600.0 340050.0 118800.0 341850.0 ;
      RECT  117600.0 330750.0 118800.0 327150.0 ;
      RECT  120300.0 340050.0 121200.0 330750.0 ;
      RECT  117600.0 330750.0 118800.0 329550.0 ;
      RECT  120000.0 330750.0 121200.0 329550.0 ;
      RECT  120000.0 330750.0 121200.0 329550.0 ;
      RECT  117600.0 330750.0 118800.0 329550.0 ;
      RECT  117600.0 340050.0 118800.0 338850.0 ;
      RECT  120000.0 340050.0 121200.0 338850.0 ;
      RECT  120000.0 340050.0 121200.0 338850.0 ;
      RECT  117600.0 340050.0 118800.0 338850.0 ;
      RECT  122400.0 330150.0 123600.0 328950.0 ;
      RECT  122400.0 340050.0 123600.0 338850.0 ;
      RECT  118200.0 335400.0 119400.0 334200.0 ;
      RECT  118200.0 335400.0 119400.0 334200.0 ;
      RECT  120750.0 335250.0 121650.0 334350.0 ;
      RECT  115800.0 328050.0 125400.0 327150.0 ;
      RECT  115800.0 341850.0 125400.0 340950.0 ;
      RECT  127200.0 339450.0 128400.0 341850.0 ;
      RECT  127200.0 330750.0 128400.0 327150.0 ;
      RECT  132000.0 330750.0 133200.0 327150.0 ;
      RECT  134400.0 329550.0 135600.0 327600.0 ;
      RECT  134400.0 341400.0 135600.0 339450.0 ;
      RECT  127200.0 330750.0 128400.0 329550.0 ;
      RECT  129600.0 330750.0 130800.0 329550.0 ;
      RECT  129600.0 330750.0 130800.0 329550.0 ;
      RECT  127200.0 330750.0 128400.0 329550.0 ;
      RECT  129600.0 330750.0 130800.0 329550.0 ;
      RECT  132000.0 330750.0 133200.0 329550.0 ;
      RECT  132000.0 330750.0 133200.0 329550.0 ;
      RECT  129600.0 330750.0 130800.0 329550.0 ;
      RECT  127200.0 339450.0 128400.0 338250.0 ;
      RECT  129600.0 339450.0 130800.0 338250.0 ;
      RECT  129600.0 339450.0 130800.0 338250.0 ;
      RECT  127200.0 339450.0 128400.0 338250.0 ;
      RECT  129600.0 339450.0 130800.0 338250.0 ;
      RECT  132000.0 339450.0 133200.0 338250.0 ;
      RECT  132000.0 339450.0 133200.0 338250.0 ;
      RECT  129600.0 339450.0 130800.0 338250.0 ;
      RECT  134400.0 330150.0 135600.0 328950.0 ;
      RECT  134400.0 340050.0 135600.0 338850.0 ;
      RECT  132000.0 336900.0 130800.0 335700.0 ;
      RECT  129000.0 334200.0 127800.0 333000.0 ;
      RECT  129600.0 330750.0 130800.0 329550.0 ;
      RECT  132000.0 339450.0 133200.0 338250.0 ;
      RECT  133200.0 334200.0 132000.0 333000.0 ;
      RECT  127800.0 334200.0 129000.0 333000.0 ;
      RECT  130800.0 336900.0 132000.0 335700.0 ;
      RECT  132000.0 334200.0 133200.0 333000.0 ;
      RECT  125400.0 328050.0 139800.0 327150.0 ;
      RECT  125400.0 341850.0 139800.0 340950.0 ;
      RECT  146400.0 329550.0 147600.0 327600.0 ;
      RECT  146400.0 341400.0 147600.0 339450.0 ;
      RECT  141600.0 340050.0 142800.0 341850.0 ;
      RECT  141600.0 330750.0 142800.0 327150.0 ;
      RECT  144300.0 340050.0 145200.0 330750.0 ;
      RECT  141600.0 330750.0 142800.0 329550.0 ;
      RECT  144000.0 330750.0 145200.0 329550.0 ;
      RECT  144000.0 330750.0 145200.0 329550.0 ;
      RECT  141600.0 330750.0 142800.0 329550.0 ;
      RECT  141600.0 340050.0 142800.0 338850.0 ;
      RECT  144000.0 340050.0 145200.0 338850.0 ;
      RECT  144000.0 340050.0 145200.0 338850.0 ;
      RECT  141600.0 340050.0 142800.0 338850.0 ;
      RECT  146400.0 330150.0 147600.0 328950.0 ;
      RECT  146400.0 340050.0 147600.0 338850.0 ;
      RECT  142200.0 335400.0 143400.0 334200.0 ;
      RECT  142200.0 335400.0 143400.0 334200.0 ;
      RECT  144750.0 335250.0 145650.0 334350.0 ;
      RECT  139800.0 328050.0 149400.0 327150.0 ;
      RECT  139800.0 341850.0 149400.0 340950.0 ;
      RECT  112050.0 334200.0 113250.0 335400.0 ;
      RECT  114000.0 336600.0 115200.0 337800.0 ;
      RECT  130800.0 335700.0 129600.0 336900.0 ;
      RECT  122400.0 353250.0 123600.0 355200.0 ;
      RECT  122400.0 341400.0 123600.0 343350.0 ;
      RECT  117600.0 342750.0 118800.0 340950.0 ;
      RECT  117600.0 352050.0 118800.0 355650.0 ;
      RECT  120300.0 342750.0 121200.0 352050.0 ;
      RECT  117600.0 352050.0 118800.0 353250.0 ;
      RECT  120000.0 352050.0 121200.0 353250.0 ;
      RECT  120000.0 352050.0 121200.0 353250.0 ;
      RECT  117600.0 352050.0 118800.0 353250.0 ;
      RECT  117600.0 342750.0 118800.0 343950.0 ;
      RECT  120000.0 342750.0 121200.0 343950.0 ;
      RECT  120000.0 342750.0 121200.0 343950.0 ;
      RECT  117600.0 342750.0 118800.0 343950.0 ;
      RECT  122400.0 352650.0 123600.0 353850.0 ;
      RECT  122400.0 342750.0 123600.0 343950.0 ;
      RECT  118200.0 347400.0 119400.0 348600.0 ;
      RECT  118200.0 347400.0 119400.0 348600.0 ;
      RECT  120750.0 347550.0 121650.0 348450.0 ;
      RECT  115800.0 354750.0 125400.0 355650.0 ;
      RECT  115800.0 340950.0 125400.0 341850.0 ;
      RECT  127200.0 343350.0 128400.0 340950.0 ;
      RECT  127200.0 352050.0 128400.0 355650.0 ;
      RECT  132000.0 352050.0 133200.0 355650.0 ;
      RECT  134400.0 353250.0 135600.0 355200.0 ;
      RECT  134400.0 341400.0 135600.0 343350.0 ;
      RECT  127200.0 352050.0 128400.0 353250.0 ;
      RECT  129600.0 352050.0 130800.0 353250.0 ;
      RECT  129600.0 352050.0 130800.0 353250.0 ;
      RECT  127200.0 352050.0 128400.0 353250.0 ;
      RECT  129600.0 352050.0 130800.0 353250.0 ;
      RECT  132000.0 352050.0 133200.0 353250.0 ;
      RECT  132000.0 352050.0 133200.0 353250.0 ;
      RECT  129600.0 352050.0 130800.0 353250.0 ;
      RECT  127200.0 343350.0 128400.0 344550.0 ;
      RECT  129600.0 343350.0 130800.0 344550.0 ;
      RECT  129600.0 343350.0 130800.0 344550.0 ;
      RECT  127200.0 343350.0 128400.0 344550.0 ;
      RECT  129600.0 343350.0 130800.0 344550.0 ;
      RECT  132000.0 343350.0 133200.0 344550.0 ;
      RECT  132000.0 343350.0 133200.0 344550.0 ;
      RECT  129600.0 343350.0 130800.0 344550.0 ;
      RECT  134400.0 352650.0 135600.0 353850.0 ;
      RECT  134400.0 342750.0 135600.0 343950.0 ;
      RECT  132000.0 345900.0 130800.0 347100.0 ;
      RECT  129000.0 348600.0 127800.0 349800.0 ;
      RECT  129600.0 352050.0 130800.0 353250.0 ;
      RECT  132000.0 343350.0 133200.0 344550.0 ;
      RECT  133200.0 348600.0 132000.0 349800.0 ;
      RECT  127800.0 348600.0 129000.0 349800.0 ;
      RECT  130800.0 345900.0 132000.0 347100.0 ;
      RECT  132000.0 348600.0 133200.0 349800.0 ;
      RECT  125400.0 354750.0 139800.0 355650.0 ;
      RECT  125400.0 340950.0 139800.0 341850.0 ;
      RECT  146400.0 353250.0 147600.0 355200.0 ;
      RECT  146400.0 341400.0 147600.0 343350.0 ;
      RECT  141600.0 342750.0 142800.0 340950.0 ;
      RECT  141600.0 352050.0 142800.0 355650.0 ;
      RECT  144300.0 342750.0 145200.0 352050.0 ;
      RECT  141600.0 352050.0 142800.0 353250.0 ;
      RECT  144000.0 352050.0 145200.0 353250.0 ;
      RECT  144000.0 352050.0 145200.0 353250.0 ;
      RECT  141600.0 352050.0 142800.0 353250.0 ;
      RECT  141600.0 342750.0 142800.0 343950.0 ;
      RECT  144000.0 342750.0 145200.0 343950.0 ;
      RECT  144000.0 342750.0 145200.0 343950.0 ;
      RECT  141600.0 342750.0 142800.0 343950.0 ;
      RECT  146400.0 352650.0 147600.0 353850.0 ;
      RECT  146400.0 342750.0 147600.0 343950.0 ;
      RECT  142200.0 347400.0 143400.0 348600.0 ;
      RECT  142200.0 347400.0 143400.0 348600.0 ;
      RECT  144750.0 347550.0 145650.0 348450.0 ;
      RECT  139800.0 354750.0 149400.0 355650.0 ;
      RECT  139800.0 340950.0 149400.0 341850.0 ;
      RECT  112050.0 347400.0 113250.0 348600.0 ;
      RECT  114000.0 345000.0 115200.0 346200.0 ;
      RECT  130800.0 345900.0 129600.0 347100.0 ;
      RECT  122400.0 357150.0 123600.0 355200.0 ;
      RECT  122400.0 369000.0 123600.0 367050.0 ;
      RECT  117600.0 367650.0 118800.0 369450.0 ;
      RECT  117600.0 358350.0 118800.0 354750.0 ;
      RECT  120300.0 367650.0 121200.0 358350.0 ;
      RECT  117600.0 358350.0 118800.0 357150.0 ;
      RECT  120000.0 358350.0 121200.0 357150.0 ;
      RECT  120000.0 358350.0 121200.0 357150.0 ;
      RECT  117600.0 358350.0 118800.0 357150.0 ;
      RECT  117600.0 367650.0 118800.0 366450.0 ;
      RECT  120000.0 367650.0 121200.0 366450.0 ;
      RECT  120000.0 367650.0 121200.0 366450.0 ;
      RECT  117600.0 367650.0 118800.0 366450.0 ;
      RECT  122400.0 357750.0 123600.0 356550.0 ;
      RECT  122400.0 367650.0 123600.0 366450.0 ;
      RECT  118200.0 363000.0 119400.0 361800.0 ;
      RECT  118200.0 363000.0 119400.0 361800.0 ;
      RECT  120750.0 362850.0 121650.0 361950.0 ;
      RECT  115800.0 355650.0 125400.0 354750.0 ;
      RECT  115800.0 369450.0 125400.0 368550.0 ;
      RECT  127200.0 367050.0 128400.0 369450.0 ;
      RECT  127200.0 358350.0 128400.0 354750.0 ;
      RECT  132000.0 358350.0 133200.0 354750.0 ;
      RECT  134400.0 357150.0 135600.0 355200.0 ;
      RECT  134400.0 369000.0 135600.0 367050.0 ;
      RECT  127200.0 358350.0 128400.0 357150.0 ;
      RECT  129600.0 358350.0 130800.0 357150.0 ;
      RECT  129600.0 358350.0 130800.0 357150.0 ;
      RECT  127200.0 358350.0 128400.0 357150.0 ;
      RECT  129600.0 358350.0 130800.0 357150.0 ;
      RECT  132000.0 358350.0 133200.0 357150.0 ;
      RECT  132000.0 358350.0 133200.0 357150.0 ;
      RECT  129600.0 358350.0 130800.0 357150.0 ;
      RECT  127200.0 367050.0 128400.0 365850.0 ;
      RECT  129600.0 367050.0 130800.0 365850.0 ;
      RECT  129600.0 367050.0 130800.0 365850.0 ;
      RECT  127200.0 367050.0 128400.0 365850.0 ;
      RECT  129600.0 367050.0 130800.0 365850.0 ;
      RECT  132000.0 367050.0 133200.0 365850.0 ;
      RECT  132000.0 367050.0 133200.0 365850.0 ;
      RECT  129600.0 367050.0 130800.0 365850.0 ;
      RECT  134400.0 357750.0 135600.0 356550.0 ;
      RECT  134400.0 367650.0 135600.0 366450.0 ;
      RECT  132000.0 364500.0 130800.0 363300.0 ;
      RECT  129000.0 361800.0 127800.0 360600.0 ;
      RECT  129600.0 358350.0 130800.0 357150.0 ;
      RECT  132000.0 367050.0 133200.0 365850.0 ;
      RECT  133200.0 361800.0 132000.0 360600.0 ;
      RECT  127800.0 361800.0 129000.0 360600.0 ;
      RECT  130800.0 364500.0 132000.0 363300.0 ;
      RECT  132000.0 361800.0 133200.0 360600.0 ;
      RECT  125400.0 355650.0 139800.0 354750.0 ;
      RECT  125400.0 369450.0 139800.0 368550.0 ;
      RECT  146400.0 357150.0 147600.0 355200.0 ;
      RECT  146400.0 369000.0 147600.0 367050.0 ;
      RECT  141600.0 367650.0 142800.0 369450.0 ;
      RECT  141600.0 358350.0 142800.0 354750.0 ;
      RECT  144300.0 367650.0 145200.0 358350.0 ;
      RECT  141600.0 358350.0 142800.0 357150.0 ;
      RECT  144000.0 358350.0 145200.0 357150.0 ;
      RECT  144000.0 358350.0 145200.0 357150.0 ;
      RECT  141600.0 358350.0 142800.0 357150.0 ;
      RECT  141600.0 367650.0 142800.0 366450.0 ;
      RECT  144000.0 367650.0 145200.0 366450.0 ;
      RECT  144000.0 367650.0 145200.0 366450.0 ;
      RECT  141600.0 367650.0 142800.0 366450.0 ;
      RECT  146400.0 357750.0 147600.0 356550.0 ;
      RECT  146400.0 367650.0 147600.0 366450.0 ;
      RECT  142200.0 363000.0 143400.0 361800.0 ;
      RECT  142200.0 363000.0 143400.0 361800.0 ;
      RECT  144750.0 362850.0 145650.0 361950.0 ;
      RECT  139800.0 355650.0 149400.0 354750.0 ;
      RECT  139800.0 369450.0 149400.0 368550.0 ;
      RECT  112050.0 361800.0 113250.0 363000.0 ;
      RECT  114000.0 364200.0 115200.0 365400.0 ;
      RECT  130800.0 363300.0 129600.0 364500.0 ;
      RECT  122400.0 380850.0 123600.0 382800.0 ;
      RECT  122400.0 369000.0 123600.0 370950.0 ;
      RECT  117600.0 370350.0 118800.0 368550.0 ;
      RECT  117600.0 379650.0 118800.0 383250.0 ;
      RECT  120300.0 370350.0 121200.0 379650.0 ;
      RECT  117600.0 379650.0 118800.0 380850.0 ;
      RECT  120000.0 379650.0 121200.0 380850.0 ;
      RECT  120000.0 379650.0 121200.0 380850.0 ;
      RECT  117600.0 379650.0 118800.0 380850.0 ;
      RECT  117600.0 370350.0 118800.0 371550.0 ;
      RECT  120000.0 370350.0 121200.0 371550.0 ;
      RECT  120000.0 370350.0 121200.0 371550.0 ;
      RECT  117600.0 370350.0 118800.0 371550.0 ;
      RECT  122400.0 380250.0 123600.0 381450.0 ;
      RECT  122400.0 370350.0 123600.0 371550.0 ;
      RECT  118200.0 375000.0 119400.0 376200.0 ;
      RECT  118200.0 375000.0 119400.0 376200.0 ;
      RECT  120750.0 375150.0 121650.0 376050.0 ;
      RECT  115800.0 382350.0 125400.0 383250.0 ;
      RECT  115800.0 368550.0 125400.0 369450.0 ;
      RECT  127200.0 370950.0 128400.0 368550.0 ;
      RECT  127200.0 379650.0 128400.0 383250.0 ;
      RECT  132000.0 379650.0 133200.0 383250.0 ;
      RECT  134400.0 380850.0 135600.0 382800.0 ;
      RECT  134400.0 369000.0 135600.0 370950.0 ;
      RECT  127200.0 379650.0 128400.0 380850.0 ;
      RECT  129600.0 379650.0 130800.0 380850.0 ;
      RECT  129600.0 379650.0 130800.0 380850.0 ;
      RECT  127200.0 379650.0 128400.0 380850.0 ;
      RECT  129600.0 379650.0 130800.0 380850.0 ;
      RECT  132000.0 379650.0 133200.0 380850.0 ;
      RECT  132000.0 379650.0 133200.0 380850.0 ;
      RECT  129600.0 379650.0 130800.0 380850.0 ;
      RECT  127200.0 370950.0 128400.0 372150.0 ;
      RECT  129600.0 370950.0 130800.0 372150.0 ;
      RECT  129600.0 370950.0 130800.0 372150.0 ;
      RECT  127200.0 370950.0 128400.0 372150.0 ;
      RECT  129600.0 370950.0 130800.0 372150.0 ;
      RECT  132000.0 370950.0 133200.0 372150.0 ;
      RECT  132000.0 370950.0 133200.0 372150.0 ;
      RECT  129600.0 370950.0 130800.0 372150.0 ;
      RECT  134400.0 380250.0 135600.0 381450.0 ;
      RECT  134400.0 370350.0 135600.0 371550.0 ;
      RECT  132000.0 373500.0 130800.0 374700.0 ;
      RECT  129000.0 376200.0 127800.0 377400.0 ;
      RECT  129600.0 379650.0 130800.0 380850.0 ;
      RECT  132000.0 370950.0 133200.0 372150.0 ;
      RECT  133200.0 376200.0 132000.0 377400.0 ;
      RECT  127800.0 376200.0 129000.0 377400.0 ;
      RECT  130800.0 373500.0 132000.0 374700.0 ;
      RECT  132000.0 376200.0 133200.0 377400.0 ;
      RECT  125400.0 382350.0 139800.0 383250.0 ;
      RECT  125400.0 368550.0 139800.0 369450.0 ;
      RECT  146400.0 380850.0 147600.0 382800.0 ;
      RECT  146400.0 369000.0 147600.0 370950.0 ;
      RECT  141600.0 370350.0 142800.0 368550.0 ;
      RECT  141600.0 379650.0 142800.0 383250.0 ;
      RECT  144300.0 370350.0 145200.0 379650.0 ;
      RECT  141600.0 379650.0 142800.0 380850.0 ;
      RECT  144000.0 379650.0 145200.0 380850.0 ;
      RECT  144000.0 379650.0 145200.0 380850.0 ;
      RECT  141600.0 379650.0 142800.0 380850.0 ;
      RECT  141600.0 370350.0 142800.0 371550.0 ;
      RECT  144000.0 370350.0 145200.0 371550.0 ;
      RECT  144000.0 370350.0 145200.0 371550.0 ;
      RECT  141600.0 370350.0 142800.0 371550.0 ;
      RECT  146400.0 380250.0 147600.0 381450.0 ;
      RECT  146400.0 370350.0 147600.0 371550.0 ;
      RECT  142200.0 375000.0 143400.0 376200.0 ;
      RECT  142200.0 375000.0 143400.0 376200.0 ;
      RECT  144750.0 375150.0 145650.0 376050.0 ;
      RECT  139800.0 382350.0 149400.0 383250.0 ;
      RECT  139800.0 368550.0 149400.0 369450.0 ;
      RECT  112050.0 375000.0 113250.0 376200.0 ;
      RECT  114000.0 372600.0 115200.0 373800.0 ;
      RECT  130800.0 373500.0 129600.0 374700.0 ;
      RECT  122400.0 384750.0 123600.0 382800.0 ;
      RECT  122400.0 396600.0 123600.0 394650.0 ;
      RECT  117600.0 395250.0 118800.0 397050.0 ;
      RECT  117600.0 385950.0 118800.0 382350.0 ;
      RECT  120300.0 395250.0 121200.0 385950.0 ;
      RECT  117600.0 385950.0 118800.0 384750.0 ;
      RECT  120000.0 385950.0 121200.0 384750.0 ;
      RECT  120000.0 385950.0 121200.0 384750.0 ;
      RECT  117600.0 385950.0 118800.0 384750.0 ;
      RECT  117600.0 395250.0 118800.0 394050.0 ;
      RECT  120000.0 395250.0 121200.0 394050.0 ;
      RECT  120000.0 395250.0 121200.0 394050.0 ;
      RECT  117600.0 395250.0 118800.0 394050.0 ;
      RECT  122400.0 385350.0 123600.0 384150.0 ;
      RECT  122400.0 395250.0 123600.0 394050.0 ;
      RECT  118200.0 390600.0 119400.0 389400.0 ;
      RECT  118200.0 390600.0 119400.0 389400.0 ;
      RECT  120750.0 390450.0 121650.0 389550.0 ;
      RECT  115800.0 383250.0 125400.0 382350.0 ;
      RECT  115800.0 397050.0 125400.0 396150.0 ;
      RECT  127200.0 394650.0 128400.0 397050.0 ;
      RECT  127200.0 385950.0 128400.0 382350.0 ;
      RECT  132000.0 385950.0 133200.0 382350.0 ;
      RECT  134400.0 384750.0 135600.0 382800.0 ;
      RECT  134400.0 396600.0 135600.0 394650.0 ;
      RECT  127200.0 385950.0 128400.0 384750.0 ;
      RECT  129600.0 385950.0 130800.0 384750.0 ;
      RECT  129600.0 385950.0 130800.0 384750.0 ;
      RECT  127200.0 385950.0 128400.0 384750.0 ;
      RECT  129600.0 385950.0 130800.0 384750.0 ;
      RECT  132000.0 385950.0 133200.0 384750.0 ;
      RECT  132000.0 385950.0 133200.0 384750.0 ;
      RECT  129600.0 385950.0 130800.0 384750.0 ;
      RECT  127200.0 394650.0 128400.0 393450.0 ;
      RECT  129600.0 394650.0 130800.0 393450.0 ;
      RECT  129600.0 394650.0 130800.0 393450.0 ;
      RECT  127200.0 394650.0 128400.0 393450.0 ;
      RECT  129600.0 394650.0 130800.0 393450.0 ;
      RECT  132000.0 394650.0 133200.0 393450.0 ;
      RECT  132000.0 394650.0 133200.0 393450.0 ;
      RECT  129600.0 394650.0 130800.0 393450.0 ;
      RECT  134400.0 385350.0 135600.0 384150.0 ;
      RECT  134400.0 395250.0 135600.0 394050.0 ;
      RECT  132000.0 392100.0 130800.0 390900.0 ;
      RECT  129000.0 389400.0 127800.0 388200.0 ;
      RECT  129600.0 385950.0 130800.0 384750.0 ;
      RECT  132000.0 394650.0 133200.0 393450.0 ;
      RECT  133200.0 389400.0 132000.0 388200.0 ;
      RECT  127800.0 389400.0 129000.0 388200.0 ;
      RECT  130800.0 392100.0 132000.0 390900.0 ;
      RECT  132000.0 389400.0 133200.0 388200.0 ;
      RECT  125400.0 383250.0 139800.0 382350.0 ;
      RECT  125400.0 397050.0 139800.0 396150.0 ;
      RECT  146400.0 384750.0 147600.0 382800.0 ;
      RECT  146400.0 396600.0 147600.0 394650.0 ;
      RECT  141600.0 395250.0 142800.0 397050.0 ;
      RECT  141600.0 385950.0 142800.0 382350.0 ;
      RECT  144300.0 395250.0 145200.0 385950.0 ;
      RECT  141600.0 385950.0 142800.0 384750.0 ;
      RECT  144000.0 385950.0 145200.0 384750.0 ;
      RECT  144000.0 385950.0 145200.0 384750.0 ;
      RECT  141600.0 385950.0 142800.0 384750.0 ;
      RECT  141600.0 395250.0 142800.0 394050.0 ;
      RECT  144000.0 395250.0 145200.0 394050.0 ;
      RECT  144000.0 395250.0 145200.0 394050.0 ;
      RECT  141600.0 395250.0 142800.0 394050.0 ;
      RECT  146400.0 385350.0 147600.0 384150.0 ;
      RECT  146400.0 395250.0 147600.0 394050.0 ;
      RECT  142200.0 390600.0 143400.0 389400.0 ;
      RECT  142200.0 390600.0 143400.0 389400.0 ;
      RECT  144750.0 390450.0 145650.0 389550.0 ;
      RECT  139800.0 383250.0 149400.0 382350.0 ;
      RECT  139800.0 397050.0 149400.0 396150.0 ;
      RECT  112050.0 389400.0 113250.0 390600.0 ;
      RECT  114000.0 391800.0 115200.0 393000.0 ;
      RECT  130800.0 390900.0 129600.0 392100.0 ;
      RECT  122400.0 408450.0 123600.0 410400.0 ;
      RECT  122400.0 396600.0 123600.0 398550.0 ;
      RECT  117600.0 397950.0 118800.0 396150.0 ;
      RECT  117600.0 407250.0 118800.0 410850.0 ;
      RECT  120300.0 397950.0 121200.0 407250.0 ;
      RECT  117600.0 407250.0 118800.0 408450.0 ;
      RECT  120000.0 407250.0 121200.0 408450.0 ;
      RECT  120000.0 407250.0 121200.0 408450.0 ;
      RECT  117600.0 407250.0 118800.0 408450.0 ;
      RECT  117600.0 397950.0 118800.0 399150.0 ;
      RECT  120000.0 397950.0 121200.0 399150.0 ;
      RECT  120000.0 397950.0 121200.0 399150.0 ;
      RECT  117600.0 397950.0 118800.0 399150.0 ;
      RECT  122400.0 407850.0 123600.0 409050.0 ;
      RECT  122400.0 397950.0 123600.0 399150.0 ;
      RECT  118200.0 402600.0 119400.0 403800.0 ;
      RECT  118200.0 402600.0 119400.0 403800.0 ;
      RECT  120750.0 402750.0 121650.0 403650.0 ;
      RECT  115800.0 409950.0 125400.0 410850.0 ;
      RECT  115800.0 396150.0 125400.0 397050.0 ;
      RECT  127200.0 398550.0 128400.0 396150.0 ;
      RECT  127200.0 407250.0 128400.0 410850.0 ;
      RECT  132000.0 407250.0 133200.0 410850.0 ;
      RECT  134400.0 408450.0 135600.0 410400.0 ;
      RECT  134400.0 396600.0 135600.0 398550.0 ;
      RECT  127200.0 407250.0 128400.0 408450.0 ;
      RECT  129600.0 407250.0 130800.0 408450.0 ;
      RECT  129600.0 407250.0 130800.0 408450.0 ;
      RECT  127200.0 407250.0 128400.0 408450.0 ;
      RECT  129600.0 407250.0 130800.0 408450.0 ;
      RECT  132000.0 407250.0 133200.0 408450.0 ;
      RECT  132000.0 407250.0 133200.0 408450.0 ;
      RECT  129600.0 407250.0 130800.0 408450.0 ;
      RECT  127200.0 398550.0 128400.0 399750.0 ;
      RECT  129600.0 398550.0 130800.0 399750.0 ;
      RECT  129600.0 398550.0 130800.0 399750.0 ;
      RECT  127200.0 398550.0 128400.0 399750.0 ;
      RECT  129600.0 398550.0 130800.0 399750.0 ;
      RECT  132000.0 398550.0 133200.0 399750.0 ;
      RECT  132000.0 398550.0 133200.0 399750.0 ;
      RECT  129600.0 398550.0 130800.0 399750.0 ;
      RECT  134400.0 407850.0 135600.0 409050.0 ;
      RECT  134400.0 397950.0 135600.0 399150.0 ;
      RECT  132000.0 401100.0 130800.0 402300.0 ;
      RECT  129000.0 403800.0 127800.0 405000.0 ;
      RECT  129600.0 407250.0 130800.0 408450.0 ;
      RECT  132000.0 398550.0 133200.0 399750.0 ;
      RECT  133200.0 403800.0 132000.0 405000.0 ;
      RECT  127800.0 403800.0 129000.0 405000.0 ;
      RECT  130800.0 401100.0 132000.0 402300.0 ;
      RECT  132000.0 403800.0 133200.0 405000.0 ;
      RECT  125400.0 409950.0 139800.0 410850.0 ;
      RECT  125400.0 396150.0 139800.0 397050.0 ;
      RECT  146400.0 408450.0 147600.0 410400.0 ;
      RECT  146400.0 396600.0 147600.0 398550.0 ;
      RECT  141600.0 397950.0 142800.0 396150.0 ;
      RECT  141600.0 407250.0 142800.0 410850.0 ;
      RECT  144300.0 397950.0 145200.0 407250.0 ;
      RECT  141600.0 407250.0 142800.0 408450.0 ;
      RECT  144000.0 407250.0 145200.0 408450.0 ;
      RECT  144000.0 407250.0 145200.0 408450.0 ;
      RECT  141600.0 407250.0 142800.0 408450.0 ;
      RECT  141600.0 397950.0 142800.0 399150.0 ;
      RECT  144000.0 397950.0 145200.0 399150.0 ;
      RECT  144000.0 397950.0 145200.0 399150.0 ;
      RECT  141600.0 397950.0 142800.0 399150.0 ;
      RECT  146400.0 407850.0 147600.0 409050.0 ;
      RECT  146400.0 397950.0 147600.0 399150.0 ;
      RECT  142200.0 402600.0 143400.0 403800.0 ;
      RECT  142200.0 402600.0 143400.0 403800.0 ;
      RECT  144750.0 402750.0 145650.0 403650.0 ;
      RECT  139800.0 409950.0 149400.0 410850.0 ;
      RECT  139800.0 396150.0 149400.0 397050.0 ;
      RECT  112050.0 402600.0 113250.0 403800.0 ;
      RECT  114000.0 400200.0 115200.0 401400.0 ;
      RECT  130800.0 401100.0 129600.0 402300.0 ;
      RECT  122400.0 412350.0 123600.0 410400.0 ;
      RECT  122400.0 424200.0 123600.0 422250.0 ;
      RECT  117600.0 422850.0 118800.0 424650.0 ;
      RECT  117600.0 413550.0 118800.0 409950.0 ;
      RECT  120300.0 422850.0 121200.0 413550.0 ;
      RECT  117600.0 413550.0 118800.0 412350.0 ;
      RECT  120000.0 413550.0 121200.0 412350.0 ;
      RECT  120000.0 413550.0 121200.0 412350.0 ;
      RECT  117600.0 413550.0 118800.0 412350.0 ;
      RECT  117600.0 422850.0 118800.0 421650.0 ;
      RECT  120000.0 422850.0 121200.0 421650.0 ;
      RECT  120000.0 422850.0 121200.0 421650.0 ;
      RECT  117600.0 422850.0 118800.0 421650.0 ;
      RECT  122400.0 412950.0 123600.0 411750.0 ;
      RECT  122400.0 422850.0 123600.0 421650.0 ;
      RECT  118200.0 418200.0 119400.0 417000.0 ;
      RECT  118200.0 418200.0 119400.0 417000.0 ;
      RECT  120750.0 418050.0 121650.0 417150.0 ;
      RECT  115800.0 410850.0 125400.0 409950.0 ;
      RECT  115800.0 424650.0 125400.0 423750.0 ;
      RECT  127200.0 422250.0 128400.0 424650.0 ;
      RECT  127200.0 413550.0 128400.0 409950.0 ;
      RECT  132000.0 413550.0 133200.0 409950.0 ;
      RECT  134400.0 412350.0 135600.0 410400.0 ;
      RECT  134400.0 424200.0 135600.0 422250.0 ;
      RECT  127200.0 413550.0 128400.0 412350.0 ;
      RECT  129600.0 413550.0 130800.0 412350.0 ;
      RECT  129600.0 413550.0 130800.0 412350.0 ;
      RECT  127200.0 413550.0 128400.0 412350.0 ;
      RECT  129600.0 413550.0 130800.0 412350.0 ;
      RECT  132000.0 413550.0 133200.0 412350.0 ;
      RECT  132000.0 413550.0 133200.0 412350.0 ;
      RECT  129600.0 413550.0 130800.0 412350.0 ;
      RECT  127200.0 422250.0 128400.0 421050.0 ;
      RECT  129600.0 422250.0 130800.0 421050.0 ;
      RECT  129600.0 422250.0 130800.0 421050.0 ;
      RECT  127200.0 422250.0 128400.0 421050.0 ;
      RECT  129600.0 422250.0 130800.0 421050.0 ;
      RECT  132000.0 422250.0 133200.0 421050.0 ;
      RECT  132000.0 422250.0 133200.0 421050.0 ;
      RECT  129600.0 422250.0 130800.0 421050.0 ;
      RECT  134400.0 412950.0 135600.0 411750.0 ;
      RECT  134400.0 422850.0 135600.0 421650.0 ;
      RECT  132000.0 419700.0 130800.0 418500.0 ;
      RECT  129000.0 417000.0 127800.0 415800.0 ;
      RECT  129600.0 413550.0 130800.0 412350.0 ;
      RECT  132000.0 422250.0 133200.0 421050.0 ;
      RECT  133200.0 417000.0 132000.0 415800.0 ;
      RECT  127800.0 417000.0 129000.0 415800.0 ;
      RECT  130800.0 419700.0 132000.0 418500.0 ;
      RECT  132000.0 417000.0 133200.0 415800.0 ;
      RECT  125400.0 410850.0 139800.0 409950.0 ;
      RECT  125400.0 424650.0 139800.0 423750.0 ;
      RECT  146400.0 412350.0 147600.0 410400.0 ;
      RECT  146400.0 424200.0 147600.0 422250.0 ;
      RECT  141600.0 422850.0 142800.0 424650.0 ;
      RECT  141600.0 413550.0 142800.0 409950.0 ;
      RECT  144300.0 422850.0 145200.0 413550.0 ;
      RECT  141600.0 413550.0 142800.0 412350.0 ;
      RECT  144000.0 413550.0 145200.0 412350.0 ;
      RECT  144000.0 413550.0 145200.0 412350.0 ;
      RECT  141600.0 413550.0 142800.0 412350.0 ;
      RECT  141600.0 422850.0 142800.0 421650.0 ;
      RECT  144000.0 422850.0 145200.0 421650.0 ;
      RECT  144000.0 422850.0 145200.0 421650.0 ;
      RECT  141600.0 422850.0 142800.0 421650.0 ;
      RECT  146400.0 412950.0 147600.0 411750.0 ;
      RECT  146400.0 422850.0 147600.0 421650.0 ;
      RECT  142200.0 418200.0 143400.0 417000.0 ;
      RECT  142200.0 418200.0 143400.0 417000.0 ;
      RECT  144750.0 418050.0 145650.0 417150.0 ;
      RECT  139800.0 410850.0 149400.0 409950.0 ;
      RECT  139800.0 424650.0 149400.0 423750.0 ;
      RECT  112050.0 417000.0 113250.0 418200.0 ;
      RECT  114000.0 419400.0 115200.0 420600.0 ;
      RECT  130800.0 418500.0 129600.0 419700.0 ;
      RECT  122400.0 436050.0 123600.0 438000.0 ;
      RECT  122400.0 424200.0 123600.0 426150.0 ;
      RECT  117600.0 425550.0 118800.0 423750.0 ;
      RECT  117600.0 434850.0 118800.0 438450.0 ;
      RECT  120300.0 425550.0 121200.0 434850.0 ;
      RECT  117600.0 434850.0 118800.0 436050.0 ;
      RECT  120000.0 434850.0 121200.0 436050.0 ;
      RECT  120000.0 434850.0 121200.0 436050.0 ;
      RECT  117600.0 434850.0 118800.0 436050.0 ;
      RECT  117600.0 425550.0 118800.0 426750.0 ;
      RECT  120000.0 425550.0 121200.0 426750.0 ;
      RECT  120000.0 425550.0 121200.0 426750.0 ;
      RECT  117600.0 425550.0 118800.0 426750.0 ;
      RECT  122400.0 435450.0 123600.0 436650.0 ;
      RECT  122400.0 425550.0 123600.0 426750.0 ;
      RECT  118200.0 430200.0 119400.0 431400.0 ;
      RECT  118200.0 430200.0 119400.0 431400.0 ;
      RECT  120750.0 430350.0 121650.0 431250.0 ;
      RECT  115800.0 437550.0 125400.0 438450.0 ;
      RECT  115800.0 423750.0 125400.0 424650.0 ;
      RECT  127200.0 426150.0 128400.0 423750.0 ;
      RECT  127200.0 434850.0 128400.0 438450.0 ;
      RECT  132000.0 434850.0 133200.0 438450.0 ;
      RECT  134400.0 436050.0 135600.0 438000.0 ;
      RECT  134400.0 424200.0 135600.0 426150.0 ;
      RECT  127200.0 434850.0 128400.0 436050.0 ;
      RECT  129600.0 434850.0 130800.0 436050.0 ;
      RECT  129600.0 434850.0 130800.0 436050.0 ;
      RECT  127200.0 434850.0 128400.0 436050.0 ;
      RECT  129600.0 434850.0 130800.0 436050.0 ;
      RECT  132000.0 434850.0 133200.0 436050.0 ;
      RECT  132000.0 434850.0 133200.0 436050.0 ;
      RECT  129600.0 434850.0 130800.0 436050.0 ;
      RECT  127200.0 426150.0 128400.0 427350.0 ;
      RECT  129600.0 426150.0 130800.0 427350.0 ;
      RECT  129600.0 426150.0 130800.0 427350.0 ;
      RECT  127200.0 426150.0 128400.0 427350.0 ;
      RECT  129600.0 426150.0 130800.0 427350.0 ;
      RECT  132000.0 426150.0 133200.0 427350.0 ;
      RECT  132000.0 426150.0 133200.0 427350.0 ;
      RECT  129600.0 426150.0 130800.0 427350.0 ;
      RECT  134400.0 435450.0 135600.0 436650.0 ;
      RECT  134400.0 425550.0 135600.0 426750.0 ;
      RECT  132000.0 428700.0 130800.0 429900.0 ;
      RECT  129000.0 431400.0 127800.0 432600.0 ;
      RECT  129600.0 434850.0 130800.0 436050.0 ;
      RECT  132000.0 426150.0 133200.0 427350.0 ;
      RECT  133200.0 431400.0 132000.0 432600.0 ;
      RECT  127800.0 431400.0 129000.0 432600.0 ;
      RECT  130800.0 428700.0 132000.0 429900.0 ;
      RECT  132000.0 431400.0 133200.0 432600.0 ;
      RECT  125400.0 437550.0 139800.0 438450.0 ;
      RECT  125400.0 423750.0 139800.0 424650.0 ;
      RECT  146400.0 436050.0 147600.0 438000.0 ;
      RECT  146400.0 424200.0 147600.0 426150.0 ;
      RECT  141600.0 425550.0 142800.0 423750.0 ;
      RECT  141600.0 434850.0 142800.0 438450.0 ;
      RECT  144300.0 425550.0 145200.0 434850.0 ;
      RECT  141600.0 434850.0 142800.0 436050.0 ;
      RECT  144000.0 434850.0 145200.0 436050.0 ;
      RECT  144000.0 434850.0 145200.0 436050.0 ;
      RECT  141600.0 434850.0 142800.0 436050.0 ;
      RECT  141600.0 425550.0 142800.0 426750.0 ;
      RECT  144000.0 425550.0 145200.0 426750.0 ;
      RECT  144000.0 425550.0 145200.0 426750.0 ;
      RECT  141600.0 425550.0 142800.0 426750.0 ;
      RECT  146400.0 435450.0 147600.0 436650.0 ;
      RECT  146400.0 425550.0 147600.0 426750.0 ;
      RECT  142200.0 430200.0 143400.0 431400.0 ;
      RECT  142200.0 430200.0 143400.0 431400.0 ;
      RECT  144750.0 430350.0 145650.0 431250.0 ;
      RECT  139800.0 437550.0 149400.0 438450.0 ;
      RECT  139800.0 423750.0 149400.0 424650.0 ;
      RECT  112050.0 430200.0 113250.0 431400.0 ;
      RECT  114000.0 427800.0 115200.0 429000.0 ;
      RECT  130800.0 428700.0 129600.0 429900.0 ;
      RECT  122400.0 439950.0 123600.0 438000.0 ;
      RECT  122400.0 451800.0 123600.0 449850.0 ;
      RECT  117600.0 450450.0 118800.0 452250.0 ;
      RECT  117600.0 441150.0 118800.0 437550.0 ;
      RECT  120300.0 450450.0 121200.0 441150.0 ;
      RECT  117600.0 441150.0 118800.0 439950.0 ;
      RECT  120000.0 441150.0 121200.0 439950.0 ;
      RECT  120000.0 441150.0 121200.0 439950.0 ;
      RECT  117600.0 441150.0 118800.0 439950.0 ;
      RECT  117600.0 450450.0 118800.0 449250.0 ;
      RECT  120000.0 450450.0 121200.0 449250.0 ;
      RECT  120000.0 450450.0 121200.0 449250.0 ;
      RECT  117600.0 450450.0 118800.0 449250.0 ;
      RECT  122400.0 440550.0 123600.0 439350.0 ;
      RECT  122400.0 450450.0 123600.0 449250.0 ;
      RECT  118200.0 445800.0 119400.0 444600.0 ;
      RECT  118200.0 445800.0 119400.0 444600.0 ;
      RECT  120750.0 445650.0 121650.0 444750.0 ;
      RECT  115800.0 438450.0 125400.0 437550.0 ;
      RECT  115800.0 452250.0 125400.0 451350.0 ;
      RECT  127200.0 449850.0 128400.0 452250.0 ;
      RECT  127200.0 441150.0 128400.0 437550.0 ;
      RECT  132000.0 441150.0 133200.0 437550.0 ;
      RECT  134400.0 439950.0 135600.0 438000.0 ;
      RECT  134400.0 451800.0 135600.0 449850.0 ;
      RECT  127200.0 441150.0 128400.0 439950.0 ;
      RECT  129600.0 441150.0 130800.0 439950.0 ;
      RECT  129600.0 441150.0 130800.0 439950.0 ;
      RECT  127200.0 441150.0 128400.0 439950.0 ;
      RECT  129600.0 441150.0 130800.0 439950.0 ;
      RECT  132000.0 441150.0 133200.0 439950.0 ;
      RECT  132000.0 441150.0 133200.0 439950.0 ;
      RECT  129600.0 441150.0 130800.0 439950.0 ;
      RECT  127200.0 449850.0 128400.0 448650.0 ;
      RECT  129600.0 449850.0 130800.0 448650.0 ;
      RECT  129600.0 449850.0 130800.0 448650.0 ;
      RECT  127200.0 449850.0 128400.0 448650.0 ;
      RECT  129600.0 449850.0 130800.0 448650.0 ;
      RECT  132000.0 449850.0 133200.0 448650.0 ;
      RECT  132000.0 449850.0 133200.0 448650.0 ;
      RECT  129600.0 449850.0 130800.0 448650.0 ;
      RECT  134400.0 440550.0 135600.0 439350.0 ;
      RECT  134400.0 450450.0 135600.0 449250.0 ;
      RECT  132000.0 447300.0 130800.0 446100.0 ;
      RECT  129000.0 444600.0 127800.0 443400.0 ;
      RECT  129600.0 441150.0 130800.0 439950.0 ;
      RECT  132000.0 449850.0 133200.0 448650.0 ;
      RECT  133200.0 444600.0 132000.0 443400.0 ;
      RECT  127800.0 444600.0 129000.0 443400.0 ;
      RECT  130800.0 447300.0 132000.0 446100.0 ;
      RECT  132000.0 444600.0 133200.0 443400.0 ;
      RECT  125400.0 438450.0 139800.0 437550.0 ;
      RECT  125400.0 452250.0 139800.0 451350.0 ;
      RECT  146400.0 439950.0 147600.0 438000.0 ;
      RECT  146400.0 451800.0 147600.0 449850.0 ;
      RECT  141600.0 450450.0 142800.0 452250.0 ;
      RECT  141600.0 441150.0 142800.0 437550.0 ;
      RECT  144300.0 450450.0 145200.0 441150.0 ;
      RECT  141600.0 441150.0 142800.0 439950.0 ;
      RECT  144000.0 441150.0 145200.0 439950.0 ;
      RECT  144000.0 441150.0 145200.0 439950.0 ;
      RECT  141600.0 441150.0 142800.0 439950.0 ;
      RECT  141600.0 450450.0 142800.0 449250.0 ;
      RECT  144000.0 450450.0 145200.0 449250.0 ;
      RECT  144000.0 450450.0 145200.0 449250.0 ;
      RECT  141600.0 450450.0 142800.0 449250.0 ;
      RECT  146400.0 440550.0 147600.0 439350.0 ;
      RECT  146400.0 450450.0 147600.0 449250.0 ;
      RECT  142200.0 445800.0 143400.0 444600.0 ;
      RECT  142200.0 445800.0 143400.0 444600.0 ;
      RECT  144750.0 445650.0 145650.0 444750.0 ;
      RECT  139800.0 438450.0 149400.0 437550.0 ;
      RECT  139800.0 452250.0 149400.0 451350.0 ;
      RECT  112050.0 444600.0 113250.0 445800.0 ;
      RECT  114000.0 447000.0 115200.0 448200.0 ;
      RECT  130800.0 446100.0 129600.0 447300.0 ;
      RECT  122400.0 463650.0 123600.0 465600.0 ;
      RECT  122400.0 451800.0 123600.0 453750.0 ;
      RECT  117600.0 453150.0 118800.0 451350.0 ;
      RECT  117600.0 462450.0 118800.0 466050.0 ;
      RECT  120300.0 453150.0 121200.0 462450.0 ;
      RECT  117600.0 462450.0 118800.0 463650.0 ;
      RECT  120000.0 462450.0 121200.0 463650.0 ;
      RECT  120000.0 462450.0 121200.0 463650.0 ;
      RECT  117600.0 462450.0 118800.0 463650.0 ;
      RECT  117600.0 453150.0 118800.0 454350.0 ;
      RECT  120000.0 453150.0 121200.0 454350.0 ;
      RECT  120000.0 453150.0 121200.0 454350.0 ;
      RECT  117600.0 453150.0 118800.0 454350.0 ;
      RECT  122400.0 463050.0 123600.0 464250.0 ;
      RECT  122400.0 453150.0 123600.0 454350.0 ;
      RECT  118200.0 457800.0 119400.0 459000.0 ;
      RECT  118200.0 457800.0 119400.0 459000.0 ;
      RECT  120750.0 457950.0 121650.0 458850.0 ;
      RECT  115800.0 465150.0 125400.0 466050.0 ;
      RECT  115800.0 451350.0 125400.0 452250.0 ;
      RECT  127200.0 453750.0 128400.0 451350.0 ;
      RECT  127200.0 462450.0 128400.0 466050.0 ;
      RECT  132000.0 462450.0 133200.0 466050.0 ;
      RECT  134400.0 463650.0 135600.0 465600.0 ;
      RECT  134400.0 451800.0 135600.0 453750.0 ;
      RECT  127200.0 462450.0 128400.0 463650.0 ;
      RECT  129600.0 462450.0 130800.0 463650.0 ;
      RECT  129600.0 462450.0 130800.0 463650.0 ;
      RECT  127200.0 462450.0 128400.0 463650.0 ;
      RECT  129600.0 462450.0 130800.0 463650.0 ;
      RECT  132000.0 462450.0 133200.0 463650.0 ;
      RECT  132000.0 462450.0 133200.0 463650.0 ;
      RECT  129600.0 462450.0 130800.0 463650.0 ;
      RECT  127200.0 453750.0 128400.0 454950.0 ;
      RECT  129600.0 453750.0 130800.0 454950.0 ;
      RECT  129600.0 453750.0 130800.0 454950.0 ;
      RECT  127200.0 453750.0 128400.0 454950.0 ;
      RECT  129600.0 453750.0 130800.0 454950.0 ;
      RECT  132000.0 453750.0 133200.0 454950.0 ;
      RECT  132000.0 453750.0 133200.0 454950.0 ;
      RECT  129600.0 453750.0 130800.0 454950.0 ;
      RECT  134400.0 463050.0 135600.0 464250.0 ;
      RECT  134400.0 453150.0 135600.0 454350.0 ;
      RECT  132000.0 456300.0 130800.0 457500.0 ;
      RECT  129000.0 459000.0 127800.0 460200.0 ;
      RECT  129600.0 462450.0 130800.0 463650.0 ;
      RECT  132000.0 453750.0 133200.0 454950.0 ;
      RECT  133200.0 459000.0 132000.0 460200.0 ;
      RECT  127800.0 459000.0 129000.0 460200.0 ;
      RECT  130800.0 456300.0 132000.0 457500.0 ;
      RECT  132000.0 459000.0 133200.0 460200.0 ;
      RECT  125400.0 465150.0 139800.0 466050.0 ;
      RECT  125400.0 451350.0 139800.0 452250.0 ;
      RECT  146400.0 463650.0 147600.0 465600.0 ;
      RECT  146400.0 451800.0 147600.0 453750.0 ;
      RECT  141600.0 453150.0 142800.0 451350.0 ;
      RECT  141600.0 462450.0 142800.0 466050.0 ;
      RECT  144300.0 453150.0 145200.0 462450.0 ;
      RECT  141600.0 462450.0 142800.0 463650.0 ;
      RECT  144000.0 462450.0 145200.0 463650.0 ;
      RECT  144000.0 462450.0 145200.0 463650.0 ;
      RECT  141600.0 462450.0 142800.0 463650.0 ;
      RECT  141600.0 453150.0 142800.0 454350.0 ;
      RECT  144000.0 453150.0 145200.0 454350.0 ;
      RECT  144000.0 453150.0 145200.0 454350.0 ;
      RECT  141600.0 453150.0 142800.0 454350.0 ;
      RECT  146400.0 463050.0 147600.0 464250.0 ;
      RECT  146400.0 453150.0 147600.0 454350.0 ;
      RECT  142200.0 457800.0 143400.0 459000.0 ;
      RECT  142200.0 457800.0 143400.0 459000.0 ;
      RECT  144750.0 457950.0 145650.0 458850.0 ;
      RECT  139800.0 465150.0 149400.0 466050.0 ;
      RECT  139800.0 451350.0 149400.0 452250.0 ;
      RECT  112050.0 457800.0 113250.0 459000.0 ;
      RECT  114000.0 455400.0 115200.0 456600.0 ;
      RECT  130800.0 456300.0 129600.0 457500.0 ;
      RECT  122400.0 467550.0 123600.0 465600.0 ;
      RECT  122400.0 479400.0 123600.0 477450.0 ;
      RECT  117600.0 478050.0 118800.0 479850.0 ;
      RECT  117600.0 468750.0 118800.0 465150.0 ;
      RECT  120300.0 478050.0 121200.0 468750.0 ;
      RECT  117600.0 468750.0 118800.0 467550.0 ;
      RECT  120000.0 468750.0 121200.0 467550.0 ;
      RECT  120000.0 468750.0 121200.0 467550.0 ;
      RECT  117600.0 468750.0 118800.0 467550.0 ;
      RECT  117600.0 478050.0 118800.0 476850.0 ;
      RECT  120000.0 478050.0 121200.0 476850.0 ;
      RECT  120000.0 478050.0 121200.0 476850.0 ;
      RECT  117600.0 478050.0 118800.0 476850.0 ;
      RECT  122400.0 468150.0 123600.0 466950.0 ;
      RECT  122400.0 478050.0 123600.0 476850.0 ;
      RECT  118200.0 473400.0 119400.0 472200.0 ;
      RECT  118200.0 473400.0 119400.0 472200.0 ;
      RECT  120750.0 473250.0 121650.0 472350.0 ;
      RECT  115800.0 466050.0 125400.0 465150.0 ;
      RECT  115800.0 479850.0 125400.0 478950.0 ;
      RECT  127200.0 477450.0 128400.0 479850.0 ;
      RECT  127200.0 468750.0 128400.0 465150.0 ;
      RECT  132000.0 468750.0 133200.0 465150.0 ;
      RECT  134400.0 467550.0 135600.0 465600.0 ;
      RECT  134400.0 479400.0 135600.0 477450.0 ;
      RECT  127200.0 468750.0 128400.0 467550.0 ;
      RECT  129600.0 468750.0 130800.0 467550.0 ;
      RECT  129600.0 468750.0 130800.0 467550.0 ;
      RECT  127200.0 468750.0 128400.0 467550.0 ;
      RECT  129600.0 468750.0 130800.0 467550.0 ;
      RECT  132000.0 468750.0 133200.0 467550.0 ;
      RECT  132000.0 468750.0 133200.0 467550.0 ;
      RECT  129600.0 468750.0 130800.0 467550.0 ;
      RECT  127200.0 477450.0 128400.0 476250.0 ;
      RECT  129600.0 477450.0 130800.0 476250.0 ;
      RECT  129600.0 477450.0 130800.0 476250.0 ;
      RECT  127200.0 477450.0 128400.0 476250.0 ;
      RECT  129600.0 477450.0 130800.0 476250.0 ;
      RECT  132000.0 477450.0 133200.0 476250.0 ;
      RECT  132000.0 477450.0 133200.0 476250.0 ;
      RECT  129600.0 477450.0 130800.0 476250.0 ;
      RECT  134400.0 468150.0 135600.0 466950.0 ;
      RECT  134400.0 478050.0 135600.0 476850.0 ;
      RECT  132000.0 474900.0 130800.0 473700.0 ;
      RECT  129000.0 472200.0 127800.0 471000.0 ;
      RECT  129600.0 468750.0 130800.0 467550.0 ;
      RECT  132000.0 477450.0 133200.0 476250.0 ;
      RECT  133200.0 472200.0 132000.0 471000.0 ;
      RECT  127800.0 472200.0 129000.0 471000.0 ;
      RECT  130800.0 474900.0 132000.0 473700.0 ;
      RECT  132000.0 472200.0 133200.0 471000.0 ;
      RECT  125400.0 466050.0 139800.0 465150.0 ;
      RECT  125400.0 479850.0 139800.0 478950.0 ;
      RECT  146400.0 467550.0 147600.0 465600.0 ;
      RECT  146400.0 479400.0 147600.0 477450.0 ;
      RECT  141600.0 478050.0 142800.0 479850.0 ;
      RECT  141600.0 468750.0 142800.0 465150.0 ;
      RECT  144300.0 478050.0 145200.0 468750.0 ;
      RECT  141600.0 468750.0 142800.0 467550.0 ;
      RECT  144000.0 468750.0 145200.0 467550.0 ;
      RECT  144000.0 468750.0 145200.0 467550.0 ;
      RECT  141600.0 468750.0 142800.0 467550.0 ;
      RECT  141600.0 478050.0 142800.0 476850.0 ;
      RECT  144000.0 478050.0 145200.0 476850.0 ;
      RECT  144000.0 478050.0 145200.0 476850.0 ;
      RECT  141600.0 478050.0 142800.0 476850.0 ;
      RECT  146400.0 468150.0 147600.0 466950.0 ;
      RECT  146400.0 478050.0 147600.0 476850.0 ;
      RECT  142200.0 473400.0 143400.0 472200.0 ;
      RECT  142200.0 473400.0 143400.0 472200.0 ;
      RECT  144750.0 473250.0 145650.0 472350.0 ;
      RECT  139800.0 466050.0 149400.0 465150.0 ;
      RECT  139800.0 479850.0 149400.0 478950.0 ;
      RECT  112050.0 472200.0 113250.0 473400.0 ;
      RECT  114000.0 474600.0 115200.0 475800.0 ;
      RECT  130800.0 473700.0 129600.0 474900.0 ;
      RECT  122400.0 491250.0 123600.0 493200.0 ;
      RECT  122400.0 479400.0 123600.0 481350.0 ;
      RECT  117600.0 480750.0 118800.0 478950.0 ;
      RECT  117600.0 490050.0 118800.0 493650.0 ;
      RECT  120300.0 480750.0 121200.0 490050.0 ;
      RECT  117600.0 490050.0 118800.0 491250.0 ;
      RECT  120000.0 490050.0 121200.0 491250.0 ;
      RECT  120000.0 490050.0 121200.0 491250.0 ;
      RECT  117600.0 490050.0 118800.0 491250.0 ;
      RECT  117600.0 480750.0 118800.0 481950.0 ;
      RECT  120000.0 480750.0 121200.0 481950.0 ;
      RECT  120000.0 480750.0 121200.0 481950.0 ;
      RECT  117600.0 480750.0 118800.0 481950.0 ;
      RECT  122400.0 490650.0 123600.0 491850.0 ;
      RECT  122400.0 480750.0 123600.0 481950.0 ;
      RECT  118200.0 485400.0 119400.0 486600.0 ;
      RECT  118200.0 485400.0 119400.0 486600.0 ;
      RECT  120750.0 485550.0 121650.0 486450.0 ;
      RECT  115800.0 492750.0 125400.0 493650.0 ;
      RECT  115800.0 478950.0 125400.0 479850.0 ;
      RECT  127200.0 481350.0 128400.0 478950.0 ;
      RECT  127200.0 490050.0 128400.0 493650.0 ;
      RECT  132000.0 490050.0 133200.0 493650.0 ;
      RECT  134400.0 491250.0 135600.0 493200.0 ;
      RECT  134400.0 479400.0 135600.0 481350.0 ;
      RECT  127200.0 490050.0 128400.0 491250.0 ;
      RECT  129600.0 490050.0 130800.0 491250.0 ;
      RECT  129600.0 490050.0 130800.0 491250.0 ;
      RECT  127200.0 490050.0 128400.0 491250.0 ;
      RECT  129600.0 490050.0 130800.0 491250.0 ;
      RECT  132000.0 490050.0 133200.0 491250.0 ;
      RECT  132000.0 490050.0 133200.0 491250.0 ;
      RECT  129600.0 490050.0 130800.0 491250.0 ;
      RECT  127200.0 481350.0 128400.0 482550.0 ;
      RECT  129600.0 481350.0 130800.0 482550.0 ;
      RECT  129600.0 481350.0 130800.0 482550.0 ;
      RECT  127200.0 481350.0 128400.0 482550.0 ;
      RECT  129600.0 481350.0 130800.0 482550.0 ;
      RECT  132000.0 481350.0 133200.0 482550.0 ;
      RECT  132000.0 481350.0 133200.0 482550.0 ;
      RECT  129600.0 481350.0 130800.0 482550.0 ;
      RECT  134400.0 490650.0 135600.0 491850.0 ;
      RECT  134400.0 480750.0 135600.0 481950.0 ;
      RECT  132000.0 483900.0 130800.0 485100.0 ;
      RECT  129000.0 486600.0 127800.0 487800.0 ;
      RECT  129600.0 490050.0 130800.0 491250.0 ;
      RECT  132000.0 481350.0 133200.0 482550.0 ;
      RECT  133200.0 486600.0 132000.0 487800.0 ;
      RECT  127800.0 486600.0 129000.0 487800.0 ;
      RECT  130800.0 483900.0 132000.0 485100.0 ;
      RECT  132000.0 486600.0 133200.0 487800.0 ;
      RECT  125400.0 492750.0 139800.0 493650.0 ;
      RECT  125400.0 478950.0 139800.0 479850.0 ;
      RECT  146400.0 491250.0 147600.0 493200.0 ;
      RECT  146400.0 479400.0 147600.0 481350.0 ;
      RECT  141600.0 480750.0 142800.0 478950.0 ;
      RECT  141600.0 490050.0 142800.0 493650.0 ;
      RECT  144300.0 480750.0 145200.0 490050.0 ;
      RECT  141600.0 490050.0 142800.0 491250.0 ;
      RECT  144000.0 490050.0 145200.0 491250.0 ;
      RECT  144000.0 490050.0 145200.0 491250.0 ;
      RECT  141600.0 490050.0 142800.0 491250.0 ;
      RECT  141600.0 480750.0 142800.0 481950.0 ;
      RECT  144000.0 480750.0 145200.0 481950.0 ;
      RECT  144000.0 480750.0 145200.0 481950.0 ;
      RECT  141600.0 480750.0 142800.0 481950.0 ;
      RECT  146400.0 490650.0 147600.0 491850.0 ;
      RECT  146400.0 480750.0 147600.0 481950.0 ;
      RECT  142200.0 485400.0 143400.0 486600.0 ;
      RECT  142200.0 485400.0 143400.0 486600.0 ;
      RECT  144750.0 485550.0 145650.0 486450.0 ;
      RECT  139800.0 492750.0 149400.0 493650.0 ;
      RECT  139800.0 478950.0 149400.0 479850.0 ;
      RECT  112050.0 485400.0 113250.0 486600.0 ;
      RECT  114000.0 483000.0 115200.0 484200.0 ;
      RECT  130800.0 483900.0 129600.0 485100.0 ;
      RECT  122400.0 495150.0 123600.0 493200.0 ;
      RECT  122400.0 507000.0 123600.0 505050.0 ;
      RECT  117600.0 505650.0 118800.0 507450.0 ;
      RECT  117600.0 496350.0 118800.0 492750.0 ;
      RECT  120300.0 505650.0 121200.0 496350.0 ;
      RECT  117600.0 496350.0 118800.0 495150.0 ;
      RECT  120000.0 496350.0 121200.0 495150.0 ;
      RECT  120000.0 496350.0 121200.0 495150.0 ;
      RECT  117600.0 496350.0 118800.0 495150.0 ;
      RECT  117600.0 505650.0 118800.0 504450.0 ;
      RECT  120000.0 505650.0 121200.0 504450.0 ;
      RECT  120000.0 505650.0 121200.0 504450.0 ;
      RECT  117600.0 505650.0 118800.0 504450.0 ;
      RECT  122400.0 495750.0 123600.0 494550.0 ;
      RECT  122400.0 505650.0 123600.0 504450.0 ;
      RECT  118200.0 501000.0 119400.0 499800.0 ;
      RECT  118200.0 501000.0 119400.0 499800.0 ;
      RECT  120750.0 500850.0 121650.0 499950.0 ;
      RECT  115800.0 493650.0 125400.0 492750.0 ;
      RECT  115800.0 507450.0 125400.0 506550.0 ;
      RECT  127200.0 505050.0 128400.0 507450.0 ;
      RECT  127200.0 496350.0 128400.0 492750.0 ;
      RECT  132000.0 496350.0 133200.0 492750.0 ;
      RECT  134400.0 495150.0 135600.0 493200.0 ;
      RECT  134400.0 507000.0 135600.0 505050.0 ;
      RECT  127200.0 496350.0 128400.0 495150.0 ;
      RECT  129600.0 496350.0 130800.0 495150.0 ;
      RECT  129600.0 496350.0 130800.0 495150.0 ;
      RECT  127200.0 496350.0 128400.0 495150.0 ;
      RECT  129600.0 496350.0 130800.0 495150.0 ;
      RECT  132000.0 496350.0 133200.0 495150.0 ;
      RECT  132000.0 496350.0 133200.0 495150.0 ;
      RECT  129600.0 496350.0 130800.0 495150.0 ;
      RECT  127200.0 505050.0 128400.0 503850.0 ;
      RECT  129600.0 505050.0 130800.0 503850.0 ;
      RECT  129600.0 505050.0 130800.0 503850.0 ;
      RECT  127200.0 505050.0 128400.0 503850.0 ;
      RECT  129600.0 505050.0 130800.0 503850.0 ;
      RECT  132000.0 505050.0 133200.0 503850.0 ;
      RECT  132000.0 505050.0 133200.0 503850.0 ;
      RECT  129600.0 505050.0 130800.0 503850.0 ;
      RECT  134400.0 495750.0 135600.0 494550.0 ;
      RECT  134400.0 505650.0 135600.0 504450.0 ;
      RECT  132000.0 502500.0 130800.0 501300.0 ;
      RECT  129000.0 499800.0 127800.0 498600.0 ;
      RECT  129600.0 496350.0 130800.0 495150.0 ;
      RECT  132000.0 505050.0 133200.0 503850.0 ;
      RECT  133200.0 499800.0 132000.0 498600.0 ;
      RECT  127800.0 499800.0 129000.0 498600.0 ;
      RECT  130800.0 502500.0 132000.0 501300.0 ;
      RECT  132000.0 499800.0 133200.0 498600.0 ;
      RECT  125400.0 493650.0 139800.0 492750.0 ;
      RECT  125400.0 507450.0 139800.0 506550.0 ;
      RECT  146400.0 495150.0 147600.0 493200.0 ;
      RECT  146400.0 507000.0 147600.0 505050.0 ;
      RECT  141600.0 505650.0 142800.0 507450.0 ;
      RECT  141600.0 496350.0 142800.0 492750.0 ;
      RECT  144300.0 505650.0 145200.0 496350.0 ;
      RECT  141600.0 496350.0 142800.0 495150.0 ;
      RECT  144000.0 496350.0 145200.0 495150.0 ;
      RECT  144000.0 496350.0 145200.0 495150.0 ;
      RECT  141600.0 496350.0 142800.0 495150.0 ;
      RECT  141600.0 505650.0 142800.0 504450.0 ;
      RECT  144000.0 505650.0 145200.0 504450.0 ;
      RECT  144000.0 505650.0 145200.0 504450.0 ;
      RECT  141600.0 505650.0 142800.0 504450.0 ;
      RECT  146400.0 495750.0 147600.0 494550.0 ;
      RECT  146400.0 505650.0 147600.0 504450.0 ;
      RECT  142200.0 501000.0 143400.0 499800.0 ;
      RECT  142200.0 501000.0 143400.0 499800.0 ;
      RECT  144750.0 500850.0 145650.0 499950.0 ;
      RECT  139800.0 493650.0 149400.0 492750.0 ;
      RECT  139800.0 507450.0 149400.0 506550.0 ;
      RECT  112050.0 499800.0 113250.0 501000.0 ;
      RECT  114000.0 502200.0 115200.0 503400.0 ;
      RECT  130800.0 501300.0 129600.0 502500.0 ;
      RECT  122400.0 518850.0 123600.0 520800.0 ;
      RECT  122400.0 507000.0 123600.0 508950.0 ;
      RECT  117600.0 508350.0 118800.0 506550.0 ;
      RECT  117600.0 517650.0 118800.0 521250.0 ;
      RECT  120300.0 508350.0 121200.0 517650.0 ;
      RECT  117600.0 517650.0 118800.0 518850.0 ;
      RECT  120000.0 517650.0 121200.0 518850.0 ;
      RECT  120000.0 517650.0 121200.0 518850.0 ;
      RECT  117600.0 517650.0 118800.0 518850.0 ;
      RECT  117600.0 508350.0 118800.0 509550.0 ;
      RECT  120000.0 508350.0 121200.0 509550.0 ;
      RECT  120000.0 508350.0 121200.0 509550.0 ;
      RECT  117600.0 508350.0 118800.0 509550.0 ;
      RECT  122400.0 518250.0 123600.0 519450.0 ;
      RECT  122400.0 508350.0 123600.0 509550.0 ;
      RECT  118200.0 513000.0 119400.0 514200.0 ;
      RECT  118200.0 513000.0 119400.0 514200.0 ;
      RECT  120750.0 513150.0 121650.0 514050.0 ;
      RECT  115800.0 520350.0 125400.0 521250.0 ;
      RECT  115800.0 506550.0 125400.0 507450.0 ;
      RECT  127200.0 508950.0 128400.0 506550.0 ;
      RECT  127200.0 517650.0 128400.0 521250.0 ;
      RECT  132000.0 517650.0 133200.0 521250.0 ;
      RECT  134400.0 518850.0 135600.0 520800.0 ;
      RECT  134400.0 507000.0 135600.0 508950.0 ;
      RECT  127200.0 517650.0 128400.0 518850.0 ;
      RECT  129600.0 517650.0 130800.0 518850.0 ;
      RECT  129600.0 517650.0 130800.0 518850.0 ;
      RECT  127200.0 517650.0 128400.0 518850.0 ;
      RECT  129600.0 517650.0 130800.0 518850.0 ;
      RECT  132000.0 517650.0 133200.0 518850.0 ;
      RECT  132000.0 517650.0 133200.0 518850.0 ;
      RECT  129600.0 517650.0 130800.0 518850.0 ;
      RECT  127200.0 508950.0 128400.0 510150.0 ;
      RECT  129600.0 508950.0 130800.0 510150.0 ;
      RECT  129600.0 508950.0 130800.0 510150.0 ;
      RECT  127200.0 508950.0 128400.0 510150.0 ;
      RECT  129600.0 508950.0 130800.0 510150.0 ;
      RECT  132000.0 508950.0 133200.0 510150.0 ;
      RECT  132000.0 508950.0 133200.0 510150.0 ;
      RECT  129600.0 508950.0 130800.0 510150.0 ;
      RECT  134400.0 518250.0 135600.0 519450.0 ;
      RECT  134400.0 508350.0 135600.0 509550.0 ;
      RECT  132000.0 511500.0 130800.0 512700.0 ;
      RECT  129000.0 514200.0 127800.0 515400.0 ;
      RECT  129600.0 517650.0 130800.0 518850.0 ;
      RECT  132000.0 508950.0 133200.0 510150.0 ;
      RECT  133200.0 514200.0 132000.0 515400.0 ;
      RECT  127800.0 514200.0 129000.0 515400.0 ;
      RECT  130800.0 511500.0 132000.0 512700.0 ;
      RECT  132000.0 514200.0 133200.0 515400.0 ;
      RECT  125400.0 520350.0 139800.0 521250.0 ;
      RECT  125400.0 506550.0 139800.0 507450.0 ;
      RECT  146400.0 518850.0 147600.0 520800.0 ;
      RECT  146400.0 507000.0 147600.0 508950.0 ;
      RECT  141600.0 508350.0 142800.0 506550.0 ;
      RECT  141600.0 517650.0 142800.0 521250.0 ;
      RECT  144300.0 508350.0 145200.0 517650.0 ;
      RECT  141600.0 517650.0 142800.0 518850.0 ;
      RECT  144000.0 517650.0 145200.0 518850.0 ;
      RECT  144000.0 517650.0 145200.0 518850.0 ;
      RECT  141600.0 517650.0 142800.0 518850.0 ;
      RECT  141600.0 508350.0 142800.0 509550.0 ;
      RECT  144000.0 508350.0 145200.0 509550.0 ;
      RECT  144000.0 508350.0 145200.0 509550.0 ;
      RECT  141600.0 508350.0 142800.0 509550.0 ;
      RECT  146400.0 518250.0 147600.0 519450.0 ;
      RECT  146400.0 508350.0 147600.0 509550.0 ;
      RECT  142200.0 513000.0 143400.0 514200.0 ;
      RECT  142200.0 513000.0 143400.0 514200.0 ;
      RECT  144750.0 513150.0 145650.0 514050.0 ;
      RECT  139800.0 520350.0 149400.0 521250.0 ;
      RECT  139800.0 506550.0 149400.0 507450.0 ;
      RECT  112050.0 513000.0 113250.0 514200.0 ;
      RECT  114000.0 510600.0 115200.0 511800.0 ;
      RECT  130800.0 511500.0 129600.0 512700.0 ;
      RECT  122400.0 522750.0 123600.0 520800.0 ;
      RECT  122400.0 534600.0 123600.0 532650.0 ;
      RECT  117600.0 533250.0 118800.0 535050.0 ;
      RECT  117600.0 523950.0 118800.0 520350.0 ;
      RECT  120300.0 533250.0 121200.0 523950.0 ;
      RECT  117600.0 523950.0 118800.0 522750.0 ;
      RECT  120000.0 523950.0 121200.0 522750.0 ;
      RECT  120000.0 523950.0 121200.0 522750.0 ;
      RECT  117600.0 523950.0 118800.0 522750.0 ;
      RECT  117600.0 533250.0 118800.0 532050.0 ;
      RECT  120000.0 533250.0 121200.0 532050.0 ;
      RECT  120000.0 533250.0 121200.0 532050.0 ;
      RECT  117600.0 533250.0 118800.0 532050.0 ;
      RECT  122400.0 523350.0 123600.0 522150.0 ;
      RECT  122400.0 533250.0 123600.0 532050.0 ;
      RECT  118200.0 528600.0 119400.0 527400.0 ;
      RECT  118200.0 528600.0 119400.0 527400.0 ;
      RECT  120750.0 528450.0 121650.0 527550.0 ;
      RECT  115800.0 521250.0 125400.0 520350.0 ;
      RECT  115800.0 535050.0 125400.0 534150.0 ;
      RECT  127200.0 532650.0 128400.0 535050.0 ;
      RECT  127200.0 523950.0 128400.0 520350.0 ;
      RECT  132000.0 523950.0 133200.0 520350.0 ;
      RECT  134400.0 522750.0 135600.0 520800.0 ;
      RECT  134400.0 534600.0 135600.0 532650.0 ;
      RECT  127200.0 523950.0 128400.0 522750.0 ;
      RECT  129600.0 523950.0 130800.0 522750.0 ;
      RECT  129600.0 523950.0 130800.0 522750.0 ;
      RECT  127200.0 523950.0 128400.0 522750.0 ;
      RECT  129600.0 523950.0 130800.0 522750.0 ;
      RECT  132000.0 523950.0 133200.0 522750.0 ;
      RECT  132000.0 523950.0 133200.0 522750.0 ;
      RECT  129600.0 523950.0 130800.0 522750.0 ;
      RECT  127200.0 532650.0 128400.0 531450.0 ;
      RECT  129600.0 532650.0 130800.0 531450.0 ;
      RECT  129600.0 532650.0 130800.0 531450.0 ;
      RECT  127200.0 532650.0 128400.0 531450.0 ;
      RECT  129600.0 532650.0 130800.0 531450.0 ;
      RECT  132000.0 532650.0 133200.0 531450.0 ;
      RECT  132000.0 532650.0 133200.0 531450.0 ;
      RECT  129600.0 532650.0 130800.0 531450.0 ;
      RECT  134400.0 523350.0 135600.0 522150.0 ;
      RECT  134400.0 533250.0 135600.0 532050.0 ;
      RECT  132000.0 530100.0 130800.0 528900.0 ;
      RECT  129000.0 527400.0 127800.0 526200.0 ;
      RECT  129600.0 523950.0 130800.0 522750.0 ;
      RECT  132000.0 532650.0 133200.0 531450.0 ;
      RECT  133200.0 527400.0 132000.0 526200.0 ;
      RECT  127800.0 527400.0 129000.0 526200.0 ;
      RECT  130800.0 530100.0 132000.0 528900.0 ;
      RECT  132000.0 527400.0 133200.0 526200.0 ;
      RECT  125400.0 521250.0 139800.0 520350.0 ;
      RECT  125400.0 535050.0 139800.0 534150.0 ;
      RECT  146400.0 522750.0 147600.0 520800.0 ;
      RECT  146400.0 534600.0 147600.0 532650.0 ;
      RECT  141600.0 533250.0 142800.0 535050.0 ;
      RECT  141600.0 523950.0 142800.0 520350.0 ;
      RECT  144300.0 533250.0 145200.0 523950.0 ;
      RECT  141600.0 523950.0 142800.0 522750.0 ;
      RECT  144000.0 523950.0 145200.0 522750.0 ;
      RECT  144000.0 523950.0 145200.0 522750.0 ;
      RECT  141600.0 523950.0 142800.0 522750.0 ;
      RECT  141600.0 533250.0 142800.0 532050.0 ;
      RECT  144000.0 533250.0 145200.0 532050.0 ;
      RECT  144000.0 533250.0 145200.0 532050.0 ;
      RECT  141600.0 533250.0 142800.0 532050.0 ;
      RECT  146400.0 523350.0 147600.0 522150.0 ;
      RECT  146400.0 533250.0 147600.0 532050.0 ;
      RECT  142200.0 528600.0 143400.0 527400.0 ;
      RECT  142200.0 528600.0 143400.0 527400.0 ;
      RECT  144750.0 528450.0 145650.0 527550.0 ;
      RECT  139800.0 521250.0 149400.0 520350.0 ;
      RECT  139800.0 535050.0 149400.0 534150.0 ;
      RECT  112050.0 527400.0 113250.0 528600.0 ;
      RECT  114000.0 529800.0 115200.0 531000.0 ;
      RECT  130800.0 528900.0 129600.0 530100.0 ;
      RECT  122400.0 546450.0 123600.0 548400.0 ;
      RECT  122400.0 534600.0 123600.0 536550.0 ;
      RECT  117600.0 535950.0 118800.0 534150.0 ;
      RECT  117600.0 545250.0 118800.0 548850.0 ;
      RECT  120300.0 535950.0 121200.0 545250.0 ;
      RECT  117600.0 545250.0 118800.0 546450.0 ;
      RECT  120000.0 545250.0 121200.0 546450.0 ;
      RECT  120000.0 545250.0 121200.0 546450.0 ;
      RECT  117600.0 545250.0 118800.0 546450.0 ;
      RECT  117600.0 535950.0 118800.0 537150.0 ;
      RECT  120000.0 535950.0 121200.0 537150.0 ;
      RECT  120000.0 535950.0 121200.0 537150.0 ;
      RECT  117600.0 535950.0 118800.0 537150.0 ;
      RECT  122400.0 545850.0 123600.0 547050.0 ;
      RECT  122400.0 535950.0 123600.0 537150.0 ;
      RECT  118200.0 540600.0 119400.0 541800.0 ;
      RECT  118200.0 540600.0 119400.0 541800.0 ;
      RECT  120750.0 540750.0 121650.0 541650.0 ;
      RECT  115800.0 547950.0 125400.0 548850.0 ;
      RECT  115800.0 534150.0 125400.0 535050.0 ;
      RECT  127200.0 536550.0 128400.0 534150.0 ;
      RECT  127200.0 545250.0 128400.0 548850.0 ;
      RECT  132000.0 545250.0 133200.0 548850.0 ;
      RECT  134400.0 546450.0 135600.0 548400.0 ;
      RECT  134400.0 534600.0 135600.0 536550.0 ;
      RECT  127200.0 545250.0 128400.0 546450.0 ;
      RECT  129600.0 545250.0 130800.0 546450.0 ;
      RECT  129600.0 545250.0 130800.0 546450.0 ;
      RECT  127200.0 545250.0 128400.0 546450.0 ;
      RECT  129600.0 545250.0 130800.0 546450.0 ;
      RECT  132000.0 545250.0 133200.0 546450.0 ;
      RECT  132000.0 545250.0 133200.0 546450.0 ;
      RECT  129600.0 545250.0 130800.0 546450.0 ;
      RECT  127200.0 536550.0 128400.0 537750.0 ;
      RECT  129600.0 536550.0 130800.0 537750.0 ;
      RECT  129600.0 536550.0 130800.0 537750.0 ;
      RECT  127200.0 536550.0 128400.0 537750.0 ;
      RECT  129600.0 536550.0 130800.0 537750.0 ;
      RECT  132000.0 536550.0 133200.0 537750.0 ;
      RECT  132000.0 536550.0 133200.0 537750.0 ;
      RECT  129600.0 536550.0 130800.0 537750.0 ;
      RECT  134400.0 545850.0 135600.0 547050.0 ;
      RECT  134400.0 535950.0 135600.0 537150.0 ;
      RECT  132000.0 539100.0 130800.0 540300.0 ;
      RECT  129000.0 541800.0 127800.0 543000.0 ;
      RECT  129600.0 545250.0 130800.0 546450.0 ;
      RECT  132000.0 536550.0 133200.0 537750.0 ;
      RECT  133200.0 541800.0 132000.0 543000.0 ;
      RECT  127800.0 541800.0 129000.0 543000.0 ;
      RECT  130800.0 539100.0 132000.0 540300.0 ;
      RECT  132000.0 541800.0 133200.0 543000.0 ;
      RECT  125400.0 547950.0 139800.0 548850.0 ;
      RECT  125400.0 534150.0 139800.0 535050.0 ;
      RECT  146400.0 546450.0 147600.0 548400.0 ;
      RECT  146400.0 534600.0 147600.0 536550.0 ;
      RECT  141600.0 535950.0 142800.0 534150.0 ;
      RECT  141600.0 545250.0 142800.0 548850.0 ;
      RECT  144300.0 535950.0 145200.0 545250.0 ;
      RECT  141600.0 545250.0 142800.0 546450.0 ;
      RECT  144000.0 545250.0 145200.0 546450.0 ;
      RECT  144000.0 545250.0 145200.0 546450.0 ;
      RECT  141600.0 545250.0 142800.0 546450.0 ;
      RECT  141600.0 535950.0 142800.0 537150.0 ;
      RECT  144000.0 535950.0 145200.0 537150.0 ;
      RECT  144000.0 535950.0 145200.0 537150.0 ;
      RECT  141600.0 535950.0 142800.0 537150.0 ;
      RECT  146400.0 545850.0 147600.0 547050.0 ;
      RECT  146400.0 535950.0 147600.0 537150.0 ;
      RECT  142200.0 540600.0 143400.0 541800.0 ;
      RECT  142200.0 540600.0 143400.0 541800.0 ;
      RECT  144750.0 540750.0 145650.0 541650.0 ;
      RECT  139800.0 547950.0 149400.0 548850.0 ;
      RECT  139800.0 534150.0 149400.0 535050.0 ;
      RECT  112050.0 540600.0 113250.0 541800.0 ;
      RECT  114000.0 538200.0 115200.0 539400.0 ;
      RECT  130800.0 539100.0 129600.0 540300.0 ;
      RECT  122400.0 550350.0 123600.0 548400.0 ;
      RECT  122400.0 562200.0 123600.0 560250.0 ;
      RECT  117600.0 560850.0 118800.0 562650.0 ;
      RECT  117600.0 551550.0 118800.0 547950.0 ;
      RECT  120300.0 560850.0 121200.0 551550.0 ;
      RECT  117600.0 551550.0 118800.0 550350.0 ;
      RECT  120000.0 551550.0 121200.0 550350.0 ;
      RECT  120000.0 551550.0 121200.0 550350.0 ;
      RECT  117600.0 551550.0 118800.0 550350.0 ;
      RECT  117600.0 560850.0 118800.0 559650.0 ;
      RECT  120000.0 560850.0 121200.0 559650.0 ;
      RECT  120000.0 560850.0 121200.0 559650.0 ;
      RECT  117600.0 560850.0 118800.0 559650.0 ;
      RECT  122400.0 550950.0 123600.0 549750.0 ;
      RECT  122400.0 560850.0 123600.0 559650.0 ;
      RECT  118200.0 556200.0 119400.0 555000.0 ;
      RECT  118200.0 556200.0 119400.0 555000.0 ;
      RECT  120750.0 556050.0 121650.0 555150.0 ;
      RECT  115800.0 548850.0 125400.0 547950.0 ;
      RECT  115800.0 562650.0 125400.0 561750.0 ;
      RECT  127200.0 560250.0 128400.0 562650.0 ;
      RECT  127200.0 551550.0 128400.0 547950.0 ;
      RECT  132000.0 551550.0 133200.0 547950.0 ;
      RECT  134400.0 550350.0 135600.0 548400.0 ;
      RECT  134400.0 562200.0 135600.0 560250.0 ;
      RECT  127200.0 551550.0 128400.0 550350.0 ;
      RECT  129600.0 551550.0 130800.0 550350.0 ;
      RECT  129600.0 551550.0 130800.0 550350.0 ;
      RECT  127200.0 551550.0 128400.0 550350.0 ;
      RECT  129600.0 551550.0 130800.0 550350.0 ;
      RECT  132000.0 551550.0 133200.0 550350.0 ;
      RECT  132000.0 551550.0 133200.0 550350.0 ;
      RECT  129600.0 551550.0 130800.0 550350.0 ;
      RECT  127200.0 560250.0 128400.0 559050.0 ;
      RECT  129600.0 560250.0 130800.0 559050.0 ;
      RECT  129600.0 560250.0 130800.0 559050.0 ;
      RECT  127200.0 560250.0 128400.0 559050.0 ;
      RECT  129600.0 560250.0 130800.0 559050.0 ;
      RECT  132000.0 560250.0 133200.0 559050.0 ;
      RECT  132000.0 560250.0 133200.0 559050.0 ;
      RECT  129600.0 560250.0 130800.0 559050.0 ;
      RECT  134400.0 550950.0 135600.0 549750.0 ;
      RECT  134400.0 560850.0 135600.0 559650.0 ;
      RECT  132000.0 557700.0 130800.0 556500.0 ;
      RECT  129000.0 555000.0 127800.0 553800.0 ;
      RECT  129600.0 551550.0 130800.0 550350.0 ;
      RECT  132000.0 560250.0 133200.0 559050.0 ;
      RECT  133200.0 555000.0 132000.0 553800.0 ;
      RECT  127800.0 555000.0 129000.0 553800.0 ;
      RECT  130800.0 557700.0 132000.0 556500.0 ;
      RECT  132000.0 555000.0 133200.0 553800.0 ;
      RECT  125400.0 548850.0 139800.0 547950.0 ;
      RECT  125400.0 562650.0 139800.0 561750.0 ;
      RECT  146400.0 550350.0 147600.0 548400.0 ;
      RECT  146400.0 562200.0 147600.0 560250.0 ;
      RECT  141600.0 560850.0 142800.0 562650.0 ;
      RECT  141600.0 551550.0 142800.0 547950.0 ;
      RECT  144300.0 560850.0 145200.0 551550.0 ;
      RECT  141600.0 551550.0 142800.0 550350.0 ;
      RECT  144000.0 551550.0 145200.0 550350.0 ;
      RECT  144000.0 551550.0 145200.0 550350.0 ;
      RECT  141600.0 551550.0 142800.0 550350.0 ;
      RECT  141600.0 560850.0 142800.0 559650.0 ;
      RECT  144000.0 560850.0 145200.0 559650.0 ;
      RECT  144000.0 560850.0 145200.0 559650.0 ;
      RECT  141600.0 560850.0 142800.0 559650.0 ;
      RECT  146400.0 550950.0 147600.0 549750.0 ;
      RECT  146400.0 560850.0 147600.0 559650.0 ;
      RECT  142200.0 556200.0 143400.0 555000.0 ;
      RECT  142200.0 556200.0 143400.0 555000.0 ;
      RECT  144750.0 556050.0 145650.0 555150.0 ;
      RECT  139800.0 548850.0 149400.0 547950.0 ;
      RECT  139800.0 562650.0 149400.0 561750.0 ;
      RECT  112050.0 555000.0 113250.0 556200.0 ;
      RECT  114000.0 557400.0 115200.0 558600.0 ;
      RECT  130800.0 556500.0 129600.0 557700.0 ;
      RECT  122400.0 574050.0 123600.0 576000.0 ;
      RECT  122400.0 562200.0 123600.0 564150.0 ;
      RECT  117600.0 563550.0 118800.0 561750.0 ;
      RECT  117600.0 572850.0 118800.0 576450.0 ;
      RECT  120300.0 563550.0 121200.0 572850.0 ;
      RECT  117600.0 572850.0 118800.0 574050.0 ;
      RECT  120000.0 572850.0 121200.0 574050.0 ;
      RECT  120000.0 572850.0 121200.0 574050.0 ;
      RECT  117600.0 572850.0 118800.0 574050.0 ;
      RECT  117600.0 563550.0 118800.0 564750.0 ;
      RECT  120000.0 563550.0 121200.0 564750.0 ;
      RECT  120000.0 563550.0 121200.0 564750.0 ;
      RECT  117600.0 563550.0 118800.0 564750.0 ;
      RECT  122400.0 573450.0 123600.0 574650.0 ;
      RECT  122400.0 563550.0 123600.0 564750.0 ;
      RECT  118200.0 568200.0 119400.0 569400.0 ;
      RECT  118200.0 568200.0 119400.0 569400.0 ;
      RECT  120750.0 568350.0 121650.0 569250.0 ;
      RECT  115800.0 575550.0 125400.0 576450.0 ;
      RECT  115800.0 561750.0 125400.0 562650.0 ;
      RECT  127200.0 564150.0 128400.0 561750.0 ;
      RECT  127200.0 572850.0 128400.0 576450.0 ;
      RECT  132000.0 572850.0 133200.0 576450.0 ;
      RECT  134400.0 574050.0 135600.0 576000.0 ;
      RECT  134400.0 562200.0 135600.0 564150.0 ;
      RECT  127200.0 572850.0 128400.0 574050.0 ;
      RECT  129600.0 572850.0 130800.0 574050.0 ;
      RECT  129600.0 572850.0 130800.0 574050.0 ;
      RECT  127200.0 572850.0 128400.0 574050.0 ;
      RECT  129600.0 572850.0 130800.0 574050.0 ;
      RECT  132000.0 572850.0 133200.0 574050.0 ;
      RECT  132000.0 572850.0 133200.0 574050.0 ;
      RECT  129600.0 572850.0 130800.0 574050.0 ;
      RECT  127200.0 564150.0 128400.0 565350.0 ;
      RECT  129600.0 564150.0 130800.0 565350.0 ;
      RECT  129600.0 564150.0 130800.0 565350.0 ;
      RECT  127200.0 564150.0 128400.0 565350.0 ;
      RECT  129600.0 564150.0 130800.0 565350.0 ;
      RECT  132000.0 564150.0 133200.0 565350.0 ;
      RECT  132000.0 564150.0 133200.0 565350.0 ;
      RECT  129600.0 564150.0 130800.0 565350.0 ;
      RECT  134400.0 573450.0 135600.0 574650.0 ;
      RECT  134400.0 563550.0 135600.0 564750.0 ;
      RECT  132000.0 566700.0 130800.0 567900.0 ;
      RECT  129000.0 569400.0 127800.0 570600.0 ;
      RECT  129600.0 572850.0 130800.0 574050.0 ;
      RECT  132000.0 564150.0 133200.0 565350.0 ;
      RECT  133200.0 569400.0 132000.0 570600.0 ;
      RECT  127800.0 569400.0 129000.0 570600.0 ;
      RECT  130800.0 566700.0 132000.0 567900.0 ;
      RECT  132000.0 569400.0 133200.0 570600.0 ;
      RECT  125400.0 575550.0 139800.0 576450.0 ;
      RECT  125400.0 561750.0 139800.0 562650.0 ;
      RECT  146400.0 574050.0 147600.0 576000.0 ;
      RECT  146400.0 562200.0 147600.0 564150.0 ;
      RECT  141600.0 563550.0 142800.0 561750.0 ;
      RECT  141600.0 572850.0 142800.0 576450.0 ;
      RECT  144300.0 563550.0 145200.0 572850.0 ;
      RECT  141600.0 572850.0 142800.0 574050.0 ;
      RECT  144000.0 572850.0 145200.0 574050.0 ;
      RECT  144000.0 572850.0 145200.0 574050.0 ;
      RECT  141600.0 572850.0 142800.0 574050.0 ;
      RECT  141600.0 563550.0 142800.0 564750.0 ;
      RECT  144000.0 563550.0 145200.0 564750.0 ;
      RECT  144000.0 563550.0 145200.0 564750.0 ;
      RECT  141600.0 563550.0 142800.0 564750.0 ;
      RECT  146400.0 573450.0 147600.0 574650.0 ;
      RECT  146400.0 563550.0 147600.0 564750.0 ;
      RECT  142200.0 568200.0 143400.0 569400.0 ;
      RECT  142200.0 568200.0 143400.0 569400.0 ;
      RECT  144750.0 568350.0 145650.0 569250.0 ;
      RECT  139800.0 575550.0 149400.0 576450.0 ;
      RECT  139800.0 561750.0 149400.0 562650.0 ;
      RECT  112050.0 568200.0 113250.0 569400.0 ;
      RECT  114000.0 565800.0 115200.0 567000.0 ;
      RECT  130800.0 566700.0 129600.0 567900.0 ;
      RECT  122400.0 577950.0 123600.0 576000.0 ;
      RECT  122400.0 589800.0 123600.0 587850.0 ;
      RECT  117600.0 588450.0 118800.0 590250.0 ;
      RECT  117600.0 579150.0 118800.0 575550.0 ;
      RECT  120300.0 588450.0 121200.0 579150.0 ;
      RECT  117600.0 579150.0 118800.0 577950.0 ;
      RECT  120000.0 579150.0 121200.0 577950.0 ;
      RECT  120000.0 579150.0 121200.0 577950.0 ;
      RECT  117600.0 579150.0 118800.0 577950.0 ;
      RECT  117600.0 588450.0 118800.0 587250.0 ;
      RECT  120000.0 588450.0 121200.0 587250.0 ;
      RECT  120000.0 588450.0 121200.0 587250.0 ;
      RECT  117600.0 588450.0 118800.0 587250.0 ;
      RECT  122400.0 578550.0 123600.0 577350.0 ;
      RECT  122400.0 588450.0 123600.0 587250.0 ;
      RECT  118200.0 583800.0 119400.0 582600.0 ;
      RECT  118200.0 583800.0 119400.0 582600.0 ;
      RECT  120750.0 583650.0 121650.0 582750.0 ;
      RECT  115800.0 576450.0 125400.0 575550.0 ;
      RECT  115800.0 590250.0 125400.0 589350.0 ;
      RECT  127200.0 587850.0 128400.0 590250.0 ;
      RECT  127200.0 579150.0 128400.0 575550.0 ;
      RECT  132000.0 579150.0 133200.0 575550.0 ;
      RECT  134400.0 577950.0 135600.0 576000.0 ;
      RECT  134400.0 589800.0 135600.0 587850.0 ;
      RECT  127200.0 579150.0 128400.0 577950.0 ;
      RECT  129600.0 579150.0 130800.0 577950.0 ;
      RECT  129600.0 579150.0 130800.0 577950.0 ;
      RECT  127200.0 579150.0 128400.0 577950.0 ;
      RECT  129600.0 579150.0 130800.0 577950.0 ;
      RECT  132000.0 579150.0 133200.0 577950.0 ;
      RECT  132000.0 579150.0 133200.0 577950.0 ;
      RECT  129600.0 579150.0 130800.0 577950.0 ;
      RECT  127200.0 587850.0 128400.0 586650.0 ;
      RECT  129600.0 587850.0 130800.0 586650.0 ;
      RECT  129600.0 587850.0 130800.0 586650.0 ;
      RECT  127200.0 587850.0 128400.0 586650.0 ;
      RECT  129600.0 587850.0 130800.0 586650.0 ;
      RECT  132000.0 587850.0 133200.0 586650.0 ;
      RECT  132000.0 587850.0 133200.0 586650.0 ;
      RECT  129600.0 587850.0 130800.0 586650.0 ;
      RECT  134400.0 578550.0 135600.0 577350.0 ;
      RECT  134400.0 588450.0 135600.0 587250.0 ;
      RECT  132000.0 585300.0 130800.0 584100.0 ;
      RECT  129000.0 582600.0 127800.0 581400.0 ;
      RECT  129600.0 579150.0 130800.0 577950.0 ;
      RECT  132000.0 587850.0 133200.0 586650.0 ;
      RECT  133200.0 582600.0 132000.0 581400.0 ;
      RECT  127800.0 582600.0 129000.0 581400.0 ;
      RECT  130800.0 585300.0 132000.0 584100.0 ;
      RECT  132000.0 582600.0 133200.0 581400.0 ;
      RECT  125400.0 576450.0 139800.0 575550.0 ;
      RECT  125400.0 590250.0 139800.0 589350.0 ;
      RECT  146400.0 577950.0 147600.0 576000.0 ;
      RECT  146400.0 589800.0 147600.0 587850.0 ;
      RECT  141600.0 588450.0 142800.0 590250.0 ;
      RECT  141600.0 579150.0 142800.0 575550.0 ;
      RECT  144300.0 588450.0 145200.0 579150.0 ;
      RECT  141600.0 579150.0 142800.0 577950.0 ;
      RECT  144000.0 579150.0 145200.0 577950.0 ;
      RECT  144000.0 579150.0 145200.0 577950.0 ;
      RECT  141600.0 579150.0 142800.0 577950.0 ;
      RECT  141600.0 588450.0 142800.0 587250.0 ;
      RECT  144000.0 588450.0 145200.0 587250.0 ;
      RECT  144000.0 588450.0 145200.0 587250.0 ;
      RECT  141600.0 588450.0 142800.0 587250.0 ;
      RECT  146400.0 578550.0 147600.0 577350.0 ;
      RECT  146400.0 588450.0 147600.0 587250.0 ;
      RECT  142200.0 583800.0 143400.0 582600.0 ;
      RECT  142200.0 583800.0 143400.0 582600.0 ;
      RECT  144750.0 583650.0 145650.0 582750.0 ;
      RECT  139800.0 576450.0 149400.0 575550.0 ;
      RECT  139800.0 590250.0 149400.0 589350.0 ;
      RECT  112050.0 582600.0 113250.0 583800.0 ;
      RECT  114000.0 585000.0 115200.0 586200.0 ;
      RECT  130800.0 584100.0 129600.0 585300.0 ;
      RECT  122400.0 601650.0 123600.0 603600.0 ;
      RECT  122400.0 589800.0 123600.0 591750.0 ;
      RECT  117600.0 591150.0 118800.0 589350.0 ;
      RECT  117600.0 600450.0 118800.0 604050.0 ;
      RECT  120300.0 591150.0 121200.0 600450.0 ;
      RECT  117600.0 600450.0 118800.0 601650.0 ;
      RECT  120000.0 600450.0 121200.0 601650.0 ;
      RECT  120000.0 600450.0 121200.0 601650.0 ;
      RECT  117600.0 600450.0 118800.0 601650.0 ;
      RECT  117600.0 591150.0 118800.0 592350.0 ;
      RECT  120000.0 591150.0 121200.0 592350.0 ;
      RECT  120000.0 591150.0 121200.0 592350.0 ;
      RECT  117600.0 591150.0 118800.0 592350.0 ;
      RECT  122400.0 601050.0 123600.0 602250.0 ;
      RECT  122400.0 591150.0 123600.0 592350.0 ;
      RECT  118200.0 595800.0 119400.0 597000.0 ;
      RECT  118200.0 595800.0 119400.0 597000.0 ;
      RECT  120750.0 595950.0 121650.0 596850.0 ;
      RECT  115800.0 603150.0 125400.0 604050.0 ;
      RECT  115800.0 589350.0 125400.0 590250.0 ;
      RECT  127200.0 591750.0 128400.0 589350.0 ;
      RECT  127200.0 600450.0 128400.0 604050.0 ;
      RECT  132000.0 600450.0 133200.0 604050.0 ;
      RECT  134400.0 601650.0 135600.0 603600.0 ;
      RECT  134400.0 589800.0 135600.0 591750.0 ;
      RECT  127200.0 600450.0 128400.0 601650.0 ;
      RECT  129600.0 600450.0 130800.0 601650.0 ;
      RECT  129600.0 600450.0 130800.0 601650.0 ;
      RECT  127200.0 600450.0 128400.0 601650.0 ;
      RECT  129600.0 600450.0 130800.0 601650.0 ;
      RECT  132000.0 600450.0 133200.0 601650.0 ;
      RECT  132000.0 600450.0 133200.0 601650.0 ;
      RECT  129600.0 600450.0 130800.0 601650.0 ;
      RECT  127200.0 591750.0 128400.0 592950.0 ;
      RECT  129600.0 591750.0 130800.0 592950.0 ;
      RECT  129600.0 591750.0 130800.0 592950.0 ;
      RECT  127200.0 591750.0 128400.0 592950.0 ;
      RECT  129600.0 591750.0 130800.0 592950.0 ;
      RECT  132000.0 591750.0 133200.0 592950.0 ;
      RECT  132000.0 591750.0 133200.0 592950.0 ;
      RECT  129600.0 591750.0 130800.0 592950.0 ;
      RECT  134400.0 601050.0 135600.0 602250.0 ;
      RECT  134400.0 591150.0 135600.0 592350.0 ;
      RECT  132000.0 594300.0 130800.0 595500.0 ;
      RECT  129000.0 597000.0 127800.0 598200.0 ;
      RECT  129600.0 600450.0 130800.0 601650.0 ;
      RECT  132000.0 591750.0 133200.0 592950.0 ;
      RECT  133200.0 597000.0 132000.0 598200.0 ;
      RECT  127800.0 597000.0 129000.0 598200.0 ;
      RECT  130800.0 594300.0 132000.0 595500.0 ;
      RECT  132000.0 597000.0 133200.0 598200.0 ;
      RECT  125400.0 603150.0 139800.0 604050.0 ;
      RECT  125400.0 589350.0 139800.0 590250.0 ;
      RECT  146400.0 601650.0 147600.0 603600.0 ;
      RECT  146400.0 589800.0 147600.0 591750.0 ;
      RECT  141600.0 591150.0 142800.0 589350.0 ;
      RECT  141600.0 600450.0 142800.0 604050.0 ;
      RECT  144300.0 591150.0 145200.0 600450.0 ;
      RECT  141600.0 600450.0 142800.0 601650.0 ;
      RECT  144000.0 600450.0 145200.0 601650.0 ;
      RECT  144000.0 600450.0 145200.0 601650.0 ;
      RECT  141600.0 600450.0 142800.0 601650.0 ;
      RECT  141600.0 591150.0 142800.0 592350.0 ;
      RECT  144000.0 591150.0 145200.0 592350.0 ;
      RECT  144000.0 591150.0 145200.0 592350.0 ;
      RECT  141600.0 591150.0 142800.0 592350.0 ;
      RECT  146400.0 601050.0 147600.0 602250.0 ;
      RECT  146400.0 591150.0 147600.0 592350.0 ;
      RECT  142200.0 595800.0 143400.0 597000.0 ;
      RECT  142200.0 595800.0 143400.0 597000.0 ;
      RECT  144750.0 595950.0 145650.0 596850.0 ;
      RECT  139800.0 603150.0 149400.0 604050.0 ;
      RECT  139800.0 589350.0 149400.0 590250.0 ;
      RECT  112050.0 595800.0 113250.0 597000.0 ;
      RECT  114000.0 593400.0 115200.0 594600.0 ;
      RECT  130800.0 594300.0 129600.0 595500.0 ;
      RECT  122400.0 605550.0 123600.0 603600.0 ;
      RECT  122400.0 617400.0 123600.0 615450.0 ;
      RECT  117600.0 616050.0 118800.0 617850.0 ;
      RECT  117600.0 606750.0 118800.0 603150.0 ;
      RECT  120300.0 616050.0 121200.0 606750.0 ;
      RECT  117600.0 606750.0 118800.0 605550.0 ;
      RECT  120000.0 606750.0 121200.0 605550.0 ;
      RECT  120000.0 606750.0 121200.0 605550.0 ;
      RECT  117600.0 606750.0 118800.0 605550.0 ;
      RECT  117600.0 616050.0 118800.0 614850.0 ;
      RECT  120000.0 616050.0 121200.0 614850.0 ;
      RECT  120000.0 616050.0 121200.0 614850.0 ;
      RECT  117600.0 616050.0 118800.0 614850.0 ;
      RECT  122400.0 606150.0 123600.0 604950.0 ;
      RECT  122400.0 616050.0 123600.0 614850.0 ;
      RECT  118200.0 611400.0 119400.0 610200.0 ;
      RECT  118200.0 611400.0 119400.0 610200.0 ;
      RECT  120750.0 611250.0 121650.0 610350.0 ;
      RECT  115800.0 604050.0 125400.0 603150.0 ;
      RECT  115800.0 617850.0 125400.0 616950.0 ;
      RECT  127200.0 615450.0 128400.0 617850.0 ;
      RECT  127200.0 606750.0 128400.0 603150.0 ;
      RECT  132000.0 606750.0 133200.0 603150.0 ;
      RECT  134400.0 605550.0 135600.0 603600.0 ;
      RECT  134400.0 617400.0 135600.0 615450.0 ;
      RECT  127200.0 606750.0 128400.0 605550.0 ;
      RECT  129600.0 606750.0 130800.0 605550.0 ;
      RECT  129600.0 606750.0 130800.0 605550.0 ;
      RECT  127200.0 606750.0 128400.0 605550.0 ;
      RECT  129600.0 606750.0 130800.0 605550.0 ;
      RECT  132000.0 606750.0 133200.0 605550.0 ;
      RECT  132000.0 606750.0 133200.0 605550.0 ;
      RECT  129600.0 606750.0 130800.0 605550.0 ;
      RECT  127200.0 615450.0 128400.0 614250.0 ;
      RECT  129600.0 615450.0 130800.0 614250.0 ;
      RECT  129600.0 615450.0 130800.0 614250.0 ;
      RECT  127200.0 615450.0 128400.0 614250.0 ;
      RECT  129600.0 615450.0 130800.0 614250.0 ;
      RECT  132000.0 615450.0 133200.0 614250.0 ;
      RECT  132000.0 615450.0 133200.0 614250.0 ;
      RECT  129600.0 615450.0 130800.0 614250.0 ;
      RECT  134400.0 606150.0 135600.0 604950.0 ;
      RECT  134400.0 616050.0 135600.0 614850.0 ;
      RECT  132000.0 612900.0 130800.0 611700.0 ;
      RECT  129000.0 610200.0 127800.0 609000.0 ;
      RECT  129600.0 606750.0 130800.0 605550.0 ;
      RECT  132000.0 615450.0 133200.0 614250.0 ;
      RECT  133200.0 610200.0 132000.0 609000.0 ;
      RECT  127800.0 610200.0 129000.0 609000.0 ;
      RECT  130800.0 612900.0 132000.0 611700.0 ;
      RECT  132000.0 610200.0 133200.0 609000.0 ;
      RECT  125400.0 604050.0 139800.0 603150.0 ;
      RECT  125400.0 617850.0 139800.0 616950.0 ;
      RECT  146400.0 605550.0 147600.0 603600.0 ;
      RECT  146400.0 617400.0 147600.0 615450.0 ;
      RECT  141600.0 616050.0 142800.0 617850.0 ;
      RECT  141600.0 606750.0 142800.0 603150.0 ;
      RECT  144300.0 616050.0 145200.0 606750.0 ;
      RECT  141600.0 606750.0 142800.0 605550.0 ;
      RECT  144000.0 606750.0 145200.0 605550.0 ;
      RECT  144000.0 606750.0 145200.0 605550.0 ;
      RECT  141600.0 606750.0 142800.0 605550.0 ;
      RECT  141600.0 616050.0 142800.0 614850.0 ;
      RECT  144000.0 616050.0 145200.0 614850.0 ;
      RECT  144000.0 616050.0 145200.0 614850.0 ;
      RECT  141600.0 616050.0 142800.0 614850.0 ;
      RECT  146400.0 606150.0 147600.0 604950.0 ;
      RECT  146400.0 616050.0 147600.0 614850.0 ;
      RECT  142200.0 611400.0 143400.0 610200.0 ;
      RECT  142200.0 611400.0 143400.0 610200.0 ;
      RECT  144750.0 611250.0 145650.0 610350.0 ;
      RECT  139800.0 604050.0 149400.0 603150.0 ;
      RECT  139800.0 617850.0 149400.0 616950.0 ;
      RECT  112050.0 610200.0 113250.0 611400.0 ;
      RECT  114000.0 612600.0 115200.0 613800.0 ;
      RECT  130800.0 611700.0 129600.0 612900.0 ;
      RECT  122400.0 629250.0 123600.0 631200.0 ;
      RECT  122400.0 617400.0 123600.0 619350.0 ;
      RECT  117600.0 618750.0 118800.0 616950.0 ;
      RECT  117600.0 628050.0 118800.0 631650.0 ;
      RECT  120300.0 618750.0 121200.0 628050.0 ;
      RECT  117600.0 628050.0 118800.0 629250.0 ;
      RECT  120000.0 628050.0 121200.0 629250.0 ;
      RECT  120000.0 628050.0 121200.0 629250.0 ;
      RECT  117600.0 628050.0 118800.0 629250.0 ;
      RECT  117600.0 618750.0 118800.0 619950.0 ;
      RECT  120000.0 618750.0 121200.0 619950.0 ;
      RECT  120000.0 618750.0 121200.0 619950.0 ;
      RECT  117600.0 618750.0 118800.0 619950.0 ;
      RECT  122400.0 628650.0 123600.0 629850.0 ;
      RECT  122400.0 618750.0 123600.0 619950.0 ;
      RECT  118200.0 623400.0 119400.0 624600.0 ;
      RECT  118200.0 623400.0 119400.0 624600.0 ;
      RECT  120750.0 623550.0 121650.0 624450.0 ;
      RECT  115800.0 630750.0 125400.0 631650.0 ;
      RECT  115800.0 616950.0 125400.0 617850.0 ;
      RECT  127200.0 619350.0 128400.0 616950.0 ;
      RECT  127200.0 628050.0 128400.0 631650.0 ;
      RECT  132000.0 628050.0 133200.0 631650.0 ;
      RECT  134400.0 629250.0 135600.0 631200.0 ;
      RECT  134400.0 617400.0 135600.0 619350.0 ;
      RECT  127200.0 628050.0 128400.0 629250.0 ;
      RECT  129600.0 628050.0 130800.0 629250.0 ;
      RECT  129600.0 628050.0 130800.0 629250.0 ;
      RECT  127200.0 628050.0 128400.0 629250.0 ;
      RECT  129600.0 628050.0 130800.0 629250.0 ;
      RECT  132000.0 628050.0 133200.0 629250.0 ;
      RECT  132000.0 628050.0 133200.0 629250.0 ;
      RECT  129600.0 628050.0 130800.0 629250.0 ;
      RECT  127200.0 619350.0 128400.0 620550.0 ;
      RECT  129600.0 619350.0 130800.0 620550.0 ;
      RECT  129600.0 619350.0 130800.0 620550.0 ;
      RECT  127200.0 619350.0 128400.0 620550.0 ;
      RECT  129600.0 619350.0 130800.0 620550.0 ;
      RECT  132000.0 619350.0 133200.0 620550.0 ;
      RECT  132000.0 619350.0 133200.0 620550.0 ;
      RECT  129600.0 619350.0 130800.0 620550.0 ;
      RECT  134400.0 628650.0 135600.0 629850.0 ;
      RECT  134400.0 618750.0 135600.0 619950.0 ;
      RECT  132000.0 621900.0 130800.0 623100.0 ;
      RECT  129000.0 624600.0 127800.0 625800.0 ;
      RECT  129600.0 628050.0 130800.0 629250.0 ;
      RECT  132000.0 619350.0 133200.0 620550.0 ;
      RECT  133200.0 624600.0 132000.0 625800.0 ;
      RECT  127800.0 624600.0 129000.0 625800.0 ;
      RECT  130800.0 621900.0 132000.0 623100.0 ;
      RECT  132000.0 624600.0 133200.0 625800.0 ;
      RECT  125400.0 630750.0 139800.0 631650.0 ;
      RECT  125400.0 616950.0 139800.0 617850.0 ;
      RECT  146400.0 629250.0 147600.0 631200.0 ;
      RECT  146400.0 617400.0 147600.0 619350.0 ;
      RECT  141600.0 618750.0 142800.0 616950.0 ;
      RECT  141600.0 628050.0 142800.0 631650.0 ;
      RECT  144300.0 618750.0 145200.0 628050.0 ;
      RECT  141600.0 628050.0 142800.0 629250.0 ;
      RECT  144000.0 628050.0 145200.0 629250.0 ;
      RECT  144000.0 628050.0 145200.0 629250.0 ;
      RECT  141600.0 628050.0 142800.0 629250.0 ;
      RECT  141600.0 618750.0 142800.0 619950.0 ;
      RECT  144000.0 618750.0 145200.0 619950.0 ;
      RECT  144000.0 618750.0 145200.0 619950.0 ;
      RECT  141600.0 618750.0 142800.0 619950.0 ;
      RECT  146400.0 628650.0 147600.0 629850.0 ;
      RECT  146400.0 618750.0 147600.0 619950.0 ;
      RECT  142200.0 623400.0 143400.0 624600.0 ;
      RECT  142200.0 623400.0 143400.0 624600.0 ;
      RECT  144750.0 623550.0 145650.0 624450.0 ;
      RECT  139800.0 630750.0 149400.0 631650.0 ;
      RECT  139800.0 616950.0 149400.0 617850.0 ;
      RECT  112050.0 623400.0 113250.0 624600.0 ;
      RECT  114000.0 621000.0 115200.0 622200.0 ;
      RECT  130800.0 621900.0 129600.0 623100.0 ;
      RECT  122400.0 633150.0 123600.0 631200.0 ;
      RECT  122400.0 645000.0 123600.0 643050.0 ;
      RECT  117600.0 643650.0 118800.0 645450.0 ;
      RECT  117600.0 634350.0 118800.0 630750.0 ;
      RECT  120300.0 643650.0 121200.0 634350.0 ;
      RECT  117600.0 634350.0 118800.0 633150.0 ;
      RECT  120000.0 634350.0 121200.0 633150.0 ;
      RECT  120000.0 634350.0 121200.0 633150.0 ;
      RECT  117600.0 634350.0 118800.0 633150.0 ;
      RECT  117600.0 643650.0 118800.0 642450.0 ;
      RECT  120000.0 643650.0 121200.0 642450.0 ;
      RECT  120000.0 643650.0 121200.0 642450.0 ;
      RECT  117600.0 643650.0 118800.0 642450.0 ;
      RECT  122400.0 633750.0 123600.0 632550.0 ;
      RECT  122400.0 643650.0 123600.0 642450.0 ;
      RECT  118200.0 639000.0 119400.0 637800.0 ;
      RECT  118200.0 639000.0 119400.0 637800.0 ;
      RECT  120750.0 638850.0 121650.0 637950.0 ;
      RECT  115800.0 631650.0 125400.0 630750.0 ;
      RECT  115800.0 645450.0 125400.0 644550.0 ;
      RECT  127200.0 643050.0 128400.0 645450.0 ;
      RECT  127200.0 634350.0 128400.0 630750.0 ;
      RECT  132000.0 634350.0 133200.0 630750.0 ;
      RECT  134400.0 633150.0 135600.0 631200.0 ;
      RECT  134400.0 645000.0 135600.0 643050.0 ;
      RECT  127200.0 634350.0 128400.0 633150.0 ;
      RECT  129600.0 634350.0 130800.0 633150.0 ;
      RECT  129600.0 634350.0 130800.0 633150.0 ;
      RECT  127200.0 634350.0 128400.0 633150.0 ;
      RECT  129600.0 634350.0 130800.0 633150.0 ;
      RECT  132000.0 634350.0 133200.0 633150.0 ;
      RECT  132000.0 634350.0 133200.0 633150.0 ;
      RECT  129600.0 634350.0 130800.0 633150.0 ;
      RECT  127200.0 643050.0 128400.0 641850.0 ;
      RECT  129600.0 643050.0 130800.0 641850.0 ;
      RECT  129600.0 643050.0 130800.0 641850.0 ;
      RECT  127200.0 643050.0 128400.0 641850.0 ;
      RECT  129600.0 643050.0 130800.0 641850.0 ;
      RECT  132000.0 643050.0 133200.0 641850.0 ;
      RECT  132000.0 643050.0 133200.0 641850.0 ;
      RECT  129600.0 643050.0 130800.0 641850.0 ;
      RECT  134400.0 633750.0 135600.0 632550.0 ;
      RECT  134400.0 643650.0 135600.0 642450.0 ;
      RECT  132000.0 640500.0 130800.0 639300.0 ;
      RECT  129000.0 637800.0 127800.0 636600.0 ;
      RECT  129600.0 634350.0 130800.0 633150.0 ;
      RECT  132000.0 643050.0 133200.0 641850.0 ;
      RECT  133200.0 637800.0 132000.0 636600.0 ;
      RECT  127800.0 637800.0 129000.0 636600.0 ;
      RECT  130800.0 640500.0 132000.0 639300.0 ;
      RECT  132000.0 637800.0 133200.0 636600.0 ;
      RECT  125400.0 631650.0 139800.0 630750.0 ;
      RECT  125400.0 645450.0 139800.0 644550.0 ;
      RECT  146400.0 633150.0 147600.0 631200.0 ;
      RECT  146400.0 645000.0 147600.0 643050.0 ;
      RECT  141600.0 643650.0 142800.0 645450.0 ;
      RECT  141600.0 634350.0 142800.0 630750.0 ;
      RECT  144300.0 643650.0 145200.0 634350.0 ;
      RECT  141600.0 634350.0 142800.0 633150.0 ;
      RECT  144000.0 634350.0 145200.0 633150.0 ;
      RECT  144000.0 634350.0 145200.0 633150.0 ;
      RECT  141600.0 634350.0 142800.0 633150.0 ;
      RECT  141600.0 643650.0 142800.0 642450.0 ;
      RECT  144000.0 643650.0 145200.0 642450.0 ;
      RECT  144000.0 643650.0 145200.0 642450.0 ;
      RECT  141600.0 643650.0 142800.0 642450.0 ;
      RECT  146400.0 633750.0 147600.0 632550.0 ;
      RECT  146400.0 643650.0 147600.0 642450.0 ;
      RECT  142200.0 639000.0 143400.0 637800.0 ;
      RECT  142200.0 639000.0 143400.0 637800.0 ;
      RECT  144750.0 638850.0 145650.0 637950.0 ;
      RECT  139800.0 631650.0 149400.0 630750.0 ;
      RECT  139800.0 645450.0 149400.0 644550.0 ;
      RECT  112050.0 637800.0 113250.0 639000.0 ;
      RECT  114000.0 640200.0 115200.0 641400.0 ;
      RECT  130800.0 639300.0 129600.0 640500.0 ;
      RECT  122400.0 656850.0 123600.0 658800.0 ;
      RECT  122400.0 645000.0 123600.0 646950.0 ;
      RECT  117600.0 646350.0 118800.0 644550.0 ;
      RECT  117600.0 655650.0 118800.0 659250.0 ;
      RECT  120300.0 646350.0 121200.0 655650.0 ;
      RECT  117600.0 655650.0 118800.0 656850.0 ;
      RECT  120000.0 655650.0 121200.0 656850.0 ;
      RECT  120000.0 655650.0 121200.0 656850.0 ;
      RECT  117600.0 655650.0 118800.0 656850.0 ;
      RECT  117600.0 646350.0 118800.0 647550.0 ;
      RECT  120000.0 646350.0 121200.0 647550.0 ;
      RECT  120000.0 646350.0 121200.0 647550.0 ;
      RECT  117600.0 646350.0 118800.0 647550.0 ;
      RECT  122400.0 656250.0 123600.0 657450.0 ;
      RECT  122400.0 646350.0 123600.0 647550.0 ;
      RECT  118200.0 651000.0 119400.0 652200.0 ;
      RECT  118200.0 651000.0 119400.0 652200.0 ;
      RECT  120750.0 651150.0 121650.0 652050.0 ;
      RECT  115800.0 658350.0 125400.0 659250.0 ;
      RECT  115800.0 644550.0 125400.0 645450.0 ;
      RECT  127200.0 646950.0 128400.0 644550.0 ;
      RECT  127200.0 655650.0 128400.0 659250.0 ;
      RECT  132000.0 655650.0 133200.0 659250.0 ;
      RECT  134400.0 656850.0 135600.0 658800.0 ;
      RECT  134400.0 645000.0 135600.0 646950.0 ;
      RECT  127200.0 655650.0 128400.0 656850.0 ;
      RECT  129600.0 655650.0 130800.0 656850.0 ;
      RECT  129600.0 655650.0 130800.0 656850.0 ;
      RECT  127200.0 655650.0 128400.0 656850.0 ;
      RECT  129600.0 655650.0 130800.0 656850.0 ;
      RECT  132000.0 655650.0 133200.0 656850.0 ;
      RECT  132000.0 655650.0 133200.0 656850.0 ;
      RECT  129600.0 655650.0 130800.0 656850.0 ;
      RECT  127200.0 646950.0 128400.0 648150.0 ;
      RECT  129600.0 646950.0 130800.0 648150.0 ;
      RECT  129600.0 646950.0 130800.0 648150.0 ;
      RECT  127200.0 646950.0 128400.0 648150.0 ;
      RECT  129600.0 646950.0 130800.0 648150.0 ;
      RECT  132000.0 646950.0 133200.0 648150.0 ;
      RECT  132000.0 646950.0 133200.0 648150.0 ;
      RECT  129600.0 646950.0 130800.0 648150.0 ;
      RECT  134400.0 656250.0 135600.0 657450.0 ;
      RECT  134400.0 646350.0 135600.0 647550.0 ;
      RECT  132000.0 649500.0 130800.0 650700.0 ;
      RECT  129000.0 652200.0 127800.0 653400.0 ;
      RECT  129600.0 655650.0 130800.0 656850.0 ;
      RECT  132000.0 646950.0 133200.0 648150.0 ;
      RECT  133200.0 652200.0 132000.0 653400.0 ;
      RECT  127800.0 652200.0 129000.0 653400.0 ;
      RECT  130800.0 649500.0 132000.0 650700.0 ;
      RECT  132000.0 652200.0 133200.0 653400.0 ;
      RECT  125400.0 658350.0 139800.0 659250.0 ;
      RECT  125400.0 644550.0 139800.0 645450.0 ;
      RECT  146400.0 656850.0 147600.0 658800.0 ;
      RECT  146400.0 645000.0 147600.0 646950.0 ;
      RECT  141600.0 646350.0 142800.0 644550.0 ;
      RECT  141600.0 655650.0 142800.0 659250.0 ;
      RECT  144300.0 646350.0 145200.0 655650.0 ;
      RECT  141600.0 655650.0 142800.0 656850.0 ;
      RECT  144000.0 655650.0 145200.0 656850.0 ;
      RECT  144000.0 655650.0 145200.0 656850.0 ;
      RECT  141600.0 655650.0 142800.0 656850.0 ;
      RECT  141600.0 646350.0 142800.0 647550.0 ;
      RECT  144000.0 646350.0 145200.0 647550.0 ;
      RECT  144000.0 646350.0 145200.0 647550.0 ;
      RECT  141600.0 646350.0 142800.0 647550.0 ;
      RECT  146400.0 656250.0 147600.0 657450.0 ;
      RECT  146400.0 646350.0 147600.0 647550.0 ;
      RECT  142200.0 651000.0 143400.0 652200.0 ;
      RECT  142200.0 651000.0 143400.0 652200.0 ;
      RECT  144750.0 651150.0 145650.0 652050.0 ;
      RECT  139800.0 658350.0 149400.0 659250.0 ;
      RECT  139800.0 644550.0 149400.0 645450.0 ;
      RECT  112050.0 651000.0 113250.0 652200.0 ;
      RECT  114000.0 648600.0 115200.0 649800.0 ;
      RECT  130800.0 649500.0 129600.0 650700.0 ;
      RECT  122400.0 660750.0 123600.0 658800.0 ;
      RECT  122400.0 672600.0 123600.0 670650.0 ;
      RECT  117600.0 671250.0 118800.0 673050.0 ;
      RECT  117600.0 661950.0 118800.0 658350.0 ;
      RECT  120300.0 671250.0 121200.0 661950.0 ;
      RECT  117600.0 661950.0 118800.0 660750.0 ;
      RECT  120000.0 661950.0 121200.0 660750.0 ;
      RECT  120000.0 661950.0 121200.0 660750.0 ;
      RECT  117600.0 661950.0 118800.0 660750.0 ;
      RECT  117600.0 671250.0 118800.0 670050.0 ;
      RECT  120000.0 671250.0 121200.0 670050.0 ;
      RECT  120000.0 671250.0 121200.0 670050.0 ;
      RECT  117600.0 671250.0 118800.0 670050.0 ;
      RECT  122400.0 661350.0 123600.0 660150.0 ;
      RECT  122400.0 671250.0 123600.0 670050.0 ;
      RECT  118200.0 666600.0 119400.0 665400.0 ;
      RECT  118200.0 666600.0 119400.0 665400.0 ;
      RECT  120750.0 666450.0 121650.0 665550.0 ;
      RECT  115800.0 659250.0 125400.0 658350.0 ;
      RECT  115800.0 673050.0 125400.0 672150.0 ;
      RECT  127200.0 670650.0 128400.0 673050.0 ;
      RECT  127200.0 661950.0 128400.0 658350.0 ;
      RECT  132000.0 661950.0 133200.0 658350.0 ;
      RECT  134400.0 660750.0 135600.0 658800.0 ;
      RECT  134400.0 672600.0 135600.0 670650.0 ;
      RECT  127200.0 661950.0 128400.0 660750.0 ;
      RECT  129600.0 661950.0 130800.0 660750.0 ;
      RECT  129600.0 661950.0 130800.0 660750.0 ;
      RECT  127200.0 661950.0 128400.0 660750.0 ;
      RECT  129600.0 661950.0 130800.0 660750.0 ;
      RECT  132000.0 661950.0 133200.0 660750.0 ;
      RECT  132000.0 661950.0 133200.0 660750.0 ;
      RECT  129600.0 661950.0 130800.0 660750.0 ;
      RECT  127200.0 670650.0 128400.0 669450.0 ;
      RECT  129600.0 670650.0 130800.0 669450.0 ;
      RECT  129600.0 670650.0 130800.0 669450.0 ;
      RECT  127200.0 670650.0 128400.0 669450.0 ;
      RECT  129600.0 670650.0 130800.0 669450.0 ;
      RECT  132000.0 670650.0 133200.0 669450.0 ;
      RECT  132000.0 670650.0 133200.0 669450.0 ;
      RECT  129600.0 670650.0 130800.0 669450.0 ;
      RECT  134400.0 661350.0 135600.0 660150.0 ;
      RECT  134400.0 671250.0 135600.0 670050.0 ;
      RECT  132000.0 668100.0 130800.0 666900.0 ;
      RECT  129000.0 665400.0 127800.0 664200.0 ;
      RECT  129600.0 661950.0 130800.0 660750.0 ;
      RECT  132000.0 670650.0 133200.0 669450.0 ;
      RECT  133200.0 665400.0 132000.0 664200.0 ;
      RECT  127800.0 665400.0 129000.0 664200.0 ;
      RECT  130800.0 668100.0 132000.0 666900.0 ;
      RECT  132000.0 665400.0 133200.0 664200.0 ;
      RECT  125400.0 659250.0 139800.0 658350.0 ;
      RECT  125400.0 673050.0 139800.0 672150.0 ;
      RECT  146400.0 660750.0 147600.0 658800.0 ;
      RECT  146400.0 672600.0 147600.0 670650.0 ;
      RECT  141600.0 671250.0 142800.0 673050.0 ;
      RECT  141600.0 661950.0 142800.0 658350.0 ;
      RECT  144300.0 671250.0 145200.0 661950.0 ;
      RECT  141600.0 661950.0 142800.0 660750.0 ;
      RECT  144000.0 661950.0 145200.0 660750.0 ;
      RECT  144000.0 661950.0 145200.0 660750.0 ;
      RECT  141600.0 661950.0 142800.0 660750.0 ;
      RECT  141600.0 671250.0 142800.0 670050.0 ;
      RECT  144000.0 671250.0 145200.0 670050.0 ;
      RECT  144000.0 671250.0 145200.0 670050.0 ;
      RECT  141600.0 671250.0 142800.0 670050.0 ;
      RECT  146400.0 661350.0 147600.0 660150.0 ;
      RECT  146400.0 671250.0 147600.0 670050.0 ;
      RECT  142200.0 666600.0 143400.0 665400.0 ;
      RECT  142200.0 666600.0 143400.0 665400.0 ;
      RECT  144750.0 666450.0 145650.0 665550.0 ;
      RECT  139800.0 659250.0 149400.0 658350.0 ;
      RECT  139800.0 673050.0 149400.0 672150.0 ;
      RECT  112050.0 665400.0 113250.0 666600.0 ;
      RECT  114000.0 667800.0 115200.0 669000.0 ;
      RECT  130800.0 666900.0 129600.0 668100.0 ;
      RECT  122400.0 684450.0 123600.0 686400.0 ;
      RECT  122400.0 672600.0 123600.0 674550.0 ;
      RECT  117600.0 673950.0 118800.0 672150.0 ;
      RECT  117600.0 683250.0 118800.0 686850.0 ;
      RECT  120300.0 673950.0 121200.0 683250.0 ;
      RECT  117600.0 683250.0 118800.0 684450.0 ;
      RECT  120000.0 683250.0 121200.0 684450.0 ;
      RECT  120000.0 683250.0 121200.0 684450.0 ;
      RECT  117600.0 683250.0 118800.0 684450.0 ;
      RECT  117600.0 673950.0 118800.0 675150.0 ;
      RECT  120000.0 673950.0 121200.0 675150.0 ;
      RECT  120000.0 673950.0 121200.0 675150.0 ;
      RECT  117600.0 673950.0 118800.0 675150.0 ;
      RECT  122400.0 683850.0 123600.0 685050.0 ;
      RECT  122400.0 673950.0 123600.0 675150.0 ;
      RECT  118200.0 678600.0 119400.0 679800.0 ;
      RECT  118200.0 678600.0 119400.0 679800.0 ;
      RECT  120750.0 678750.0 121650.0 679650.0 ;
      RECT  115800.0 685950.0 125400.0 686850.0 ;
      RECT  115800.0 672150.0 125400.0 673050.0 ;
      RECT  127200.0 674550.0 128400.0 672150.0 ;
      RECT  127200.0 683250.0 128400.0 686850.0 ;
      RECT  132000.0 683250.0 133200.0 686850.0 ;
      RECT  134400.0 684450.0 135600.0 686400.0 ;
      RECT  134400.0 672600.0 135600.0 674550.0 ;
      RECT  127200.0 683250.0 128400.0 684450.0 ;
      RECT  129600.0 683250.0 130800.0 684450.0 ;
      RECT  129600.0 683250.0 130800.0 684450.0 ;
      RECT  127200.0 683250.0 128400.0 684450.0 ;
      RECT  129600.0 683250.0 130800.0 684450.0 ;
      RECT  132000.0 683250.0 133200.0 684450.0 ;
      RECT  132000.0 683250.0 133200.0 684450.0 ;
      RECT  129600.0 683250.0 130800.0 684450.0 ;
      RECT  127200.0 674550.0 128400.0 675750.0 ;
      RECT  129600.0 674550.0 130800.0 675750.0 ;
      RECT  129600.0 674550.0 130800.0 675750.0 ;
      RECT  127200.0 674550.0 128400.0 675750.0 ;
      RECT  129600.0 674550.0 130800.0 675750.0 ;
      RECT  132000.0 674550.0 133200.0 675750.0 ;
      RECT  132000.0 674550.0 133200.0 675750.0 ;
      RECT  129600.0 674550.0 130800.0 675750.0 ;
      RECT  134400.0 683850.0 135600.0 685050.0 ;
      RECT  134400.0 673950.0 135600.0 675150.0 ;
      RECT  132000.0 677100.0 130800.0 678300.0 ;
      RECT  129000.0 679800.0 127800.0 681000.0 ;
      RECT  129600.0 683250.0 130800.0 684450.0 ;
      RECT  132000.0 674550.0 133200.0 675750.0 ;
      RECT  133200.0 679800.0 132000.0 681000.0 ;
      RECT  127800.0 679800.0 129000.0 681000.0 ;
      RECT  130800.0 677100.0 132000.0 678300.0 ;
      RECT  132000.0 679800.0 133200.0 681000.0 ;
      RECT  125400.0 685950.0 139800.0 686850.0 ;
      RECT  125400.0 672150.0 139800.0 673050.0 ;
      RECT  146400.0 684450.0 147600.0 686400.0 ;
      RECT  146400.0 672600.0 147600.0 674550.0 ;
      RECT  141600.0 673950.0 142800.0 672150.0 ;
      RECT  141600.0 683250.0 142800.0 686850.0 ;
      RECT  144300.0 673950.0 145200.0 683250.0 ;
      RECT  141600.0 683250.0 142800.0 684450.0 ;
      RECT  144000.0 683250.0 145200.0 684450.0 ;
      RECT  144000.0 683250.0 145200.0 684450.0 ;
      RECT  141600.0 683250.0 142800.0 684450.0 ;
      RECT  141600.0 673950.0 142800.0 675150.0 ;
      RECT  144000.0 673950.0 145200.0 675150.0 ;
      RECT  144000.0 673950.0 145200.0 675150.0 ;
      RECT  141600.0 673950.0 142800.0 675150.0 ;
      RECT  146400.0 683850.0 147600.0 685050.0 ;
      RECT  146400.0 673950.0 147600.0 675150.0 ;
      RECT  142200.0 678600.0 143400.0 679800.0 ;
      RECT  142200.0 678600.0 143400.0 679800.0 ;
      RECT  144750.0 678750.0 145650.0 679650.0 ;
      RECT  139800.0 685950.0 149400.0 686850.0 ;
      RECT  139800.0 672150.0 149400.0 673050.0 ;
      RECT  112050.0 678600.0 113250.0 679800.0 ;
      RECT  114000.0 676200.0 115200.0 677400.0 ;
      RECT  130800.0 677100.0 129600.0 678300.0 ;
      RECT  122400.0 688350.0 123600.0 686400.0 ;
      RECT  122400.0 700200.0 123600.0 698250.0 ;
      RECT  117600.0 698850.0 118800.0 700650.0 ;
      RECT  117600.0 689550.0 118800.0 685950.0 ;
      RECT  120300.0 698850.0 121200.0 689550.0 ;
      RECT  117600.0 689550.0 118800.0 688350.0 ;
      RECT  120000.0 689550.0 121200.0 688350.0 ;
      RECT  120000.0 689550.0 121200.0 688350.0 ;
      RECT  117600.0 689550.0 118800.0 688350.0 ;
      RECT  117600.0 698850.0 118800.0 697650.0 ;
      RECT  120000.0 698850.0 121200.0 697650.0 ;
      RECT  120000.0 698850.0 121200.0 697650.0 ;
      RECT  117600.0 698850.0 118800.0 697650.0 ;
      RECT  122400.0 688950.0 123600.0 687750.0 ;
      RECT  122400.0 698850.0 123600.0 697650.0 ;
      RECT  118200.0 694200.0 119400.0 693000.0 ;
      RECT  118200.0 694200.0 119400.0 693000.0 ;
      RECT  120750.0 694050.0 121650.0 693150.0 ;
      RECT  115800.0 686850.0 125400.0 685950.0 ;
      RECT  115800.0 700650.0 125400.0 699750.0 ;
      RECT  127200.0 698250.0 128400.0 700650.0 ;
      RECT  127200.0 689550.0 128400.0 685950.0 ;
      RECT  132000.0 689550.0 133200.0 685950.0 ;
      RECT  134400.0 688350.0 135600.0 686400.0 ;
      RECT  134400.0 700200.0 135600.0 698250.0 ;
      RECT  127200.0 689550.0 128400.0 688350.0 ;
      RECT  129600.0 689550.0 130800.0 688350.0 ;
      RECT  129600.0 689550.0 130800.0 688350.0 ;
      RECT  127200.0 689550.0 128400.0 688350.0 ;
      RECT  129600.0 689550.0 130800.0 688350.0 ;
      RECT  132000.0 689550.0 133200.0 688350.0 ;
      RECT  132000.0 689550.0 133200.0 688350.0 ;
      RECT  129600.0 689550.0 130800.0 688350.0 ;
      RECT  127200.0 698250.0 128400.0 697050.0 ;
      RECT  129600.0 698250.0 130800.0 697050.0 ;
      RECT  129600.0 698250.0 130800.0 697050.0 ;
      RECT  127200.0 698250.0 128400.0 697050.0 ;
      RECT  129600.0 698250.0 130800.0 697050.0 ;
      RECT  132000.0 698250.0 133200.0 697050.0 ;
      RECT  132000.0 698250.0 133200.0 697050.0 ;
      RECT  129600.0 698250.0 130800.0 697050.0 ;
      RECT  134400.0 688950.0 135600.0 687750.0 ;
      RECT  134400.0 698850.0 135600.0 697650.0 ;
      RECT  132000.0 695700.0 130800.0 694500.0 ;
      RECT  129000.0 693000.0 127800.0 691800.0 ;
      RECT  129600.0 689550.0 130800.0 688350.0 ;
      RECT  132000.0 698250.0 133200.0 697050.0 ;
      RECT  133200.0 693000.0 132000.0 691800.0 ;
      RECT  127800.0 693000.0 129000.0 691800.0 ;
      RECT  130800.0 695700.0 132000.0 694500.0 ;
      RECT  132000.0 693000.0 133200.0 691800.0 ;
      RECT  125400.0 686850.0 139800.0 685950.0 ;
      RECT  125400.0 700650.0 139800.0 699750.0 ;
      RECT  146400.0 688350.0 147600.0 686400.0 ;
      RECT  146400.0 700200.0 147600.0 698250.0 ;
      RECT  141600.0 698850.0 142800.0 700650.0 ;
      RECT  141600.0 689550.0 142800.0 685950.0 ;
      RECT  144300.0 698850.0 145200.0 689550.0 ;
      RECT  141600.0 689550.0 142800.0 688350.0 ;
      RECT  144000.0 689550.0 145200.0 688350.0 ;
      RECT  144000.0 689550.0 145200.0 688350.0 ;
      RECT  141600.0 689550.0 142800.0 688350.0 ;
      RECT  141600.0 698850.0 142800.0 697650.0 ;
      RECT  144000.0 698850.0 145200.0 697650.0 ;
      RECT  144000.0 698850.0 145200.0 697650.0 ;
      RECT  141600.0 698850.0 142800.0 697650.0 ;
      RECT  146400.0 688950.0 147600.0 687750.0 ;
      RECT  146400.0 698850.0 147600.0 697650.0 ;
      RECT  142200.0 694200.0 143400.0 693000.0 ;
      RECT  142200.0 694200.0 143400.0 693000.0 ;
      RECT  144750.0 694050.0 145650.0 693150.0 ;
      RECT  139800.0 686850.0 149400.0 685950.0 ;
      RECT  139800.0 700650.0 149400.0 699750.0 ;
      RECT  112050.0 693000.0 113250.0 694200.0 ;
      RECT  114000.0 695400.0 115200.0 696600.0 ;
      RECT  130800.0 694500.0 129600.0 695700.0 ;
      RECT  122400.0 712050.0 123600.0 714000.0 ;
      RECT  122400.0 700200.0 123600.0 702150.0 ;
      RECT  117600.0 701550.0 118800.0 699750.0 ;
      RECT  117600.0 710850.0 118800.0 714450.0 ;
      RECT  120300.0 701550.0 121200.0 710850.0 ;
      RECT  117600.0 710850.0 118800.0 712050.0 ;
      RECT  120000.0 710850.0 121200.0 712050.0 ;
      RECT  120000.0 710850.0 121200.0 712050.0 ;
      RECT  117600.0 710850.0 118800.0 712050.0 ;
      RECT  117600.0 701550.0 118800.0 702750.0 ;
      RECT  120000.0 701550.0 121200.0 702750.0 ;
      RECT  120000.0 701550.0 121200.0 702750.0 ;
      RECT  117600.0 701550.0 118800.0 702750.0 ;
      RECT  122400.0 711450.0 123600.0 712650.0 ;
      RECT  122400.0 701550.0 123600.0 702750.0 ;
      RECT  118200.0 706200.0 119400.0 707400.0 ;
      RECT  118200.0 706200.0 119400.0 707400.0 ;
      RECT  120750.0 706350.0 121650.0 707250.0 ;
      RECT  115800.0 713550.0 125400.0 714450.0 ;
      RECT  115800.0 699750.0 125400.0 700650.0 ;
      RECT  127200.0 702150.0 128400.0 699750.0 ;
      RECT  127200.0 710850.0 128400.0 714450.0 ;
      RECT  132000.0 710850.0 133200.0 714450.0 ;
      RECT  134400.0 712050.0 135600.0 714000.0 ;
      RECT  134400.0 700200.0 135600.0 702150.0 ;
      RECT  127200.0 710850.0 128400.0 712050.0 ;
      RECT  129600.0 710850.0 130800.0 712050.0 ;
      RECT  129600.0 710850.0 130800.0 712050.0 ;
      RECT  127200.0 710850.0 128400.0 712050.0 ;
      RECT  129600.0 710850.0 130800.0 712050.0 ;
      RECT  132000.0 710850.0 133200.0 712050.0 ;
      RECT  132000.0 710850.0 133200.0 712050.0 ;
      RECT  129600.0 710850.0 130800.0 712050.0 ;
      RECT  127200.0 702150.0 128400.0 703350.0 ;
      RECT  129600.0 702150.0 130800.0 703350.0 ;
      RECT  129600.0 702150.0 130800.0 703350.0 ;
      RECT  127200.0 702150.0 128400.0 703350.0 ;
      RECT  129600.0 702150.0 130800.0 703350.0 ;
      RECT  132000.0 702150.0 133200.0 703350.0 ;
      RECT  132000.0 702150.0 133200.0 703350.0 ;
      RECT  129600.0 702150.0 130800.0 703350.0 ;
      RECT  134400.0 711450.0 135600.0 712650.0 ;
      RECT  134400.0 701550.0 135600.0 702750.0 ;
      RECT  132000.0 704700.0 130800.0 705900.0 ;
      RECT  129000.0 707400.0 127800.0 708600.0 ;
      RECT  129600.0 710850.0 130800.0 712050.0 ;
      RECT  132000.0 702150.0 133200.0 703350.0 ;
      RECT  133200.0 707400.0 132000.0 708600.0 ;
      RECT  127800.0 707400.0 129000.0 708600.0 ;
      RECT  130800.0 704700.0 132000.0 705900.0 ;
      RECT  132000.0 707400.0 133200.0 708600.0 ;
      RECT  125400.0 713550.0 139800.0 714450.0 ;
      RECT  125400.0 699750.0 139800.0 700650.0 ;
      RECT  146400.0 712050.0 147600.0 714000.0 ;
      RECT  146400.0 700200.0 147600.0 702150.0 ;
      RECT  141600.0 701550.0 142800.0 699750.0 ;
      RECT  141600.0 710850.0 142800.0 714450.0 ;
      RECT  144300.0 701550.0 145200.0 710850.0 ;
      RECT  141600.0 710850.0 142800.0 712050.0 ;
      RECT  144000.0 710850.0 145200.0 712050.0 ;
      RECT  144000.0 710850.0 145200.0 712050.0 ;
      RECT  141600.0 710850.0 142800.0 712050.0 ;
      RECT  141600.0 701550.0 142800.0 702750.0 ;
      RECT  144000.0 701550.0 145200.0 702750.0 ;
      RECT  144000.0 701550.0 145200.0 702750.0 ;
      RECT  141600.0 701550.0 142800.0 702750.0 ;
      RECT  146400.0 711450.0 147600.0 712650.0 ;
      RECT  146400.0 701550.0 147600.0 702750.0 ;
      RECT  142200.0 706200.0 143400.0 707400.0 ;
      RECT  142200.0 706200.0 143400.0 707400.0 ;
      RECT  144750.0 706350.0 145650.0 707250.0 ;
      RECT  139800.0 713550.0 149400.0 714450.0 ;
      RECT  139800.0 699750.0 149400.0 700650.0 ;
      RECT  112050.0 706200.0 113250.0 707400.0 ;
      RECT  114000.0 703800.0 115200.0 705000.0 ;
      RECT  130800.0 704700.0 129600.0 705900.0 ;
      RECT  122400.0 715950.0 123600.0 714000.0 ;
      RECT  122400.0 727800.0 123600.0 725850.0 ;
      RECT  117600.0 726450.0 118800.0 728250.0 ;
      RECT  117600.0 717150.0 118800.0 713550.0 ;
      RECT  120300.0 726450.0 121200.0 717150.0 ;
      RECT  117600.0 717150.0 118800.0 715950.0 ;
      RECT  120000.0 717150.0 121200.0 715950.0 ;
      RECT  120000.0 717150.0 121200.0 715950.0 ;
      RECT  117600.0 717150.0 118800.0 715950.0 ;
      RECT  117600.0 726450.0 118800.0 725250.0 ;
      RECT  120000.0 726450.0 121200.0 725250.0 ;
      RECT  120000.0 726450.0 121200.0 725250.0 ;
      RECT  117600.0 726450.0 118800.0 725250.0 ;
      RECT  122400.0 716550.0 123600.0 715350.0 ;
      RECT  122400.0 726450.0 123600.0 725250.0 ;
      RECT  118200.0 721800.0 119400.0 720600.0 ;
      RECT  118200.0 721800.0 119400.0 720600.0 ;
      RECT  120750.0 721650.0 121650.0 720750.0 ;
      RECT  115800.0 714450.0 125400.0 713550.0 ;
      RECT  115800.0 728250.0 125400.0 727350.0 ;
      RECT  127200.0 725850.0 128400.0 728250.0 ;
      RECT  127200.0 717150.0 128400.0 713550.0 ;
      RECT  132000.0 717150.0 133200.0 713550.0 ;
      RECT  134400.0 715950.0 135600.0 714000.0 ;
      RECT  134400.0 727800.0 135600.0 725850.0 ;
      RECT  127200.0 717150.0 128400.0 715950.0 ;
      RECT  129600.0 717150.0 130800.0 715950.0 ;
      RECT  129600.0 717150.0 130800.0 715950.0 ;
      RECT  127200.0 717150.0 128400.0 715950.0 ;
      RECT  129600.0 717150.0 130800.0 715950.0 ;
      RECT  132000.0 717150.0 133200.0 715950.0 ;
      RECT  132000.0 717150.0 133200.0 715950.0 ;
      RECT  129600.0 717150.0 130800.0 715950.0 ;
      RECT  127200.0 725850.0 128400.0 724650.0 ;
      RECT  129600.0 725850.0 130800.0 724650.0 ;
      RECT  129600.0 725850.0 130800.0 724650.0 ;
      RECT  127200.0 725850.0 128400.0 724650.0 ;
      RECT  129600.0 725850.0 130800.0 724650.0 ;
      RECT  132000.0 725850.0 133200.0 724650.0 ;
      RECT  132000.0 725850.0 133200.0 724650.0 ;
      RECT  129600.0 725850.0 130800.0 724650.0 ;
      RECT  134400.0 716550.0 135600.0 715350.0 ;
      RECT  134400.0 726450.0 135600.0 725250.0 ;
      RECT  132000.0 723300.0 130800.0 722100.0 ;
      RECT  129000.0 720600.0 127800.0 719400.0 ;
      RECT  129600.0 717150.0 130800.0 715950.0 ;
      RECT  132000.0 725850.0 133200.0 724650.0 ;
      RECT  133200.0 720600.0 132000.0 719400.0 ;
      RECT  127800.0 720600.0 129000.0 719400.0 ;
      RECT  130800.0 723300.0 132000.0 722100.0 ;
      RECT  132000.0 720600.0 133200.0 719400.0 ;
      RECT  125400.0 714450.0 139800.0 713550.0 ;
      RECT  125400.0 728250.0 139800.0 727350.0 ;
      RECT  146400.0 715950.0 147600.0 714000.0 ;
      RECT  146400.0 727800.0 147600.0 725850.0 ;
      RECT  141600.0 726450.0 142800.0 728250.0 ;
      RECT  141600.0 717150.0 142800.0 713550.0 ;
      RECT  144300.0 726450.0 145200.0 717150.0 ;
      RECT  141600.0 717150.0 142800.0 715950.0 ;
      RECT  144000.0 717150.0 145200.0 715950.0 ;
      RECT  144000.0 717150.0 145200.0 715950.0 ;
      RECT  141600.0 717150.0 142800.0 715950.0 ;
      RECT  141600.0 726450.0 142800.0 725250.0 ;
      RECT  144000.0 726450.0 145200.0 725250.0 ;
      RECT  144000.0 726450.0 145200.0 725250.0 ;
      RECT  141600.0 726450.0 142800.0 725250.0 ;
      RECT  146400.0 716550.0 147600.0 715350.0 ;
      RECT  146400.0 726450.0 147600.0 725250.0 ;
      RECT  142200.0 721800.0 143400.0 720600.0 ;
      RECT  142200.0 721800.0 143400.0 720600.0 ;
      RECT  144750.0 721650.0 145650.0 720750.0 ;
      RECT  139800.0 714450.0 149400.0 713550.0 ;
      RECT  139800.0 728250.0 149400.0 727350.0 ;
      RECT  112050.0 720600.0 113250.0 721800.0 ;
      RECT  114000.0 723000.0 115200.0 724200.0 ;
      RECT  130800.0 722100.0 129600.0 723300.0 ;
      RECT  122400.0 739650.0 123600.0 741600.0 ;
      RECT  122400.0 727800.0 123600.0 729750.0 ;
      RECT  117600.0 729150.0 118800.0 727350.0 ;
      RECT  117600.0 738450.0 118800.0 742050.0 ;
      RECT  120300.0 729150.0 121200.0 738450.0 ;
      RECT  117600.0 738450.0 118800.0 739650.0 ;
      RECT  120000.0 738450.0 121200.0 739650.0 ;
      RECT  120000.0 738450.0 121200.0 739650.0 ;
      RECT  117600.0 738450.0 118800.0 739650.0 ;
      RECT  117600.0 729150.0 118800.0 730350.0 ;
      RECT  120000.0 729150.0 121200.0 730350.0 ;
      RECT  120000.0 729150.0 121200.0 730350.0 ;
      RECT  117600.0 729150.0 118800.0 730350.0 ;
      RECT  122400.0 739050.0 123600.0 740250.0 ;
      RECT  122400.0 729150.0 123600.0 730350.0 ;
      RECT  118200.0 733800.0 119400.0 735000.0 ;
      RECT  118200.0 733800.0 119400.0 735000.0 ;
      RECT  120750.0 733950.0 121650.0 734850.0 ;
      RECT  115800.0 741150.0 125400.0 742050.0 ;
      RECT  115800.0 727350.0 125400.0 728250.0 ;
      RECT  127200.0 729750.0 128400.0 727350.0 ;
      RECT  127200.0 738450.0 128400.0 742050.0 ;
      RECT  132000.0 738450.0 133200.0 742050.0 ;
      RECT  134400.0 739650.0 135600.0 741600.0 ;
      RECT  134400.0 727800.0 135600.0 729750.0 ;
      RECT  127200.0 738450.0 128400.0 739650.0 ;
      RECT  129600.0 738450.0 130800.0 739650.0 ;
      RECT  129600.0 738450.0 130800.0 739650.0 ;
      RECT  127200.0 738450.0 128400.0 739650.0 ;
      RECT  129600.0 738450.0 130800.0 739650.0 ;
      RECT  132000.0 738450.0 133200.0 739650.0 ;
      RECT  132000.0 738450.0 133200.0 739650.0 ;
      RECT  129600.0 738450.0 130800.0 739650.0 ;
      RECT  127200.0 729750.0 128400.0 730950.0 ;
      RECT  129600.0 729750.0 130800.0 730950.0 ;
      RECT  129600.0 729750.0 130800.0 730950.0 ;
      RECT  127200.0 729750.0 128400.0 730950.0 ;
      RECT  129600.0 729750.0 130800.0 730950.0 ;
      RECT  132000.0 729750.0 133200.0 730950.0 ;
      RECT  132000.0 729750.0 133200.0 730950.0 ;
      RECT  129600.0 729750.0 130800.0 730950.0 ;
      RECT  134400.0 739050.0 135600.0 740250.0 ;
      RECT  134400.0 729150.0 135600.0 730350.0 ;
      RECT  132000.0 732300.0 130800.0 733500.0 ;
      RECT  129000.0 735000.0 127800.0 736200.0 ;
      RECT  129600.0 738450.0 130800.0 739650.0 ;
      RECT  132000.0 729750.0 133200.0 730950.0 ;
      RECT  133200.0 735000.0 132000.0 736200.0 ;
      RECT  127800.0 735000.0 129000.0 736200.0 ;
      RECT  130800.0 732300.0 132000.0 733500.0 ;
      RECT  132000.0 735000.0 133200.0 736200.0 ;
      RECT  125400.0 741150.0 139800.0 742050.0 ;
      RECT  125400.0 727350.0 139800.0 728250.0 ;
      RECT  146400.0 739650.0 147600.0 741600.0 ;
      RECT  146400.0 727800.0 147600.0 729750.0 ;
      RECT  141600.0 729150.0 142800.0 727350.0 ;
      RECT  141600.0 738450.0 142800.0 742050.0 ;
      RECT  144300.0 729150.0 145200.0 738450.0 ;
      RECT  141600.0 738450.0 142800.0 739650.0 ;
      RECT  144000.0 738450.0 145200.0 739650.0 ;
      RECT  144000.0 738450.0 145200.0 739650.0 ;
      RECT  141600.0 738450.0 142800.0 739650.0 ;
      RECT  141600.0 729150.0 142800.0 730350.0 ;
      RECT  144000.0 729150.0 145200.0 730350.0 ;
      RECT  144000.0 729150.0 145200.0 730350.0 ;
      RECT  141600.0 729150.0 142800.0 730350.0 ;
      RECT  146400.0 739050.0 147600.0 740250.0 ;
      RECT  146400.0 729150.0 147600.0 730350.0 ;
      RECT  142200.0 733800.0 143400.0 735000.0 ;
      RECT  142200.0 733800.0 143400.0 735000.0 ;
      RECT  144750.0 733950.0 145650.0 734850.0 ;
      RECT  139800.0 741150.0 149400.0 742050.0 ;
      RECT  139800.0 727350.0 149400.0 728250.0 ;
      RECT  112050.0 733800.0 113250.0 735000.0 ;
      RECT  114000.0 731400.0 115200.0 732600.0 ;
      RECT  130800.0 732300.0 129600.0 733500.0 ;
      RECT  122400.0 743550.0 123600.0 741600.0 ;
      RECT  122400.0 755400.0 123600.0 753450.0 ;
      RECT  117600.0 754050.0 118800.0 755850.0 ;
      RECT  117600.0 744750.0 118800.0 741150.0 ;
      RECT  120300.0 754050.0 121200.0 744750.0 ;
      RECT  117600.0 744750.0 118800.0 743550.0 ;
      RECT  120000.0 744750.0 121200.0 743550.0 ;
      RECT  120000.0 744750.0 121200.0 743550.0 ;
      RECT  117600.0 744750.0 118800.0 743550.0 ;
      RECT  117600.0 754050.0 118800.0 752850.0 ;
      RECT  120000.0 754050.0 121200.0 752850.0 ;
      RECT  120000.0 754050.0 121200.0 752850.0 ;
      RECT  117600.0 754050.0 118800.0 752850.0 ;
      RECT  122400.0 744150.0 123600.0 742950.0 ;
      RECT  122400.0 754050.0 123600.0 752850.0 ;
      RECT  118200.0 749400.0 119400.0 748200.0 ;
      RECT  118200.0 749400.0 119400.0 748200.0 ;
      RECT  120750.0 749250.0 121650.0 748350.0 ;
      RECT  115800.0 742050.0 125400.0 741150.0 ;
      RECT  115800.0 755850.0 125400.0 754950.0 ;
      RECT  127200.0 753450.0 128400.0 755850.0 ;
      RECT  127200.0 744750.0 128400.0 741150.0 ;
      RECT  132000.0 744750.0 133200.0 741150.0 ;
      RECT  134400.0 743550.0 135600.0 741600.0 ;
      RECT  134400.0 755400.0 135600.0 753450.0 ;
      RECT  127200.0 744750.0 128400.0 743550.0 ;
      RECT  129600.0 744750.0 130800.0 743550.0 ;
      RECT  129600.0 744750.0 130800.0 743550.0 ;
      RECT  127200.0 744750.0 128400.0 743550.0 ;
      RECT  129600.0 744750.0 130800.0 743550.0 ;
      RECT  132000.0 744750.0 133200.0 743550.0 ;
      RECT  132000.0 744750.0 133200.0 743550.0 ;
      RECT  129600.0 744750.0 130800.0 743550.0 ;
      RECT  127200.0 753450.0 128400.0 752250.0 ;
      RECT  129600.0 753450.0 130800.0 752250.0 ;
      RECT  129600.0 753450.0 130800.0 752250.0 ;
      RECT  127200.0 753450.0 128400.0 752250.0 ;
      RECT  129600.0 753450.0 130800.0 752250.0 ;
      RECT  132000.0 753450.0 133200.0 752250.0 ;
      RECT  132000.0 753450.0 133200.0 752250.0 ;
      RECT  129600.0 753450.0 130800.0 752250.0 ;
      RECT  134400.0 744150.0 135600.0 742950.0 ;
      RECT  134400.0 754050.0 135600.0 752850.0 ;
      RECT  132000.0 750900.0 130800.0 749700.0 ;
      RECT  129000.0 748200.0 127800.0 747000.0 ;
      RECT  129600.0 744750.0 130800.0 743550.0 ;
      RECT  132000.0 753450.0 133200.0 752250.0 ;
      RECT  133200.0 748200.0 132000.0 747000.0 ;
      RECT  127800.0 748200.0 129000.0 747000.0 ;
      RECT  130800.0 750900.0 132000.0 749700.0 ;
      RECT  132000.0 748200.0 133200.0 747000.0 ;
      RECT  125400.0 742050.0 139800.0 741150.0 ;
      RECT  125400.0 755850.0 139800.0 754950.0 ;
      RECT  146400.0 743550.0 147600.0 741600.0 ;
      RECT  146400.0 755400.0 147600.0 753450.0 ;
      RECT  141600.0 754050.0 142800.0 755850.0 ;
      RECT  141600.0 744750.0 142800.0 741150.0 ;
      RECT  144300.0 754050.0 145200.0 744750.0 ;
      RECT  141600.0 744750.0 142800.0 743550.0 ;
      RECT  144000.0 744750.0 145200.0 743550.0 ;
      RECT  144000.0 744750.0 145200.0 743550.0 ;
      RECT  141600.0 744750.0 142800.0 743550.0 ;
      RECT  141600.0 754050.0 142800.0 752850.0 ;
      RECT  144000.0 754050.0 145200.0 752850.0 ;
      RECT  144000.0 754050.0 145200.0 752850.0 ;
      RECT  141600.0 754050.0 142800.0 752850.0 ;
      RECT  146400.0 744150.0 147600.0 742950.0 ;
      RECT  146400.0 754050.0 147600.0 752850.0 ;
      RECT  142200.0 749400.0 143400.0 748200.0 ;
      RECT  142200.0 749400.0 143400.0 748200.0 ;
      RECT  144750.0 749250.0 145650.0 748350.0 ;
      RECT  139800.0 742050.0 149400.0 741150.0 ;
      RECT  139800.0 755850.0 149400.0 754950.0 ;
      RECT  112050.0 748200.0 113250.0 749400.0 ;
      RECT  114000.0 750600.0 115200.0 751800.0 ;
      RECT  130800.0 749700.0 129600.0 750900.0 ;
      RECT  122400.0 767250.0 123600.0 769200.0 ;
      RECT  122400.0 755400.0 123600.0 757350.0 ;
      RECT  117600.0 756750.0 118800.0 754950.0 ;
      RECT  117600.0 766050.0 118800.0 769650.0 ;
      RECT  120300.0 756750.0 121200.0 766050.0 ;
      RECT  117600.0 766050.0 118800.0 767250.0 ;
      RECT  120000.0 766050.0 121200.0 767250.0 ;
      RECT  120000.0 766050.0 121200.0 767250.0 ;
      RECT  117600.0 766050.0 118800.0 767250.0 ;
      RECT  117600.0 756750.0 118800.0 757950.0 ;
      RECT  120000.0 756750.0 121200.0 757950.0 ;
      RECT  120000.0 756750.0 121200.0 757950.0 ;
      RECT  117600.0 756750.0 118800.0 757950.0 ;
      RECT  122400.0 766650.0 123600.0 767850.0 ;
      RECT  122400.0 756750.0 123600.0 757950.0 ;
      RECT  118200.0 761400.0 119400.0 762600.0 ;
      RECT  118200.0 761400.0 119400.0 762600.0 ;
      RECT  120750.0 761550.0 121650.0 762450.0 ;
      RECT  115800.0 768750.0 125400.0 769650.0 ;
      RECT  115800.0 754950.0 125400.0 755850.0 ;
      RECT  127200.0 757350.0 128400.0 754950.0 ;
      RECT  127200.0 766050.0 128400.0 769650.0 ;
      RECT  132000.0 766050.0 133200.0 769650.0 ;
      RECT  134400.0 767250.0 135600.0 769200.0 ;
      RECT  134400.0 755400.0 135600.0 757350.0 ;
      RECT  127200.0 766050.0 128400.0 767250.0 ;
      RECT  129600.0 766050.0 130800.0 767250.0 ;
      RECT  129600.0 766050.0 130800.0 767250.0 ;
      RECT  127200.0 766050.0 128400.0 767250.0 ;
      RECT  129600.0 766050.0 130800.0 767250.0 ;
      RECT  132000.0 766050.0 133200.0 767250.0 ;
      RECT  132000.0 766050.0 133200.0 767250.0 ;
      RECT  129600.0 766050.0 130800.0 767250.0 ;
      RECT  127200.0 757350.0 128400.0 758550.0 ;
      RECT  129600.0 757350.0 130800.0 758550.0 ;
      RECT  129600.0 757350.0 130800.0 758550.0 ;
      RECT  127200.0 757350.0 128400.0 758550.0 ;
      RECT  129600.0 757350.0 130800.0 758550.0 ;
      RECT  132000.0 757350.0 133200.0 758550.0 ;
      RECT  132000.0 757350.0 133200.0 758550.0 ;
      RECT  129600.0 757350.0 130800.0 758550.0 ;
      RECT  134400.0 766650.0 135600.0 767850.0 ;
      RECT  134400.0 756750.0 135600.0 757950.0 ;
      RECT  132000.0 759900.0 130800.0 761100.0 ;
      RECT  129000.0 762600.0 127800.0 763800.0 ;
      RECT  129600.0 766050.0 130800.0 767250.0 ;
      RECT  132000.0 757350.0 133200.0 758550.0 ;
      RECT  133200.0 762600.0 132000.0 763800.0 ;
      RECT  127800.0 762600.0 129000.0 763800.0 ;
      RECT  130800.0 759900.0 132000.0 761100.0 ;
      RECT  132000.0 762600.0 133200.0 763800.0 ;
      RECT  125400.0 768750.0 139800.0 769650.0 ;
      RECT  125400.0 754950.0 139800.0 755850.0 ;
      RECT  146400.0 767250.0 147600.0 769200.0 ;
      RECT  146400.0 755400.0 147600.0 757350.0 ;
      RECT  141600.0 756750.0 142800.0 754950.0 ;
      RECT  141600.0 766050.0 142800.0 769650.0 ;
      RECT  144300.0 756750.0 145200.0 766050.0 ;
      RECT  141600.0 766050.0 142800.0 767250.0 ;
      RECT  144000.0 766050.0 145200.0 767250.0 ;
      RECT  144000.0 766050.0 145200.0 767250.0 ;
      RECT  141600.0 766050.0 142800.0 767250.0 ;
      RECT  141600.0 756750.0 142800.0 757950.0 ;
      RECT  144000.0 756750.0 145200.0 757950.0 ;
      RECT  144000.0 756750.0 145200.0 757950.0 ;
      RECT  141600.0 756750.0 142800.0 757950.0 ;
      RECT  146400.0 766650.0 147600.0 767850.0 ;
      RECT  146400.0 756750.0 147600.0 757950.0 ;
      RECT  142200.0 761400.0 143400.0 762600.0 ;
      RECT  142200.0 761400.0 143400.0 762600.0 ;
      RECT  144750.0 761550.0 145650.0 762450.0 ;
      RECT  139800.0 768750.0 149400.0 769650.0 ;
      RECT  139800.0 754950.0 149400.0 755850.0 ;
      RECT  112050.0 761400.0 113250.0 762600.0 ;
      RECT  114000.0 759000.0 115200.0 760200.0 ;
      RECT  130800.0 759900.0 129600.0 761100.0 ;
      RECT  122400.0 771150.0 123600.0 769200.0 ;
      RECT  122400.0 783000.0 123600.0 781050.0 ;
      RECT  117600.0 781650.0 118800.0 783450.0 ;
      RECT  117600.0 772350.0 118800.0 768750.0 ;
      RECT  120300.0 781650.0 121200.0 772350.0 ;
      RECT  117600.0 772350.0 118800.0 771150.0 ;
      RECT  120000.0 772350.0 121200.0 771150.0 ;
      RECT  120000.0 772350.0 121200.0 771150.0 ;
      RECT  117600.0 772350.0 118800.0 771150.0 ;
      RECT  117600.0 781650.0 118800.0 780450.0 ;
      RECT  120000.0 781650.0 121200.0 780450.0 ;
      RECT  120000.0 781650.0 121200.0 780450.0 ;
      RECT  117600.0 781650.0 118800.0 780450.0 ;
      RECT  122400.0 771750.0 123600.0 770550.0 ;
      RECT  122400.0 781650.0 123600.0 780450.0 ;
      RECT  118200.0 777000.0 119400.0 775800.0 ;
      RECT  118200.0 777000.0 119400.0 775800.0 ;
      RECT  120750.0 776850.0 121650.0 775950.0 ;
      RECT  115800.0 769650.0 125400.0 768750.0 ;
      RECT  115800.0 783450.0 125400.0 782550.0 ;
      RECT  127200.0 781050.0 128400.0 783450.0 ;
      RECT  127200.0 772350.0 128400.0 768750.0 ;
      RECT  132000.0 772350.0 133200.0 768750.0 ;
      RECT  134400.0 771150.0 135600.0 769200.0 ;
      RECT  134400.0 783000.0 135600.0 781050.0 ;
      RECT  127200.0 772350.0 128400.0 771150.0 ;
      RECT  129600.0 772350.0 130800.0 771150.0 ;
      RECT  129600.0 772350.0 130800.0 771150.0 ;
      RECT  127200.0 772350.0 128400.0 771150.0 ;
      RECT  129600.0 772350.0 130800.0 771150.0 ;
      RECT  132000.0 772350.0 133200.0 771150.0 ;
      RECT  132000.0 772350.0 133200.0 771150.0 ;
      RECT  129600.0 772350.0 130800.0 771150.0 ;
      RECT  127200.0 781050.0 128400.0 779850.0 ;
      RECT  129600.0 781050.0 130800.0 779850.0 ;
      RECT  129600.0 781050.0 130800.0 779850.0 ;
      RECT  127200.0 781050.0 128400.0 779850.0 ;
      RECT  129600.0 781050.0 130800.0 779850.0 ;
      RECT  132000.0 781050.0 133200.0 779850.0 ;
      RECT  132000.0 781050.0 133200.0 779850.0 ;
      RECT  129600.0 781050.0 130800.0 779850.0 ;
      RECT  134400.0 771750.0 135600.0 770550.0 ;
      RECT  134400.0 781650.0 135600.0 780450.0 ;
      RECT  132000.0 778500.0 130800.0 777300.0 ;
      RECT  129000.0 775800.0 127800.0 774600.0 ;
      RECT  129600.0 772350.0 130800.0 771150.0 ;
      RECT  132000.0 781050.0 133200.0 779850.0 ;
      RECT  133200.0 775800.0 132000.0 774600.0 ;
      RECT  127800.0 775800.0 129000.0 774600.0 ;
      RECT  130800.0 778500.0 132000.0 777300.0 ;
      RECT  132000.0 775800.0 133200.0 774600.0 ;
      RECT  125400.0 769650.0 139800.0 768750.0 ;
      RECT  125400.0 783450.0 139800.0 782550.0 ;
      RECT  146400.0 771150.0 147600.0 769200.0 ;
      RECT  146400.0 783000.0 147600.0 781050.0 ;
      RECT  141600.0 781650.0 142800.0 783450.0 ;
      RECT  141600.0 772350.0 142800.0 768750.0 ;
      RECT  144300.0 781650.0 145200.0 772350.0 ;
      RECT  141600.0 772350.0 142800.0 771150.0 ;
      RECT  144000.0 772350.0 145200.0 771150.0 ;
      RECT  144000.0 772350.0 145200.0 771150.0 ;
      RECT  141600.0 772350.0 142800.0 771150.0 ;
      RECT  141600.0 781650.0 142800.0 780450.0 ;
      RECT  144000.0 781650.0 145200.0 780450.0 ;
      RECT  144000.0 781650.0 145200.0 780450.0 ;
      RECT  141600.0 781650.0 142800.0 780450.0 ;
      RECT  146400.0 771750.0 147600.0 770550.0 ;
      RECT  146400.0 781650.0 147600.0 780450.0 ;
      RECT  142200.0 777000.0 143400.0 775800.0 ;
      RECT  142200.0 777000.0 143400.0 775800.0 ;
      RECT  144750.0 776850.0 145650.0 775950.0 ;
      RECT  139800.0 769650.0 149400.0 768750.0 ;
      RECT  139800.0 783450.0 149400.0 782550.0 ;
      RECT  112050.0 775800.0 113250.0 777000.0 ;
      RECT  114000.0 778200.0 115200.0 779400.0 ;
      RECT  130800.0 777300.0 129600.0 778500.0 ;
      RECT  122400.0 794850.0 123600.0 796800.0 ;
      RECT  122400.0 783000.0 123600.0 784950.0 ;
      RECT  117600.0 784350.0 118800.0 782550.0 ;
      RECT  117600.0 793650.0 118800.0 797250.0 ;
      RECT  120300.0 784350.0 121200.0 793650.0 ;
      RECT  117600.0 793650.0 118800.0 794850.0 ;
      RECT  120000.0 793650.0 121200.0 794850.0 ;
      RECT  120000.0 793650.0 121200.0 794850.0 ;
      RECT  117600.0 793650.0 118800.0 794850.0 ;
      RECT  117600.0 784350.0 118800.0 785550.0 ;
      RECT  120000.0 784350.0 121200.0 785550.0 ;
      RECT  120000.0 784350.0 121200.0 785550.0 ;
      RECT  117600.0 784350.0 118800.0 785550.0 ;
      RECT  122400.0 794250.0 123600.0 795450.0 ;
      RECT  122400.0 784350.0 123600.0 785550.0 ;
      RECT  118200.0 789000.0 119400.0 790200.0 ;
      RECT  118200.0 789000.0 119400.0 790200.0 ;
      RECT  120750.0 789150.0 121650.0 790050.0 ;
      RECT  115800.0 796350.0 125400.0 797250.0 ;
      RECT  115800.0 782550.0 125400.0 783450.0 ;
      RECT  127200.0 784950.0 128400.0 782550.0 ;
      RECT  127200.0 793650.0 128400.0 797250.0 ;
      RECT  132000.0 793650.0 133200.0 797250.0 ;
      RECT  134400.0 794850.0 135600.0 796800.0 ;
      RECT  134400.0 783000.0 135600.0 784950.0 ;
      RECT  127200.0 793650.0 128400.0 794850.0 ;
      RECT  129600.0 793650.0 130800.0 794850.0 ;
      RECT  129600.0 793650.0 130800.0 794850.0 ;
      RECT  127200.0 793650.0 128400.0 794850.0 ;
      RECT  129600.0 793650.0 130800.0 794850.0 ;
      RECT  132000.0 793650.0 133200.0 794850.0 ;
      RECT  132000.0 793650.0 133200.0 794850.0 ;
      RECT  129600.0 793650.0 130800.0 794850.0 ;
      RECT  127200.0 784950.0 128400.0 786150.0 ;
      RECT  129600.0 784950.0 130800.0 786150.0 ;
      RECT  129600.0 784950.0 130800.0 786150.0 ;
      RECT  127200.0 784950.0 128400.0 786150.0 ;
      RECT  129600.0 784950.0 130800.0 786150.0 ;
      RECT  132000.0 784950.0 133200.0 786150.0 ;
      RECT  132000.0 784950.0 133200.0 786150.0 ;
      RECT  129600.0 784950.0 130800.0 786150.0 ;
      RECT  134400.0 794250.0 135600.0 795450.0 ;
      RECT  134400.0 784350.0 135600.0 785550.0 ;
      RECT  132000.0 787500.0 130800.0 788700.0 ;
      RECT  129000.0 790200.0 127800.0 791400.0 ;
      RECT  129600.0 793650.0 130800.0 794850.0 ;
      RECT  132000.0 784950.0 133200.0 786150.0 ;
      RECT  133200.0 790200.0 132000.0 791400.0 ;
      RECT  127800.0 790200.0 129000.0 791400.0 ;
      RECT  130800.0 787500.0 132000.0 788700.0 ;
      RECT  132000.0 790200.0 133200.0 791400.0 ;
      RECT  125400.0 796350.0 139800.0 797250.0 ;
      RECT  125400.0 782550.0 139800.0 783450.0 ;
      RECT  146400.0 794850.0 147600.0 796800.0 ;
      RECT  146400.0 783000.0 147600.0 784950.0 ;
      RECT  141600.0 784350.0 142800.0 782550.0 ;
      RECT  141600.0 793650.0 142800.0 797250.0 ;
      RECT  144300.0 784350.0 145200.0 793650.0 ;
      RECT  141600.0 793650.0 142800.0 794850.0 ;
      RECT  144000.0 793650.0 145200.0 794850.0 ;
      RECT  144000.0 793650.0 145200.0 794850.0 ;
      RECT  141600.0 793650.0 142800.0 794850.0 ;
      RECT  141600.0 784350.0 142800.0 785550.0 ;
      RECT  144000.0 784350.0 145200.0 785550.0 ;
      RECT  144000.0 784350.0 145200.0 785550.0 ;
      RECT  141600.0 784350.0 142800.0 785550.0 ;
      RECT  146400.0 794250.0 147600.0 795450.0 ;
      RECT  146400.0 784350.0 147600.0 785550.0 ;
      RECT  142200.0 789000.0 143400.0 790200.0 ;
      RECT  142200.0 789000.0 143400.0 790200.0 ;
      RECT  144750.0 789150.0 145650.0 790050.0 ;
      RECT  139800.0 796350.0 149400.0 797250.0 ;
      RECT  139800.0 782550.0 149400.0 783450.0 ;
      RECT  112050.0 789000.0 113250.0 790200.0 ;
      RECT  114000.0 786600.0 115200.0 787800.0 ;
      RECT  130800.0 787500.0 129600.0 788700.0 ;
      RECT  122400.0 798750.0 123600.0 796800.0 ;
      RECT  122400.0 810600.0 123600.0 808650.0 ;
      RECT  117600.0 809250.0 118800.0 811050.0 ;
      RECT  117600.0 799950.0 118800.0 796350.0 ;
      RECT  120300.0 809250.0 121200.0 799950.0 ;
      RECT  117600.0 799950.0 118800.0 798750.0 ;
      RECT  120000.0 799950.0 121200.0 798750.0 ;
      RECT  120000.0 799950.0 121200.0 798750.0 ;
      RECT  117600.0 799950.0 118800.0 798750.0 ;
      RECT  117600.0 809250.0 118800.0 808050.0 ;
      RECT  120000.0 809250.0 121200.0 808050.0 ;
      RECT  120000.0 809250.0 121200.0 808050.0 ;
      RECT  117600.0 809250.0 118800.0 808050.0 ;
      RECT  122400.0 799350.0 123600.0 798150.0 ;
      RECT  122400.0 809250.0 123600.0 808050.0 ;
      RECT  118200.0 804600.0 119400.0 803400.0 ;
      RECT  118200.0 804600.0 119400.0 803400.0 ;
      RECT  120750.0 804450.0 121650.0 803550.0 ;
      RECT  115800.0 797250.0 125400.0 796350.0 ;
      RECT  115800.0 811050.0 125400.0 810150.0 ;
      RECT  127200.0 808650.0 128400.0 811050.0 ;
      RECT  127200.0 799950.0 128400.0 796350.0 ;
      RECT  132000.0 799950.0 133200.0 796350.0 ;
      RECT  134400.0 798750.0 135600.0 796800.0 ;
      RECT  134400.0 810600.0 135600.0 808650.0 ;
      RECT  127200.0 799950.0 128400.0 798750.0 ;
      RECT  129600.0 799950.0 130800.0 798750.0 ;
      RECT  129600.0 799950.0 130800.0 798750.0 ;
      RECT  127200.0 799950.0 128400.0 798750.0 ;
      RECT  129600.0 799950.0 130800.0 798750.0 ;
      RECT  132000.0 799950.0 133200.0 798750.0 ;
      RECT  132000.0 799950.0 133200.0 798750.0 ;
      RECT  129600.0 799950.0 130800.0 798750.0 ;
      RECT  127200.0 808650.0 128400.0 807450.0 ;
      RECT  129600.0 808650.0 130800.0 807450.0 ;
      RECT  129600.0 808650.0 130800.0 807450.0 ;
      RECT  127200.0 808650.0 128400.0 807450.0 ;
      RECT  129600.0 808650.0 130800.0 807450.0 ;
      RECT  132000.0 808650.0 133200.0 807450.0 ;
      RECT  132000.0 808650.0 133200.0 807450.0 ;
      RECT  129600.0 808650.0 130800.0 807450.0 ;
      RECT  134400.0 799350.0 135600.0 798150.0 ;
      RECT  134400.0 809250.0 135600.0 808050.0 ;
      RECT  132000.0 806100.0 130800.0 804900.0 ;
      RECT  129000.0 803400.0 127800.0 802200.0 ;
      RECT  129600.0 799950.0 130800.0 798750.0 ;
      RECT  132000.0 808650.0 133200.0 807450.0 ;
      RECT  133200.0 803400.0 132000.0 802200.0 ;
      RECT  127800.0 803400.0 129000.0 802200.0 ;
      RECT  130800.0 806100.0 132000.0 804900.0 ;
      RECT  132000.0 803400.0 133200.0 802200.0 ;
      RECT  125400.0 797250.0 139800.0 796350.0 ;
      RECT  125400.0 811050.0 139800.0 810150.0 ;
      RECT  146400.0 798750.0 147600.0 796800.0 ;
      RECT  146400.0 810600.0 147600.0 808650.0 ;
      RECT  141600.0 809250.0 142800.0 811050.0 ;
      RECT  141600.0 799950.0 142800.0 796350.0 ;
      RECT  144300.0 809250.0 145200.0 799950.0 ;
      RECT  141600.0 799950.0 142800.0 798750.0 ;
      RECT  144000.0 799950.0 145200.0 798750.0 ;
      RECT  144000.0 799950.0 145200.0 798750.0 ;
      RECT  141600.0 799950.0 142800.0 798750.0 ;
      RECT  141600.0 809250.0 142800.0 808050.0 ;
      RECT  144000.0 809250.0 145200.0 808050.0 ;
      RECT  144000.0 809250.0 145200.0 808050.0 ;
      RECT  141600.0 809250.0 142800.0 808050.0 ;
      RECT  146400.0 799350.0 147600.0 798150.0 ;
      RECT  146400.0 809250.0 147600.0 808050.0 ;
      RECT  142200.0 804600.0 143400.0 803400.0 ;
      RECT  142200.0 804600.0 143400.0 803400.0 ;
      RECT  144750.0 804450.0 145650.0 803550.0 ;
      RECT  139800.0 797250.0 149400.0 796350.0 ;
      RECT  139800.0 811050.0 149400.0 810150.0 ;
      RECT  112050.0 803400.0 113250.0 804600.0 ;
      RECT  114000.0 805800.0 115200.0 807000.0 ;
      RECT  130800.0 804900.0 129600.0 806100.0 ;
      RECT  122400.0 822450.0 123600.0 824400.0 ;
      RECT  122400.0 810600.0 123600.0 812550.0 ;
      RECT  117600.0 811950.0 118800.0 810150.0 ;
      RECT  117600.0 821250.0 118800.0 824850.0 ;
      RECT  120300.0 811950.0 121200.0 821250.0 ;
      RECT  117600.0 821250.0 118800.0 822450.0 ;
      RECT  120000.0 821250.0 121200.0 822450.0 ;
      RECT  120000.0 821250.0 121200.0 822450.0 ;
      RECT  117600.0 821250.0 118800.0 822450.0 ;
      RECT  117600.0 811950.0 118800.0 813150.0 ;
      RECT  120000.0 811950.0 121200.0 813150.0 ;
      RECT  120000.0 811950.0 121200.0 813150.0 ;
      RECT  117600.0 811950.0 118800.0 813150.0 ;
      RECT  122400.0 821850.0 123600.0 823050.0 ;
      RECT  122400.0 811950.0 123600.0 813150.0 ;
      RECT  118200.0 816600.0 119400.0 817800.0 ;
      RECT  118200.0 816600.0 119400.0 817800.0 ;
      RECT  120750.0 816750.0 121650.0 817650.0 ;
      RECT  115800.0 823950.0 125400.0 824850.0 ;
      RECT  115800.0 810150.0 125400.0 811050.0 ;
      RECT  127200.0 812550.0 128400.0 810150.0 ;
      RECT  127200.0 821250.0 128400.0 824850.0 ;
      RECT  132000.0 821250.0 133200.0 824850.0 ;
      RECT  134400.0 822450.0 135600.0 824400.0 ;
      RECT  134400.0 810600.0 135600.0 812550.0 ;
      RECT  127200.0 821250.0 128400.0 822450.0 ;
      RECT  129600.0 821250.0 130800.0 822450.0 ;
      RECT  129600.0 821250.0 130800.0 822450.0 ;
      RECT  127200.0 821250.0 128400.0 822450.0 ;
      RECT  129600.0 821250.0 130800.0 822450.0 ;
      RECT  132000.0 821250.0 133200.0 822450.0 ;
      RECT  132000.0 821250.0 133200.0 822450.0 ;
      RECT  129600.0 821250.0 130800.0 822450.0 ;
      RECT  127200.0 812550.0 128400.0 813750.0 ;
      RECT  129600.0 812550.0 130800.0 813750.0 ;
      RECT  129600.0 812550.0 130800.0 813750.0 ;
      RECT  127200.0 812550.0 128400.0 813750.0 ;
      RECT  129600.0 812550.0 130800.0 813750.0 ;
      RECT  132000.0 812550.0 133200.0 813750.0 ;
      RECT  132000.0 812550.0 133200.0 813750.0 ;
      RECT  129600.0 812550.0 130800.0 813750.0 ;
      RECT  134400.0 821850.0 135600.0 823050.0 ;
      RECT  134400.0 811950.0 135600.0 813150.0 ;
      RECT  132000.0 815100.0 130800.0 816300.0 ;
      RECT  129000.0 817800.0 127800.0 819000.0 ;
      RECT  129600.0 821250.0 130800.0 822450.0 ;
      RECT  132000.0 812550.0 133200.0 813750.0 ;
      RECT  133200.0 817800.0 132000.0 819000.0 ;
      RECT  127800.0 817800.0 129000.0 819000.0 ;
      RECT  130800.0 815100.0 132000.0 816300.0 ;
      RECT  132000.0 817800.0 133200.0 819000.0 ;
      RECT  125400.0 823950.0 139800.0 824850.0 ;
      RECT  125400.0 810150.0 139800.0 811050.0 ;
      RECT  146400.0 822450.0 147600.0 824400.0 ;
      RECT  146400.0 810600.0 147600.0 812550.0 ;
      RECT  141600.0 811950.0 142800.0 810150.0 ;
      RECT  141600.0 821250.0 142800.0 824850.0 ;
      RECT  144300.0 811950.0 145200.0 821250.0 ;
      RECT  141600.0 821250.0 142800.0 822450.0 ;
      RECT  144000.0 821250.0 145200.0 822450.0 ;
      RECT  144000.0 821250.0 145200.0 822450.0 ;
      RECT  141600.0 821250.0 142800.0 822450.0 ;
      RECT  141600.0 811950.0 142800.0 813150.0 ;
      RECT  144000.0 811950.0 145200.0 813150.0 ;
      RECT  144000.0 811950.0 145200.0 813150.0 ;
      RECT  141600.0 811950.0 142800.0 813150.0 ;
      RECT  146400.0 821850.0 147600.0 823050.0 ;
      RECT  146400.0 811950.0 147600.0 813150.0 ;
      RECT  142200.0 816600.0 143400.0 817800.0 ;
      RECT  142200.0 816600.0 143400.0 817800.0 ;
      RECT  144750.0 816750.0 145650.0 817650.0 ;
      RECT  139800.0 823950.0 149400.0 824850.0 ;
      RECT  139800.0 810150.0 149400.0 811050.0 ;
      RECT  112050.0 816600.0 113250.0 817800.0 ;
      RECT  114000.0 814200.0 115200.0 815400.0 ;
      RECT  130800.0 815100.0 129600.0 816300.0 ;
      RECT  122400.0 826350.0 123600.0 824400.0 ;
      RECT  122400.0 838200.0 123600.0 836250.0 ;
      RECT  117600.0 836850.0 118800.0 838650.0 ;
      RECT  117600.0 827550.0 118800.0 823950.0 ;
      RECT  120300.0 836850.0 121200.0 827550.0 ;
      RECT  117600.0 827550.0 118800.0 826350.0 ;
      RECT  120000.0 827550.0 121200.0 826350.0 ;
      RECT  120000.0 827550.0 121200.0 826350.0 ;
      RECT  117600.0 827550.0 118800.0 826350.0 ;
      RECT  117600.0 836850.0 118800.0 835650.0 ;
      RECT  120000.0 836850.0 121200.0 835650.0 ;
      RECT  120000.0 836850.0 121200.0 835650.0 ;
      RECT  117600.0 836850.0 118800.0 835650.0 ;
      RECT  122400.0 826950.0 123600.0 825750.0 ;
      RECT  122400.0 836850.0 123600.0 835650.0 ;
      RECT  118200.0 832200.0 119400.0 831000.0 ;
      RECT  118200.0 832200.0 119400.0 831000.0 ;
      RECT  120750.0 832050.0 121650.0 831150.0 ;
      RECT  115800.0 824850.0 125400.0 823950.0 ;
      RECT  115800.0 838650.0 125400.0 837750.0 ;
      RECT  127200.0 836250.0 128400.0 838650.0 ;
      RECT  127200.0 827550.0 128400.0 823950.0 ;
      RECT  132000.0 827550.0 133200.0 823950.0 ;
      RECT  134400.0 826350.0 135600.0 824400.0 ;
      RECT  134400.0 838200.0 135600.0 836250.0 ;
      RECT  127200.0 827550.0 128400.0 826350.0 ;
      RECT  129600.0 827550.0 130800.0 826350.0 ;
      RECT  129600.0 827550.0 130800.0 826350.0 ;
      RECT  127200.0 827550.0 128400.0 826350.0 ;
      RECT  129600.0 827550.0 130800.0 826350.0 ;
      RECT  132000.0 827550.0 133200.0 826350.0 ;
      RECT  132000.0 827550.0 133200.0 826350.0 ;
      RECT  129600.0 827550.0 130800.0 826350.0 ;
      RECT  127200.0 836250.0 128400.0 835050.0 ;
      RECT  129600.0 836250.0 130800.0 835050.0 ;
      RECT  129600.0 836250.0 130800.0 835050.0 ;
      RECT  127200.0 836250.0 128400.0 835050.0 ;
      RECT  129600.0 836250.0 130800.0 835050.0 ;
      RECT  132000.0 836250.0 133200.0 835050.0 ;
      RECT  132000.0 836250.0 133200.0 835050.0 ;
      RECT  129600.0 836250.0 130800.0 835050.0 ;
      RECT  134400.0 826950.0 135600.0 825750.0 ;
      RECT  134400.0 836850.0 135600.0 835650.0 ;
      RECT  132000.0 833700.0 130800.0 832500.0 ;
      RECT  129000.0 831000.0 127800.0 829800.0 ;
      RECT  129600.0 827550.0 130800.0 826350.0 ;
      RECT  132000.0 836250.0 133200.0 835050.0 ;
      RECT  133200.0 831000.0 132000.0 829800.0 ;
      RECT  127800.0 831000.0 129000.0 829800.0 ;
      RECT  130800.0 833700.0 132000.0 832500.0 ;
      RECT  132000.0 831000.0 133200.0 829800.0 ;
      RECT  125400.0 824850.0 139800.0 823950.0 ;
      RECT  125400.0 838650.0 139800.0 837750.0 ;
      RECT  146400.0 826350.0 147600.0 824400.0 ;
      RECT  146400.0 838200.0 147600.0 836250.0 ;
      RECT  141600.0 836850.0 142800.0 838650.0 ;
      RECT  141600.0 827550.0 142800.0 823950.0 ;
      RECT  144300.0 836850.0 145200.0 827550.0 ;
      RECT  141600.0 827550.0 142800.0 826350.0 ;
      RECT  144000.0 827550.0 145200.0 826350.0 ;
      RECT  144000.0 827550.0 145200.0 826350.0 ;
      RECT  141600.0 827550.0 142800.0 826350.0 ;
      RECT  141600.0 836850.0 142800.0 835650.0 ;
      RECT  144000.0 836850.0 145200.0 835650.0 ;
      RECT  144000.0 836850.0 145200.0 835650.0 ;
      RECT  141600.0 836850.0 142800.0 835650.0 ;
      RECT  146400.0 826950.0 147600.0 825750.0 ;
      RECT  146400.0 836850.0 147600.0 835650.0 ;
      RECT  142200.0 832200.0 143400.0 831000.0 ;
      RECT  142200.0 832200.0 143400.0 831000.0 ;
      RECT  144750.0 832050.0 145650.0 831150.0 ;
      RECT  139800.0 824850.0 149400.0 823950.0 ;
      RECT  139800.0 838650.0 149400.0 837750.0 ;
      RECT  112050.0 831000.0 113250.0 832200.0 ;
      RECT  114000.0 833400.0 115200.0 834600.0 ;
      RECT  130800.0 832500.0 129600.0 833700.0 ;
      RECT  122400.0 850050.0 123600.0 852000.0 ;
      RECT  122400.0 838200.0 123600.0 840150.0 ;
      RECT  117600.0 839550.0 118800.0 837750.0 ;
      RECT  117600.0 848850.0 118800.0 852450.0 ;
      RECT  120300.0 839550.0 121200.0 848850.0 ;
      RECT  117600.0 848850.0 118800.0 850050.0 ;
      RECT  120000.0 848850.0 121200.0 850050.0 ;
      RECT  120000.0 848850.0 121200.0 850050.0 ;
      RECT  117600.0 848850.0 118800.0 850050.0 ;
      RECT  117600.0 839550.0 118800.0 840750.0 ;
      RECT  120000.0 839550.0 121200.0 840750.0 ;
      RECT  120000.0 839550.0 121200.0 840750.0 ;
      RECT  117600.0 839550.0 118800.0 840750.0 ;
      RECT  122400.0 849450.0 123600.0 850650.0 ;
      RECT  122400.0 839550.0 123600.0 840750.0 ;
      RECT  118200.0 844200.0 119400.0 845400.0 ;
      RECT  118200.0 844200.0 119400.0 845400.0 ;
      RECT  120750.0 844350.0 121650.0 845250.0 ;
      RECT  115800.0 851550.0 125400.0 852450.0 ;
      RECT  115800.0 837750.0 125400.0 838650.0 ;
      RECT  127200.0 840150.0 128400.0 837750.0 ;
      RECT  127200.0 848850.0 128400.0 852450.0 ;
      RECT  132000.0 848850.0 133200.0 852450.0 ;
      RECT  134400.0 850050.0 135600.0 852000.0 ;
      RECT  134400.0 838200.0 135600.0 840150.0 ;
      RECT  127200.0 848850.0 128400.0 850050.0 ;
      RECT  129600.0 848850.0 130800.0 850050.0 ;
      RECT  129600.0 848850.0 130800.0 850050.0 ;
      RECT  127200.0 848850.0 128400.0 850050.0 ;
      RECT  129600.0 848850.0 130800.0 850050.0 ;
      RECT  132000.0 848850.0 133200.0 850050.0 ;
      RECT  132000.0 848850.0 133200.0 850050.0 ;
      RECT  129600.0 848850.0 130800.0 850050.0 ;
      RECT  127200.0 840150.0 128400.0 841350.0 ;
      RECT  129600.0 840150.0 130800.0 841350.0 ;
      RECT  129600.0 840150.0 130800.0 841350.0 ;
      RECT  127200.0 840150.0 128400.0 841350.0 ;
      RECT  129600.0 840150.0 130800.0 841350.0 ;
      RECT  132000.0 840150.0 133200.0 841350.0 ;
      RECT  132000.0 840150.0 133200.0 841350.0 ;
      RECT  129600.0 840150.0 130800.0 841350.0 ;
      RECT  134400.0 849450.0 135600.0 850650.0 ;
      RECT  134400.0 839550.0 135600.0 840750.0 ;
      RECT  132000.0 842700.0 130800.0 843900.0 ;
      RECT  129000.0 845400.0 127800.0 846600.0 ;
      RECT  129600.0 848850.0 130800.0 850050.0 ;
      RECT  132000.0 840150.0 133200.0 841350.0 ;
      RECT  133200.0 845400.0 132000.0 846600.0 ;
      RECT  127800.0 845400.0 129000.0 846600.0 ;
      RECT  130800.0 842700.0 132000.0 843900.0 ;
      RECT  132000.0 845400.0 133200.0 846600.0 ;
      RECT  125400.0 851550.0 139800.0 852450.0 ;
      RECT  125400.0 837750.0 139800.0 838650.0 ;
      RECT  146400.0 850050.0 147600.0 852000.0 ;
      RECT  146400.0 838200.0 147600.0 840150.0 ;
      RECT  141600.0 839550.0 142800.0 837750.0 ;
      RECT  141600.0 848850.0 142800.0 852450.0 ;
      RECT  144300.0 839550.0 145200.0 848850.0 ;
      RECT  141600.0 848850.0 142800.0 850050.0 ;
      RECT  144000.0 848850.0 145200.0 850050.0 ;
      RECT  144000.0 848850.0 145200.0 850050.0 ;
      RECT  141600.0 848850.0 142800.0 850050.0 ;
      RECT  141600.0 839550.0 142800.0 840750.0 ;
      RECT  144000.0 839550.0 145200.0 840750.0 ;
      RECT  144000.0 839550.0 145200.0 840750.0 ;
      RECT  141600.0 839550.0 142800.0 840750.0 ;
      RECT  146400.0 849450.0 147600.0 850650.0 ;
      RECT  146400.0 839550.0 147600.0 840750.0 ;
      RECT  142200.0 844200.0 143400.0 845400.0 ;
      RECT  142200.0 844200.0 143400.0 845400.0 ;
      RECT  144750.0 844350.0 145650.0 845250.0 ;
      RECT  139800.0 851550.0 149400.0 852450.0 ;
      RECT  139800.0 837750.0 149400.0 838650.0 ;
      RECT  112050.0 844200.0 113250.0 845400.0 ;
      RECT  114000.0 841800.0 115200.0 843000.0 ;
      RECT  130800.0 842700.0 129600.0 843900.0 ;
      RECT  122400.0 853950.0 123600.0 852000.0 ;
      RECT  122400.0 865800.0 123600.0 863850.0 ;
      RECT  117600.0 864450.0 118800.0 866250.0 ;
      RECT  117600.0 855150.0 118800.0 851550.0 ;
      RECT  120300.0 864450.0 121200.0 855150.0 ;
      RECT  117600.0 855150.0 118800.0 853950.0 ;
      RECT  120000.0 855150.0 121200.0 853950.0 ;
      RECT  120000.0 855150.0 121200.0 853950.0 ;
      RECT  117600.0 855150.0 118800.0 853950.0 ;
      RECT  117600.0 864450.0 118800.0 863250.0 ;
      RECT  120000.0 864450.0 121200.0 863250.0 ;
      RECT  120000.0 864450.0 121200.0 863250.0 ;
      RECT  117600.0 864450.0 118800.0 863250.0 ;
      RECT  122400.0 854550.0 123600.0 853350.0 ;
      RECT  122400.0 864450.0 123600.0 863250.0 ;
      RECT  118200.0 859800.0 119400.0 858600.0 ;
      RECT  118200.0 859800.0 119400.0 858600.0 ;
      RECT  120750.0 859650.0 121650.0 858750.0 ;
      RECT  115800.0 852450.0 125400.0 851550.0 ;
      RECT  115800.0 866250.0 125400.0 865350.0 ;
      RECT  127200.0 863850.0 128400.0 866250.0 ;
      RECT  127200.0 855150.0 128400.0 851550.0 ;
      RECT  132000.0 855150.0 133200.0 851550.0 ;
      RECT  134400.0 853950.0 135600.0 852000.0 ;
      RECT  134400.0 865800.0 135600.0 863850.0 ;
      RECT  127200.0 855150.0 128400.0 853950.0 ;
      RECT  129600.0 855150.0 130800.0 853950.0 ;
      RECT  129600.0 855150.0 130800.0 853950.0 ;
      RECT  127200.0 855150.0 128400.0 853950.0 ;
      RECT  129600.0 855150.0 130800.0 853950.0 ;
      RECT  132000.0 855150.0 133200.0 853950.0 ;
      RECT  132000.0 855150.0 133200.0 853950.0 ;
      RECT  129600.0 855150.0 130800.0 853950.0 ;
      RECT  127200.0 863850.0 128400.0 862650.0 ;
      RECT  129600.0 863850.0 130800.0 862650.0 ;
      RECT  129600.0 863850.0 130800.0 862650.0 ;
      RECT  127200.0 863850.0 128400.0 862650.0 ;
      RECT  129600.0 863850.0 130800.0 862650.0 ;
      RECT  132000.0 863850.0 133200.0 862650.0 ;
      RECT  132000.0 863850.0 133200.0 862650.0 ;
      RECT  129600.0 863850.0 130800.0 862650.0 ;
      RECT  134400.0 854550.0 135600.0 853350.0 ;
      RECT  134400.0 864450.0 135600.0 863250.0 ;
      RECT  132000.0 861300.0 130800.0 860100.0 ;
      RECT  129000.0 858600.0 127800.0 857400.0 ;
      RECT  129600.0 855150.0 130800.0 853950.0 ;
      RECT  132000.0 863850.0 133200.0 862650.0 ;
      RECT  133200.0 858600.0 132000.0 857400.0 ;
      RECT  127800.0 858600.0 129000.0 857400.0 ;
      RECT  130800.0 861300.0 132000.0 860100.0 ;
      RECT  132000.0 858600.0 133200.0 857400.0 ;
      RECT  125400.0 852450.0 139800.0 851550.0 ;
      RECT  125400.0 866250.0 139800.0 865350.0 ;
      RECT  146400.0 853950.0 147600.0 852000.0 ;
      RECT  146400.0 865800.0 147600.0 863850.0 ;
      RECT  141600.0 864450.0 142800.0 866250.0 ;
      RECT  141600.0 855150.0 142800.0 851550.0 ;
      RECT  144300.0 864450.0 145200.0 855150.0 ;
      RECT  141600.0 855150.0 142800.0 853950.0 ;
      RECT  144000.0 855150.0 145200.0 853950.0 ;
      RECT  144000.0 855150.0 145200.0 853950.0 ;
      RECT  141600.0 855150.0 142800.0 853950.0 ;
      RECT  141600.0 864450.0 142800.0 863250.0 ;
      RECT  144000.0 864450.0 145200.0 863250.0 ;
      RECT  144000.0 864450.0 145200.0 863250.0 ;
      RECT  141600.0 864450.0 142800.0 863250.0 ;
      RECT  146400.0 854550.0 147600.0 853350.0 ;
      RECT  146400.0 864450.0 147600.0 863250.0 ;
      RECT  142200.0 859800.0 143400.0 858600.0 ;
      RECT  142200.0 859800.0 143400.0 858600.0 ;
      RECT  144750.0 859650.0 145650.0 858750.0 ;
      RECT  139800.0 852450.0 149400.0 851550.0 ;
      RECT  139800.0 866250.0 149400.0 865350.0 ;
      RECT  112050.0 858600.0 113250.0 859800.0 ;
      RECT  114000.0 861000.0 115200.0 862200.0 ;
      RECT  130800.0 860100.0 129600.0 861300.0 ;
      RECT  122400.0 877650.0 123600.0 879600.0 ;
      RECT  122400.0 865800.0 123600.0 867750.0 ;
      RECT  117600.0 867150.0 118800.0 865350.0 ;
      RECT  117600.0 876450.0 118800.0 880050.0 ;
      RECT  120300.0 867150.0 121200.0 876450.0 ;
      RECT  117600.0 876450.0 118800.0 877650.0 ;
      RECT  120000.0 876450.0 121200.0 877650.0 ;
      RECT  120000.0 876450.0 121200.0 877650.0 ;
      RECT  117600.0 876450.0 118800.0 877650.0 ;
      RECT  117600.0 867150.0 118800.0 868350.0 ;
      RECT  120000.0 867150.0 121200.0 868350.0 ;
      RECT  120000.0 867150.0 121200.0 868350.0 ;
      RECT  117600.0 867150.0 118800.0 868350.0 ;
      RECT  122400.0 877050.0 123600.0 878250.0 ;
      RECT  122400.0 867150.0 123600.0 868350.0 ;
      RECT  118200.0 871800.0 119400.0 873000.0 ;
      RECT  118200.0 871800.0 119400.0 873000.0 ;
      RECT  120750.0 871950.0 121650.0 872850.0 ;
      RECT  115800.0 879150.0 125400.0 880050.0 ;
      RECT  115800.0 865350.0 125400.0 866250.0 ;
      RECT  127200.0 867750.0 128400.0 865350.0 ;
      RECT  127200.0 876450.0 128400.0 880050.0 ;
      RECT  132000.0 876450.0 133200.0 880050.0 ;
      RECT  134400.0 877650.0 135600.0 879600.0 ;
      RECT  134400.0 865800.0 135600.0 867750.0 ;
      RECT  127200.0 876450.0 128400.0 877650.0 ;
      RECT  129600.0 876450.0 130800.0 877650.0 ;
      RECT  129600.0 876450.0 130800.0 877650.0 ;
      RECT  127200.0 876450.0 128400.0 877650.0 ;
      RECT  129600.0 876450.0 130800.0 877650.0 ;
      RECT  132000.0 876450.0 133200.0 877650.0 ;
      RECT  132000.0 876450.0 133200.0 877650.0 ;
      RECT  129600.0 876450.0 130800.0 877650.0 ;
      RECT  127200.0 867750.0 128400.0 868950.0 ;
      RECT  129600.0 867750.0 130800.0 868950.0 ;
      RECT  129600.0 867750.0 130800.0 868950.0 ;
      RECT  127200.0 867750.0 128400.0 868950.0 ;
      RECT  129600.0 867750.0 130800.0 868950.0 ;
      RECT  132000.0 867750.0 133200.0 868950.0 ;
      RECT  132000.0 867750.0 133200.0 868950.0 ;
      RECT  129600.0 867750.0 130800.0 868950.0 ;
      RECT  134400.0 877050.0 135600.0 878250.0 ;
      RECT  134400.0 867150.0 135600.0 868350.0 ;
      RECT  132000.0 870300.0 130800.0 871500.0 ;
      RECT  129000.0 873000.0 127800.0 874200.0 ;
      RECT  129600.0 876450.0 130800.0 877650.0 ;
      RECT  132000.0 867750.0 133200.0 868950.0 ;
      RECT  133200.0 873000.0 132000.0 874200.0 ;
      RECT  127800.0 873000.0 129000.0 874200.0 ;
      RECT  130800.0 870300.0 132000.0 871500.0 ;
      RECT  132000.0 873000.0 133200.0 874200.0 ;
      RECT  125400.0 879150.0 139800.0 880050.0 ;
      RECT  125400.0 865350.0 139800.0 866250.0 ;
      RECT  146400.0 877650.0 147600.0 879600.0 ;
      RECT  146400.0 865800.0 147600.0 867750.0 ;
      RECT  141600.0 867150.0 142800.0 865350.0 ;
      RECT  141600.0 876450.0 142800.0 880050.0 ;
      RECT  144300.0 867150.0 145200.0 876450.0 ;
      RECT  141600.0 876450.0 142800.0 877650.0 ;
      RECT  144000.0 876450.0 145200.0 877650.0 ;
      RECT  144000.0 876450.0 145200.0 877650.0 ;
      RECT  141600.0 876450.0 142800.0 877650.0 ;
      RECT  141600.0 867150.0 142800.0 868350.0 ;
      RECT  144000.0 867150.0 145200.0 868350.0 ;
      RECT  144000.0 867150.0 145200.0 868350.0 ;
      RECT  141600.0 867150.0 142800.0 868350.0 ;
      RECT  146400.0 877050.0 147600.0 878250.0 ;
      RECT  146400.0 867150.0 147600.0 868350.0 ;
      RECT  142200.0 871800.0 143400.0 873000.0 ;
      RECT  142200.0 871800.0 143400.0 873000.0 ;
      RECT  144750.0 871950.0 145650.0 872850.0 ;
      RECT  139800.0 879150.0 149400.0 880050.0 ;
      RECT  139800.0 865350.0 149400.0 866250.0 ;
      RECT  112050.0 871800.0 113250.0 873000.0 ;
      RECT  114000.0 869400.0 115200.0 870600.0 ;
      RECT  130800.0 870300.0 129600.0 871500.0 ;
      RECT  122400.0 881550.0 123600.0 879600.0 ;
      RECT  122400.0 893400.0 123600.0 891450.0 ;
      RECT  117600.0 892050.0 118800.0 893850.0 ;
      RECT  117600.0 882750.0 118800.0 879150.0 ;
      RECT  120300.0 892050.0 121200.0 882750.0 ;
      RECT  117600.0 882750.0 118800.0 881550.0 ;
      RECT  120000.0 882750.0 121200.0 881550.0 ;
      RECT  120000.0 882750.0 121200.0 881550.0 ;
      RECT  117600.0 882750.0 118800.0 881550.0 ;
      RECT  117600.0 892050.0 118800.0 890850.0 ;
      RECT  120000.0 892050.0 121200.0 890850.0 ;
      RECT  120000.0 892050.0 121200.0 890850.0 ;
      RECT  117600.0 892050.0 118800.0 890850.0 ;
      RECT  122400.0 882150.0 123600.0 880950.0 ;
      RECT  122400.0 892050.0 123600.0 890850.0 ;
      RECT  118200.0 887400.0 119400.0 886200.0 ;
      RECT  118200.0 887400.0 119400.0 886200.0 ;
      RECT  120750.0 887250.0 121650.0 886350.0 ;
      RECT  115800.0 880050.0 125400.0 879150.0 ;
      RECT  115800.0 893850.0 125400.0 892950.0 ;
      RECT  127200.0 891450.0 128400.0 893850.0 ;
      RECT  127200.0 882750.0 128400.0 879150.0 ;
      RECT  132000.0 882750.0 133200.0 879150.0 ;
      RECT  134400.0 881550.0 135600.0 879600.0 ;
      RECT  134400.0 893400.0 135600.0 891450.0 ;
      RECT  127200.0 882750.0 128400.0 881550.0 ;
      RECT  129600.0 882750.0 130800.0 881550.0 ;
      RECT  129600.0 882750.0 130800.0 881550.0 ;
      RECT  127200.0 882750.0 128400.0 881550.0 ;
      RECT  129600.0 882750.0 130800.0 881550.0 ;
      RECT  132000.0 882750.0 133200.0 881550.0 ;
      RECT  132000.0 882750.0 133200.0 881550.0 ;
      RECT  129600.0 882750.0 130800.0 881550.0 ;
      RECT  127200.0 891450.0 128400.0 890250.0 ;
      RECT  129600.0 891450.0 130800.0 890250.0 ;
      RECT  129600.0 891450.0 130800.0 890250.0 ;
      RECT  127200.0 891450.0 128400.0 890250.0 ;
      RECT  129600.0 891450.0 130800.0 890250.0 ;
      RECT  132000.0 891450.0 133200.0 890250.0 ;
      RECT  132000.0 891450.0 133200.0 890250.0 ;
      RECT  129600.0 891450.0 130800.0 890250.0 ;
      RECT  134400.0 882150.0 135600.0 880950.0 ;
      RECT  134400.0 892050.0 135600.0 890850.0 ;
      RECT  132000.0 888900.0 130800.0 887700.0 ;
      RECT  129000.0 886200.0 127800.0 885000.0 ;
      RECT  129600.0 882750.0 130800.0 881550.0 ;
      RECT  132000.0 891450.0 133200.0 890250.0 ;
      RECT  133200.0 886200.0 132000.0 885000.0 ;
      RECT  127800.0 886200.0 129000.0 885000.0 ;
      RECT  130800.0 888900.0 132000.0 887700.0 ;
      RECT  132000.0 886200.0 133200.0 885000.0 ;
      RECT  125400.0 880050.0 139800.0 879150.0 ;
      RECT  125400.0 893850.0 139800.0 892950.0 ;
      RECT  146400.0 881550.0 147600.0 879600.0 ;
      RECT  146400.0 893400.0 147600.0 891450.0 ;
      RECT  141600.0 892050.0 142800.0 893850.0 ;
      RECT  141600.0 882750.0 142800.0 879150.0 ;
      RECT  144300.0 892050.0 145200.0 882750.0 ;
      RECT  141600.0 882750.0 142800.0 881550.0 ;
      RECT  144000.0 882750.0 145200.0 881550.0 ;
      RECT  144000.0 882750.0 145200.0 881550.0 ;
      RECT  141600.0 882750.0 142800.0 881550.0 ;
      RECT  141600.0 892050.0 142800.0 890850.0 ;
      RECT  144000.0 892050.0 145200.0 890850.0 ;
      RECT  144000.0 892050.0 145200.0 890850.0 ;
      RECT  141600.0 892050.0 142800.0 890850.0 ;
      RECT  146400.0 882150.0 147600.0 880950.0 ;
      RECT  146400.0 892050.0 147600.0 890850.0 ;
      RECT  142200.0 887400.0 143400.0 886200.0 ;
      RECT  142200.0 887400.0 143400.0 886200.0 ;
      RECT  144750.0 887250.0 145650.0 886350.0 ;
      RECT  139800.0 880050.0 149400.0 879150.0 ;
      RECT  139800.0 893850.0 149400.0 892950.0 ;
      RECT  112050.0 886200.0 113250.0 887400.0 ;
      RECT  114000.0 888600.0 115200.0 889800.0 ;
      RECT  130800.0 887700.0 129600.0 888900.0 ;
      RECT  122400.0 905250.0 123600.0 907200.0 ;
      RECT  122400.0 893400.0 123600.0 895350.0 ;
      RECT  117600.0 894750.0 118800.0 892950.0 ;
      RECT  117600.0 904050.0 118800.0 907650.0 ;
      RECT  120300.0 894750.0 121200.0 904050.0 ;
      RECT  117600.0 904050.0 118800.0 905250.0 ;
      RECT  120000.0 904050.0 121200.0 905250.0 ;
      RECT  120000.0 904050.0 121200.0 905250.0 ;
      RECT  117600.0 904050.0 118800.0 905250.0 ;
      RECT  117600.0 894750.0 118800.0 895950.0 ;
      RECT  120000.0 894750.0 121200.0 895950.0 ;
      RECT  120000.0 894750.0 121200.0 895950.0 ;
      RECT  117600.0 894750.0 118800.0 895950.0 ;
      RECT  122400.0 904650.0 123600.0 905850.0 ;
      RECT  122400.0 894750.0 123600.0 895950.0 ;
      RECT  118200.0 899400.0 119400.0 900600.0 ;
      RECT  118200.0 899400.0 119400.0 900600.0 ;
      RECT  120750.0 899550.0 121650.0 900450.0 ;
      RECT  115800.0 906750.0 125400.0 907650.0 ;
      RECT  115800.0 892950.0 125400.0 893850.0 ;
      RECT  127200.0 895350.0 128400.0 892950.0 ;
      RECT  127200.0 904050.0 128400.0 907650.0 ;
      RECT  132000.0 904050.0 133200.0 907650.0 ;
      RECT  134400.0 905250.0 135600.0 907200.0 ;
      RECT  134400.0 893400.0 135600.0 895350.0 ;
      RECT  127200.0 904050.0 128400.0 905250.0 ;
      RECT  129600.0 904050.0 130800.0 905250.0 ;
      RECT  129600.0 904050.0 130800.0 905250.0 ;
      RECT  127200.0 904050.0 128400.0 905250.0 ;
      RECT  129600.0 904050.0 130800.0 905250.0 ;
      RECT  132000.0 904050.0 133200.0 905250.0 ;
      RECT  132000.0 904050.0 133200.0 905250.0 ;
      RECT  129600.0 904050.0 130800.0 905250.0 ;
      RECT  127200.0 895350.0 128400.0 896550.0 ;
      RECT  129600.0 895350.0 130800.0 896550.0 ;
      RECT  129600.0 895350.0 130800.0 896550.0 ;
      RECT  127200.0 895350.0 128400.0 896550.0 ;
      RECT  129600.0 895350.0 130800.0 896550.0 ;
      RECT  132000.0 895350.0 133200.0 896550.0 ;
      RECT  132000.0 895350.0 133200.0 896550.0 ;
      RECT  129600.0 895350.0 130800.0 896550.0 ;
      RECT  134400.0 904650.0 135600.0 905850.0 ;
      RECT  134400.0 894750.0 135600.0 895950.0 ;
      RECT  132000.0 897900.0 130800.0 899100.0 ;
      RECT  129000.0 900600.0 127800.0 901800.0 ;
      RECT  129600.0 904050.0 130800.0 905250.0 ;
      RECT  132000.0 895350.0 133200.0 896550.0 ;
      RECT  133200.0 900600.0 132000.0 901800.0 ;
      RECT  127800.0 900600.0 129000.0 901800.0 ;
      RECT  130800.0 897900.0 132000.0 899100.0 ;
      RECT  132000.0 900600.0 133200.0 901800.0 ;
      RECT  125400.0 906750.0 139800.0 907650.0 ;
      RECT  125400.0 892950.0 139800.0 893850.0 ;
      RECT  146400.0 905250.0 147600.0 907200.0 ;
      RECT  146400.0 893400.0 147600.0 895350.0 ;
      RECT  141600.0 894750.0 142800.0 892950.0 ;
      RECT  141600.0 904050.0 142800.0 907650.0 ;
      RECT  144300.0 894750.0 145200.0 904050.0 ;
      RECT  141600.0 904050.0 142800.0 905250.0 ;
      RECT  144000.0 904050.0 145200.0 905250.0 ;
      RECT  144000.0 904050.0 145200.0 905250.0 ;
      RECT  141600.0 904050.0 142800.0 905250.0 ;
      RECT  141600.0 894750.0 142800.0 895950.0 ;
      RECT  144000.0 894750.0 145200.0 895950.0 ;
      RECT  144000.0 894750.0 145200.0 895950.0 ;
      RECT  141600.0 894750.0 142800.0 895950.0 ;
      RECT  146400.0 904650.0 147600.0 905850.0 ;
      RECT  146400.0 894750.0 147600.0 895950.0 ;
      RECT  142200.0 899400.0 143400.0 900600.0 ;
      RECT  142200.0 899400.0 143400.0 900600.0 ;
      RECT  144750.0 899550.0 145650.0 900450.0 ;
      RECT  139800.0 906750.0 149400.0 907650.0 ;
      RECT  139800.0 892950.0 149400.0 893850.0 ;
      RECT  112050.0 899400.0 113250.0 900600.0 ;
      RECT  114000.0 897000.0 115200.0 898200.0 ;
      RECT  130800.0 897900.0 129600.0 899100.0 ;
      RECT  122400.0 909150.0 123600.0 907200.0 ;
      RECT  122400.0 921000.0 123600.0 919050.0 ;
      RECT  117600.0 919650.0 118800.0 921450.0 ;
      RECT  117600.0 910350.0 118800.0 906750.0 ;
      RECT  120300.0 919650.0 121200.0 910350.0 ;
      RECT  117600.0 910350.0 118800.0 909150.0 ;
      RECT  120000.0 910350.0 121200.0 909150.0 ;
      RECT  120000.0 910350.0 121200.0 909150.0 ;
      RECT  117600.0 910350.0 118800.0 909150.0 ;
      RECT  117600.0 919650.0 118800.0 918450.0 ;
      RECT  120000.0 919650.0 121200.0 918450.0 ;
      RECT  120000.0 919650.0 121200.0 918450.0 ;
      RECT  117600.0 919650.0 118800.0 918450.0 ;
      RECT  122400.0 909750.0 123600.0 908550.0 ;
      RECT  122400.0 919650.0 123600.0 918450.0 ;
      RECT  118200.0 915000.0 119400.0 913800.0 ;
      RECT  118200.0 915000.0 119400.0 913800.0 ;
      RECT  120750.0 914850.0 121650.0 913950.0 ;
      RECT  115800.0 907650.0 125400.0 906750.0 ;
      RECT  115800.0 921450.0 125400.0 920550.0 ;
      RECT  127200.0 919050.0 128400.0 921450.0 ;
      RECT  127200.0 910350.0 128400.0 906750.0 ;
      RECT  132000.0 910350.0 133200.0 906750.0 ;
      RECT  134400.0 909150.0 135600.0 907200.0 ;
      RECT  134400.0 921000.0 135600.0 919050.0 ;
      RECT  127200.0 910350.0 128400.0 909150.0 ;
      RECT  129600.0 910350.0 130800.0 909150.0 ;
      RECT  129600.0 910350.0 130800.0 909150.0 ;
      RECT  127200.0 910350.0 128400.0 909150.0 ;
      RECT  129600.0 910350.0 130800.0 909150.0 ;
      RECT  132000.0 910350.0 133200.0 909150.0 ;
      RECT  132000.0 910350.0 133200.0 909150.0 ;
      RECT  129600.0 910350.0 130800.0 909150.0 ;
      RECT  127200.0 919050.0 128400.0 917850.0 ;
      RECT  129600.0 919050.0 130800.0 917850.0 ;
      RECT  129600.0 919050.0 130800.0 917850.0 ;
      RECT  127200.0 919050.0 128400.0 917850.0 ;
      RECT  129600.0 919050.0 130800.0 917850.0 ;
      RECT  132000.0 919050.0 133200.0 917850.0 ;
      RECT  132000.0 919050.0 133200.0 917850.0 ;
      RECT  129600.0 919050.0 130800.0 917850.0 ;
      RECT  134400.0 909750.0 135600.0 908550.0 ;
      RECT  134400.0 919650.0 135600.0 918450.0 ;
      RECT  132000.0 916500.0 130800.0 915300.0 ;
      RECT  129000.0 913800.0 127800.0 912600.0 ;
      RECT  129600.0 910350.0 130800.0 909150.0 ;
      RECT  132000.0 919050.0 133200.0 917850.0 ;
      RECT  133200.0 913800.0 132000.0 912600.0 ;
      RECT  127800.0 913800.0 129000.0 912600.0 ;
      RECT  130800.0 916500.0 132000.0 915300.0 ;
      RECT  132000.0 913800.0 133200.0 912600.0 ;
      RECT  125400.0 907650.0 139800.0 906750.0 ;
      RECT  125400.0 921450.0 139800.0 920550.0 ;
      RECT  146400.0 909150.0 147600.0 907200.0 ;
      RECT  146400.0 921000.0 147600.0 919050.0 ;
      RECT  141600.0 919650.0 142800.0 921450.0 ;
      RECT  141600.0 910350.0 142800.0 906750.0 ;
      RECT  144300.0 919650.0 145200.0 910350.0 ;
      RECT  141600.0 910350.0 142800.0 909150.0 ;
      RECT  144000.0 910350.0 145200.0 909150.0 ;
      RECT  144000.0 910350.0 145200.0 909150.0 ;
      RECT  141600.0 910350.0 142800.0 909150.0 ;
      RECT  141600.0 919650.0 142800.0 918450.0 ;
      RECT  144000.0 919650.0 145200.0 918450.0 ;
      RECT  144000.0 919650.0 145200.0 918450.0 ;
      RECT  141600.0 919650.0 142800.0 918450.0 ;
      RECT  146400.0 909750.0 147600.0 908550.0 ;
      RECT  146400.0 919650.0 147600.0 918450.0 ;
      RECT  142200.0 915000.0 143400.0 913800.0 ;
      RECT  142200.0 915000.0 143400.0 913800.0 ;
      RECT  144750.0 914850.0 145650.0 913950.0 ;
      RECT  139800.0 907650.0 149400.0 906750.0 ;
      RECT  139800.0 921450.0 149400.0 920550.0 ;
      RECT  112050.0 913800.0 113250.0 915000.0 ;
      RECT  114000.0 916200.0 115200.0 917400.0 ;
      RECT  130800.0 915300.0 129600.0 916500.0 ;
      RECT  122400.0 932850.0 123600.0 934800.0 ;
      RECT  122400.0 921000.0 123600.0 922950.0 ;
      RECT  117600.0 922350.0 118800.0 920550.0 ;
      RECT  117600.0 931650.0 118800.0 935250.0 ;
      RECT  120300.0 922350.0 121200.0 931650.0 ;
      RECT  117600.0 931650.0 118800.0 932850.0 ;
      RECT  120000.0 931650.0 121200.0 932850.0 ;
      RECT  120000.0 931650.0 121200.0 932850.0 ;
      RECT  117600.0 931650.0 118800.0 932850.0 ;
      RECT  117600.0 922350.0 118800.0 923550.0 ;
      RECT  120000.0 922350.0 121200.0 923550.0 ;
      RECT  120000.0 922350.0 121200.0 923550.0 ;
      RECT  117600.0 922350.0 118800.0 923550.0 ;
      RECT  122400.0 932250.0 123600.0 933450.0 ;
      RECT  122400.0 922350.0 123600.0 923550.0 ;
      RECT  118200.0 927000.0 119400.0 928200.0 ;
      RECT  118200.0 927000.0 119400.0 928200.0 ;
      RECT  120750.0 927150.0 121650.0 928050.0 ;
      RECT  115800.0 934350.0 125400.0 935250.0 ;
      RECT  115800.0 920550.0 125400.0 921450.0 ;
      RECT  127200.0 922950.0 128400.0 920550.0 ;
      RECT  127200.0 931650.0 128400.0 935250.0 ;
      RECT  132000.0 931650.0 133200.0 935250.0 ;
      RECT  134400.0 932850.0 135600.0 934800.0 ;
      RECT  134400.0 921000.0 135600.0 922950.0 ;
      RECT  127200.0 931650.0 128400.0 932850.0 ;
      RECT  129600.0 931650.0 130800.0 932850.0 ;
      RECT  129600.0 931650.0 130800.0 932850.0 ;
      RECT  127200.0 931650.0 128400.0 932850.0 ;
      RECT  129600.0 931650.0 130800.0 932850.0 ;
      RECT  132000.0 931650.0 133200.0 932850.0 ;
      RECT  132000.0 931650.0 133200.0 932850.0 ;
      RECT  129600.0 931650.0 130800.0 932850.0 ;
      RECT  127200.0 922950.0 128400.0 924150.0 ;
      RECT  129600.0 922950.0 130800.0 924150.0 ;
      RECT  129600.0 922950.0 130800.0 924150.0 ;
      RECT  127200.0 922950.0 128400.0 924150.0 ;
      RECT  129600.0 922950.0 130800.0 924150.0 ;
      RECT  132000.0 922950.0 133200.0 924150.0 ;
      RECT  132000.0 922950.0 133200.0 924150.0 ;
      RECT  129600.0 922950.0 130800.0 924150.0 ;
      RECT  134400.0 932250.0 135600.0 933450.0 ;
      RECT  134400.0 922350.0 135600.0 923550.0 ;
      RECT  132000.0 925500.0 130800.0 926700.0 ;
      RECT  129000.0 928200.0 127800.0 929400.0 ;
      RECT  129600.0 931650.0 130800.0 932850.0 ;
      RECT  132000.0 922950.0 133200.0 924150.0 ;
      RECT  133200.0 928200.0 132000.0 929400.0 ;
      RECT  127800.0 928200.0 129000.0 929400.0 ;
      RECT  130800.0 925500.0 132000.0 926700.0 ;
      RECT  132000.0 928200.0 133200.0 929400.0 ;
      RECT  125400.0 934350.0 139800.0 935250.0 ;
      RECT  125400.0 920550.0 139800.0 921450.0 ;
      RECT  146400.0 932850.0 147600.0 934800.0 ;
      RECT  146400.0 921000.0 147600.0 922950.0 ;
      RECT  141600.0 922350.0 142800.0 920550.0 ;
      RECT  141600.0 931650.0 142800.0 935250.0 ;
      RECT  144300.0 922350.0 145200.0 931650.0 ;
      RECT  141600.0 931650.0 142800.0 932850.0 ;
      RECT  144000.0 931650.0 145200.0 932850.0 ;
      RECT  144000.0 931650.0 145200.0 932850.0 ;
      RECT  141600.0 931650.0 142800.0 932850.0 ;
      RECT  141600.0 922350.0 142800.0 923550.0 ;
      RECT  144000.0 922350.0 145200.0 923550.0 ;
      RECT  144000.0 922350.0 145200.0 923550.0 ;
      RECT  141600.0 922350.0 142800.0 923550.0 ;
      RECT  146400.0 932250.0 147600.0 933450.0 ;
      RECT  146400.0 922350.0 147600.0 923550.0 ;
      RECT  142200.0 927000.0 143400.0 928200.0 ;
      RECT  142200.0 927000.0 143400.0 928200.0 ;
      RECT  144750.0 927150.0 145650.0 928050.0 ;
      RECT  139800.0 934350.0 149400.0 935250.0 ;
      RECT  139800.0 920550.0 149400.0 921450.0 ;
      RECT  112050.0 927000.0 113250.0 928200.0 ;
      RECT  114000.0 924600.0 115200.0 925800.0 ;
      RECT  130800.0 925500.0 129600.0 926700.0 ;
      RECT  122400.0 936750.0 123600.0 934800.0 ;
      RECT  122400.0 948600.0 123600.0 946650.0 ;
      RECT  117600.0 947250.0 118800.0 949050.0 ;
      RECT  117600.0 937950.0 118800.0 934350.0 ;
      RECT  120300.0 947250.0 121200.0 937950.0 ;
      RECT  117600.0 937950.0 118800.0 936750.0 ;
      RECT  120000.0 937950.0 121200.0 936750.0 ;
      RECT  120000.0 937950.0 121200.0 936750.0 ;
      RECT  117600.0 937950.0 118800.0 936750.0 ;
      RECT  117600.0 947250.0 118800.0 946050.0 ;
      RECT  120000.0 947250.0 121200.0 946050.0 ;
      RECT  120000.0 947250.0 121200.0 946050.0 ;
      RECT  117600.0 947250.0 118800.0 946050.0 ;
      RECT  122400.0 937350.0 123600.0 936150.0 ;
      RECT  122400.0 947250.0 123600.0 946050.0 ;
      RECT  118200.0 942600.0 119400.0 941400.0 ;
      RECT  118200.0 942600.0 119400.0 941400.0 ;
      RECT  120750.0 942450.0 121650.0 941550.0 ;
      RECT  115800.0 935250.0 125400.0 934350.0 ;
      RECT  115800.0 949050.0 125400.0 948150.0 ;
      RECT  127200.0 946650.0 128400.0 949050.0 ;
      RECT  127200.0 937950.0 128400.0 934350.0 ;
      RECT  132000.0 937950.0 133200.0 934350.0 ;
      RECT  134400.0 936750.0 135600.0 934800.0 ;
      RECT  134400.0 948600.0 135600.0 946650.0 ;
      RECT  127200.0 937950.0 128400.0 936750.0 ;
      RECT  129600.0 937950.0 130800.0 936750.0 ;
      RECT  129600.0 937950.0 130800.0 936750.0 ;
      RECT  127200.0 937950.0 128400.0 936750.0 ;
      RECT  129600.0 937950.0 130800.0 936750.0 ;
      RECT  132000.0 937950.0 133200.0 936750.0 ;
      RECT  132000.0 937950.0 133200.0 936750.0 ;
      RECT  129600.0 937950.0 130800.0 936750.0 ;
      RECT  127200.0 946650.0 128400.0 945450.0 ;
      RECT  129600.0 946650.0 130800.0 945450.0 ;
      RECT  129600.0 946650.0 130800.0 945450.0 ;
      RECT  127200.0 946650.0 128400.0 945450.0 ;
      RECT  129600.0 946650.0 130800.0 945450.0 ;
      RECT  132000.0 946650.0 133200.0 945450.0 ;
      RECT  132000.0 946650.0 133200.0 945450.0 ;
      RECT  129600.0 946650.0 130800.0 945450.0 ;
      RECT  134400.0 937350.0 135600.0 936150.0 ;
      RECT  134400.0 947250.0 135600.0 946050.0 ;
      RECT  132000.0 944100.0 130800.0 942900.0 ;
      RECT  129000.0 941400.0 127800.0 940200.0 ;
      RECT  129600.0 937950.0 130800.0 936750.0 ;
      RECT  132000.0 946650.0 133200.0 945450.0 ;
      RECT  133200.0 941400.0 132000.0 940200.0 ;
      RECT  127800.0 941400.0 129000.0 940200.0 ;
      RECT  130800.0 944100.0 132000.0 942900.0 ;
      RECT  132000.0 941400.0 133200.0 940200.0 ;
      RECT  125400.0 935250.0 139800.0 934350.0 ;
      RECT  125400.0 949050.0 139800.0 948150.0 ;
      RECT  146400.0 936750.0 147600.0 934800.0 ;
      RECT  146400.0 948600.0 147600.0 946650.0 ;
      RECT  141600.0 947250.0 142800.0 949050.0 ;
      RECT  141600.0 937950.0 142800.0 934350.0 ;
      RECT  144300.0 947250.0 145200.0 937950.0 ;
      RECT  141600.0 937950.0 142800.0 936750.0 ;
      RECT  144000.0 937950.0 145200.0 936750.0 ;
      RECT  144000.0 937950.0 145200.0 936750.0 ;
      RECT  141600.0 937950.0 142800.0 936750.0 ;
      RECT  141600.0 947250.0 142800.0 946050.0 ;
      RECT  144000.0 947250.0 145200.0 946050.0 ;
      RECT  144000.0 947250.0 145200.0 946050.0 ;
      RECT  141600.0 947250.0 142800.0 946050.0 ;
      RECT  146400.0 937350.0 147600.0 936150.0 ;
      RECT  146400.0 947250.0 147600.0 946050.0 ;
      RECT  142200.0 942600.0 143400.0 941400.0 ;
      RECT  142200.0 942600.0 143400.0 941400.0 ;
      RECT  144750.0 942450.0 145650.0 941550.0 ;
      RECT  139800.0 935250.0 149400.0 934350.0 ;
      RECT  139800.0 949050.0 149400.0 948150.0 ;
      RECT  112050.0 941400.0 113250.0 942600.0 ;
      RECT  114000.0 943800.0 115200.0 945000.0 ;
      RECT  130800.0 942900.0 129600.0 944100.0 ;
      RECT  122400.0 960450.0 123600.0 962400.0 ;
      RECT  122400.0 948600.0 123600.0 950550.0 ;
      RECT  117600.0 949950.0 118800.0 948150.0 ;
      RECT  117600.0 959250.0 118800.0 962850.0 ;
      RECT  120300.0 949950.0 121200.0 959250.0 ;
      RECT  117600.0 959250.0 118800.0 960450.0 ;
      RECT  120000.0 959250.0 121200.0 960450.0 ;
      RECT  120000.0 959250.0 121200.0 960450.0 ;
      RECT  117600.0 959250.0 118800.0 960450.0 ;
      RECT  117600.0 949950.0 118800.0 951150.0 ;
      RECT  120000.0 949950.0 121200.0 951150.0 ;
      RECT  120000.0 949950.0 121200.0 951150.0 ;
      RECT  117600.0 949950.0 118800.0 951150.0 ;
      RECT  122400.0 959850.0 123600.0 961050.0 ;
      RECT  122400.0 949950.0 123600.0 951150.0 ;
      RECT  118200.0 954600.0 119400.0 955800.0 ;
      RECT  118200.0 954600.0 119400.0 955800.0 ;
      RECT  120750.0 954750.0 121650.0 955650.0 ;
      RECT  115800.0 961950.0 125400.0 962850.0 ;
      RECT  115800.0 948150.0 125400.0 949050.0 ;
      RECT  127200.0 950550.0 128400.0 948150.0 ;
      RECT  127200.0 959250.0 128400.0 962850.0 ;
      RECT  132000.0 959250.0 133200.0 962850.0 ;
      RECT  134400.0 960450.0 135600.0 962400.0 ;
      RECT  134400.0 948600.0 135600.0 950550.0 ;
      RECT  127200.0 959250.0 128400.0 960450.0 ;
      RECT  129600.0 959250.0 130800.0 960450.0 ;
      RECT  129600.0 959250.0 130800.0 960450.0 ;
      RECT  127200.0 959250.0 128400.0 960450.0 ;
      RECT  129600.0 959250.0 130800.0 960450.0 ;
      RECT  132000.0 959250.0 133200.0 960450.0 ;
      RECT  132000.0 959250.0 133200.0 960450.0 ;
      RECT  129600.0 959250.0 130800.0 960450.0 ;
      RECT  127200.0 950550.0 128400.0 951750.0 ;
      RECT  129600.0 950550.0 130800.0 951750.0 ;
      RECT  129600.0 950550.0 130800.0 951750.0 ;
      RECT  127200.0 950550.0 128400.0 951750.0 ;
      RECT  129600.0 950550.0 130800.0 951750.0 ;
      RECT  132000.0 950550.0 133200.0 951750.0 ;
      RECT  132000.0 950550.0 133200.0 951750.0 ;
      RECT  129600.0 950550.0 130800.0 951750.0 ;
      RECT  134400.0 959850.0 135600.0 961050.0 ;
      RECT  134400.0 949950.0 135600.0 951150.0 ;
      RECT  132000.0 953100.0 130800.0 954300.0 ;
      RECT  129000.0 955800.0 127800.0 957000.0 ;
      RECT  129600.0 959250.0 130800.0 960450.0 ;
      RECT  132000.0 950550.0 133200.0 951750.0 ;
      RECT  133200.0 955800.0 132000.0 957000.0 ;
      RECT  127800.0 955800.0 129000.0 957000.0 ;
      RECT  130800.0 953100.0 132000.0 954300.0 ;
      RECT  132000.0 955800.0 133200.0 957000.0 ;
      RECT  125400.0 961950.0 139800.0 962850.0 ;
      RECT  125400.0 948150.0 139800.0 949050.0 ;
      RECT  146400.0 960450.0 147600.0 962400.0 ;
      RECT  146400.0 948600.0 147600.0 950550.0 ;
      RECT  141600.0 949950.0 142800.0 948150.0 ;
      RECT  141600.0 959250.0 142800.0 962850.0 ;
      RECT  144300.0 949950.0 145200.0 959250.0 ;
      RECT  141600.0 959250.0 142800.0 960450.0 ;
      RECT  144000.0 959250.0 145200.0 960450.0 ;
      RECT  144000.0 959250.0 145200.0 960450.0 ;
      RECT  141600.0 959250.0 142800.0 960450.0 ;
      RECT  141600.0 949950.0 142800.0 951150.0 ;
      RECT  144000.0 949950.0 145200.0 951150.0 ;
      RECT  144000.0 949950.0 145200.0 951150.0 ;
      RECT  141600.0 949950.0 142800.0 951150.0 ;
      RECT  146400.0 959850.0 147600.0 961050.0 ;
      RECT  146400.0 949950.0 147600.0 951150.0 ;
      RECT  142200.0 954600.0 143400.0 955800.0 ;
      RECT  142200.0 954600.0 143400.0 955800.0 ;
      RECT  144750.0 954750.0 145650.0 955650.0 ;
      RECT  139800.0 961950.0 149400.0 962850.0 ;
      RECT  139800.0 948150.0 149400.0 949050.0 ;
      RECT  112050.0 954600.0 113250.0 955800.0 ;
      RECT  114000.0 952200.0 115200.0 953400.0 ;
      RECT  130800.0 953100.0 129600.0 954300.0 ;
      RECT  122400.0 964350.0 123600.0 962400.0 ;
      RECT  122400.0 976200.0 123600.0 974250.0 ;
      RECT  117600.0 974850.0 118800.0 976650.0 ;
      RECT  117600.0 965550.0 118800.0 961950.0 ;
      RECT  120300.0 974850.0 121200.0 965550.0 ;
      RECT  117600.0 965550.0 118800.0 964350.0 ;
      RECT  120000.0 965550.0 121200.0 964350.0 ;
      RECT  120000.0 965550.0 121200.0 964350.0 ;
      RECT  117600.0 965550.0 118800.0 964350.0 ;
      RECT  117600.0 974850.0 118800.0 973650.0 ;
      RECT  120000.0 974850.0 121200.0 973650.0 ;
      RECT  120000.0 974850.0 121200.0 973650.0 ;
      RECT  117600.0 974850.0 118800.0 973650.0 ;
      RECT  122400.0 964950.0 123600.0 963750.0 ;
      RECT  122400.0 974850.0 123600.0 973650.0 ;
      RECT  118200.0 970200.0 119400.0 969000.0 ;
      RECT  118200.0 970200.0 119400.0 969000.0 ;
      RECT  120750.0 970050.0 121650.0 969150.0 ;
      RECT  115800.0 962850.0 125400.0 961950.0 ;
      RECT  115800.0 976650.0 125400.0 975750.0 ;
      RECT  127200.0 974250.0 128400.0 976650.0 ;
      RECT  127200.0 965550.0 128400.0 961950.0 ;
      RECT  132000.0 965550.0 133200.0 961950.0 ;
      RECT  134400.0 964350.0 135600.0 962400.0 ;
      RECT  134400.0 976200.0 135600.0 974250.0 ;
      RECT  127200.0 965550.0 128400.0 964350.0 ;
      RECT  129600.0 965550.0 130800.0 964350.0 ;
      RECT  129600.0 965550.0 130800.0 964350.0 ;
      RECT  127200.0 965550.0 128400.0 964350.0 ;
      RECT  129600.0 965550.0 130800.0 964350.0 ;
      RECT  132000.0 965550.0 133200.0 964350.0 ;
      RECT  132000.0 965550.0 133200.0 964350.0 ;
      RECT  129600.0 965550.0 130800.0 964350.0 ;
      RECT  127200.0 974250.0 128400.0 973050.0 ;
      RECT  129600.0 974250.0 130800.0 973050.0 ;
      RECT  129600.0 974250.0 130800.0 973050.0 ;
      RECT  127200.0 974250.0 128400.0 973050.0 ;
      RECT  129600.0 974250.0 130800.0 973050.0 ;
      RECT  132000.0 974250.0 133200.0 973050.0 ;
      RECT  132000.0 974250.0 133200.0 973050.0 ;
      RECT  129600.0 974250.0 130800.0 973050.0 ;
      RECT  134400.0 964950.0 135600.0 963750.0 ;
      RECT  134400.0 974850.0 135600.0 973650.0 ;
      RECT  132000.0 971700.0 130800.0 970500.0 ;
      RECT  129000.0 969000.0 127800.0 967800.0 ;
      RECT  129600.0 965550.0 130800.0 964350.0 ;
      RECT  132000.0 974250.0 133200.0 973050.0 ;
      RECT  133200.0 969000.0 132000.0 967800.0 ;
      RECT  127800.0 969000.0 129000.0 967800.0 ;
      RECT  130800.0 971700.0 132000.0 970500.0 ;
      RECT  132000.0 969000.0 133200.0 967800.0 ;
      RECT  125400.0 962850.0 139800.0 961950.0 ;
      RECT  125400.0 976650.0 139800.0 975750.0 ;
      RECT  146400.0 964350.0 147600.0 962400.0 ;
      RECT  146400.0 976200.0 147600.0 974250.0 ;
      RECT  141600.0 974850.0 142800.0 976650.0 ;
      RECT  141600.0 965550.0 142800.0 961950.0 ;
      RECT  144300.0 974850.0 145200.0 965550.0 ;
      RECT  141600.0 965550.0 142800.0 964350.0 ;
      RECT  144000.0 965550.0 145200.0 964350.0 ;
      RECT  144000.0 965550.0 145200.0 964350.0 ;
      RECT  141600.0 965550.0 142800.0 964350.0 ;
      RECT  141600.0 974850.0 142800.0 973650.0 ;
      RECT  144000.0 974850.0 145200.0 973650.0 ;
      RECT  144000.0 974850.0 145200.0 973650.0 ;
      RECT  141600.0 974850.0 142800.0 973650.0 ;
      RECT  146400.0 964950.0 147600.0 963750.0 ;
      RECT  146400.0 974850.0 147600.0 973650.0 ;
      RECT  142200.0 970200.0 143400.0 969000.0 ;
      RECT  142200.0 970200.0 143400.0 969000.0 ;
      RECT  144750.0 970050.0 145650.0 969150.0 ;
      RECT  139800.0 962850.0 149400.0 961950.0 ;
      RECT  139800.0 976650.0 149400.0 975750.0 ;
      RECT  112050.0 969000.0 113250.0 970200.0 ;
      RECT  114000.0 971400.0 115200.0 972600.0 ;
      RECT  130800.0 970500.0 129600.0 971700.0 ;
      RECT  122400.0 988050.0 123600.0 990000.0 ;
      RECT  122400.0 976200.0 123600.0 978150.0 ;
      RECT  117600.0 977550.0 118800.0 975750.0 ;
      RECT  117600.0 986850.0 118800.0 990450.0 ;
      RECT  120300.0 977550.0 121200.0 986850.0 ;
      RECT  117600.0 986850.0 118800.0 988050.0 ;
      RECT  120000.0 986850.0 121200.0 988050.0 ;
      RECT  120000.0 986850.0 121200.0 988050.0 ;
      RECT  117600.0 986850.0 118800.0 988050.0 ;
      RECT  117600.0 977550.0 118800.0 978750.0 ;
      RECT  120000.0 977550.0 121200.0 978750.0 ;
      RECT  120000.0 977550.0 121200.0 978750.0 ;
      RECT  117600.0 977550.0 118800.0 978750.0 ;
      RECT  122400.0 987450.0 123600.0 988650.0 ;
      RECT  122400.0 977550.0 123600.0 978750.0 ;
      RECT  118200.0 982200.0 119400.0 983400.0 ;
      RECT  118200.0 982200.0 119400.0 983400.0 ;
      RECT  120750.0 982350.0 121650.0 983250.0 ;
      RECT  115800.0 989550.0 125400.0 990450.0 ;
      RECT  115800.0 975750.0 125400.0 976650.0 ;
      RECT  127200.0 978150.0 128400.0 975750.0 ;
      RECT  127200.0 986850.0 128400.0 990450.0 ;
      RECT  132000.0 986850.0 133200.0 990450.0 ;
      RECT  134400.0 988050.0 135600.0 990000.0 ;
      RECT  134400.0 976200.0 135600.0 978150.0 ;
      RECT  127200.0 986850.0 128400.0 988050.0 ;
      RECT  129600.0 986850.0 130800.0 988050.0 ;
      RECT  129600.0 986850.0 130800.0 988050.0 ;
      RECT  127200.0 986850.0 128400.0 988050.0 ;
      RECT  129600.0 986850.0 130800.0 988050.0 ;
      RECT  132000.0 986850.0 133200.0 988050.0 ;
      RECT  132000.0 986850.0 133200.0 988050.0 ;
      RECT  129600.0 986850.0 130800.0 988050.0 ;
      RECT  127200.0 978150.0 128400.0 979350.0 ;
      RECT  129600.0 978150.0 130800.0 979350.0 ;
      RECT  129600.0 978150.0 130800.0 979350.0 ;
      RECT  127200.0 978150.0 128400.0 979350.0 ;
      RECT  129600.0 978150.0 130800.0 979350.0 ;
      RECT  132000.0 978150.0 133200.0 979350.0 ;
      RECT  132000.0 978150.0 133200.0 979350.0 ;
      RECT  129600.0 978150.0 130800.0 979350.0 ;
      RECT  134400.0 987450.0 135600.0 988650.0 ;
      RECT  134400.0 977550.0 135600.0 978750.0 ;
      RECT  132000.0 980700.0 130800.0 981900.0 ;
      RECT  129000.0 983400.0 127800.0 984600.0 ;
      RECT  129600.0 986850.0 130800.0 988050.0 ;
      RECT  132000.0 978150.0 133200.0 979350.0 ;
      RECT  133200.0 983400.0 132000.0 984600.0 ;
      RECT  127800.0 983400.0 129000.0 984600.0 ;
      RECT  130800.0 980700.0 132000.0 981900.0 ;
      RECT  132000.0 983400.0 133200.0 984600.0 ;
      RECT  125400.0 989550.0 139800.0 990450.0 ;
      RECT  125400.0 975750.0 139800.0 976650.0 ;
      RECT  146400.0 988050.0 147600.0 990000.0 ;
      RECT  146400.0 976200.0 147600.0 978150.0 ;
      RECT  141600.0 977550.0 142800.0 975750.0 ;
      RECT  141600.0 986850.0 142800.0 990450.0 ;
      RECT  144300.0 977550.0 145200.0 986850.0 ;
      RECT  141600.0 986850.0 142800.0 988050.0 ;
      RECT  144000.0 986850.0 145200.0 988050.0 ;
      RECT  144000.0 986850.0 145200.0 988050.0 ;
      RECT  141600.0 986850.0 142800.0 988050.0 ;
      RECT  141600.0 977550.0 142800.0 978750.0 ;
      RECT  144000.0 977550.0 145200.0 978750.0 ;
      RECT  144000.0 977550.0 145200.0 978750.0 ;
      RECT  141600.0 977550.0 142800.0 978750.0 ;
      RECT  146400.0 987450.0 147600.0 988650.0 ;
      RECT  146400.0 977550.0 147600.0 978750.0 ;
      RECT  142200.0 982200.0 143400.0 983400.0 ;
      RECT  142200.0 982200.0 143400.0 983400.0 ;
      RECT  144750.0 982350.0 145650.0 983250.0 ;
      RECT  139800.0 989550.0 149400.0 990450.0 ;
      RECT  139800.0 975750.0 149400.0 976650.0 ;
      RECT  112050.0 982200.0 113250.0 983400.0 ;
      RECT  114000.0 979800.0 115200.0 981000.0 ;
      RECT  130800.0 980700.0 129600.0 981900.0 ;
      RECT  122400.0 991950.0 123600.0 990000.0 ;
      RECT  122400.0 1003800.0 123600.0 1001850.0 ;
      RECT  117600.0 1002450.0 118800.0 1004250.0 ;
      RECT  117600.0 993150.0 118800.0 989550.0 ;
      RECT  120300.0 1002450.0 121200.0 993150.0 ;
      RECT  117600.0 993150.0 118800.0 991950.0 ;
      RECT  120000.0 993150.0 121200.0 991950.0 ;
      RECT  120000.0 993150.0 121200.0 991950.0 ;
      RECT  117600.0 993150.0 118800.0 991950.0 ;
      RECT  117600.0 1002450.0 118800.0 1001250.0 ;
      RECT  120000.0 1002450.0 121200.0 1001250.0 ;
      RECT  120000.0 1002450.0 121200.0 1001250.0 ;
      RECT  117600.0 1002450.0 118800.0 1001250.0 ;
      RECT  122400.0 992550.0 123600.0 991350.0 ;
      RECT  122400.0 1002450.0 123600.0 1001250.0 ;
      RECT  118200.0 997800.0 119400.0 996600.0 ;
      RECT  118200.0 997800.0 119400.0 996600.0 ;
      RECT  120750.0 997650.0 121650.0 996750.0 ;
      RECT  115800.0 990450.0 125400.0 989550.0 ;
      RECT  115800.0 1004250.0 125400.0 1003350.0 ;
      RECT  127200.0 1001850.0 128400.0 1004250.0 ;
      RECT  127200.0 993150.0 128400.0 989550.0 ;
      RECT  132000.0 993150.0 133200.0 989550.0 ;
      RECT  134400.0 991950.0 135600.0 990000.0 ;
      RECT  134400.0 1003800.0 135600.0 1001850.0 ;
      RECT  127200.0 993150.0 128400.0 991950.0 ;
      RECT  129600.0 993150.0 130800.0 991950.0 ;
      RECT  129600.0 993150.0 130800.0 991950.0 ;
      RECT  127200.0 993150.0 128400.0 991950.0 ;
      RECT  129600.0 993150.0 130800.0 991950.0 ;
      RECT  132000.0 993150.0 133200.0 991950.0 ;
      RECT  132000.0 993150.0 133200.0 991950.0 ;
      RECT  129600.0 993150.0 130800.0 991950.0 ;
      RECT  127200.0 1001850.0 128400.0 1000650.0 ;
      RECT  129600.0 1001850.0 130800.0 1000650.0 ;
      RECT  129600.0 1001850.0 130800.0 1000650.0 ;
      RECT  127200.0 1001850.0 128400.0 1000650.0 ;
      RECT  129600.0 1001850.0 130800.0 1000650.0 ;
      RECT  132000.0 1001850.0 133200.0 1000650.0 ;
      RECT  132000.0 1001850.0 133200.0 1000650.0 ;
      RECT  129600.0 1001850.0 130800.0 1000650.0 ;
      RECT  134400.0 992550.0 135600.0 991350.0 ;
      RECT  134400.0 1002450.0 135600.0 1001250.0 ;
      RECT  132000.0 999300.0 130800.0 998100.0 ;
      RECT  129000.0 996600.0 127800.0 995400.0 ;
      RECT  129600.0 993150.0 130800.0 991950.0 ;
      RECT  132000.0 1001850.0 133200.0 1000650.0 ;
      RECT  133200.0 996600.0 132000.0 995400.0 ;
      RECT  127800.0 996600.0 129000.0 995400.0 ;
      RECT  130800.0 999300.0 132000.0 998100.0 ;
      RECT  132000.0 996600.0 133200.0 995400.0 ;
      RECT  125400.0 990450.0 139800.0 989550.0 ;
      RECT  125400.0 1004250.0 139800.0 1003350.0 ;
      RECT  146400.0 991950.0 147600.0 990000.0 ;
      RECT  146400.0 1003800.0 147600.0 1001850.0 ;
      RECT  141600.0 1002450.0 142800.0 1004250.0 ;
      RECT  141600.0 993150.0 142800.0 989550.0 ;
      RECT  144300.0 1002450.0 145200.0 993150.0 ;
      RECT  141600.0 993150.0 142800.0 991950.0 ;
      RECT  144000.0 993150.0 145200.0 991950.0 ;
      RECT  144000.0 993150.0 145200.0 991950.0 ;
      RECT  141600.0 993150.0 142800.0 991950.0 ;
      RECT  141600.0 1002450.0 142800.0 1001250.0 ;
      RECT  144000.0 1002450.0 145200.0 1001250.0 ;
      RECT  144000.0 1002450.0 145200.0 1001250.0 ;
      RECT  141600.0 1002450.0 142800.0 1001250.0 ;
      RECT  146400.0 992550.0 147600.0 991350.0 ;
      RECT  146400.0 1002450.0 147600.0 1001250.0 ;
      RECT  142200.0 997800.0 143400.0 996600.0 ;
      RECT  142200.0 997800.0 143400.0 996600.0 ;
      RECT  144750.0 997650.0 145650.0 996750.0 ;
      RECT  139800.0 990450.0 149400.0 989550.0 ;
      RECT  139800.0 1004250.0 149400.0 1003350.0 ;
      RECT  112050.0 996600.0 113250.0 997800.0 ;
      RECT  114000.0 999000.0 115200.0 1000200.0 ;
      RECT  130800.0 998100.0 129600.0 999300.0 ;
      RECT  122400.0 1015650.0 123600.0 1017600.0 ;
      RECT  122400.0 1003800.0 123600.0 1005750.0 ;
      RECT  117600.0 1005150.0 118800.0 1003350.0 ;
      RECT  117600.0 1014450.0 118800.0 1018050.0 ;
      RECT  120300.0 1005150.0 121200.0 1014450.0 ;
      RECT  117600.0 1014450.0 118800.0 1015650.0 ;
      RECT  120000.0 1014450.0 121200.0 1015650.0 ;
      RECT  120000.0 1014450.0 121200.0 1015650.0 ;
      RECT  117600.0 1014450.0 118800.0 1015650.0 ;
      RECT  117600.0 1005150.0 118800.0 1006350.0 ;
      RECT  120000.0 1005150.0 121200.0 1006350.0 ;
      RECT  120000.0 1005150.0 121200.0 1006350.0 ;
      RECT  117600.0 1005150.0 118800.0 1006350.0 ;
      RECT  122400.0 1015050.0 123600.0 1016250.0 ;
      RECT  122400.0 1005150.0 123600.0 1006350.0 ;
      RECT  118200.0 1009800.0 119400.0 1011000.0 ;
      RECT  118200.0 1009800.0 119400.0 1011000.0 ;
      RECT  120750.0 1009950.0 121650.0 1010850.0 ;
      RECT  115800.0 1017150.0 125400.0 1018050.0 ;
      RECT  115800.0 1003350.0 125400.0 1004250.0 ;
      RECT  127200.0 1005750.0 128400.0 1003350.0 ;
      RECT  127200.0 1014450.0 128400.0 1018050.0 ;
      RECT  132000.0 1014450.0 133200.0 1018050.0 ;
      RECT  134400.0 1015650.0 135600.0 1017600.0 ;
      RECT  134400.0 1003800.0 135600.0 1005750.0 ;
      RECT  127200.0 1014450.0 128400.0 1015650.0 ;
      RECT  129600.0 1014450.0 130800.0 1015650.0 ;
      RECT  129600.0 1014450.0 130800.0 1015650.0 ;
      RECT  127200.0 1014450.0 128400.0 1015650.0 ;
      RECT  129600.0 1014450.0 130800.0 1015650.0 ;
      RECT  132000.0 1014450.0 133200.0 1015650.0 ;
      RECT  132000.0 1014450.0 133200.0 1015650.0 ;
      RECT  129600.0 1014450.0 130800.0 1015650.0 ;
      RECT  127200.0 1005750.0 128400.0 1006950.0 ;
      RECT  129600.0 1005750.0 130800.0 1006950.0 ;
      RECT  129600.0 1005750.0 130800.0 1006950.0 ;
      RECT  127200.0 1005750.0 128400.0 1006950.0 ;
      RECT  129600.0 1005750.0 130800.0 1006950.0 ;
      RECT  132000.0 1005750.0 133200.0 1006950.0 ;
      RECT  132000.0 1005750.0 133200.0 1006950.0 ;
      RECT  129600.0 1005750.0 130800.0 1006950.0 ;
      RECT  134400.0 1015050.0 135600.0 1016250.0 ;
      RECT  134400.0 1005150.0 135600.0 1006350.0 ;
      RECT  132000.0 1008300.0 130800.0 1009500.0 ;
      RECT  129000.0 1011000.0 127800.0 1012200.0 ;
      RECT  129600.0 1014450.0 130800.0 1015650.0 ;
      RECT  132000.0 1005750.0 133200.0 1006950.0 ;
      RECT  133200.0 1011000.0 132000.0 1012200.0 ;
      RECT  127800.0 1011000.0 129000.0 1012200.0 ;
      RECT  130800.0 1008300.0 132000.0 1009500.0 ;
      RECT  132000.0 1011000.0 133200.0 1012200.0 ;
      RECT  125400.0 1017150.0 139800.0 1018050.0 ;
      RECT  125400.0 1003350.0 139800.0 1004250.0 ;
      RECT  146400.0 1015650.0 147600.0 1017600.0 ;
      RECT  146400.0 1003800.0 147600.0 1005750.0 ;
      RECT  141600.0 1005150.0 142800.0 1003350.0 ;
      RECT  141600.0 1014450.0 142800.0 1018050.0 ;
      RECT  144300.0 1005150.0 145200.0 1014450.0 ;
      RECT  141600.0 1014450.0 142800.0 1015650.0 ;
      RECT  144000.0 1014450.0 145200.0 1015650.0 ;
      RECT  144000.0 1014450.0 145200.0 1015650.0 ;
      RECT  141600.0 1014450.0 142800.0 1015650.0 ;
      RECT  141600.0 1005150.0 142800.0 1006350.0 ;
      RECT  144000.0 1005150.0 145200.0 1006350.0 ;
      RECT  144000.0 1005150.0 145200.0 1006350.0 ;
      RECT  141600.0 1005150.0 142800.0 1006350.0 ;
      RECT  146400.0 1015050.0 147600.0 1016250.0 ;
      RECT  146400.0 1005150.0 147600.0 1006350.0 ;
      RECT  142200.0 1009800.0 143400.0 1011000.0 ;
      RECT  142200.0 1009800.0 143400.0 1011000.0 ;
      RECT  144750.0 1009950.0 145650.0 1010850.0 ;
      RECT  139800.0 1017150.0 149400.0 1018050.0 ;
      RECT  139800.0 1003350.0 149400.0 1004250.0 ;
      RECT  112050.0 1009800.0 113250.0 1011000.0 ;
      RECT  114000.0 1007400.0 115200.0 1008600.0 ;
      RECT  130800.0 1008300.0 129600.0 1009500.0 ;
      RECT  122400.0 1019550.0 123600.0 1017600.0 ;
      RECT  122400.0 1031400.0 123600.0 1029450.0 ;
      RECT  117600.0 1030050.0 118800.0 1031850.0 ;
      RECT  117600.0 1020750.0 118800.0 1017150.0 ;
      RECT  120300.0 1030050.0 121200.0 1020750.0 ;
      RECT  117600.0 1020750.0 118800.0 1019550.0 ;
      RECT  120000.0 1020750.0 121200.0 1019550.0 ;
      RECT  120000.0 1020750.0 121200.0 1019550.0 ;
      RECT  117600.0 1020750.0 118800.0 1019550.0 ;
      RECT  117600.0 1030050.0 118800.0 1028850.0 ;
      RECT  120000.0 1030050.0 121200.0 1028850.0 ;
      RECT  120000.0 1030050.0 121200.0 1028850.0 ;
      RECT  117600.0 1030050.0 118800.0 1028850.0 ;
      RECT  122400.0 1020150.0 123600.0 1018950.0 ;
      RECT  122400.0 1030050.0 123600.0 1028850.0 ;
      RECT  118200.0 1025400.0 119400.0 1024200.0 ;
      RECT  118200.0 1025400.0 119400.0 1024200.0 ;
      RECT  120750.0 1025250.0 121650.0 1024350.0 ;
      RECT  115800.0 1018050.0 125400.0 1017150.0 ;
      RECT  115800.0 1031850.0 125400.0 1030950.0 ;
      RECT  127200.0 1029450.0 128400.0 1031850.0 ;
      RECT  127200.0 1020750.0 128400.0 1017150.0 ;
      RECT  132000.0 1020750.0 133200.0 1017150.0 ;
      RECT  134400.0 1019550.0 135600.0 1017600.0 ;
      RECT  134400.0 1031400.0 135600.0 1029450.0 ;
      RECT  127200.0 1020750.0 128400.0 1019550.0 ;
      RECT  129600.0 1020750.0 130800.0 1019550.0 ;
      RECT  129600.0 1020750.0 130800.0 1019550.0 ;
      RECT  127200.0 1020750.0 128400.0 1019550.0 ;
      RECT  129600.0 1020750.0 130800.0 1019550.0 ;
      RECT  132000.0 1020750.0 133200.0 1019550.0 ;
      RECT  132000.0 1020750.0 133200.0 1019550.0 ;
      RECT  129600.0 1020750.0 130800.0 1019550.0 ;
      RECT  127200.0 1029450.0 128400.0 1028250.0 ;
      RECT  129600.0 1029450.0 130800.0 1028250.0 ;
      RECT  129600.0 1029450.0 130800.0 1028250.0 ;
      RECT  127200.0 1029450.0 128400.0 1028250.0 ;
      RECT  129600.0 1029450.0 130800.0 1028250.0 ;
      RECT  132000.0 1029450.0 133200.0 1028250.0 ;
      RECT  132000.0 1029450.0 133200.0 1028250.0 ;
      RECT  129600.0 1029450.0 130800.0 1028250.0 ;
      RECT  134400.0 1020150.0 135600.0 1018950.0 ;
      RECT  134400.0 1030050.0 135600.0 1028850.0 ;
      RECT  132000.0 1026900.0 130800.0 1025700.0 ;
      RECT  129000.0 1024200.0 127800.0 1023000.0 ;
      RECT  129600.0 1020750.0 130800.0 1019550.0 ;
      RECT  132000.0 1029450.0 133200.0 1028250.0 ;
      RECT  133200.0 1024200.0 132000.0 1023000.0 ;
      RECT  127800.0 1024200.0 129000.0 1023000.0 ;
      RECT  130800.0 1026900.0 132000.0 1025700.0 ;
      RECT  132000.0 1024200.0 133200.0 1023000.0 ;
      RECT  125400.0 1018050.0 139800.0 1017150.0 ;
      RECT  125400.0 1031850.0 139800.0 1030950.0 ;
      RECT  146400.0 1019550.0 147600.0 1017600.0 ;
      RECT  146400.0 1031400.0 147600.0 1029450.0 ;
      RECT  141600.0 1030050.0 142800.0 1031850.0 ;
      RECT  141600.0 1020750.0 142800.0 1017150.0 ;
      RECT  144300.0 1030050.0 145200.0 1020750.0 ;
      RECT  141600.0 1020750.0 142800.0 1019550.0 ;
      RECT  144000.0 1020750.0 145200.0 1019550.0 ;
      RECT  144000.0 1020750.0 145200.0 1019550.0 ;
      RECT  141600.0 1020750.0 142800.0 1019550.0 ;
      RECT  141600.0 1030050.0 142800.0 1028850.0 ;
      RECT  144000.0 1030050.0 145200.0 1028850.0 ;
      RECT  144000.0 1030050.0 145200.0 1028850.0 ;
      RECT  141600.0 1030050.0 142800.0 1028850.0 ;
      RECT  146400.0 1020150.0 147600.0 1018950.0 ;
      RECT  146400.0 1030050.0 147600.0 1028850.0 ;
      RECT  142200.0 1025400.0 143400.0 1024200.0 ;
      RECT  142200.0 1025400.0 143400.0 1024200.0 ;
      RECT  144750.0 1025250.0 145650.0 1024350.0 ;
      RECT  139800.0 1018050.0 149400.0 1017150.0 ;
      RECT  139800.0 1031850.0 149400.0 1030950.0 ;
      RECT  112050.0 1024200.0 113250.0 1025400.0 ;
      RECT  114000.0 1026600.0 115200.0 1027800.0 ;
      RECT  130800.0 1025700.0 129600.0 1026900.0 ;
      RECT  122400.0 1043250.0 123600.0 1045200.0 ;
      RECT  122400.0 1031400.0 123600.0 1033350.0 ;
      RECT  117600.0 1032750.0 118800.0 1030950.0 ;
      RECT  117600.0 1042050.0 118800.0 1045650.0 ;
      RECT  120300.0 1032750.0 121200.0 1042050.0 ;
      RECT  117600.0 1042050.0 118800.0 1043250.0 ;
      RECT  120000.0 1042050.0 121200.0 1043250.0 ;
      RECT  120000.0 1042050.0 121200.0 1043250.0 ;
      RECT  117600.0 1042050.0 118800.0 1043250.0 ;
      RECT  117600.0 1032750.0 118800.0 1033950.0 ;
      RECT  120000.0 1032750.0 121200.0 1033950.0 ;
      RECT  120000.0 1032750.0 121200.0 1033950.0 ;
      RECT  117600.0 1032750.0 118800.0 1033950.0 ;
      RECT  122400.0 1042650.0 123600.0 1043850.0 ;
      RECT  122400.0 1032750.0 123600.0 1033950.0 ;
      RECT  118200.0 1037400.0 119400.0 1038600.0 ;
      RECT  118200.0 1037400.0 119400.0 1038600.0 ;
      RECT  120750.0 1037550.0 121650.0 1038450.0 ;
      RECT  115800.0 1044750.0 125400.0 1045650.0 ;
      RECT  115800.0 1030950.0 125400.0 1031850.0 ;
      RECT  127200.0 1033350.0 128400.0 1030950.0 ;
      RECT  127200.0 1042050.0 128400.0 1045650.0 ;
      RECT  132000.0 1042050.0 133200.0 1045650.0 ;
      RECT  134400.0 1043250.0 135600.0 1045200.0 ;
      RECT  134400.0 1031400.0 135600.0 1033350.0 ;
      RECT  127200.0 1042050.0 128400.0 1043250.0 ;
      RECT  129600.0 1042050.0 130800.0 1043250.0 ;
      RECT  129600.0 1042050.0 130800.0 1043250.0 ;
      RECT  127200.0 1042050.0 128400.0 1043250.0 ;
      RECT  129600.0 1042050.0 130800.0 1043250.0 ;
      RECT  132000.0 1042050.0 133200.0 1043250.0 ;
      RECT  132000.0 1042050.0 133200.0 1043250.0 ;
      RECT  129600.0 1042050.0 130800.0 1043250.0 ;
      RECT  127200.0 1033350.0 128400.0 1034550.0 ;
      RECT  129600.0 1033350.0 130800.0 1034550.0 ;
      RECT  129600.0 1033350.0 130800.0 1034550.0 ;
      RECT  127200.0 1033350.0 128400.0 1034550.0 ;
      RECT  129600.0 1033350.0 130800.0 1034550.0 ;
      RECT  132000.0 1033350.0 133200.0 1034550.0 ;
      RECT  132000.0 1033350.0 133200.0 1034550.0 ;
      RECT  129600.0 1033350.0 130800.0 1034550.0 ;
      RECT  134400.0 1042650.0 135600.0 1043850.0 ;
      RECT  134400.0 1032750.0 135600.0 1033950.0 ;
      RECT  132000.0 1035900.0 130800.0 1037100.0 ;
      RECT  129000.0 1038600.0 127800.0 1039800.0 ;
      RECT  129600.0 1042050.0 130800.0 1043250.0 ;
      RECT  132000.0 1033350.0 133200.0 1034550.0 ;
      RECT  133200.0 1038600.0 132000.0 1039800.0 ;
      RECT  127800.0 1038600.0 129000.0 1039800.0 ;
      RECT  130800.0 1035900.0 132000.0 1037100.0 ;
      RECT  132000.0 1038600.0 133200.0 1039800.0 ;
      RECT  125400.0 1044750.0 139800.0 1045650.0 ;
      RECT  125400.0 1030950.0 139800.0 1031850.0 ;
      RECT  146400.0 1043250.0 147600.0 1045200.0 ;
      RECT  146400.0 1031400.0 147600.0 1033350.0 ;
      RECT  141600.0 1032750.0 142800.0 1030950.0 ;
      RECT  141600.0 1042050.0 142800.0 1045650.0 ;
      RECT  144300.0 1032750.0 145200.0 1042050.0 ;
      RECT  141600.0 1042050.0 142800.0 1043250.0 ;
      RECT  144000.0 1042050.0 145200.0 1043250.0 ;
      RECT  144000.0 1042050.0 145200.0 1043250.0 ;
      RECT  141600.0 1042050.0 142800.0 1043250.0 ;
      RECT  141600.0 1032750.0 142800.0 1033950.0 ;
      RECT  144000.0 1032750.0 145200.0 1033950.0 ;
      RECT  144000.0 1032750.0 145200.0 1033950.0 ;
      RECT  141600.0 1032750.0 142800.0 1033950.0 ;
      RECT  146400.0 1042650.0 147600.0 1043850.0 ;
      RECT  146400.0 1032750.0 147600.0 1033950.0 ;
      RECT  142200.0 1037400.0 143400.0 1038600.0 ;
      RECT  142200.0 1037400.0 143400.0 1038600.0 ;
      RECT  144750.0 1037550.0 145650.0 1038450.0 ;
      RECT  139800.0 1044750.0 149400.0 1045650.0 ;
      RECT  139800.0 1030950.0 149400.0 1031850.0 ;
      RECT  112050.0 1037400.0 113250.0 1038600.0 ;
      RECT  114000.0 1035000.0 115200.0 1036200.0 ;
      RECT  130800.0 1035900.0 129600.0 1037100.0 ;
      RECT  122400.0 1047150.0 123600.0 1045200.0 ;
      RECT  122400.0 1059000.0 123600.0 1057050.0 ;
      RECT  117600.0 1057650.0 118800.0 1059450.0 ;
      RECT  117600.0 1048350.0 118800.0 1044750.0 ;
      RECT  120300.0 1057650.0 121200.0 1048350.0 ;
      RECT  117600.0 1048350.0 118800.0 1047150.0 ;
      RECT  120000.0 1048350.0 121200.0 1047150.0 ;
      RECT  120000.0 1048350.0 121200.0 1047150.0 ;
      RECT  117600.0 1048350.0 118800.0 1047150.0 ;
      RECT  117600.0 1057650.0 118800.0 1056450.0 ;
      RECT  120000.0 1057650.0 121200.0 1056450.0 ;
      RECT  120000.0 1057650.0 121200.0 1056450.0 ;
      RECT  117600.0 1057650.0 118800.0 1056450.0 ;
      RECT  122400.0 1047750.0 123600.0 1046550.0 ;
      RECT  122400.0 1057650.0 123600.0 1056450.0 ;
      RECT  118200.0 1053000.0 119400.0 1051800.0 ;
      RECT  118200.0 1053000.0 119400.0 1051800.0 ;
      RECT  120750.0 1052850.0 121650.0 1051950.0 ;
      RECT  115800.0 1045650.0 125400.0 1044750.0 ;
      RECT  115800.0 1059450.0 125400.0 1058550.0 ;
      RECT  127200.0 1057050.0 128400.0 1059450.0 ;
      RECT  127200.0 1048350.0 128400.0 1044750.0 ;
      RECT  132000.0 1048350.0 133200.0 1044750.0 ;
      RECT  134400.0 1047150.0 135600.0 1045200.0 ;
      RECT  134400.0 1059000.0 135600.0 1057050.0 ;
      RECT  127200.0 1048350.0 128400.0 1047150.0 ;
      RECT  129600.0 1048350.0 130800.0 1047150.0 ;
      RECT  129600.0 1048350.0 130800.0 1047150.0 ;
      RECT  127200.0 1048350.0 128400.0 1047150.0 ;
      RECT  129600.0 1048350.0 130800.0 1047150.0 ;
      RECT  132000.0 1048350.0 133200.0 1047150.0 ;
      RECT  132000.0 1048350.0 133200.0 1047150.0 ;
      RECT  129600.0 1048350.0 130800.0 1047150.0 ;
      RECT  127200.0 1057050.0 128400.0 1055850.0 ;
      RECT  129600.0 1057050.0 130800.0 1055850.0 ;
      RECT  129600.0 1057050.0 130800.0 1055850.0 ;
      RECT  127200.0 1057050.0 128400.0 1055850.0 ;
      RECT  129600.0 1057050.0 130800.0 1055850.0 ;
      RECT  132000.0 1057050.0 133200.0 1055850.0 ;
      RECT  132000.0 1057050.0 133200.0 1055850.0 ;
      RECT  129600.0 1057050.0 130800.0 1055850.0 ;
      RECT  134400.0 1047750.0 135600.0 1046550.0 ;
      RECT  134400.0 1057650.0 135600.0 1056450.0 ;
      RECT  132000.0 1054500.0 130800.0 1053300.0 ;
      RECT  129000.0 1051800.0 127800.0 1050600.0 ;
      RECT  129600.0 1048350.0 130800.0 1047150.0 ;
      RECT  132000.0 1057050.0 133200.0 1055850.0 ;
      RECT  133200.0 1051800.0 132000.0 1050600.0 ;
      RECT  127800.0 1051800.0 129000.0 1050600.0 ;
      RECT  130800.0 1054500.0 132000.0 1053300.0 ;
      RECT  132000.0 1051800.0 133200.0 1050600.0 ;
      RECT  125400.0 1045650.0 139800.0 1044750.0 ;
      RECT  125400.0 1059450.0 139800.0 1058550.0 ;
      RECT  146400.0 1047150.0 147600.0 1045200.0 ;
      RECT  146400.0 1059000.0 147600.0 1057050.0 ;
      RECT  141600.0 1057650.0 142800.0 1059450.0 ;
      RECT  141600.0 1048350.0 142800.0 1044750.0 ;
      RECT  144300.0 1057650.0 145200.0 1048350.0 ;
      RECT  141600.0 1048350.0 142800.0 1047150.0 ;
      RECT  144000.0 1048350.0 145200.0 1047150.0 ;
      RECT  144000.0 1048350.0 145200.0 1047150.0 ;
      RECT  141600.0 1048350.0 142800.0 1047150.0 ;
      RECT  141600.0 1057650.0 142800.0 1056450.0 ;
      RECT  144000.0 1057650.0 145200.0 1056450.0 ;
      RECT  144000.0 1057650.0 145200.0 1056450.0 ;
      RECT  141600.0 1057650.0 142800.0 1056450.0 ;
      RECT  146400.0 1047750.0 147600.0 1046550.0 ;
      RECT  146400.0 1057650.0 147600.0 1056450.0 ;
      RECT  142200.0 1053000.0 143400.0 1051800.0 ;
      RECT  142200.0 1053000.0 143400.0 1051800.0 ;
      RECT  144750.0 1052850.0 145650.0 1051950.0 ;
      RECT  139800.0 1045650.0 149400.0 1044750.0 ;
      RECT  139800.0 1059450.0 149400.0 1058550.0 ;
      RECT  112050.0 1051800.0 113250.0 1053000.0 ;
      RECT  114000.0 1054200.0 115200.0 1055400.0 ;
      RECT  130800.0 1053300.0 129600.0 1054500.0 ;
      RECT  122400.0 1070850.0 123600.0 1072800.0 ;
      RECT  122400.0 1059000.0 123600.0 1060950.0 ;
      RECT  117600.0 1060350.0 118800.0 1058550.0 ;
      RECT  117600.0 1069650.0 118800.0 1073250.0 ;
      RECT  120300.0 1060350.0 121200.0 1069650.0 ;
      RECT  117600.0 1069650.0 118800.0 1070850.0 ;
      RECT  120000.0 1069650.0 121200.0 1070850.0 ;
      RECT  120000.0 1069650.0 121200.0 1070850.0 ;
      RECT  117600.0 1069650.0 118800.0 1070850.0 ;
      RECT  117600.0 1060350.0 118800.0 1061550.0 ;
      RECT  120000.0 1060350.0 121200.0 1061550.0 ;
      RECT  120000.0 1060350.0 121200.0 1061550.0 ;
      RECT  117600.0 1060350.0 118800.0 1061550.0 ;
      RECT  122400.0 1070250.0 123600.0 1071450.0 ;
      RECT  122400.0 1060350.0 123600.0 1061550.0 ;
      RECT  118200.0 1065000.0 119400.0 1066200.0 ;
      RECT  118200.0 1065000.0 119400.0 1066200.0 ;
      RECT  120750.0 1065150.0 121650.0 1066050.0 ;
      RECT  115800.0 1072350.0 125400.0 1073250.0 ;
      RECT  115800.0 1058550.0 125400.0 1059450.0 ;
      RECT  127200.0 1060950.0 128400.0 1058550.0 ;
      RECT  127200.0 1069650.0 128400.0 1073250.0 ;
      RECT  132000.0 1069650.0 133200.0 1073250.0 ;
      RECT  134400.0 1070850.0 135600.0 1072800.0 ;
      RECT  134400.0 1059000.0 135600.0 1060950.0 ;
      RECT  127200.0 1069650.0 128400.0 1070850.0 ;
      RECT  129600.0 1069650.0 130800.0 1070850.0 ;
      RECT  129600.0 1069650.0 130800.0 1070850.0 ;
      RECT  127200.0 1069650.0 128400.0 1070850.0 ;
      RECT  129600.0 1069650.0 130800.0 1070850.0 ;
      RECT  132000.0 1069650.0 133200.0 1070850.0 ;
      RECT  132000.0 1069650.0 133200.0 1070850.0 ;
      RECT  129600.0 1069650.0 130800.0 1070850.0 ;
      RECT  127200.0 1060950.0 128400.0 1062150.0 ;
      RECT  129600.0 1060950.0 130800.0 1062150.0 ;
      RECT  129600.0 1060950.0 130800.0 1062150.0 ;
      RECT  127200.0 1060950.0 128400.0 1062150.0 ;
      RECT  129600.0 1060950.0 130800.0 1062150.0 ;
      RECT  132000.0 1060950.0 133200.0 1062150.0 ;
      RECT  132000.0 1060950.0 133200.0 1062150.0 ;
      RECT  129600.0 1060950.0 130800.0 1062150.0 ;
      RECT  134400.0 1070250.0 135600.0 1071450.0 ;
      RECT  134400.0 1060350.0 135600.0 1061550.0 ;
      RECT  132000.0 1063500.0 130800.0 1064700.0 ;
      RECT  129000.0 1066200.0 127800.0 1067400.0 ;
      RECT  129600.0 1069650.0 130800.0 1070850.0 ;
      RECT  132000.0 1060950.0 133200.0 1062150.0 ;
      RECT  133200.0 1066200.0 132000.0 1067400.0 ;
      RECT  127800.0 1066200.0 129000.0 1067400.0 ;
      RECT  130800.0 1063500.0 132000.0 1064700.0 ;
      RECT  132000.0 1066200.0 133200.0 1067400.0 ;
      RECT  125400.0 1072350.0 139800.0 1073250.0 ;
      RECT  125400.0 1058550.0 139800.0 1059450.0 ;
      RECT  146400.0 1070850.0 147600.0 1072800.0 ;
      RECT  146400.0 1059000.0 147600.0 1060950.0 ;
      RECT  141600.0 1060350.0 142800.0 1058550.0 ;
      RECT  141600.0 1069650.0 142800.0 1073250.0 ;
      RECT  144300.0 1060350.0 145200.0 1069650.0 ;
      RECT  141600.0 1069650.0 142800.0 1070850.0 ;
      RECT  144000.0 1069650.0 145200.0 1070850.0 ;
      RECT  144000.0 1069650.0 145200.0 1070850.0 ;
      RECT  141600.0 1069650.0 142800.0 1070850.0 ;
      RECT  141600.0 1060350.0 142800.0 1061550.0 ;
      RECT  144000.0 1060350.0 145200.0 1061550.0 ;
      RECT  144000.0 1060350.0 145200.0 1061550.0 ;
      RECT  141600.0 1060350.0 142800.0 1061550.0 ;
      RECT  146400.0 1070250.0 147600.0 1071450.0 ;
      RECT  146400.0 1060350.0 147600.0 1061550.0 ;
      RECT  142200.0 1065000.0 143400.0 1066200.0 ;
      RECT  142200.0 1065000.0 143400.0 1066200.0 ;
      RECT  144750.0 1065150.0 145650.0 1066050.0 ;
      RECT  139800.0 1072350.0 149400.0 1073250.0 ;
      RECT  139800.0 1058550.0 149400.0 1059450.0 ;
      RECT  112050.0 1065000.0 113250.0 1066200.0 ;
      RECT  114000.0 1062600.0 115200.0 1063800.0 ;
      RECT  130800.0 1063500.0 129600.0 1064700.0 ;
      RECT  122400.0 1074750.0 123600.0 1072800.0 ;
      RECT  122400.0 1086600.0 123600.0 1084650.0 ;
      RECT  117600.0 1085250.0 118800.0 1087050.0 ;
      RECT  117600.0 1075950.0 118800.0 1072350.0 ;
      RECT  120300.0 1085250.0 121200.0 1075950.0 ;
      RECT  117600.0 1075950.0 118800.0 1074750.0 ;
      RECT  120000.0 1075950.0 121200.0 1074750.0 ;
      RECT  120000.0 1075950.0 121200.0 1074750.0 ;
      RECT  117600.0 1075950.0 118800.0 1074750.0 ;
      RECT  117600.0 1085250.0 118800.0 1084050.0 ;
      RECT  120000.0 1085250.0 121200.0 1084050.0 ;
      RECT  120000.0 1085250.0 121200.0 1084050.0 ;
      RECT  117600.0 1085250.0 118800.0 1084050.0 ;
      RECT  122400.0 1075350.0 123600.0 1074150.0 ;
      RECT  122400.0 1085250.0 123600.0 1084050.0 ;
      RECT  118200.0 1080600.0 119400.0 1079400.0 ;
      RECT  118200.0 1080600.0 119400.0 1079400.0 ;
      RECT  120750.0 1080450.0 121650.0 1079550.0 ;
      RECT  115800.0 1073250.0 125400.0 1072350.0 ;
      RECT  115800.0 1087050.0 125400.0 1086150.0 ;
      RECT  127200.0 1084650.0 128400.0 1087050.0 ;
      RECT  127200.0 1075950.0 128400.0 1072350.0 ;
      RECT  132000.0 1075950.0 133200.0 1072350.0 ;
      RECT  134400.0 1074750.0 135600.0 1072800.0 ;
      RECT  134400.0 1086600.0 135600.0 1084650.0 ;
      RECT  127200.0 1075950.0 128400.0 1074750.0 ;
      RECT  129600.0 1075950.0 130800.0 1074750.0 ;
      RECT  129600.0 1075950.0 130800.0 1074750.0 ;
      RECT  127200.0 1075950.0 128400.0 1074750.0 ;
      RECT  129600.0 1075950.0 130800.0 1074750.0 ;
      RECT  132000.0 1075950.0 133200.0 1074750.0 ;
      RECT  132000.0 1075950.0 133200.0 1074750.0 ;
      RECT  129600.0 1075950.0 130800.0 1074750.0 ;
      RECT  127200.0 1084650.0 128400.0 1083450.0 ;
      RECT  129600.0 1084650.0 130800.0 1083450.0 ;
      RECT  129600.0 1084650.0 130800.0 1083450.0 ;
      RECT  127200.0 1084650.0 128400.0 1083450.0 ;
      RECT  129600.0 1084650.0 130800.0 1083450.0 ;
      RECT  132000.0 1084650.0 133200.0 1083450.0 ;
      RECT  132000.0 1084650.0 133200.0 1083450.0 ;
      RECT  129600.0 1084650.0 130800.0 1083450.0 ;
      RECT  134400.0 1075350.0 135600.0 1074150.0 ;
      RECT  134400.0 1085250.0 135600.0 1084050.0 ;
      RECT  132000.0 1082100.0 130800.0 1080900.0 ;
      RECT  129000.0 1079400.0 127800.0 1078200.0 ;
      RECT  129600.0 1075950.0 130800.0 1074750.0 ;
      RECT  132000.0 1084650.0 133200.0 1083450.0 ;
      RECT  133200.0 1079400.0 132000.0 1078200.0 ;
      RECT  127800.0 1079400.0 129000.0 1078200.0 ;
      RECT  130800.0 1082100.0 132000.0 1080900.0 ;
      RECT  132000.0 1079400.0 133200.0 1078200.0 ;
      RECT  125400.0 1073250.0 139800.0 1072350.0 ;
      RECT  125400.0 1087050.0 139800.0 1086150.0 ;
      RECT  146400.0 1074750.0 147600.0 1072800.0 ;
      RECT  146400.0 1086600.0 147600.0 1084650.0 ;
      RECT  141600.0 1085250.0 142800.0 1087050.0 ;
      RECT  141600.0 1075950.0 142800.0 1072350.0 ;
      RECT  144300.0 1085250.0 145200.0 1075950.0 ;
      RECT  141600.0 1075950.0 142800.0 1074750.0 ;
      RECT  144000.0 1075950.0 145200.0 1074750.0 ;
      RECT  144000.0 1075950.0 145200.0 1074750.0 ;
      RECT  141600.0 1075950.0 142800.0 1074750.0 ;
      RECT  141600.0 1085250.0 142800.0 1084050.0 ;
      RECT  144000.0 1085250.0 145200.0 1084050.0 ;
      RECT  144000.0 1085250.0 145200.0 1084050.0 ;
      RECT  141600.0 1085250.0 142800.0 1084050.0 ;
      RECT  146400.0 1075350.0 147600.0 1074150.0 ;
      RECT  146400.0 1085250.0 147600.0 1084050.0 ;
      RECT  142200.0 1080600.0 143400.0 1079400.0 ;
      RECT  142200.0 1080600.0 143400.0 1079400.0 ;
      RECT  144750.0 1080450.0 145650.0 1079550.0 ;
      RECT  139800.0 1073250.0 149400.0 1072350.0 ;
      RECT  139800.0 1087050.0 149400.0 1086150.0 ;
      RECT  112050.0 1079400.0 113250.0 1080600.0 ;
      RECT  114000.0 1081800.0 115200.0 1083000.0 ;
      RECT  130800.0 1080900.0 129600.0 1082100.0 ;
      RECT  122400.0 1098450.0 123600.0 1100400.0 ;
      RECT  122400.0 1086600.0 123600.0 1088550.0 ;
      RECT  117600.0 1087950.0 118800.0 1086150.0 ;
      RECT  117600.0 1097250.0 118800.0 1100850.0 ;
      RECT  120300.0 1087950.0 121200.0 1097250.0 ;
      RECT  117600.0 1097250.0 118800.0 1098450.0 ;
      RECT  120000.0 1097250.0 121200.0 1098450.0 ;
      RECT  120000.0 1097250.0 121200.0 1098450.0 ;
      RECT  117600.0 1097250.0 118800.0 1098450.0 ;
      RECT  117600.0 1087950.0 118800.0 1089150.0 ;
      RECT  120000.0 1087950.0 121200.0 1089150.0 ;
      RECT  120000.0 1087950.0 121200.0 1089150.0 ;
      RECT  117600.0 1087950.0 118800.0 1089150.0 ;
      RECT  122400.0 1097850.0 123600.0 1099050.0 ;
      RECT  122400.0 1087950.0 123600.0 1089150.0 ;
      RECT  118200.0 1092600.0 119400.0 1093800.0 ;
      RECT  118200.0 1092600.0 119400.0 1093800.0 ;
      RECT  120750.0 1092750.0 121650.0 1093650.0 ;
      RECT  115800.0 1099950.0 125400.0 1100850.0 ;
      RECT  115800.0 1086150.0 125400.0 1087050.0 ;
      RECT  127200.0 1088550.0 128400.0 1086150.0 ;
      RECT  127200.0 1097250.0 128400.0 1100850.0 ;
      RECT  132000.0 1097250.0 133200.0 1100850.0 ;
      RECT  134400.0 1098450.0 135600.0 1100400.0 ;
      RECT  134400.0 1086600.0 135600.0 1088550.0 ;
      RECT  127200.0 1097250.0 128400.0 1098450.0 ;
      RECT  129600.0 1097250.0 130800.0 1098450.0 ;
      RECT  129600.0 1097250.0 130800.0 1098450.0 ;
      RECT  127200.0 1097250.0 128400.0 1098450.0 ;
      RECT  129600.0 1097250.0 130800.0 1098450.0 ;
      RECT  132000.0 1097250.0 133200.0 1098450.0 ;
      RECT  132000.0 1097250.0 133200.0 1098450.0 ;
      RECT  129600.0 1097250.0 130800.0 1098450.0 ;
      RECT  127200.0 1088550.0 128400.0 1089750.0 ;
      RECT  129600.0 1088550.0 130800.0 1089750.0 ;
      RECT  129600.0 1088550.0 130800.0 1089750.0 ;
      RECT  127200.0 1088550.0 128400.0 1089750.0 ;
      RECT  129600.0 1088550.0 130800.0 1089750.0 ;
      RECT  132000.0 1088550.0 133200.0 1089750.0 ;
      RECT  132000.0 1088550.0 133200.0 1089750.0 ;
      RECT  129600.0 1088550.0 130800.0 1089750.0 ;
      RECT  134400.0 1097850.0 135600.0 1099050.0 ;
      RECT  134400.0 1087950.0 135600.0 1089150.0 ;
      RECT  132000.0 1091100.0 130800.0 1092300.0 ;
      RECT  129000.0 1093800.0 127800.0 1095000.0 ;
      RECT  129600.0 1097250.0 130800.0 1098450.0 ;
      RECT  132000.0 1088550.0 133200.0 1089750.0 ;
      RECT  133200.0 1093800.0 132000.0 1095000.0 ;
      RECT  127800.0 1093800.0 129000.0 1095000.0 ;
      RECT  130800.0 1091100.0 132000.0 1092300.0 ;
      RECT  132000.0 1093800.0 133200.0 1095000.0 ;
      RECT  125400.0 1099950.0 139800.0 1100850.0 ;
      RECT  125400.0 1086150.0 139800.0 1087050.0 ;
      RECT  146400.0 1098450.0 147600.0 1100400.0 ;
      RECT  146400.0 1086600.0 147600.0 1088550.0 ;
      RECT  141600.0 1087950.0 142800.0 1086150.0 ;
      RECT  141600.0 1097250.0 142800.0 1100850.0 ;
      RECT  144300.0 1087950.0 145200.0 1097250.0 ;
      RECT  141600.0 1097250.0 142800.0 1098450.0 ;
      RECT  144000.0 1097250.0 145200.0 1098450.0 ;
      RECT  144000.0 1097250.0 145200.0 1098450.0 ;
      RECT  141600.0 1097250.0 142800.0 1098450.0 ;
      RECT  141600.0 1087950.0 142800.0 1089150.0 ;
      RECT  144000.0 1087950.0 145200.0 1089150.0 ;
      RECT  144000.0 1087950.0 145200.0 1089150.0 ;
      RECT  141600.0 1087950.0 142800.0 1089150.0 ;
      RECT  146400.0 1097850.0 147600.0 1099050.0 ;
      RECT  146400.0 1087950.0 147600.0 1089150.0 ;
      RECT  142200.0 1092600.0 143400.0 1093800.0 ;
      RECT  142200.0 1092600.0 143400.0 1093800.0 ;
      RECT  144750.0 1092750.0 145650.0 1093650.0 ;
      RECT  139800.0 1099950.0 149400.0 1100850.0 ;
      RECT  139800.0 1086150.0 149400.0 1087050.0 ;
      RECT  112050.0 1092600.0 113250.0 1093800.0 ;
      RECT  114000.0 1090200.0 115200.0 1091400.0 ;
      RECT  130800.0 1091100.0 129600.0 1092300.0 ;
      RECT  122400.0 1102350.0 123600.0 1100400.0 ;
      RECT  122400.0 1114200.0 123600.0 1112250.0 ;
      RECT  117600.0 1112850.0 118800.0 1114650.0 ;
      RECT  117600.0 1103550.0 118800.0 1099950.0 ;
      RECT  120300.0 1112850.0 121200.0 1103550.0 ;
      RECT  117600.0 1103550.0 118800.0 1102350.0 ;
      RECT  120000.0 1103550.0 121200.0 1102350.0 ;
      RECT  120000.0 1103550.0 121200.0 1102350.0 ;
      RECT  117600.0 1103550.0 118800.0 1102350.0 ;
      RECT  117600.0 1112850.0 118800.0 1111650.0 ;
      RECT  120000.0 1112850.0 121200.0 1111650.0 ;
      RECT  120000.0 1112850.0 121200.0 1111650.0 ;
      RECT  117600.0 1112850.0 118800.0 1111650.0 ;
      RECT  122400.0 1102950.0 123600.0 1101750.0 ;
      RECT  122400.0 1112850.0 123600.0 1111650.0 ;
      RECT  118200.0 1108200.0 119400.0 1107000.0 ;
      RECT  118200.0 1108200.0 119400.0 1107000.0 ;
      RECT  120750.0 1108050.0 121650.0 1107150.0 ;
      RECT  115800.0 1100850.0 125400.0 1099950.0 ;
      RECT  115800.0 1114650.0 125400.0 1113750.0 ;
      RECT  127200.0 1112250.0 128400.0 1114650.0 ;
      RECT  127200.0 1103550.0 128400.0 1099950.0 ;
      RECT  132000.0 1103550.0 133200.0 1099950.0 ;
      RECT  134400.0 1102350.0 135600.0 1100400.0 ;
      RECT  134400.0 1114200.0 135600.0 1112250.0 ;
      RECT  127200.0 1103550.0 128400.0 1102350.0 ;
      RECT  129600.0 1103550.0 130800.0 1102350.0 ;
      RECT  129600.0 1103550.0 130800.0 1102350.0 ;
      RECT  127200.0 1103550.0 128400.0 1102350.0 ;
      RECT  129600.0 1103550.0 130800.0 1102350.0 ;
      RECT  132000.0 1103550.0 133200.0 1102350.0 ;
      RECT  132000.0 1103550.0 133200.0 1102350.0 ;
      RECT  129600.0 1103550.0 130800.0 1102350.0 ;
      RECT  127200.0 1112250.0 128400.0 1111050.0 ;
      RECT  129600.0 1112250.0 130800.0 1111050.0 ;
      RECT  129600.0 1112250.0 130800.0 1111050.0 ;
      RECT  127200.0 1112250.0 128400.0 1111050.0 ;
      RECT  129600.0 1112250.0 130800.0 1111050.0 ;
      RECT  132000.0 1112250.0 133200.0 1111050.0 ;
      RECT  132000.0 1112250.0 133200.0 1111050.0 ;
      RECT  129600.0 1112250.0 130800.0 1111050.0 ;
      RECT  134400.0 1102950.0 135600.0 1101750.0 ;
      RECT  134400.0 1112850.0 135600.0 1111650.0 ;
      RECT  132000.0 1109700.0 130800.0 1108500.0 ;
      RECT  129000.0 1107000.0 127800.0 1105800.0 ;
      RECT  129600.0 1103550.0 130800.0 1102350.0 ;
      RECT  132000.0 1112250.0 133200.0 1111050.0 ;
      RECT  133200.0 1107000.0 132000.0 1105800.0 ;
      RECT  127800.0 1107000.0 129000.0 1105800.0 ;
      RECT  130800.0 1109700.0 132000.0 1108500.0 ;
      RECT  132000.0 1107000.0 133200.0 1105800.0 ;
      RECT  125400.0 1100850.0 139800.0 1099950.0 ;
      RECT  125400.0 1114650.0 139800.0 1113750.0 ;
      RECT  146400.0 1102350.0 147600.0 1100400.0 ;
      RECT  146400.0 1114200.0 147600.0 1112250.0 ;
      RECT  141600.0 1112850.0 142800.0 1114650.0 ;
      RECT  141600.0 1103550.0 142800.0 1099950.0 ;
      RECT  144300.0 1112850.0 145200.0 1103550.0 ;
      RECT  141600.0 1103550.0 142800.0 1102350.0 ;
      RECT  144000.0 1103550.0 145200.0 1102350.0 ;
      RECT  144000.0 1103550.0 145200.0 1102350.0 ;
      RECT  141600.0 1103550.0 142800.0 1102350.0 ;
      RECT  141600.0 1112850.0 142800.0 1111650.0 ;
      RECT  144000.0 1112850.0 145200.0 1111650.0 ;
      RECT  144000.0 1112850.0 145200.0 1111650.0 ;
      RECT  141600.0 1112850.0 142800.0 1111650.0 ;
      RECT  146400.0 1102950.0 147600.0 1101750.0 ;
      RECT  146400.0 1112850.0 147600.0 1111650.0 ;
      RECT  142200.0 1108200.0 143400.0 1107000.0 ;
      RECT  142200.0 1108200.0 143400.0 1107000.0 ;
      RECT  144750.0 1108050.0 145650.0 1107150.0 ;
      RECT  139800.0 1100850.0 149400.0 1099950.0 ;
      RECT  139800.0 1114650.0 149400.0 1113750.0 ;
      RECT  112050.0 1107000.0 113250.0 1108200.0 ;
      RECT  114000.0 1109400.0 115200.0 1110600.0 ;
      RECT  130800.0 1108500.0 129600.0 1109700.0 ;
      RECT  122400.0 1126050.0 123600.0 1128000.0 ;
      RECT  122400.0 1114200.0 123600.0 1116150.0 ;
      RECT  117600.0 1115550.0 118800.0 1113750.0 ;
      RECT  117600.0 1124850.0 118800.0 1128450.0 ;
      RECT  120300.0 1115550.0 121200.0 1124850.0 ;
      RECT  117600.0 1124850.0 118800.0 1126050.0 ;
      RECT  120000.0 1124850.0 121200.0 1126050.0 ;
      RECT  120000.0 1124850.0 121200.0 1126050.0 ;
      RECT  117600.0 1124850.0 118800.0 1126050.0 ;
      RECT  117600.0 1115550.0 118800.0 1116750.0 ;
      RECT  120000.0 1115550.0 121200.0 1116750.0 ;
      RECT  120000.0 1115550.0 121200.0 1116750.0 ;
      RECT  117600.0 1115550.0 118800.0 1116750.0 ;
      RECT  122400.0 1125450.0 123600.0 1126650.0 ;
      RECT  122400.0 1115550.0 123600.0 1116750.0 ;
      RECT  118200.0 1120200.0 119400.0 1121400.0 ;
      RECT  118200.0 1120200.0 119400.0 1121400.0 ;
      RECT  120750.0 1120350.0 121650.0 1121250.0 ;
      RECT  115800.0 1127550.0 125400.0 1128450.0 ;
      RECT  115800.0 1113750.0 125400.0 1114650.0 ;
      RECT  127200.0 1116150.0 128400.0 1113750.0 ;
      RECT  127200.0 1124850.0 128400.0 1128450.0 ;
      RECT  132000.0 1124850.0 133200.0 1128450.0 ;
      RECT  134400.0 1126050.0 135600.0 1128000.0 ;
      RECT  134400.0 1114200.0 135600.0 1116150.0 ;
      RECT  127200.0 1124850.0 128400.0 1126050.0 ;
      RECT  129600.0 1124850.0 130800.0 1126050.0 ;
      RECT  129600.0 1124850.0 130800.0 1126050.0 ;
      RECT  127200.0 1124850.0 128400.0 1126050.0 ;
      RECT  129600.0 1124850.0 130800.0 1126050.0 ;
      RECT  132000.0 1124850.0 133200.0 1126050.0 ;
      RECT  132000.0 1124850.0 133200.0 1126050.0 ;
      RECT  129600.0 1124850.0 130800.0 1126050.0 ;
      RECT  127200.0 1116150.0 128400.0 1117350.0 ;
      RECT  129600.0 1116150.0 130800.0 1117350.0 ;
      RECT  129600.0 1116150.0 130800.0 1117350.0 ;
      RECT  127200.0 1116150.0 128400.0 1117350.0 ;
      RECT  129600.0 1116150.0 130800.0 1117350.0 ;
      RECT  132000.0 1116150.0 133200.0 1117350.0 ;
      RECT  132000.0 1116150.0 133200.0 1117350.0 ;
      RECT  129600.0 1116150.0 130800.0 1117350.0 ;
      RECT  134400.0 1125450.0 135600.0 1126650.0 ;
      RECT  134400.0 1115550.0 135600.0 1116750.0 ;
      RECT  132000.0 1118700.0 130800.0 1119900.0 ;
      RECT  129000.0 1121400.0 127800.0 1122600.0 ;
      RECT  129600.0 1124850.0 130800.0 1126050.0 ;
      RECT  132000.0 1116150.0 133200.0 1117350.0 ;
      RECT  133200.0 1121400.0 132000.0 1122600.0 ;
      RECT  127800.0 1121400.0 129000.0 1122600.0 ;
      RECT  130800.0 1118700.0 132000.0 1119900.0 ;
      RECT  132000.0 1121400.0 133200.0 1122600.0 ;
      RECT  125400.0 1127550.0 139800.0 1128450.0 ;
      RECT  125400.0 1113750.0 139800.0 1114650.0 ;
      RECT  146400.0 1126050.0 147600.0 1128000.0 ;
      RECT  146400.0 1114200.0 147600.0 1116150.0 ;
      RECT  141600.0 1115550.0 142800.0 1113750.0 ;
      RECT  141600.0 1124850.0 142800.0 1128450.0 ;
      RECT  144300.0 1115550.0 145200.0 1124850.0 ;
      RECT  141600.0 1124850.0 142800.0 1126050.0 ;
      RECT  144000.0 1124850.0 145200.0 1126050.0 ;
      RECT  144000.0 1124850.0 145200.0 1126050.0 ;
      RECT  141600.0 1124850.0 142800.0 1126050.0 ;
      RECT  141600.0 1115550.0 142800.0 1116750.0 ;
      RECT  144000.0 1115550.0 145200.0 1116750.0 ;
      RECT  144000.0 1115550.0 145200.0 1116750.0 ;
      RECT  141600.0 1115550.0 142800.0 1116750.0 ;
      RECT  146400.0 1125450.0 147600.0 1126650.0 ;
      RECT  146400.0 1115550.0 147600.0 1116750.0 ;
      RECT  142200.0 1120200.0 143400.0 1121400.0 ;
      RECT  142200.0 1120200.0 143400.0 1121400.0 ;
      RECT  144750.0 1120350.0 145650.0 1121250.0 ;
      RECT  139800.0 1127550.0 149400.0 1128450.0 ;
      RECT  139800.0 1113750.0 149400.0 1114650.0 ;
      RECT  112050.0 1120200.0 113250.0 1121400.0 ;
      RECT  114000.0 1117800.0 115200.0 1119000.0 ;
      RECT  130800.0 1118700.0 129600.0 1119900.0 ;
      RECT  122400.0 1129950.0 123600.0 1128000.0 ;
      RECT  122400.0 1141800.0 123600.0 1139850.0 ;
      RECT  117600.0 1140450.0 118800.0 1142250.0 ;
      RECT  117600.0 1131150.0 118800.0 1127550.0 ;
      RECT  120300.0 1140450.0 121200.0 1131150.0 ;
      RECT  117600.0 1131150.0 118800.0 1129950.0 ;
      RECT  120000.0 1131150.0 121200.0 1129950.0 ;
      RECT  120000.0 1131150.0 121200.0 1129950.0 ;
      RECT  117600.0 1131150.0 118800.0 1129950.0 ;
      RECT  117600.0 1140450.0 118800.0 1139250.0 ;
      RECT  120000.0 1140450.0 121200.0 1139250.0 ;
      RECT  120000.0 1140450.0 121200.0 1139250.0 ;
      RECT  117600.0 1140450.0 118800.0 1139250.0 ;
      RECT  122400.0 1130550.0 123600.0 1129350.0 ;
      RECT  122400.0 1140450.0 123600.0 1139250.0 ;
      RECT  118200.0 1135800.0 119400.0 1134600.0 ;
      RECT  118200.0 1135800.0 119400.0 1134600.0 ;
      RECT  120750.0 1135650.0 121650.0 1134750.0 ;
      RECT  115800.0 1128450.0 125400.0 1127550.0 ;
      RECT  115800.0 1142250.0 125400.0 1141350.0 ;
      RECT  127200.0 1139850.0 128400.0 1142250.0 ;
      RECT  127200.0 1131150.0 128400.0 1127550.0 ;
      RECT  132000.0 1131150.0 133200.0 1127550.0 ;
      RECT  134400.0 1129950.0 135600.0 1128000.0 ;
      RECT  134400.0 1141800.0 135600.0 1139850.0 ;
      RECT  127200.0 1131150.0 128400.0 1129950.0 ;
      RECT  129600.0 1131150.0 130800.0 1129950.0 ;
      RECT  129600.0 1131150.0 130800.0 1129950.0 ;
      RECT  127200.0 1131150.0 128400.0 1129950.0 ;
      RECT  129600.0 1131150.0 130800.0 1129950.0 ;
      RECT  132000.0 1131150.0 133200.0 1129950.0 ;
      RECT  132000.0 1131150.0 133200.0 1129950.0 ;
      RECT  129600.0 1131150.0 130800.0 1129950.0 ;
      RECT  127200.0 1139850.0 128400.0 1138650.0 ;
      RECT  129600.0 1139850.0 130800.0 1138650.0 ;
      RECT  129600.0 1139850.0 130800.0 1138650.0 ;
      RECT  127200.0 1139850.0 128400.0 1138650.0 ;
      RECT  129600.0 1139850.0 130800.0 1138650.0 ;
      RECT  132000.0 1139850.0 133200.0 1138650.0 ;
      RECT  132000.0 1139850.0 133200.0 1138650.0 ;
      RECT  129600.0 1139850.0 130800.0 1138650.0 ;
      RECT  134400.0 1130550.0 135600.0 1129350.0 ;
      RECT  134400.0 1140450.0 135600.0 1139250.0 ;
      RECT  132000.0 1137300.0 130800.0 1136100.0 ;
      RECT  129000.0 1134600.0 127800.0 1133400.0 ;
      RECT  129600.0 1131150.0 130800.0 1129950.0 ;
      RECT  132000.0 1139850.0 133200.0 1138650.0 ;
      RECT  133200.0 1134600.0 132000.0 1133400.0 ;
      RECT  127800.0 1134600.0 129000.0 1133400.0 ;
      RECT  130800.0 1137300.0 132000.0 1136100.0 ;
      RECT  132000.0 1134600.0 133200.0 1133400.0 ;
      RECT  125400.0 1128450.0 139800.0 1127550.0 ;
      RECT  125400.0 1142250.0 139800.0 1141350.0 ;
      RECT  146400.0 1129950.0 147600.0 1128000.0 ;
      RECT  146400.0 1141800.0 147600.0 1139850.0 ;
      RECT  141600.0 1140450.0 142800.0 1142250.0 ;
      RECT  141600.0 1131150.0 142800.0 1127550.0 ;
      RECT  144300.0 1140450.0 145200.0 1131150.0 ;
      RECT  141600.0 1131150.0 142800.0 1129950.0 ;
      RECT  144000.0 1131150.0 145200.0 1129950.0 ;
      RECT  144000.0 1131150.0 145200.0 1129950.0 ;
      RECT  141600.0 1131150.0 142800.0 1129950.0 ;
      RECT  141600.0 1140450.0 142800.0 1139250.0 ;
      RECT  144000.0 1140450.0 145200.0 1139250.0 ;
      RECT  144000.0 1140450.0 145200.0 1139250.0 ;
      RECT  141600.0 1140450.0 142800.0 1139250.0 ;
      RECT  146400.0 1130550.0 147600.0 1129350.0 ;
      RECT  146400.0 1140450.0 147600.0 1139250.0 ;
      RECT  142200.0 1135800.0 143400.0 1134600.0 ;
      RECT  142200.0 1135800.0 143400.0 1134600.0 ;
      RECT  144750.0 1135650.0 145650.0 1134750.0 ;
      RECT  139800.0 1128450.0 149400.0 1127550.0 ;
      RECT  139800.0 1142250.0 149400.0 1141350.0 ;
      RECT  112050.0 1134600.0 113250.0 1135800.0 ;
      RECT  114000.0 1137000.0 115200.0 1138200.0 ;
      RECT  130800.0 1136100.0 129600.0 1137300.0 ;
      RECT  122400.0 1153650.0 123600.0 1155600.0 ;
      RECT  122400.0 1141800.0 123600.0 1143750.0 ;
      RECT  117600.0 1143150.0 118800.0 1141350.0 ;
      RECT  117600.0 1152450.0 118800.0 1156050.0 ;
      RECT  120300.0 1143150.0 121200.0 1152450.0 ;
      RECT  117600.0 1152450.0 118800.0 1153650.0 ;
      RECT  120000.0 1152450.0 121200.0 1153650.0 ;
      RECT  120000.0 1152450.0 121200.0 1153650.0 ;
      RECT  117600.0 1152450.0 118800.0 1153650.0 ;
      RECT  117600.0 1143150.0 118800.0 1144350.0 ;
      RECT  120000.0 1143150.0 121200.0 1144350.0 ;
      RECT  120000.0 1143150.0 121200.0 1144350.0 ;
      RECT  117600.0 1143150.0 118800.0 1144350.0 ;
      RECT  122400.0 1153050.0 123600.0 1154250.0 ;
      RECT  122400.0 1143150.0 123600.0 1144350.0 ;
      RECT  118200.0 1147800.0 119400.0 1149000.0 ;
      RECT  118200.0 1147800.0 119400.0 1149000.0 ;
      RECT  120750.0 1147950.0 121650.0 1148850.0 ;
      RECT  115800.0 1155150.0 125400.0 1156050.0 ;
      RECT  115800.0 1141350.0 125400.0 1142250.0 ;
      RECT  127200.0 1143750.0 128400.0 1141350.0 ;
      RECT  127200.0 1152450.0 128400.0 1156050.0 ;
      RECT  132000.0 1152450.0 133200.0 1156050.0 ;
      RECT  134400.0 1153650.0 135600.0 1155600.0 ;
      RECT  134400.0 1141800.0 135600.0 1143750.0 ;
      RECT  127200.0 1152450.0 128400.0 1153650.0 ;
      RECT  129600.0 1152450.0 130800.0 1153650.0 ;
      RECT  129600.0 1152450.0 130800.0 1153650.0 ;
      RECT  127200.0 1152450.0 128400.0 1153650.0 ;
      RECT  129600.0 1152450.0 130800.0 1153650.0 ;
      RECT  132000.0 1152450.0 133200.0 1153650.0 ;
      RECT  132000.0 1152450.0 133200.0 1153650.0 ;
      RECT  129600.0 1152450.0 130800.0 1153650.0 ;
      RECT  127200.0 1143750.0 128400.0 1144950.0 ;
      RECT  129600.0 1143750.0 130800.0 1144950.0 ;
      RECT  129600.0 1143750.0 130800.0 1144950.0 ;
      RECT  127200.0 1143750.0 128400.0 1144950.0 ;
      RECT  129600.0 1143750.0 130800.0 1144950.0 ;
      RECT  132000.0 1143750.0 133200.0 1144950.0 ;
      RECT  132000.0 1143750.0 133200.0 1144950.0 ;
      RECT  129600.0 1143750.0 130800.0 1144950.0 ;
      RECT  134400.0 1153050.0 135600.0 1154250.0 ;
      RECT  134400.0 1143150.0 135600.0 1144350.0 ;
      RECT  132000.0 1146300.0 130800.0 1147500.0 ;
      RECT  129000.0 1149000.0 127800.0 1150200.0 ;
      RECT  129600.0 1152450.0 130800.0 1153650.0 ;
      RECT  132000.0 1143750.0 133200.0 1144950.0 ;
      RECT  133200.0 1149000.0 132000.0 1150200.0 ;
      RECT  127800.0 1149000.0 129000.0 1150200.0 ;
      RECT  130800.0 1146300.0 132000.0 1147500.0 ;
      RECT  132000.0 1149000.0 133200.0 1150200.0 ;
      RECT  125400.0 1155150.0 139800.0 1156050.0 ;
      RECT  125400.0 1141350.0 139800.0 1142250.0 ;
      RECT  146400.0 1153650.0 147600.0 1155600.0 ;
      RECT  146400.0 1141800.0 147600.0 1143750.0 ;
      RECT  141600.0 1143150.0 142800.0 1141350.0 ;
      RECT  141600.0 1152450.0 142800.0 1156050.0 ;
      RECT  144300.0 1143150.0 145200.0 1152450.0 ;
      RECT  141600.0 1152450.0 142800.0 1153650.0 ;
      RECT  144000.0 1152450.0 145200.0 1153650.0 ;
      RECT  144000.0 1152450.0 145200.0 1153650.0 ;
      RECT  141600.0 1152450.0 142800.0 1153650.0 ;
      RECT  141600.0 1143150.0 142800.0 1144350.0 ;
      RECT  144000.0 1143150.0 145200.0 1144350.0 ;
      RECT  144000.0 1143150.0 145200.0 1144350.0 ;
      RECT  141600.0 1143150.0 142800.0 1144350.0 ;
      RECT  146400.0 1153050.0 147600.0 1154250.0 ;
      RECT  146400.0 1143150.0 147600.0 1144350.0 ;
      RECT  142200.0 1147800.0 143400.0 1149000.0 ;
      RECT  142200.0 1147800.0 143400.0 1149000.0 ;
      RECT  144750.0 1147950.0 145650.0 1148850.0 ;
      RECT  139800.0 1155150.0 149400.0 1156050.0 ;
      RECT  139800.0 1141350.0 149400.0 1142250.0 ;
      RECT  112050.0 1147800.0 113250.0 1149000.0 ;
      RECT  114000.0 1145400.0 115200.0 1146600.0 ;
      RECT  130800.0 1146300.0 129600.0 1147500.0 ;
      RECT  122400.0 1157550.0 123600.0 1155600.0 ;
      RECT  122400.0 1169400.0 123600.0 1167450.0 ;
      RECT  117600.0 1168050.0 118800.0 1169850.0 ;
      RECT  117600.0 1158750.0 118800.0 1155150.0 ;
      RECT  120300.0 1168050.0 121200.0 1158750.0 ;
      RECT  117600.0 1158750.0 118800.0 1157550.0 ;
      RECT  120000.0 1158750.0 121200.0 1157550.0 ;
      RECT  120000.0 1158750.0 121200.0 1157550.0 ;
      RECT  117600.0 1158750.0 118800.0 1157550.0 ;
      RECT  117600.0 1168050.0 118800.0 1166850.0 ;
      RECT  120000.0 1168050.0 121200.0 1166850.0 ;
      RECT  120000.0 1168050.0 121200.0 1166850.0 ;
      RECT  117600.0 1168050.0 118800.0 1166850.0 ;
      RECT  122400.0 1158150.0 123600.0 1156950.0 ;
      RECT  122400.0 1168050.0 123600.0 1166850.0 ;
      RECT  118200.0 1163400.0 119400.0 1162200.0 ;
      RECT  118200.0 1163400.0 119400.0 1162200.0 ;
      RECT  120750.0 1163250.0 121650.0 1162350.0 ;
      RECT  115800.0 1156050.0 125400.0 1155150.0 ;
      RECT  115800.0 1169850.0 125400.0 1168950.0 ;
      RECT  127200.0 1167450.0 128400.0 1169850.0 ;
      RECT  127200.0 1158750.0 128400.0 1155150.0 ;
      RECT  132000.0 1158750.0 133200.0 1155150.0 ;
      RECT  134400.0 1157550.0 135600.0 1155600.0 ;
      RECT  134400.0 1169400.0 135600.0 1167450.0 ;
      RECT  127200.0 1158750.0 128400.0 1157550.0 ;
      RECT  129600.0 1158750.0 130800.0 1157550.0 ;
      RECT  129600.0 1158750.0 130800.0 1157550.0 ;
      RECT  127200.0 1158750.0 128400.0 1157550.0 ;
      RECT  129600.0 1158750.0 130800.0 1157550.0 ;
      RECT  132000.0 1158750.0 133200.0 1157550.0 ;
      RECT  132000.0 1158750.0 133200.0 1157550.0 ;
      RECT  129600.0 1158750.0 130800.0 1157550.0 ;
      RECT  127200.0 1167450.0 128400.0 1166250.0 ;
      RECT  129600.0 1167450.0 130800.0 1166250.0 ;
      RECT  129600.0 1167450.0 130800.0 1166250.0 ;
      RECT  127200.0 1167450.0 128400.0 1166250.0 ;
      RECT  129600.0 1167450.0 130800.0 1166250.0 ;
      RECT  132000.0 1167450.0 133200.0 1166250.0 ;
      RECT  132000.0 1167450.0 133200.0 1166250.0 ;
      RECT  129600.0 1167450.0 130800.0 1166250.0 ;
      RECT  134400.0 1158150.0 135600.0 1156950.0 ;
      RECT  134400.0 1168050.0 135600.0 1166850.0 ;
      RECT  132000.0 1164900.0 130800.0 1163700.0 ;
      RECT  129000.0 1162200.0 127800.0 1161000.0 ;
      RECT  129600.0 1158750.0 130800.0 1157550.0 ;
      RECT  132000.0 1167450.0 133200.0 1166250.0 ;
      RECT  133200.0 1162200.0 132000.0 1161000.0 ;
      RECT  127800.0 1162200.0 129000.0 1161000.0 ;
      RECT  130800.0 1164900.0 132000.0 1163700.0 ;
      RECT  132000.0 1162200.0 133200.0 1161000.0 ;
      RECT  125400.0 1156050.0 139800.0 1155150.0 ;
      RECT  125400.0 1169850.0 139800.0 1168950.0 ;
      RECT  146400.0 1157550.0 147600.0 1155600.0 ;
      RECT  146400.0 1169400.0 147600.0 1167450.0 ;
      RECT  141600.0 1168050.0 142800.0 1169850.0 ;
      RECT  141600.0 1158750.0 142800.0 1155150.0 ;
      RECT  144300.0 1168050.0 145200.0 1158750.0 ;
      RECT  141600.0 1158750.0 142800.0 1157550.0 ;
      RECT  144000.0 1158750.0 145200.0 1157550.0 ;
      RECT  144000.0 1158750.0 145200.0 1157550.0 ;
      RECT  141600.0 1158750.0 142800.0 1157550.0 ;
      RECT  141600.0 1168050.0 142800.0 1166850.0 ;
      RECT  144000.0 1168050.0 145200.0 1166850.0 ;
      RECT  144000.0 1168050.0 145200.0 1166850.0 ;
      RECT  141600.0 1168050.0 142800.0 1166850.0 ;
      RECT  146400.0 1158150.0 147600.0 1156950.0 ;
      RECT  146400.0 1168050.0 147600.0 1166850.0 ;
      RECT  142200.0 1163400.0 143400.0 1162200.0 ;
      RECT  142200.0 1163400.0 143400.0 1162200.0 ;
      RECT  144750.0 1163250.0 145650.0 1162350.0 ;
      RECT  139800.0 1156050.0 149400.0 1155150.0 ;
      RECT  139800.0 1169850.0 149400.0 1168950.0 ;
      RECT  112050.0 1162200.0 113250.0 1163400.0 ;
      RECT  114000.0 1164600.0 115200.0 1165800.0 ;
      RECT  130800.0 1163700.0 129600.0 1164900.0 ;
      RECT  122400.0 1181250.0 123600.0 1183200.0 ;
      RECT  122400.0 1169400.0 123600.0 1171350.0 ;
      RECT  117600.0 1170750.0 118800.0 1168950.0 ;
      RECT  117600.0 1180050.0 118800.0 1183650.0 ;
      RECT  120300.0 1170750.0 121200.0 1180050.0 ;
      RECT  117600.0 1180050.0 118800.0 1181250.0 ;
      RECT  120000.0 1180050.0 121200.0 1181250.0 ;
      RECT  120000.0 1180050.0 121200.0 1181250.0 ;
      RECT  117600.0 1180050.0 118800.0 1181250.0 ;
      RECT  117600.0 1170750.0 118800.0 1171950.0 ;
      RECT  120000.0 1170750.0 121200.0 1171950.0 ;
      RECT  120000.0 1170750.0 121200.0 1171950.0 ;
      RECT  117600.0 1170750.0 118800.0 1171950.0 ;
      RECT  122400.0 1180650.0 123600.0 1181850.0 ;
      RECT  122400.0 1170750.0 123600.0 1171950.0 ;
      RECT  118200.0 1175400.0 119400.0 1176600.0 ;
      RECT  118200.0 1175400.0 119400.0 1176600.0 ;
      RECT  120750.0 1175550.0 121650.0 1176450.0 ;
      RECT  115800.0 1182750.0 125400.0 1183650.0 ;
      RECT  115800.0 1168950.0 125400.0 1169850.0 ;
      RECT  127200.0 1171350.0 128400.0 1168950.0 ;
      RECT  127200.0 1180050.0 128400.0 1183650.0 ;
      RECT  132000.0 1180050.0 133200.0 1183650.0 ;
      RECT  134400.0 1181250.0 135600.0 1183200.0 ;
      RECT  134400.0 1169400.0 135600.0 1171350.0 ;
      RECT  127200.0 1180050.0 128400.0 1181250.0 ;
      RECT  129600.0 1180050.0 130800.0 1181250.0 ;
      RECT  129600.0 1180050.0 130800.0 1181250.0 ;
      RECT  127200.0 1180050.0 128400.0 1181250.0 ;
      RECT  129600.0 1180050.0 130800.0 1181250.0 ;
      RECT  132000.0 1180050.0 133200.0 1181250.0 ;
      RECT  132000.0 1180050.0 133200.0 1181250.0 ;
      RECT  129600.0 1180050.0 130800.0 1181250.0 ;
      RECT  127200.0 1171350.0 128400.0 1172550.0 ;
      RECT  129600.0 1171350.0 130800.0 1172550.0 ;
      RECT  129600.0 1171350.0 130800.0 1172550.0 ;
      RECT  127200.0 1171350.0 128400.0 1172550.0 ;
      RECT  129600.0 1171350.0 130800.0 1172550.0 ;
      RECT  132000.0 1171350.0 133200.0 1172550.0 ;
      RECT  132000.0 1171350.0 133200.0 1172550.0 ;
      RECT  129600.0 1171350.0 130800.0 1172550.0 ;
      RECT  134400.0 1180650.0 135600.0 1181850.0 ;
      RECT  134400.0 1170750.0 135600.0 1171950.0 ;
      RECT  132000.0 1173900.0 130800.0 1175100.0 ;
      RECT  129000.0 1176600.0 127800.0 1177800.0 ;
      RECT  129600.0 1180050.0 130800.0 1181250.0 ;
      RECT  132000.0 1171350.0 133200.0 1172550.0 ;
      RECT  133200.0 1176600.0 132000.0 1177800.0 ;
      RECT  127800.0 1176600.0 129000.0 1177800.0 ;
      RECT  130800.0 1173900.0 132000.0 1175100.0 ;
      RECT  132000.0 1176600.0 133200.0 1177800.0 ;
      RECT  125400.0 1182750.0 139800.0 1183650.0 ;
      RECT  125400.0 1168950.0 139800.0 1169850.0 ;
      RECT  146400.0 1181250.0 147600.0 1183200.0 ;
      RECT  146400.0 1169400.0 147600.0 1171350.0 ;
      RECT  141600.0 1170750.0 142800.0 1168950.0 ;
      RECT  141600.0 1180050.0 142800.0 1183650.0 ;
      RECT  144300.0 1170750.0 145200.0 1180050.0 ;
      RECT  141600.0 1180050.0 142800.0 1181250.0 ;
      RECT  144000.0 1180050.0 145200.0 1181250.0 ;
      RECT  144000.0 1180050.0 145200.0 1181250.0 ;
      RECT  141600.0 1180050.0 142800.0 1181250.0 ;
      RECT  141600.0 1170750.0 142800.0 1171950.0 ;
      RECT  144000.0 1170750.0 145200.0 1171950.0 ;
      RECT  144000.0 1170750.0 145200.0 1171950.0 ;
      RECT  141600.0 1170750.0 142800.0 1171950.0 ;
      RECT  146400.0 1180650.0 147600.0 1181850.0 ;
      RECT  146400.0 1170750.0 147600.0 1171950.0 ;
      RECT  142200.0 1175400.0 143400.0 1176600.0 ;
      RECT  142200.0 1175400.0 143400.0 1176600.0 ;
      RECT  144750.0 1175550.0 145650.0 1176450.0 ;
      RECT  139800.0 1182750.0 149400.0 1183650.0 ;
      RECT  139800.0 1168950.0 149400.0 1169850.0 ;
      RECT  112050.0 1175400.0 113250.0 1176600.0 ;
      RECT  114000.0 1173000.0 115200.0 1174200.0 ;
      RECT  130800.0 1173900.0 129600.0 1175100.0 ;
      RECT  122400.0 1185150.0 123600.0 1183200.0 ;
      RECT  122400.0 1197000.0 123600.0 1195050.0 ;
      RECT  117600.0 1195650.0 118800.0 1197450.0 ;
      RECT  117600.0 1186350.0 118800.0 1182750.0 ;
      RECT  120300.0 1195650.0 121200.0 1186350.0 ;
      RECT  117600.0 1186350.0 118800.0 1185150.0 ;
      RECT  120000.0 1186350.0 121200.0 1185150.0 ;
      RECT  120000.0 1186350.0 121200.0 1185150.0 ;
      RECT  117600.0 1186350.0 118800.0 1185150.0 ;
      RECT  117600.0 1195650.0 118800.0 1194450.0 ;
      RECT  120000.0 1195650.0 121200.0 1194450.0 ;
      RECT  120000.0 1195650.0 121200.0 1194450.0 ;
      RECT  117600.0 1195650.0 118800.0 1194450.0 ;
      RECT  122400.0 1185750.0 123600.0 1184550.0 ;
      RECT  122400.0 1195650.0 123600.0 1194450.0 ;
      RECT  118200.0 1191000.0 119400.0 1189800.0 ;
      RECT  118200.0 1191000.0 119400.0 1189800.0 ;
      RECT  120750.0 1190850.0 121650.0 1189950.0 ;
      RECT  115800.0 1183650.0 125400.0 1182750.0 ;
      RECT  115800.0 1197450.0 125400.0 1196550.0 ;
      RECT  127200.0 1195050.0 128400.0 1197450.0 ;
      RECT  127200.0 1186350.0 128400.0 1182750.0 ;
      RECT  132000.0 1186350.0 133200.0 1182750.0 ;
      RECT  134400.0 1185150.0 135600.0 1183200.0 ;
      RECT  134400.0 1197000.0 135600.0 1195050.0 ;
      RECT  127200.0 1186350.0 128400.0 1185150.0 ;
      RECT  129600.0 1186350.0 130800.0 1185150.0 ;
      RECT  129600.0 1186350.0 130800.0 1185150.0 ;
      RECT  127200.0 1186350.0 128400.0 1185150.0 ;
      RECT  129600.0 1186350.0 130800.0 1185150.0 ;
      RECT  132000.0 1186350.0 133200.0 1185150.0 ;
      RECT  132000.0 1186350.0 133200.0 1185150.0 ;
      RECT  129600.0 1186350.0 130800.0 1185150.0 ;
      RECT  127200.0 1195050.0 128400.0 1193850.0 ;
      RECT  129600.0 1195050.0 130800.0 1193850.0 ;
      RECT  129600.0 1195050.0 130800.0 1193850.0 ;
      RECT  127200.0 1195050.0 128400.0 1193850.0 ;
      RECT  129600.0 1195050.0 130800.0 1193850.0 ;
      RECT  132000.0 1195050.0 133200.0 1193850.0 ;
      RECT  132000.0 1195050.0 133200.0 1193850.0 ;
      RECT  129600.0 1195050.0 130800.0 1193850.0 ;
      RECT  134400.0 1185750.0 135600.0 1184550.0 ;
      RECT  134400.0 1195650.0 135600.0 1194450.0 ;
      RECT  132000.0 1192500.0 130800.0 1191300.0 ;
      RECT  129000.0 1189800.0 127800.0 1188600.0 ;
      RECT  129600.0 1186350.0 130800.0 1185150.0 ;
      RECT  132000.0 1195050.0 133200.0 1193850.0 ;
      RECT  133200.0 1189800.0 132000.0 1188600.0 ;
      RECT  127800.0 1189800.0 129000.0 1188600.0 ;
      RECT  130800.0 1192500.0 132000.0 1191300.0 ;
      RECT  132000.0 1189800.0 133200.0 1188600.0 ;
      RECT  125400.0 1183650.0 139800.0 1182750.0 ;
      RECT  125400.0 1197450.0 139800.0 1196550.0 ;
      RECT  146400.0 1185150.0 147600.0 1183200.0 ;
      RECT  146400.0 1197000.0 147600.0 1195050.0 ;
      RECT  141600.0 1195650.0 142800.0 1197450.0 ;
      RECT  141600.0 1186350.0 142800.0 1182750.0 ;
      RECT  144300.0 1195650.0 145200.0 1186350.0 ;
      RECT  141600.0 1186350.0 142800.0 1185150.0 ;
      RECT  144000.0 1186350.0 145200.0 1185150.0 ;
      RECT  144000.0 1186350.0 145200.0 1185150.0 ;
      RECT  141600.0 1186350.0 142800.0 1185150.0 ;
      RECT  141600.0 1195650.0 142800.0 1194450.0 ;
      RECT  144000.0 1195650.0 145200.0 1194450.0 ;
      RECT  144000.0 1195650.0 145200.0 1194450.0 ;
      RECT  141600.0 1195650.0 142800.0 1194450.0 ;
      RECT  146400.0 1185750.0 147600.0 1184550.0 ;
      RECT  146400.0 1195650.0 147600.0 1194450.0 ;
      RECT  142200.0 1191000.0 143400.0 1189800.0 ;
      RECT  142200.0 1191000.0 143400.0 1189800.0 ;
      RECT  144750.0 1190850.0 145650.0 1189950.0 ;
      RECT  139800.0 1183650.0 149400.0 1182750.0 ;
      RECT  139800.0 1197450.0 149400.0 1196550.0 ;
      RECT  112050.0 1189800.0 113250.0 1191000.0 ;
      RECT  114000.0 1192200.0 115200.0 1193400.0 ;
      RECT  130800.0 1191300.0 129600.0 1192500.0 ;
      RECT  109500.0 317550.0 114600.0 318450.0 ;
      RECT  109500.0 336750.0 114600.0 337650.0 ;
      RECT  109500.0 345150.0 114600.0 346050.0 ;
      RECT  109500.0 364350.0 114600.0 365250.0 ;
      RECT  109500.0 372750.0 114600.0 373650.0 ;
      RECT  109500.0 391950.0 114600.0 392850.0 ;
      RECT  109500.0 400350.0 114600.0 401250.0 ;
      RECT  109500.0 419550.0 114600.0 420450.0 ;
      RECT  109500.0 427950.0 114600.0 428850.0 ;
      RECT  109500.0 447150.0 114600.0 448050.0 ;
      RECT  109500.0 455550.0 114600.0 456450.0 ;
      RECT  109500.0 474750.0 114600.0 475650.0 ;
      RECT  109500.0 483150.0 114600.0 484050.0 ;
      RECT  109500.0 502350.0 114600.0 503250.0 ;
      RECT  109500.0 510750.0 114600.0 511650.0 ;
      RECT  109500.0 529950.0 114600.0 530850.0 ;
      RECT  109500.0 538350.0 114600.0 539250.0 ;
      RECT  109500.0 557550.0 114600.0 558450.0 ;
      RECT  109500.0 565950.0 114600.0 566850.0 ;
      RECT  109500.0 585150.0 114600.0 586050.0 ;
      RECT  109500.0 593550.0 114600.0 594450.0 ;
      RECT  109500.0 612750.0 114600.0 613650.0 ;
      RECT  109500.0 621150.0 114600.0 622050.0 ;
      RECT  109500.0 640350.0 114600.0 641250.0 ;
      RECT  109500.0 648750.0 114600.0 649650.0 ;
      RECT  109500.0 667950.0 114600.0 668850.0 ;
      RECT  109500.0 676350.0 114600.0 677250.0 ;
      RECT  109500.0 695550.0 114600.0 696450.0 ;
      RECT  109500.0 703950.0 114600.0 704850.0 ;
      RECT  109500.0 723150.0 114600.0 724050.0 ;
      RECT  109500.0 731550.0 114600.0 732450.0 ;
      RECT  109500.0 750750.0 114600.0 751650.0 ;
      RECT  109500.0 759150.0 114600.0 760050.0 ;
      RECT  109500.0 778350.0 114600.0 779250.0 ;
      RECT  109500.0 786750.0 114600.0 787650.0 ;
      RECT  109500.0 805950.0 114600.0 806850.0 ;
      RECT  109500.0 814350.0 114600.0 815250.0 ;
      RECT  109500.0 833550.0 114600.0 834450.0 ;
      RECT  109500.0 841950.0 114600.0 842850.0 ;
      RECT  109500.0 861150.0 114600.0 862050.0 ;
      RECT  109500.0 869550.0 114600.0 870450.0 ;
      RECT  109500.0 888750.0 114600.0 889650.0 ;
      RECT  109500.0 897150.0 114600.0 898050.0 ;
      RECT  109500.0 916350.0 114600.0 917250.0 ;
      RECT  109500.0 924750.0 114600.0 925650.0 ;
      RECT  109500.0 943950.0 114600.0 944850.0 ;
      RECT  109500.0 952350.0 114600.0 953250.0 ;
      RECT  109500.0 971550.0 114600.0 972450.0 ;
      RECT  109500.0 979950.0 114600.0 980850.0 ;
      RECT  109500.0 999150.0 114600.0 1000050.0 ;
      RECT  109500.0 1007550.0 114600.0 1008450.0 ;
      RECT  109500.0 1026750.0 114600.0 1027650.0 ;
      RECT  109500.0 1035150.0 114600.0 1036050.0 ;
      RECT  109500.0 1054350.0 114600.0 1055250.0 ;
      RECT  109500.0 1062750.0 114600.0 1063650.0 ;
      RECT  109500.0 1081950.0 114600.0 1082850.0 ;
      RECT  109500.0 1090350.0 114600.0 1091250.0 ;
      RECT  109500.0 1109550.0 114600.0 1110450.0 ;
      RECT  109500.0 1117950.0 114600.0 1118850.0 ;
      RECT  109500.0 1137150.0 114600.0 1138050.0 ;
      RECT  109500.0 1145550.0 114600.0 1146450.0 ;
      RECT  109500.0 1164750.0 114600.0 1165650.0 ;
      RECT  109500.0 1173150.0 114600.0 1174050.0 ;
      RECT  109500.0 1192350.0 114600.0 1193250.0 ;
      RECT  144750.0 319950.0 145650.0 320850.0 ;
      RECT  144750.0 334350.0 145650.0 335250.0 ;
      RECT  144750.0 347550.0 145650.0 348450.0 ;
      RECT  144750.0 361950.0 145650.0 362850.0 ;
      RECT  144750.0 375150.0 145650.0 376050.0 ;
      RECT  144750.0 389550.0 145650.0 390450.0 ;
      RECT  144750.0 402750.0 145650.0 403650.0 ;
      RECT  144750.0 417150.0 145650.0 418050.0 ;
      RECT  144750.0 430350.0 145650.0 431250.0 ;
      RECT  144750.0 444750.0 145650.0 445650.0 ;
      RECT  144750.0 457950.0 145650.0 458850.0 ;
      RECT  144750.0 472350.0 145650.0 473250.0 ;
      RECT  144750.0 485550.0 145650.0 486450.0 ;
      RECT  144750.0 499950.0 145650.0 500850.0 ;
      RECT  144750.0 513150.0 145650.0 514050.0 ;
      RECT  144750.0 527550.0 145650.0 528450.0 ;
      RECT  144750.0 540750.0 145650.0 541650.0 ;
      RECT  144750.0 555150.0 145650.0 556050.0 ;
      RECT  144750.0 568350.0 145650.0 569250.0 ;
      RECT  144750.0 582750.0 145650.0 583650.0 ;
      RECT  144750.0 595950.0 145650.0 596850.0 ;
      RECT  144750.0 610350.0 145650.0 611250.0 ;
      RECT  144750.0 623550.0 145650.0 624450.0 ;
      RECT  144750.0 637950.0 145650.0 638850.0 ;
      RECT  144750.0 651150.0 145650.0 652050.0 ;
      RECT  144750.0 665550.0 145650.0 666450.0 ;
      RECT  144750.0 678750.0 145650.0 679650.0 ;
      RECT  144750.0 693150.0 145650.0 694050.0 ;
      RECT  144750.0 706350.0 145650.0 707250.0 ;
      RECT  144750.0 720750.0 145650.0 721650.0 ;
      RECT  144750.0 733950.0 145650.0 734850.0 ;
      RECT  144750.0 748350.0 145650.0 749250.0 ;
      RECT  144750.0 761550.0 145650.0 762450.0 ;
      RECT  144750.0 775950.0 145650.0 776850.0 ;
      RECT  144750.0 789150.0 145650.0 790050.0 ;
      RECT  144750.0 803550.0 145650.0 804450.0 ;
      RECT  144750.0 816750.0 145650.0 817650.0 ;
      RECT  144750.0 831150.0 145650.0 832050.0 ;
      RECT  144750.0 844350.0 145650.0 845250.0 ;
      RECT  144750.0 858750.0 145650.0 859650.0 ;
      RECT  144750.0 871950.0 145650.0 872850.0 ;
      RECT  144750.0 886350.0 145650.0 887250.0 ;
      RECT  144750.0 899550.0 145650.0 900450.0 ;
      RECT  144750.0 913950.0 145650.0 914850.0 ;
      RECT  144750.0 927150.0 145650.0 928050.0 ;
      RECT  144750.0 941550.0 145650.0 942450.0 ;
      RECT  144750.0 954750.0 145650.0 955650.0 ;
      RECT  144750.0 969150.0 145650.0 970050.0 ;
      RECT  144750.0 982350.0 145650.0 983250.0 ;
      RECT  144750.0 996750.0 145650.0 997650.0 ;
      RECT  144750.0 1009950.0 145650.0 1010850.0 ;
      RECT  144750.0 1024350.0 145650.0 1025250.0 ;
      RECT  144750.0 1037550.0 145650.0 1038450.0 ;
      RECT  144750.0 1051950.0 145650.0 1052850.0 ;
      RECT  144750.0 1065150.0 145650.0 1066050.0 ;
      RECT  144750.0 1079550.0 145650.0 1080450.0 ;
      RECT  144750.0 1092750.0 145650.0 1093650.0 ;
      RECT  144750.0 1107150.0 145650.0 1108050.0 ;
      RECT  144750.0 1120350.0 145650.0 1121250.0 ;
      RECT  144750.0 1134750.0 145650.0 1135650.0 ;
      RECT  144750.0 1147950.0 145650.0 1148850.0 ;
      RECT  144750.0 1162350.0 145650.0 1163250.0 ;
      RECT  144750.0 1175550.0 145650.0 1176450.0 ;
      RECT  144750.0 1189950.0 145650.0 1190850.0 ;
      RECT  109500.0 327150.0 115800.0 328050.0 ;
      RECT  109500.0 354750.0 115800.0 355650.0 ;
      RECT  109500.0 382350.0 115800.0 383250.0 ;
      RECT  109500.0 409950.0 115800.0 410850.0 ;
      RECT  109500.0 437550.0 115800.0 438450.0 ;
      RECT  109500.0 465150.0 115800.0 466050.0 ;
      RECT  109500.0 492750.0 115800.0 493650.0 ;
      RECT  109500.0 520350.0 115800.0 521250.0 ;
      RECT  109500.0 547950.0 115800.0 548850.0 ;
      RECT  109500.0 575550.0 115800.0 576450.0 ;
      RECT  109500.0 603150.0 115800.0 604050.0 ;
      RECT  109500.0 630750.0 115800.0 631650.0 ;
      RECT  109500.0 658350.0 115800.0 659250.0 ;
      RECT  109500.0 685950.0 115800.0 686850.0 ;
      RECT  109500.0 713550.0 115800.0 714450.0 ;
      RECT  109500.0 741150.0 115800.0 742050.0 ;
      RECT  109500.0 768750.0 115800.0 769650.0 ;
      RECT  109500.0 796350.0 115800.0 797250.0 ;
      RECT  109500.0 823950.0 115800.0 824850.0 ;
      RECT  109500.0 851550.0 115800.0 852450.0 ;
      RECT  109500.0 879150.0 115800.0 880050.0 ;
      RECT  109500.0 906750.0 115800.0 907650.0 ;
      RECT  109500.0 934350.0 115800.0 935250.0 ;
      RECT  109500.0 961950.0 115800.0 962850.0 ;
      RECT  109500.0 989550.0 115800.0 990450.0 ;
      RECT  109500.0 1017150.0 115800.0 1018050.0 ;
      RECT  109500.0 1044750.0 115800.0 1045650.0 ;
      RECT  109500.0 1072350.0 115800.0 1073250.0 ;
      RECT  109500.0 1099950.0 115800.0 1100850.0 ;
      RECT  109500.0 1127550.0 115800.0 1128450.0 ;
      RECT  109500.0 1155150.0 115800.0 1156050.0 ;
      RECT  109500.0 1182750.0 115800.0 1183650.0 ;
      RECT  109500.0 313350.0 115800.0 314250.0 ;
      RECT  109500.0 340950.0 115800.0 341850.0 ;
      RECT  109500.0 368550.0 115800.0 369450.0 ;
      RECT  109500.0 396150.0 115800.0 397050.0 ;
      RECT  109500.0 423750.0 115800.0 424650.0 ;
      RECT  109500.0 451350.0 115800.0 452250.0 ;
      RECT  109500.0 478950.0 115800.0 479850.0 ;
      RECT  109500.0 506550.0 115800.0 507450.0 ;
      RECT  109500.0 534150.0 115800.0 535050.0 ;
      RECT  109500.0 561750.0 115800.0 562650.0 ;
      RECT  109500.0 589350.0 115800.0 590250.0 ;
      RECT  109500.0 616950.0 115800.0 617850.0 ;
      RECT  109500.0 644550.0 115800.0 645450.0 ;
      RECT  109500.0 672150.0 115800.0 673050.0 ;
      RECT  109500.0 699750.0 115800.0 700650.0 ;
      RECT  109500.0 727350.0 115800.0 728250.0 ;
      RECT  109500.0 754950.0 115800.0 755850.0 ;
      RECT  109500.0 782550.0 115800.0 783450.0 ;
      RECT  109500.0 810150.0 115800.0 811050.0 ;
      RECT  109500.0 837750.0 115800.0 838650.0 ;
      RECT  109500.0 865350.0 115800.0 866250.0 ;
      RECT  109500.0 892950.0 115800.0 893850.0 ;
      RECT  109500.0 920550.0 115800.0 921450.0 ;
      RECT  109500.0 948150.0 115800.0 949050.0 ;
      RECT  109500.0 975750.0 115800.0 976650.0 ;
      RECT  109500.0 1003350.0 115800.0 1004250.0 ;
      RECT  109500.0 1030950.0 115800.0 1031850.0 ;
      RECT  109500.0 1058550.0 115800.0 1059450.0 ;
      RECT  109500.0 1086150.0 115800.0 1087050.0 ;
      RECT  109500.0 1113750.0 115800.0 1114650.0 ;
      RECT  109500.0 1141350.0 115800.0 1142250.0 ;
      RECT  109500.0 1168950.0 115800.0 1169850.0 ;
      RECT  109500.0 1196550.0 115800.0 1197450.0 ;
      RECT  59100.0 142800.0 119100.0 132600.0 ;
      RECT  59100.0 122400.0 119100.0 132600.0 ;
      RECT  59100.0 122400.0 119100.0 112200.0 ;
      RECT  59100.0 102000.0 119100.0 112200.0 ;
      RECT  59100.0 102000.0 119100.0 91800.0 ;
      RECT  59100.0 81600.0 119100.0 91800.0 ;
      RECT  59100.0 81600.0 119100.0 71400.0 ;
      RECT  59100.0 61200.0 119100.0 71400.0 ;
      RECT  61500.0 142800.0 62400.0 61200.0 ;
      RECT  115500.0 142800.0 116400.0 61200.0 ;
      RECT  172650.0 314400.0 173850.0 313200.0 ;
      RECT  172650.0 342000.0 173850.0 340800.0 ;
      RECT  172650.0 369600.0 173850.0 368400.0 ;
      RECT  172650.0 397200.0 173850.0 396000.0 ;
      RECT  172650.0 424800.0 173850.0 423600.0 ;
      RECT  172650.0 452400.0 173850.0 451200.0 ;
      RECT  172650.0 480000.0 173850.0 478800.0 ;
      RECT  172650.0 507600.0 173850.0 506400.0 ;
      RECT  172650.0 535200.0 173850.0 534000.0 ;
      RECT  172650.0 562800.0 173850.0 561600.0 ;
      RECT  172650.0 590400.0 173850.0 589200.0 ;
      RECT  172650.0 618000.0 173850.0 616800.0 ;
      RECT  172650.0 645600.0 173850.0 644400.0 ;
      RECT  172650.0 673200.0 173850.0 672000.0 ;
      RECT  172650.0 700800.0 173850.0 699600.0 ;
      RECT  172650.0 728400.0 173850.0 727200.0 ;
      RECT  172650.0 756000.0 173850.0 754800.0 ;
      RECT  172650.0 783600.0 173850.0 782400.0 ;
      RECT  172650.0 811200.0 173850.0 810000.0 ;
      RECT  172650.0 838800.0 173850.0 837600.0 ;
      RECT  172650.0 866400.0 173850.0 865200.0 ;
      RECT  172650.0 894000.0 173850.0 892800.0 ;
      RECT  172650.0 921600.0 173850.0 920400.0 ;
      RECT  172650.0 949200.0 173850.0 948000.0 ;
      RECT  172650.0 976800.0 173850.0 975600.0 ;
      RECT  172650.0 1004400.0 173850.0 1003200.0 ;
      RECT  172650.0 1032000.0 173850.0 1030800.0 ;
      RECT  172650.0 1059600.0 173850.0 1058400.0 ;
      RECT  172650.0 1087200.0 173850.0 1086000.0 ;
      RECT  172650.0 1114800.0 173850.0 1113600.0 ;
      RECT  172650.0 1142400.0 173850.0 1141200.0 ;
      RECT  172650.0 1170000.0 173850.0 1168800.0 ;
      RECT  172650.0 1197600.0 173850.0 1196400.0 ;
      RECT  138900.0 150450.0 137700.0 151650.0 ;
      RECT  144000.0 150300.0 142800.0 151500.0 ;
      RECT  135900.0 164250.0 134700.0 165450.0 ;
      RECT  146700.0 164100.0 145500.0 165300.0 ;
      RECT  138900.0 205650.0 137700.0 206850.0 ;
      RECT  149400.0 205500.0 148200.0 206700.0 ;
      RECT  135900.0 219450.0 134700.0 220650.0 ;
      RECT  152100.0 219300.0 150900.0 220500.0 ;
      RECT  138900.0 260850.0 137700.0 262050.0 ;
      RECT  154800.0 260700.0 153600.0 261900.0 ;
      RECT  135900.0 274650.0 134700.0 275850.0 ;
      RECT  157500.0 274500.0 156300.0 275700.0 ;
      RECT  141000.0 147600.0 139800.0 148800.0 ;
      RECT  141000.0 175200.0 139800.0 176400.0 ;
      RECT  141000.0 202800.0 139800.0 204000.0 ;
      RECT  141000.0 230400.0 139800.0 231600.0 ;
      RECT  141000.0 258000.0 139800.0 259200.0 ;
      RECT  141000.0 285600.0 139800.0 286800.0 ;
      RECT  160200.0 285750.0 159000.0 286950.0 ;
      RECT  162900.0 283650.0 161700.0 284850.0 ;
      RECT  165600.0 281550.0 164400.0 282750.0 ;
      RECT  168300.0 279450.0 167100.0 280650.0 ;
      RECT  160200.0 6600.0 159000.0 7800.0 ;
      RECT  162900.0 21000.0 161700.0 22200.0 ;
      RECT  165600.0 34200.0 164400.0 35400.0 ;
      RECT  168300.0 48600.0 167100.0 49800.0 ;
      RECT  172650.0 1200.0 173850.0 -1.15463194561e-11 ;
      RECT  172650.0 28800.0 173850.0 27600.0 ;
      RECT  172650.0 56400.0 173850.0 55200.0 ;
      RECT  118500.0 136350.0 117300.0 137550.0 ;
      RECT  144000.0 136350.0 142800.0 137550.0 ;
      RECT  118500.0 127650.0 117300.0 128850.0 ;
      RECT  146700.0 127650.0 145500.0 128850.0 ;
      RECT  118500.0 115950.0 117300.0 117150.0 ;
      RECT  149400.0 115950.0 148200.0 117150.0 ;
      RECT  118500.0 107250.0 117300.0 108450.0 ;
      RECT  152100.0 107250.0 150900.0 108450.0 ;
      RECT  118500.0 95550.0 117300.0 96750.0 ;
      RECT  154800.0 95550.0 153600.0 96750.0 ;
      RECT  118500.0 86850.0 117300.0 88050.0 ;
      RECT  157500.0 86850.0 156300.0 88050.0 ;
      RECT  120300.0 132000.0 119100.0 133200.0 ;
      RECT  173850.0 132150.0 172650.0 133350.0 ;
      RECT  120300.0 111600.0 119100.0 112800.0 ;
      RECT  173850.0 111750.0 172650.0 112950.0 ;
      RECT  120300.0 91200.0 119100.0 92400.0 ;
      RECT  173850.0 91350.0 172650.0 92550.0 ;
      RECT  120300.0 70800.0 119100.0 72000.0 ;
      RECT  173850.0 70950.0 172650.0 72150.0 ;
      RECT  189000.0 105900.0 187800.0 107100.0 ;
      RECT  183600.0 101400.0 182400.0 102600.0 ;
      RECT  186300.0 99000.0 185100.0 100200.0 ;
      RECT  189000.0 1205250.0 187800.0 1206450.0 ;
      RECT  191700.0 170700.0 190500.0 171900.0 ;
      RECT  194400.0 268800.0 193200.0 270000.0 ;
      RECT  180900.0 144300.0 179700.0 145500.0 ;
      RECT  113250.0 1198500.0 112050.0 1199700.0 ;
      RECT  180900.0 1198500.0 179700.0 1199700.0 ;
      RECT  177150.0 97050.0 175950.0 98250.0 ;
      RECT  177150.0 266850.0 175950.0 268050.0 ;
      RECT  177150.0 168750.0 175950.0 169950.0 ;
      RECT  529200.0 600.0 533700.0 1217400.0 ;
      RECT  52800.0 600.0 57300.0 1217400.0 ;
      RECT  43650.0 322200.0 42750.0 331800.0 ;
      RECT  43800.0 338400.0 42900.0 339300.0 ;
      RECT  43350.0 338400.0 43200.0 339300.0 ;
      RECT  43800.0 338850.0 42900.0 346200.0 ;
      RECT  43800.0 358050.0 42900.0 365400.0 ;
      RECT  35550.0 373200.0 30600.0 374100.0 ;
      RECT  43650.0 321750.0 42750.0 322650.0 ;
      RECT  43650.0 338400.0 42750.0 339300.0 ;
      RECT  29250.0 476700.0 28350.0 490050.0 ;
      RECT  43800.0 387300.0 42900.0 399450.0 ;
      RECT  33300.0 319200.0 30600.0 320100.0 ;
      RECT  29700.0 399450.0 28800.0 426300.0 ;
      RECT  27000.0 404850.0 26100.0 429300.0 ;
      RECT  41700.0 418350.0 40800.0 426900.0 ;
      RECT  43650.0 415650.0 42750.0 429300.0 ;
      RECT  45600.0 407550.0 44700.0 431700.0 ;
      RECT  41700.0 441450.0 40800.0 442350.0 ;
      RECT  41700.0 432900.0 40800.0 441900.0 ;
      RECT  43200.0 441450.0 41250.0 442350.0 ;
      RECT  43800.0 443850.0 42900.0 444750.0 ;
      RECT  43350.0 443850.0 43200.0 444750.0 ;
      RECT  43800.0 444300.0 42900.0 501900.0 ;
      RECT  14100.0 418350.0 13200.0 436500.0 ;
      RECT  16050.0 407550.0 15150.0 438900.0 ;
      RECT  18000.0 410250.0 17100.0 441300.0 ;
      RECT  14100.0 451050.0 13200.0 451950.0 ;
      RECT  14100.0 442500.0 13200.0 451500.0 ;
      RECT  15600.0 451050.0 13650.0 451950.0 ;
      RECT  16050.0 453900.0 15150.0 461100.0 ;
      RECT  16050.0 463500.0 15150.0 470700.0 ;
      RECT  29250.0 476250.0 28350.0 477150.0 ;
      RECT  28800.0 476250.0 28350.0 477150.0 ;
      RECT  29250.0 474300.0 28350.0 476700.0 ;
      RECT  29250.0 464100.0 28350.0 471300.0 ;
      RECT  29700.0 431400.0 28800.0 437700.0 ;
      RECT  30450.0 447600.0 29550.0 454800.0 ;
      RECT  16050.0 473100.0 15150.0 477300.0 ;
      RECT  29250.0 457500.0 28350.0 461700.0 ;
      RECT  50250.0 316800.0 49350.0 476700.0 ;
      RECT  50250.0 402150.0 49350.0 423300.0 ;
      RECT  36450.0 316800.0 35550.0 476700.0 ;
      RECT  36450.0 412950.0 35550.0 423300.0 ;
      RECT  22650.0 423300.0 21750.0 476700.0 ;
      RECT  22650.0 402150.0 21750.0 423300.0 ;
      RECT  8850.0 423300.0 7950.0 476700.0 ;
      RECT  8850.0 412950.0 7950.0 423300.0 ;
      RECT  8850.0 476250.0 7950.0 477150.0 ;
      RECT  8850.0 474600.0 7950.0 476700.0 ;
      RECT  8400.0 476250.0 3600.0 477150.0 ;
      RECT  7.1054273576e-12 316800.0 10200.0 376800.0 ;
      RECT  20400.0 316800.0 10200.0 376800.0 ;
      RECT  20400.0 316800.0 30600.0 376800.0 ;
      RECT  7.1054273576e-12 319200.0 30600.0 320100.0 ;
      RECT  1.42108547152e-11 373200.0 30600.0 374100.0 ;
      RECT  37950.0 325800.0 36000.0 327000.0 ;
      RECT  49800.0 325800.0 47850.0 327000.0 ;
      RECT  48450.0 321300.0 39150.0 322200.0 ;
      RECT  38550.0 318750.0 36600.0 319650.0 ;
      RECT  38550.0 323550.0 36600.0 324450.0 ;
      RECT  39150.0 318600.0 37950.0 319800.0 ;
      RECT  39150.0 323400.0 37950.0 324600.0 ;
      RECT  39150.0 321000.0 37950.0 322200.0 ;
      RECT  39150.0 321000.0 37950.0 322200.0 ;
      RECT  37050.0 318750.0 36150.0 324450.0 ;
      RECT  49800.0 318750.0 47850.0 319650.0 ;
      RECT  49800.0 323550.0 47850.0 324450.0 ;
      RECT  48450.0 318600.0 47250.0 319800.0 ;
      RECT  48450.0 323400.0 47250.0 324600.0 ;
      RECT  48450.0 321000.0 47250.0 322200.0 ;
      RECT  48450.0 321000.0 47250.0 322200.0 ;
      RECT  50250.0 318750.0 49350.0 324450.0 ;
      RECT  38550.0 325800.0 37350.0 327000.0 ;
      RECT  48450.0 325800.0 47250.0 327000.0 ;
      RECT  43800.0 319200.0 42600.0 320400.0 ;
      RECT  43800.0 319200.0 42600.0 320400.0 ;
      RECT  43650.0 321750.0 42750.0 322650.0 ;
      RECT  36450.0 316800.0 35550.0 328800.0 ;
      RECT  50250.0 316800.0 49350.0 328800.0 ;
      RECT  37950.0 340200.0 36000.0 341400.0 ;
      RECT  49800.0 340200.0 47850.0 341400.0 ;
      RECT  37350.0 330750.0 35550.0 336450.0 ;
      RECT  46050.0 337950.0 41250.0 338850.0 ;
      RECT  38850.0 330750.0 36900.0 331650.0 ;
      RECT  38850.0 335550.0 36900.0 336450.0 ;
      RECT  40800.0 333150.0 38850.0 334050.0 ;
      RECT  40800.0 337950.0 38850.0 338850.0 ;
      RECT  39450.0 330600.0 38250.0 331800.0 ;
      RECT  39450.0 335400.0 38250.0 336600.0 ;
      RECT  39450.0 333000.0 38250.0 334200.0 ;
      RECT  39450.0 337800.0 38250.0 339000.0 ;
      RECT  41250.0 333150.0 40350.0 338850.0 ;
      RECT  37350.0 330750.0 36450.0 336450.0 ;
      RECT  49500.0 330750.0 47550.0 331650.0 ;
      RECT  49500.0 335550.0 47550.0 336450.0 ;
      RECT  47550.0 333150.0 45600.0 334050.0 ;
      RECT  47550.0 337950.0 45600.0 338850.0 ;
      RECT  48150.0 330600.0 46950.0 331800.0 ;
      RECT  48150.0 335400.0 46950.0 336600.0 ;
      RECT  48150.0 333000.0 46950.0 334200.0 ;
      RECT  48150.0 337800.0 46950.0 339000.0 ;
      RECT  46050.0 333150.0 45150.0 338850.0 ;
      RECT  49950.0 330750.0 49050.0 336450.0 ;
      RECT  38550.0 340200.0 37350.0 341400.0 ;
      RECT  48450.0 340200.0 47250.0 341400.0 ;
      RECT  43800.0 331200.0 42600.0 332400.0 ;
      RECT  43800.0 331200.0 42600.0 332400.0 ;
      RECT  43650.0 338400.0 42750.0 339300.0 ;
      RECT  36450.0 328800.0 35550.0 343200.0 ;
      RECT  50250.0 328800.0 49350.0 343200.0 ;
      RECT  37950.0 359400.0 36000.0 360600.0 ;
      RECT  49800.0 359400.0 47850.0 360600.0 ;
      RECT  37800.0 345150.0 35550.0 355650.0 ;
      RECT  45900.0 357150.0 41700.0 358050.0 ;
      RECT  39300.0 345150.0 37350.0 346050.0 ;
      RECT  39300.0 349950.0 37350.0 350850.0 ;
      RECT  39300.0 354750.0 37350.0 355650.0 ;
      RECT  41250.0 347550.0 39300.0 348450.0 ;
      RECT  41250.0 352350.0 39300.0 353250.0 ;
      RECT  41250.0 357150.0 39300.0 358050.0 ;
      RECT  39900.0 345000.0 38700.0 346200.0 ;
      RECT  39900.0 349800.0 38700.0 351000.0 ;
      RECT  39900.0 354600.0 38700.0 355800.0 ;
      RECT  39900.0 347400.0 38700.0 348600.0 ;
      RECT  39900.0 352200.0 38700.0 353400.0 ;
      RECT  39900.0 357000.0 38700.0 358200.0 ;
      RECT  41700.0 347550.0 40800.0 358050.0 ;
      RECT  37800.0 345150.0 36900.0 355650.0 ;
      RECT  49350.0 345150.0 47400.0 346050.0 ;
      RECT  49350.0 349950.0 47400.0 350850.0 ;
      RECT  49350.0 354750.0 47400.0 355650.0 ;
      RECT  47400.0 347550.0 45450.0 348450.0 ;
      RECT  47400.0 352350.0 45450.0 353250.0 ;
      RECT  47400.0 357150.0 45450.0 358050.0 ;
      RECT  48000.0 345000.0 46800.0 346200.0 ;
      RECT  48000.0 349800.0 46800.0 351000.0 ;
      RECT  48000.0 354600.0 46800.0 355800.0 ;
      RECT  48000.0 347400.0 46800.0 348600.0 ;
      RECT  48000.0 352200.0 46800.0 353400.0 ;
      RECT  48000.0 357000.0 46800.0 358200.0 ;
      RECT  45900.0 347550.0 45000.0 358050.0 ;
      RECT  49800.0 345150.0 48900.0 355650.0 ;
      RECT  38550.0 359400.0 37350.0 360600.0 ;
      RECT  48450.0 359400.0 47250.0 360600.0 ;
      RECT  43950.0 345600.0 42750.0 346800.0 ;
      RECT  43950.0 345600.0 42750.0 346800.0 ;
      RECT  43800.0 357600.0 42900.0 358500.0 ;
      RECT  36450.0 343200.0 35550.0 362400.0 ;
      RECT  50250.0 343200.0 49350.0 362400.0 ;
      RECT  37950.0 390600.0 36000.0 391800.0 ;
      RECT  49800.0 390600.0 47850.0 391800.0 ;
      RECT  37800.0 364350.0 35550.0 389250.0 ;
      RECT  45900.0 385950.0 41700.0 386850.0 ;
      RECT  39300.0 364350.0 37350.0 365250.0 ;
      RECT  39300.0 369150.0 37350.0 370050.0 ;
      RECT  39300.0 373950.0 37350.0 374850.0 ;
      RECT  39300.0 378750.0 37350.0 379650.0 ;
      RECT  39300.0 383550.0 37350.0 384450.0 ;
      RECT  39300.0 388350.0 37350.0 389250.0 ;
      RECT  41250.0 366750.0 39300.0 367650.0 ;
      RECT  41250.0 371550.0 39300.0 372450.0 ;
      RECT  41250.0 376350.0 39300.0 377250.0 ;
      RECT  41250.0 381150.0 39300.0 382050.0 ;
      RECT  41250.0 385950.0 39300.0 386850.0 ;
      RECT  39900.0 364200.0 38700.0 365400.0 ;
      RECT  39900.0 369000.0 38700.0 370200.0 ;
      RECT  39900.0 373800.0 38700.0 375000.0 ;
      RECT  39900.0 378600.0 38700.0 379800.0 ;
      RECT  39900.0 383400.0 38700.0 384600.0 ;
      RECT  39900.0 388200.0 38700.0 389400.0 ;
      RECT  39900.0 366600.0 38700.0 367800.0 ;
      RECT  39900.0 371400.0 38700.0 372600.0 ;
      RECT  39900.0 376200.0 38700.0 377400.0 ;
      RECT  39900.0 381000.0 38700.0 382200.0 ;
      RECT  39900.0 385800.0 38700.0 387000.0 ;
      RECT  41700.0 366750.0 40800.0 386850.0 ;
      RECT  37800.0 364350.0 36900.0 389250.0 ;
      RECT  49350.0 364350.0 47400.0 365250.0 ;
      RECT  49350.0 369150.0 47400.0 370050.0 ;
      RECT  49350.0 373950.0 47400.0 374850.0 ;
      RECT  49350.0 378750.0 47400.0 379650.0 ;
      RECT  49350.0 383550.0 47400.0 384450.0 ;
      RECT  49350.0 388350.0 47400.0 389250.0 ;
      RECT  47400.0 366750.0 45450.0 367650.0 ;
      RECT  47400.0 371550.0 45450.0 372450.0 ;
      RECT  47400.0 376350.0 45450.0 377250.0 ;
      RECT  47400.0 381150.0 45450.0 382050.0 ;
      RECT  47400.0 385950.0 45450.0 386850.0 ;
      RECT  48000.0 364200.0 46800.0 365400.0 ;
      RECT  48000.0 369000.0 46800.0 370200.0 ;
      RECT  48000.0 373800.0 46800.0 375000.0 ;
      RECT  48000.0 378600.0 46800.0 379800.0 ;
      RECT  48000.0 383400.0 46800.0 384600.0 ;
      RECT  48000.0 388200.0 46800.0 389400.0 ;
      RECT  48000.0 366600.0 46800.0 367800.0 ;
      RECT  48000.0 371400.0 46800.0 372600.0 ;
      RECT  48000.0 376200.0 46800.0 377400.0 ;
      RECT  48000.0 381000.0 46800.0 382200.0 ;
      RECT  48000.0 385800.0 46800.0 387000.0 ;
      RECT  45900.0 366750.0 45000.0 386850.0 ;
      RECT  49800.0 364350.0 48900.0 389250.0 ;
      RECT  38550.0 390600.0 37350.0 391800.0 ;
      RECT  48450.0 390600.0 47250.0 391800.0 ;
      RECT  43950.0 364800.0 42750.0 366000.0 ;
      RECT  43950.0 364800.0 42750.0 366000.0 ;
      RECT  43800.0 386400.0 42900.0 387300.0 ;
      RECT  36450.0 362400.0 35550.0 393600.0 ;
      RECT  50250.0 362400.0 49350.0 393600.0 ;
      RECT  47850.0 425100.0 50250.0 426300.0 ;
      RECT  39150.0 425100.0 35550.0 426300.0 ;
      RECT  39150.0 429900.0 35550.0 431100.0 ;
      RECT  37950.0 434700.0 36000.0 435900.0 ;
      RECT  49800.0 434700.0 47850.0 435900.0 ;
      RECT  39150.0 425100.0 37950.0 426300.0 ;
      RECT  39150.0 427500.0 37950.0 428700.0 ;
      RECT  39150.0 427500.0 37950.0 428700.0 ;
      RECT  39150.0 425100.0 37950.0 426300.0 ;
      RECT  39150.0 427500.0 37950.0 428700.0 ;
      RECT  39150.0 429900.0 37950.0 431100.0 ;
      RECT  39150.0 429900.0 37950.0 431100.0 ;
      RECT  39150.0 427500.0 37950.0 428700.0 ;
      RECT  39150.0 429900.0 37950.0 431100.0 ;
      RECT  39150.0 432300.0 37950.0 433500.0 ;
      RECT  39150.0 432300.0 37950.0 433500.0 ;
      RECT  39150.0 429900.0 37950.0 431100.0 ;
      RECT  47850.0 425100.0 46650.0 426300.0 ;
      RECT  47850.0 427500.0 46650.0 428700.0 ;
      RECT  47850.0 427500.0 46650.0 428700.0 ;
      RECT  47850.0 425100.0 46650.0 426300.0 ;
      RECT  47850.0 427500.0 46650.0 428700.0 ;
      RECT  47850.0 429900.0 46650.0 431100.0 ;
      RECT  47850.0 429900.0 46650.0 431100.0 ;
      RECT  47850.0 427500.0 46650.0 428700.0 ;
      RECT  47850.0 429900.0 46650.0 431100.0 ;
      RECT  47850.0 432300.0 46650.0 433500.0 ;
      RECT  47850.0 432300.0 46650.0 433500.0 ;
      RECT  47850.0 429900.0 46650.0 431100.0 ;
      RECT  38550.0 434700.0 37350.0 435900.0 ;
      RECT  48450.0 434700.0 47250.0 435900.0 ;
      RECT  45750.0 432300.0 44550.0 431100.0 ;
      RECT  43800.0 429900.0 42600.0 428700.0 ;
      RECT  41850.0 427500.0 40650.0 426300.0 ;
      RECT  39150.0 427500.0 37950.0 428700.0 ;
      RECT  39150.0 432300.0 37950.0 433500.0 ;
      RECT  47850.0 432300.0 46650.0 433500.0 ;
      RECT  41850.0 432300.0 40650.0 433500.0 ;
      RECT  41850.0 426300.0 40650.0 427500.0 ;
      RECT  43800.0 428700.0 42600.0 429900.0 ;
      RECT  45750.0 431100.0 44550.0 432300.0 ;
      RECT  41850.0 432300.0 40650.0 433500.0 ;
      RECT  36450.0 423300.0 35550.0 438900.0 ;
      RECT  50250.0 423300.0 49350.0 438900.0 ;
      RECT  37950.0 445500.0 36000.0 446700.0 ;
      RECT  49800.0 445500.0 47850.0 446700.0 ;
      RECT  48450.0 440700.0 50250.0 441900.0 ;
      RECT  39150.0 440700.0 35550.0 441900.0 ;
      RECT  48450.0 443400.0 39150.0 444300.0 ;
      RECT  39150.0 440700.0 37950.0 441900.0 ;
      RECT  39150.0 443100.0 37950.0 444300.0 ;
      RECT  39150.0 443100.0 37950.0 444300.0 ;
      RECT  39150.0 440700.0 37950.0 441900.0 ;
      RECT  48450.0 440700.0 47250.0 441900.0 ;
      RECT  48450.0 443100.0 47250.0 444300.0 ;
      RECT  48450.0 443100.0 47250.0 444300.0 ;
      RECT  48450.0 440700.0 47250.0 441900.0 ;
      RECT  38550.0 445500.0 37350.0 446700.0 ;
      RECT  48450.0 445500.0 47250.0 446700.0 ;
      RECT  43800.0 441300.0 42600.0 442500.0 ;
      RECT  43800.0 441300.0 42600.0 442500.0 ;
      RECT  43650.0 443850.0 42750.0 444750.0 ;
      RECT  36450.0 438900.0 35550.0 448500.0 ;
      RECT  50250.0 438900.0 49350.0 448500.0 ;
      RECT  23550.0 425100.0 21750.0 426300.0 ;
      RECT  23550.0 429900.0 21750.0 431100.0 ;
      RECT  32250.0 425100.0 36450.0 426300.0 ;
      RECT  34050.0 432300.0 36000.0 433500.0 ;
      RECT  22200.0 432300.0 24150.0 433500.0 ;
      RECT  32250.0 425100.0 33450.0 426300.0 ;
      RECT  32250.0 427500.0 33450.0 428700.0 ;
      RECT  32250.0 427500.0 33450.0 428700.0 ;
      RECT  32250.0 425100.0 33450.0 426300.0 ;
      RECT  32250.0 427500.0 33450.0 428700.0 ;
      RECT  32250.0 429900.0 33450.0 431100.0 ;
      RECT  32250.0 429900.0 33450.0 431100.0 ;
      RECT  32250.0 427500.0 33450.0 428700.0 ;
      RECT  23550.0 425100.0 24750.0 426300.0 ;
      RECT  23550.0 427500.0 24750.0 428700.0 ;
      RECT  23550.0 427500.0 24750.0 428700.0 ;
      RECT  23550.0 425100.0 24750.0 426300.0 ;
      RECT  23550.0 427500.0 24750.0 428700.0 ;
      RECT  23550.0 429900.0 24750.0 431100.0 ;
      RECT  23550.0 429900.0 24750.0 431100.0 ;
      RECT  23550.0 427500.0 24750.0 428700.0 ;
      RECT  33450.0 432300.0 34650.0 433500.0 ;
      RECT  23550.0 432300.0 24750.0 433500.0 ;
      RECT  25950.0 429900.0 27150.0 428700.0 ;
      RECT  28650.0 426900.0 29850.0 425700.0 ;
      RECT  32250.0 429900.0 33450.0 431100.0 ;
      RECT  23550.0 428700.0 24750.0 427500.0 ;
      RECT  28650.0 432000.0 29850.0 430800.0 ;
      RECT  28650.0 425700.0 29850.0 426900.0 ;
      RECT  25950.0 428700.0 27150.0 429900.0 ;
      RECT  28650.0 430800.0 29850.0 432000.0 ;
      RECT  35550.0 423300.0 36450.0 437700.0 ;
      RECT  21750.0 423300.0 22650.0 437700.0 ;
      RECT  24150.0 442200.0 21750.0 443400.0 ;
      RECT  32850.0 442200.0 36450.0 443400.0 ;
      RECT  32850.0 447000.0 36450.0 448200.0 ;
      RECT  34050.0 449400.0 36000.0 450600.0 ;
      RECT  22200.0 449400.0 24150.0 450600.0 ;
      RECT  32850.0 442200.0 34050.0 443400.0 ;
      RECT  32850.0 444600.0 34050.0 445800.0 ;
      RECT  32850.0 444600.0 34050.0 445800.0 ;
      RECT  32850.0 442200.0 34050.0 443400.0 ;
      RECT  32850.0 444600.0 34050.0 445800.0 ;
      RECT  32850.0 447000.0 34050.0 448200.0 ;
      RECT  32850.0 447000.0 34050.0 448200.0 ;
      RECT  32850.0 444600.0 34050.0 445800.0 ;
      RECT  24150.0 442200.0 25350.0 443400.0 ;
      RECT  24150.0 444600.0 25350.0 445800.0 ;
      RECT  24150.0 444600.0 25350.0 445800.0 ;
      RECT  24150.0 442200.0 25350.0 443400.0 ;
      RECT  24150.0 444600.0 25350.0 445800.0 ;
      RECT  24150.0 447000.0 25350.0 448200.0 ;
      RECT  24150.0 447000.0 25350.0 448200.0 ;
      RECT  24150.0 444600.0 25350.0 445800.0 ;
      RECT  33450.0 449400.0 34650.0 450600.0 ;
      RECT  23550.0 449400.0 24750.0 450600.0 ;
      RECT  26700.0 447000.0 27900.0 445800.0 ;
      RECT  29400.0 444000.0 30600.0 442800.0 ;
      RECT  32850.0 444600.0 34050.0 445800.0 ;
      RECT  24150.0 447000.0 25350.0 448200.0 ;
      RECT  29400.0 448200.0 30600.0 447000.0 ;
      RECT  29400.0 442800.0 30600.0 444000.0 ;
      RECT  26700.0 445800.0 27900.0 447000.0 ;
      RECT  29400.0 447000.0 30600.0 448200.0 ;
      RECT  35550.0 440400.0 36450.0 454800.0 ;
      RECT  21750.0 440400.0 22650.0 454800.0 ;
      RECT  34050.0 460500.0 36000.0 459300.0 ;
      RECT  22200.0 460500.0 24150.0 459300.0 ;
      RECT  23550.0 465300.0 21750.0 464100.0 ;
      RECT  32850.0 465300.0 36450.0 464100.0 ;
      RECT  23550.0 462600.0 32850.0 461700.0 ;
      RECT  32850.0 465300.0 34050.0 464100.0 ;
      RECT  32850.0 462900.0 34050.0 461700.0 ;
      RECT  32850.0 462900.0 34050.0 461700.0 ;
      RECT  32850.0 465300.0 34050.0 464100.0 ;
      RECT  23550.0 465300.0 24750.0 464100.0 ;
      RECT  23550.0 462900.0 24750.0 461700.0 ;
      RECT  23550.0 462900.0 24750.0 461700.0 ;
      RECT  23550.0 465300.0 24750.0 464100.0 ;
      RECT  33450.0 460500.0 34650.0 459300.0 ;
      RECT  23550.0 460500.0 24750.0 459300.0 ;
      RECT  28200.0 464700.0 29400.0 463500.0 ;
      RECT  28200.0 464700.0 29400.0 463500.0 ;
      RECT  28350.0 462150.0 29250.0 461250.0 ;
      RECT  35550.0 467100.0 36450.0 457500.0 ;
      RECT  21750.0 467100.0 22650.0 457500.0 ;
      RECT  34050.0 470100.0 36000.0 468900.0 ;
      RECT  22200.0 470100.0 24150.0 468900.0 ;
      RECT  23550.0 474900.0 21750.0 473700.0 ;
      RECT  32850.0 474900.0 36450.0 473700.0 ;
      RECT  23550.0 472200.0 32850.0 471300.0 ;
      RECT  32850.0 474900.0 34050.0 473700.0 ;
      RECT  32850.0 472500.0 34050.0 471300.0 ;
      RECT  32850.0 472500.0 34050.0 471300.0 ;
      RECT  32850.0 474900.0 34050.0 473700.0 ;
      RECT  23550.0 474900.0 24750.0 473700.0 ;
      RECT  23550.0 472500.0 24750.0 471300.0 ;
      RECT  23550.0 472500.0 24750.0 471300.0 ;
      RECT  23550.0 474900.0 24750.0 473700.0 ;
      RECT  33450.0 470100.0 34650.0 468900.0 ;
      RECT  23550.0 470100.0 24750.0 468900.0 ;
      RECT  28200.0 474300.0 29400.0 473100.0 ;
      RECT  28200.0 474300.0 29400.0 473100.0 ;
      RECT  28350.0 471750.0 29250.0 470850.0 ;
      RECT  35550.0 476700.0 36450.0 467100.0 ;
      RECT  21750.0 476700.0 22650.0 467100.0 ;
      RECT  20250.0 434700.0 22650.0 435900.0 ;
      RECT  11550.0 434700.0 7950.0 435900.0 ;
      RECT  11550.0 439500.0 7950.0 440700.0 ;
      RECT  10350.0 444300.0 8400.0 445500.0 ;
      RECT  22200.0 444300.0 20250.0 445500.0 ;
      RECT  11550.0 434700.0 10350.0 435900.0 ;
      RECT  11550.0 437100.0 10350.0 438300.0 ;
      RECT  11550.0 437100.0 10350.0 438300.0 ;
      RECT  11550.0 434700.0 10350.0 435900.0 ;
      RECT  11550.0 437100.0 10350.0 438300.0 ;
      RECT  11550.0 439500.0 10350.0 440700.0 ;
      RECT  11550.0 439500.0 10350.0 440700.0 ;
      RECT  11550.0 437100.0 10350.0 438300.0 ;
      RECT  11550.0 439500.0 10350.0 440700.0 ;
      RECT  11550.0 441900.0 10350.0 443100.0 ;
      RECT  11550.0 441900.0 10350.0 443100.0 ;
      RECT  11550.0 439500.0 10350.0 440700.0 ;
      RECT  20250.0 434700.0 19050.0 435900.0 ;
      RECT  20250.0 437100.0 19050.0 438300.0 ;
      RECT  20250.0 437100.0 19050.0 438300.0 ;
      RECT  20250.0 434700.0 19050.0 435900.0 ;
      RECT  20250.0 437100.0 19050.0 438300.0 ;
      RECT  20250.0 439500.0 19050.0 440700.0 ;
      RECT  20250.0 439500.0 19050.0 440700.0 ;
      RECT  20250.0 437100.0 19050.0 438300.0 ;
      RECT  20250.0 439500.0 19050.0 440700.0 ;
      RECT  20250.0 441900.0 19050.0 443100.0 ;
      RECT  20250.0 441900.0 19050.0 443100.0 ;
      RECT  20250.0 439500.0 19050.0 440700.0 ;
      RECT  10950.0 444300.0 9750.0 445500.0 ;
      RECT  20850.0 444300.0 19650.0 445500.0 ;
      RECT  18150.0 441900.0 16950.0 440700.0 ;
      RECT  16200.0 439500.0 15000.0 438300.0 ;
      RECT  14250.0 437100.0 13050.0 435900.0 ;
      RECT  11550.0 437100.0 10350.0 438300.0 ;
      RECT  11550.0 441900.0 10350.0 443100.0 ;
      RECT  20250.0 441900.0 19050.0 443100.0 ;
      RECT  14250.0 441900.0 13050.0 443100.0 ;
      RECT  14250.0 435900.0 13050.0 437100.0 ;
      RECT  16200.0 438300.0 15000.0 439500.0 ;
      RECT  18150.0 440700.0 16950.0 441900.0 ;
      RECT  14250.0 441900.0 13050.0 443100.0 ;
      RECT  8850.0 432900.0 7950.0 448500.0 ;
      RECT  22650.0 432900.0 21750.0 448500.0 ;
      RECT  10350.0 455100.0 8400.0 456300.0 ;
      RECT  22200.0 455100.0 20250.0 456300.0 ;
      RECT  20850.0 450300.0 22650.0 451500.0 ;
      RECT  11550.0 450300.0 7950.0 451500.0 ;
      RECT  20850.0 453000.0 11550.0 453900.0 ;
      RECT  11550.0 450300.0 10350.0 451500.0 ;
      RECT  11550.0 452700.0 10350.0 453900.0 ;
      RECT  11550.0 452700.0 10350.0 453900.0 ;
      RECT  11550.0 450300.0 10350.0 451500.0 ;
      RECT  20850.0 450300.0 19650.0 451500.0 ;
      RECT  20850.0 452700.0 19650.0 453900.0 ;
      RECT  20850.0 452700.0 19650.0 453900.0 ;
      RECT  20850.0 450300.0 19650.0 451500.0 ;
      RECT  10950.0 455100.0 9750.0 456300.0 ;
      RECT  20850.0 455100.0 19650.0 456300.0 ;
      RECT  16200.0 450900.0 15000.0 452100.0 ;
      RECT  16200.0 450900.0 15000.0 452100.0 ;
      RECT  16050.0 453450.0 15150.0 454350.0 ;
      RECT  8850.0 448500.0 7950.0 458100.0 ;
      RECT  22650.0 448500.0 21750.0 458100.0 ;
      RECT  10350.0 464700.0 8400.0 465900.0 ;
      RECT  22200.0 464700.0 20250.0 465900.0 ;
      RECT  20850.0 459900.0 22650.0 461100.0 ;
      RECT  11550.0 459900.0 7950.0 461100.0 ;
      RECT  20850.0 462600.0 11550.0 463500.0 ;
      RECT  11550.0 459900.0 10350.0 461100.0 ;
      RECT  11550.0 462300.0 10350.0 463500.0 ;
      RECT  11550.0 462300.0 10350.0 463500.0 ;
      RECT  11550.0 459900.0 10350.0 461100.0 ;
      RECT  20850.0 459900.0 19650.0 461100.0 ;
      RECT  20850.0 462300.0 19650.0 463500.0 ;
      RECT  20850.0 462300.0 19650.0 463500.0 ;
      RECT  20850.0 459900.0 19650.0 461100.0 ;
      RECT  10950.0 464700.0 9750.0 465900.0 ;
      RECT  20850.0 464700.0 19650.0 465900.0 ;
      RECT  16200.0 460500.0 15000.0 461700.0 ;
      RECT  16200.0 460500.0 15000.0 461700.0 ;
      RECT  16050.0 463050.0 15150.0 463950.0 ;
      RECT  8850.0 458100.0 7950.0 467700.0 ;
      RECT  22650.0 458100.0 21750.0 467700.0 ;
      RECT  10350.0 474300.0 8400.0 475500.0 ;
      RECT  22200.0 474300.0 20250.0 475500.0 ;
      RECT  20850.0 469500.0 22650.0 470700.0 ;
      RECT  11550.0 469500.0 7950.0 470700.0 ;
      RECT  20850.0 472200.0 11550.0 473100.0 ;
      RECT  11550.0 469500.0 10350.0 470700.0 ;
      RECT  11550.0 471900.0 10350.0 473100.0 ;
      RECT  11550.0 471900.0 10350.0 473100.0 ;
      RECT  11550.0 469500.0 10350.0 470700.0 ;
      RECT  20850.0 469500.0 19650.0 470700.0 ;
      RECT  20850.0 471900.0 19650.0 473100.0 ;
      RECT  20850.0 471900.0 19650.0 473100.0 ;
      RECT  20850.0 469500.0 19650.0 470700.0 ;
      RECT  10950.0 474300.0 9750.0 475500.0 ;
      RECT  20850.0 474300.0 19650.0 475500.0 ;
      RECT  16200.0 470100.0 15000.0 471300.0 ;
      RECT  16200.0 470100.0 15000.0 471300.0 ;
      RECT  16050.0 472650.0 15150.0 473550.0 ;
      RECT  8850.0 467700.0 7950.0 477300.0 ;
      RECT  22650.0 467700.0 21750.0 477300.0 ;
      RECT  22650.0 594150.0 21750.0 696300.0 ;
      RECT  21750.0 511350.0 17400.0 512250.0 ;
      RECT  21750.0 534750.0 17400.0 535650.0 ;
      RECT  21750.0 538950.0 17400.0 539850.0 ;
      RECT  21750.0 562350.0 17400.0 563250.0 ;
      RECT  21750.0 566550.0 17400.0 567450.0 ;
      RECT  21750.0 589950.0 17400.0 590850.0 ;
      RECT  21750.0 594150.0 17400.0 595050.0 ;
      RECT  21750.0 617550.0 17400.0 618450.0 ;
      RECT  21750.0 621750.0 17400.0 622650.0 ;
      RECT  21750.0 645150.0 17400.0 646050.0 ;
      RECT  21750.0 649350.0 17400.0 650250.0 ;
      RECT  21750.0 672750.0 17400.0 673650.0 ;
      RECT  21750.0 676950.0 17400.0 677850.0 ;
      RECT  22650.0 485850.0 16800.0 486750.0 ;
      RECT  16800.0 485850.0 6600.0 486750.0 ;
      RECT  4500.0 522900.0 16800.0 523800.0 ;
      RECT  4500.0 550500.0 16800.0 551400.0 ;
      RECT  4500.0 578100.0 16800.0 579000.0 ;
      RECT  4500.0 605700.0 16800.0 606600.0 ;
      RECT  4500.0 633300.0 16800.0 634200.0 ;
      RECT  4500.0 660900.0 16800.0 661800.0 ;
      RECT  4500.0 688500.0 16800.0 689400.0 ;
      RECT  4500.0 495300.0 16800.0 496200.0 ;
      RECT  29250.0 512100.0 28350.0 524700.0 ;
      RECT  29250.0 507150.0 28350.0 508050.0 ;
      RECT  29250.0 507600.0 28350.0 512100.0 ;
      RECT  28800.0 507150.0 17400.0 508050.0 ;
      RECT  36000.0 512850.0 33750.0 513750.0 ;
      RECT  33600.0 498150.0 32700.0 499050.0 ;
      RECT  29250.0 498150.0 28350.0 499050.0 ;
      RECT  33600.0 498600.0 32700.0 510300.0 ;
      RECT  33150.0 498150.0 28800.0 499050.0 ;
      RECT  29250.0 493500.0 28350.0 498600.0 ;
      RECT  28800.0 498150.0 19950.0 499050.0 ;
      RECT  19950.0 490050.0 13200.0 490950.0 ;
      RECT  29400.0 492300.0 28200.0 493500.0 ;
      RECT  29250.0 524700.0 28350.0 528450.0 ;
      RECT  34050.0 489300.0 36000.0 488100.0 ;
      RECT  22200.0 489300.0 24150.0 488100.0 ;
      RECT  23550.0 494100.0 21750.0 492900.0 ;
      RECT  32850.0 494100.0 36450.0 492900.0 ;
      RECT  23550.0 491400.0 32850.0 490500.0 ;
      RECT  32850.0 494100.0 34050.0 492900.0 ;
      RECT  32850.0 491700.0 34050.0 490500.0 ;
      RECT  32850.0 491700.0 34050.0 490500.0 ;
      RECT  32850.0 494100.0 34050.0 492900.0 ;
      RECT  23550.0 494100.0 24750.0 492900.0 ;
      RECT  23550.0 491700.0 24750.0 490500.0 ;
      RECT  23550.0 491700.0 24750.0 490500.0 ;
      RECT  23550.0 494100.0 24750.0 492900.0 ;
      RECT  33450.0 489300.0 34650.0 488100.0 ;
      RECT  23550.0 489300.0 24750.0 488100.0 ;
      RECT  28200.0 493500.0 29400.0 492300.0 ;
      RECT  28200.0 493500.0 29400.0 492300.0 ;
      RECT  28350.0 490950.0 29250.0 490050.0 ;
      RECT  35550.0 495900.0 36450.0 486300.0 ;
      RECT  21750.0 495900.0 22650.0 486300.0 ;
      RECT  32550.0 510300.0 33750.0 511500.0 ;
      RECT  32550.0 512700.0 33750.0 513900.0 ;
      RECT  32550.0 512700.0 33750.0 513900.0 ;
      RECT  32550.0 510300.0 33750.0 511500.0 ;
      RECT  21750.0 593250.0 22650.0 594150.0 ;
      RECT  49350.0 593250.0 50250.0 594150.0 ;
      RECT  21750.0 591900.0 22650.0 593700.0 ;
      RECT  22200.0 593250.0 49800.0 594150.0 ;
      RECT  49350.0 591900.0 50250.0 593700.0 ;
      RECT  37950.0 531300.0 36000.0 532500.0 ;
      RECT  49800.0 531300.0 47850.0 532500.0 ;
      RECT  48450.0 526500.0 50250.0 527700.0 ;
      RECT  39150.0 526500.0 35550.0 527700.0 ;
      RECT  48450.0 529200.0 39150.0 530100.0 ;
      RECT  39150.0 526500.0 37950.0 527700.0 ;
      RECT  39150.0 528900.0 37950.0 530100.0 ;
      RECT  39150.0 528900.0 37950.0 530100.0 ;
      RECT  39150.0 526500.0 37950.0 527700.0 ;
      RECT  48450.0 526500.0 47250.0 527700.0 ;
      RECT  48450.0 528900.0 47250.0 530100.0 ;
      RECT  48450.0 528900.0 47250.0 530100.0 ;
      RECT  48450.0 526500.0 47250.0 527700.0 ;
      RECT  38550.0 531300.0 37350.0 532500.0 ;
      RECT  48450.0 531300.0 47250.0 532500.0 ;
      RECT  43800.0 527100.0 42600.0 528300.0 ;
      RECT  43800.0 527100.0 42600.0 528300.0 ;
      RECT  43650.0 529650.0 42750.0 530550.0 ;
      RECT  36450.0 524700.0 35550.0 534300.0 ;
      RECT  50250.0 524700.0 49350.0 534300.0 ;
      RECT  37950.0 540900.0 36000.0 542100.0 ;
      RECT  49800.0 540900.0 47850.0 542100.0 ;
      RECT  48450.0 536100.0 50250.0 537300.0 ;
      RECT  39150.0 536100.0 35550.0 537300.0 ;
      RECT  48450.0 538800.0 39150.0 539700.0 ;
      RECT  39150.0 536100.0 37950.0 537300.0 ;
      RECT  39150.0 538500.0 37950.0 539700.0 ;
      RECT  39150.0 538500.0 37950.0 539700.0 ;
      RECT  39150.0 536100.0 37950.0 537300.0 ;
      RECT  48450.0 536100.0 47250.0 537300.0 ;
      RECT  48450.0 538500.0 47250.0 539700.0 ;
      RECT  48450.0 538500.0 47250.0 539700.0 ;
      RECT  48450.0 536100.0 47250.0 537300.0 ;
      RECT  38550.0 540900.0 37350.0 542100.0 ;
      RECT  48450.0 540900.0 47250.0 542100.0 ;
      RECT  43800.0 536700.0 42600.0 537900.0 ;
      RECT  43800.0 536700.0 42600.0 537900.0 ;
      RECT  43650.0 539250.0 42750.0 540150.0 ;
      RECT  36450.0 534300.0 35550.0 543900.0 ;
      RECT  50250.0 534300.0 49350.0 543900.0 ;
      RECT  42600.0 536700.0 43800.0 537900.0 ;
      RECT  37950.0 550500.0 36000.0 551700.0 ;
      RECT  49800.0 550500.0 47850.0 551700.0 ;
      RECT  48450.0 545700.0 50250.0 546900.0 ;
      RECT  39150.0 545700.0 35550.0 546900.0 ;
      RECT  48450.0 548400.0 39150.0 549300.0 ;
      RECT  39150.0 545700.0 37950.0 546900.0 ;
      RECT  39150.0 548100.0 37950.0 549300.0 ;
      RECT  39150.0 548100.0 37950.0 549300.0 ;
      RECT  39150.0 545700.0 37950.0 546900.0 ;
      RECT  48450.0 545700.0 47250.0 546900.0 ;
      RECT  48450.0 548100.0 47250.0 549300.0 ;
      RECT  48450.0 548100.0 47250.0 549300.0 ;
      RECT  48450.0 545700.0 47250.0 546900.0 ;
      RECT  38550.0 550500.0 37350.0 551700.0 ;
      RECT  48450.0 550500.0 47250.0 551700.0 ;
      RECT  43800.0 546300.0 42600.0 547500.0 ;
      RECT  43800.0 546300.0 42600.0 547500.0 ;
      RECT  43650.0 548850.0 42750.0 549750.0 ;
      RECT  36450.0 543900.0 35550.0 553500.0 ;
      RECT  50250.0 543900.0 49350.0 553500.0 ;
      RECT  42600.0 546300.0 43800.0 547500.0 ;
      RECT  37950.0 560100.0 36000.0 561300.0 ;
      RECT  49800.0 560100.0 47850.0 561300.0 ;
      RECT  48450.0 555300.0 50250.0 556500.0 ;
      RECT  39150.0 555300.0 35550.0 556500.0 ;
      RECT  48450.0 558000.0 39150.0 558900.0 ;
      RECT  39150.0 555300.0 37950.0 556500.0 ;
      RECT  39150.0 557700.0 37950.0 558900.0 ;
      RECT  39150.0 557700.0 37950.0 558900.0 ;
      RECT  39150.0 555300.0 37950.0 556500.0 ;
      RECT  48450.0 555300.0 47250.0 556500.0 ;
      RECT  48450.0 557700.0 47250.0 558900.0 ;
      RECT  48450.0 557700.0 47250.0 558900.0 ;
      RECT  48450.0 555300.0 47250.0 556500.0 ;
      RECT  38550.0 560100.0 37350.0 561300.0 ;
      RECT  48450.0 560100.0 47250.0 561300.0 ;
      RECT  43800.0 555900.0 42600.0 557100.0 ;
      RECT  43800.0 555900.0 42600.0 557100.0 ;
      RECT  43650.0 558450.0 42750.0 559350.0 ;
      RECT  36450.0 553500.0 35550.0 563100.0 ;
      RECT  50250.0 553500.0 49350.0 563100.0 ;
      RECT  42600.0 555900.0 43800.0 557100.0 ;
      RECT  37950.0 569700.0 36000.0 570900.0 ;
      RECT  49800.0 569700.0 47850.0 570900.0 ;
      RECT  48450.0 564900.0 50250.0 566100.0 ;
      RECT  39150.0 564900.0 35550.0 566100.0 ;
      RECT  48450.0 567600.0 39150.0 568500.0 ;
      RECT  39150.0 564900.0 37950.0 566100.0 ;
      RECT  39150.0 567300.0 37950.0 568500.0 ;
      RECT  39150.0 567300.0 37950.0 568500.0 ;
      RECT  39150.0 564900.0 37950.0 566100.0 ;
      RECT  48450.0 564900.0 47250.0 566100.0 ;
      RECT  48450.0 567300.0 47250.0 568500.0 ;
      RECT  48450.0 567300.0 47250.0 568500.0 ;
      RECT  48450.0 564900.0 47250.0 566100.0 ;
      RECT  38550.0 569700.0 37350.0 570900.0 ;
      RECT  48450.0 569700.0 47250.0 570900.0 ;
      RECT  43800.0 565500.0 42600.0 566700.0 ;
      RECT  43800.0 565500.0 42600.0 566700.0 ;
      RECT  43650.0 568050.0 42750.0 568950.0 ;
      RECT  36450.0 563100.0 35550.0 572700.0 ;
      RECT  50250.0 563100.0 49350.0 572700.0 ;
      RECT  42600.0 565500.0 43800.0 566700.0 ;
      RECT  37950.0 579300.0 36000.0 580500.0 ;
      RECT  49800.0 579300.0 47850.0 580500.0 ;
      RECT  48450.0 574500.0 50250.0 575700.0 ;
      RECT  39150.0 574500.0 35550.0 575700.0 ;
      RECT  48450.0 577200.0 39150.0 578100.0 ;
      RECT  39150.0 574500.0 37950.0 575700.0 ;
      RECT  39150.0 576900.0 37950.0 578100.0 ;
      RECT  39150.0 576900.0 37950.0 578100.0 ;
      RECT  39150.0 574500.0 37950.0 575700.0 ;
      RECT  48450.0 574500.0 47250.0 575700.0 ;
      RECT  48450.0 576900.0 47250.0 578100.0 ;
      RECT  48450.0 576900.0 47250.0 578100.0 ;
      RECT  48450.0 574500.0 47250.0 575700.0 ;
      RECT  38550.0 579300.0 37350.0 580500.0 ;
      RECT  48450.0 579300.0 47250.0 580500.0 ;
      RECT  43800.0 575100.0 42600.0 576300.0 ;
      RECT  43800.0 575100.0 42600.0 576300.0 ;
      RECT  43650.0 577650.0 42750.0 578550.0 ;
      RECT  36450.0 572700.0 35550.0 582300.0 ;
      RECT  50250.0 572700.0 49350.0 582300.0 ;
      RECT  42600.0 575100.0 43800.0 576300.0 ;
      RECT  37950.0 588900.0 36000.0 590100.0 ;
      RECT  49800.0 588900.0 47850.0 590100.0 ;
      RECT  48450.0 584100.0 50250.0 585300.0 ;
      RECT  39150.0 584100.0 35550.0 585300.0 ;
      RECT  48450.0 586800.0 39150.0 587700.0 ;
      RECT  39150.0 584100.0 37950.0 585300.0 ;
      RECT  39150.0 586500.0 37950.0 587700.0 ;
      RECT  39150.0 586500.0 37950.0 587700.0 ;
      RECT  39150.0 584100.0 37950.0 585300.0 ;
      RECT  48450.0 584100.0 47250.0 585300.0 ;
      RECT  48450.0 586500.0 47250.0 587700.0 ;
      RECT  48450.0 586500.0 47250.0 587700.0 ;
      RECT  48450.0 584100.0 47250.0 585300.0 ;
      RECT  38550.0 588900.0 37350.0 590100.0 ;
      RECT  48450.0 588900.0 47250.0 590100.0 ;
      RECT  43800.0 584700.0 42600.0 585900.0 ;
      RECT  43800.0 584700.0 42600.0 585900.0 ;
      RECT  43650.0 587250.0 42750.0 588150.0 ;
      RECT  36450.0 582300.0 35550.0 591900.0 ;
      RECT  50250.0 582300.0 49350.0 591900.0 ;
      RECT  42600.0 584700.0 43800.0 585900.0 ;
      RECT  34050.0 575700.0 36000.0 574500.0 ;
      RECT  22200.0 575700.0 24150.0 574500.0 ;
      RECT  23550.0 580500.0 21750.0 579300.0 ;
      RECT  32850.0 580500.0 36450.0 579300.0 ;
      RECT  23550.0 577800.0 32850.0 576900.0 ;
      RECT  32850.0 580500.0 34050.0 579300.0 ;
      RECT  32850.0 578100.0 34050.0 576900.0 ;
      RECT  32850.0 578100.0 34050.0 576900.0 ;
      RECT  32850.0 580500.0 34050.0 579300.0 ;
      RECT  23550.0 580500.0 24750.0 579300.0 ;
      RECT  23550.0 578100.0 24750.0 576900.0 ;
      RECT  23550.0 578100.0 24750.0 576900.0 ;
      RECT  23550.0 580500.0 24750.0 579300.0 ;
      RECT  33450.0 575700.0 34650.0 574500.0 ;
      RECT  23550.0 575700.0 24750.0 574500.0 ;
      RECT  28200.0 579900.0 29400.0 578700.0 ;
      RECT  28200.0 579900.0 29400.0 578700.0 ;
      RECT  28350.0 577350.0 29250.0 576450.0 ;
      RECT  35550.0 582300.0 36450.0 572700.0 ;
      RECT  21750.0 582300.0 22650.0 572700.0 ;
      RECT  28200.0 578700.0 29400.0 579900.0 ;
      RECT  34050.0 566100.0 36000.0 564900.0 ;
      RECT  22200.0 566100.0 24150.0 564900.0 ;
      RECT  23550.0 570900.0 21750.0 569700.0 ;
      RECT  32850.0 570900.0 36450.0 569700.0 ;
      RECT  23550.0 568200.0 32850.0 567300.0 ;
      RECT  32850.0 570900.0 34050.0 569700.0 ;
      RECT  32850.0 568500.0 34050.0 567300.0 ;
      RECT  32850.0 568500.0 34050.0 567300.0 ;
      RECT  32850.0 570900.0 34050.0 569700.0 ;
      RECT  23550.0 570900.0 24750.0 569700.0 ;
      RECT  23550.0 568500.0 24750.0 567300.0 ;
      RECT  23550.0 568500.0 24750.0 567300.0 ;
      RECT  23550.0 570900.0 24750.0 569700.0 ;
      RECT  33450.0 566100.0 34650.0 564900.0 ;
      RECT  23550.0 566100.0 24750.0 564900.0 ;
      RECT  28200.0 570300.0 29400.0 569100.0 ;
      RECT  28200.0 570300.0 29400.0 569100.0 ;
      RECT  28350.0 567750.0 29250.0 566850.0 ;
      RECT  35550.0 572700.0 36450.0 563100.0 ;
      RECT  21750.0 572700.0 22650.0 563100.0 ;
      RECT  28200.0 569100.0 29400.0 570300.0 ;
      RECT  34050.0 556500.0 36000.0 555300.0 ;
      RECT  22200.0 556500.0 24150.0 555300.0 ;
      RECT  23550.0 561300.0 21750.0 560100.0 ;
      RECT  32850.0 561300.0 36450.0 560100.0 ;
      RECT  23550.0 558600.0 32850.0 557700.0 ;
      RECT  32850.0 561300.0 34050.0 560100.0 ;
      RECT  32850.0 558900.0 34050.0 557700.0 ;
      RECT  32850.0 558900.0 34050.0 557700.0 ;
      RECT  32850.0 561300.0 34050.0 560100.0 ;
      RECT  23550.0 561300.0 24750.0 560100.0 ;
      RECT  23550.0 558900.0 24750.0 557700.0 ;
      RECT  23550.0 558900.0 24750.0 557700.0 ;
      RECT  23550.0 561300.0 24750.0 560100.0 ;
      RECT  33450.0 556500.0 34650.0 555300.0 ;
      RECT  23550.0 556500.0 24750.0 555300.0 ;
      RECT  28200.0 560700.0 29400.0 559500.0 ;
      RECT  28200.0 560700.0 29400.0 559500.0 ;
      RECT  28350.0 558150.0 29250.0 557250.0 ;
      RECT  35550.0 563100.0 36450.0 553500.0 ;
      RECT  21750.0 563100.0 22650.0 553500.0 ;
      RECT  28200.0 559500.0 29400.0 560700.0 ;
      RECT  34050.0 546900.0 36000.0 545700.0 ;
      RECT  22200.0 546900.0 24150.0 545700.0 ;
      RECT  23550.0 551700.0 21750.0 550500.0 ;
      RECT  32850.0 551700.0 36450.0 550500.0 ;
      RECT  23550.0 549000.0 32850.0 548100.0 ;
      RECT  32850.0 551700.0 34050.0 550500.0 ;
      RECT  32850.0 549300.0 34050.0 548100.0 ;
      RECT  32850.0 549300.0 34050.0 548100.0 ;
      RECT  32850.0 551700.0 34050.0 550500.0 ;
      RECT  23550.0 551700.0 24750.0 550500.0 ;
      RECT  23550.0 549300.0 24750.0 548100.0 ;
      RECT  23550.0 549300.0 24750.0 548100.0 ;
      RECT  23550.0 551700.0 24750.0 550500.0 ;
      RECT  33450.0 546900.0 34650.0 545700.0 ;
      RECT  23550.0 546900.0 24750.0 545700.0 ;
      RECT  28200.0 551100.0 29400.0 549900.0 ;
      RECT  28200.0 551100.0 29400.0 549900.0 ;
      RECT  28350.0 548550.0 29250.0 547650.0 ;
      RECT  35550.0 553500.0 36450.0 543900.0 ;
      RECT  21750.0 553500.0 22650.0 543900.0 ;
      RECT  28200.0 549900.0 29400.0 551100.0 ;
      RECT  34050.0 537300.0 36000.0 536100.0 ;
      RECT  22200.0 537300.0 24150.0 536100.0 ;
      RECT  23550.0 542100.0 21750.0 540900.0 ;
      RECT  32850.0 542100.0 36450.0 540900.0 ;
      RECT  23550.0 539400.0 32850.0 538500.0 ;
      RECT  32850.0 542100.0 34050.0 540900.0 ;
      RECT  32850.0 539700.0 34050.0 538500.0 ;
      RECT  32850.0 539700.0 34050.0 538500.0 ;
      RECT  32850.0 542100.0 34050.0 540900.0 ;
      RECT  23550.0 542100.0 24750.0 540900.0 ;
      RECT  23550.0 539700.0 24750.0 538500.0 ;
      RECT  23550.0 539700.0 24750.0 538500.0 ;
      RECT  23550.0 542100.0 24750.0 540900.0 ;
      RECT  33450.0 537300.0 34650.0 536100.0 ;
      RECT  23550.0 537300.0 24750.0 536100.0 ;
      RECT  28200.0 541500.0 29400.0 540300.0 ;
      RECT  28200.0 541500.0 29400.0 540300.0 ;
      RECT  28350.0 538950.0 29250.0 538050.0 ;
      RECT  35550.0 543900.0 36450.0 534300.0 ;
      RECT  21750.0 543900.0 22650.0 534300.0 ;
      RECT  28200.0 540300.0 29400.0 541500.0 ;
      RECT  34050.0 527700.0 36000.0 526500.0 ;
      RECT  22200.0 527700.0 24150.0 526500.0 ;
      RECT  23550.0 532500.0 21750.0 531300.0 ;
      RECT  32850.0 532500.0 36450.0 531300.0 ;
      RECT  23550.0 529800.0 32850.0 528900.0 ;
      RECT  32850.0 532500.0 34050.0 531300.0 ;
      RECT  32850.0 530100.0 34050.0 528900.0 ;
      RECT  32850.0 530100.0 34050.0 528900.0 ;
      RECT  32850.0 532500.0 34050.0 531300.0 ;
      RECT  23550.0 532500.0 24750.0 531300.0 ;
      RECT  23550.0 530100.0 24750.0 528900.0 ;
      RECT  23550.0 530100.0 24750.0 528900.0 ;
      RECT  23550.0 532500.0 24750.0 531300.0 ;
      RECT  33450.0 527700.0 34650.0 526500.0 ;
      RECT  23550.0 527700.0 24750.0 526500.0 ;
      RECT  28200.0 531900.0 29400.0 530700.0 ;
      RECT  28200.0 531900.0 29400.0 530700.0 ;
      RECT  28350.0 529350.0 29250.0 528450.0 ;
      RECT  35550.0 534300.0 36450.0 524700.0 ;
      RECT  21750.0 534300.0 22650.0 524700.0 ;
      RECT  28200.0 530700.0 29400.0 531900.0 ;
      RECT  42600.0 529500.0 43800.0 530700.0 ;
      RECT  42600.0 558300.0 43800.0 559500.0 ;
      RECT  42600.0 587100.0 43800.0 588300.0 ;
      RECT  28200.0 557100.0 29400.0 558300.0 ;
      RECT  42600.0 527100.0 43800.0 528300.0 ;
      RECT  28350.0 524700.0 29250.0 528450.0 ;
      RECT  35550.0 524700.0 36450.0 591900.0 ;
      RECT  21750.0 524700.0 22650.0 591900.0 ;
      RECT  49350.0 524700.0 50250.0 591900.0 ;
      RECT  16800.0 509700.0 6600.0 495900.0 ;
      RECT  16800.0 509700.0 6600.0 523500.0 ;
      RECT  16800.0 537300.0 6600.0 523500.0 ;
      RECT  16800.0 537300.0 6600.0 551100.0 ;
      RECT  16800.0 564900.0 6600.0 551100.0 ;
      RECT  16800.0 564900.0 6600.0 578700.0 ;
      RECT  16800.0 592500.0 6600.0 578700.0 ;
      RECT  16800.0 592500.0 6600.0 606300.0 ;
      RECT  16800.0 620100.0 6600.0 606300.0 ;
      RECT  16800.0 620100.0 6600.0 633900.0 ;
      RECT  16800.0 647700.0 6600.0 633900.0 ;
      RECT  16800.0 647700.0 6600.0 661500.0 ;
      RECT  16800.0 675300.0 6600.0 661500.0 ;
      RECT  16800.0 675300.0 6600.0 689100.0 ;
      RECT  17400.0 511200.0 6000.0 512400.0 ;
      RECT  17400.0 534600.0 6000.0 535800.0 ;
      RECT  17400.0 538800.0 6000.0 540000.0 ;
      RECT  17400.0 562200.0 6000.0 563400.0 ;
      RECT  17400.0 566400.0 6000.0 567600.0 ;
      RECT  17400.0 589800.0 6000.0 591000.0 ;
      RECT  17400.0 594000.0 6000.0 595200.0 ;
      RECT  17400.0 617400.0 6000.0 618600.0 ;
      RECT  17400.0 621600.0 6000.0 622800.0 ;
      RECT  17400.0 645000.0 6000.0 646200.0 ;
      RECT  17400.0 649200.0 6000.0 650400.0 ;
      RECT  17400.0 672600.0 6000.0 673800.0 ;
      RECT  17400.0 676800.0 6000.0 678000.0 ;
      RECT  17400.0 522900.0 6000.0 523800.0 ;
      RECT  17400.0 550500.0 6000.0 551400.0 ;
      RECT  17400.0 578100.0 6000.0 579000.0 ;
      RECT  17400.0 605700.0 6000.0 606600.0 ;
      RECT  17400.0 633300.0 6000.0 634200.0 ;
      RECT  17400.0 660900.0 6000.0 661800.0 ;
      RECT  17400.0 688500.0 6000.0 689400.0 ;
      RECT  22350.0 511200.0 21150.0 512400.0 ;
      RECT  22350.0 534600.0 21150.0 535800.0 ;
      RECT  22350.0 538800.0 21150.0 540000.0 ;
      RECT  22350.0 562200.0 21150.0 563400.0 ;
      RECT  22350.0 566400.0 21150.0 567600.0 ;
      RECT  22350.0 589800.0 21150.0 591000.0 ;
      RECT  22350.0 594000.0 21150.0 595200.0 ;
      RECT  22350.0 617400.0 21150.0 618600.0 ;
      RECT  22350.0 621600.0 21150.0 622800.0 ;
      RECT  22350.0 645000.0 21150.0 646200.0 ;
      RECT  22350.0 649200.0 21150.0 650400.0 ;
      RECT  22350.0 672600.0 21150.0 673800.0 ;
      RECT  22350.0 676800.0 21150.0 678000.0 ;
      RECT  22200.0 524700.0 21000.0 525900.0 ;
      RECT  22800.0 485100.0 21600.0 486300.0 ;
      RECT  16200.0 485700.0 17400.0 486900.0 ;
      RECT  6000.0 485700.0 7200.0 486900.0 ;
      RECT  29400.0 511500.0 28200.0 512700.0 ;
      RECT  19350.0 498000.0 20550.0 499200.0 ;
      RECT  19350.0 489900.0 20550.0 491100.0 ;
      RECT  12600.0 489900.0 13800.0 491100.0 ;
      RECT  43800.0 476700.0 42900.0 527100.0 ;
      RECT  29250.0 476700.0 28350.0 490050.0 ;
      RECT  4500.0 476700.0 3600.0 691350.0 ;
      RECT  36450.0 476700.0 35550.0 524700.0 ;
      RECT  22650.0 476700.0 21750.0 486300.0 ;
      RECT  50250.0 476700.0 49350.0 524700.0 ;
      RECT  43950.0 400050.0 42750.0 398850.0 ;
      RECT  43950.0 359100.0 42750.0 357900.0 ;
      RECT  33900.0 320250.0 32700.0 319050.0 ;
      RECT  29850.0 400050.0 28650.0 398850.0 ;
      RECT  27150.0 405450.0 25950.0 404250.0 ;
      RECT  30600.0 442800.0 29400.0 441600.0 ;
      RECT  27900.0 445800.0 26700.0 444600.0 ;
      RECT  41850.0 418950.0 40650.0 417750.0 ;
      RECT  43800.0 416250.0 42600.0 415050.0 ;
      RECT  45750.0 408150.0 44550.0 406950.0 ;
      RECT  14250.0 418950.0 13050.0 417750.0 ;
      RECT  16200.0 408150.0 15000.0 406950.0 ;
      RECT  18150.0 410850.0 16950.0 409650.0 ;
      RECT  29850.0 437100.0 28650.0 438300.0 ;
      RECT  30600.0 454200.0 29400.0 455400.0 ;
      RECT  16200.0 476700.0 15000.0 477900.0 ;
      RECT  29400.0 456900.0 28200.0 458100.0 ;
      RECT  50400.0 402750.0 49200.0 401550.0 ;
      RECT  36600.0 413550.0 35400.0 412350.0 ;
      RECT  22800.0 402750.0 21600.0 401550.0 ;
      RECT  9000.0 413550.0 7800.0 412350.0 ;
      RECT  43800.0 316800.0 42600.0 320400.0 ;
      RECT  36450.0 316800.0 35550.0 317700.0 ;
      RECT  50250.0 316800.0 49350.0 317700.0 ;
      RECT  55650.0 412350.0 54450.0 413550.0 ;
   LAYER  metal2 ;
      RECT  193350.0 454800.0 194250.0 457500.0 ;
      RECT  190650.0 474600.0 191550.0 477300.0 ;
      RECT  185250.0 435000.0 186150.0 437700.0 ;
      RECT  182550.0 452100.0 183450.0 454800.0 ;
      RECT  187950.0 415650.0 188850.0 418350.0 ;
      RECT  179850.0 396750.0 180750.0 399450.0 ;
      RECT  49800.0 412500.0 55050.0 413400.0 ;
      RECT  174450.0 399450.0 175350.0 402150.0 ;
      RECT  179850.0 600.0 180750.0 1217400.0 ;
      RECT  182550.0 600.0 183450.0 1217400.0 ;
      RECT  185250.0 600.0 186150.0 1217400.0 ;
      RECT  187950.0 600.0 188850.0 1217400.0 ;
      RECT  190650.0 600.0 191550.0 1217400.0 ;
      RECT  193350.0 600.0 194250.0 1217400.0 ;
      RECT  142950.0 600.0 143850.0 313800.0 ;
      RECT  145650.0 600.0 146550.0 313800.0 ;
      RECT  148350.0 600.0 149250.0 313800.0 ;
      RECT  151050.0 600.0 151950.0 313800.0 ;
      RECT  153750.0 600.0 154650.0 313800.0 ;
      RECT  156450.0 600.0 157350.0 313800.0 ;
      RECT  159150.0 600.0 160050.0 313800.0 ;
      RECT  161850.0 600.0 162750.0 313800.0 ;
      RECT  164550.0 600.0 165450.0 313800.0 ;
      RECT  167250.0 600.0 168150.0 313800.0 ;
      RECT  206250.0 1199400.0 207150.0 1200600.0 ;
      RECT  216450.0 1199400.0 217350.0 1200600.0 ;
      RECT  226650.0 1199400.0 227550.0 1200600.0 ;
      RECT  236850.0 1199400.0 237750.0 1200600.0 ;
      RECT  247050.0 1199400.0 247950.0 1200600.0 ;
      RECT  257250.0 1199400.0 258150.0 1200600.0 ;
      RECT  267450.0 1199400.0 268350.0 1200600.0 ;
      RECT  277650.0 1199400.0 278550.0 1200600.0 ;
      RECT  287850.0 1199400.0 288750.0 1200600.0 ;
      RECT  298050.0 1199400.0 298950.0 1200600.0 ;
      RECT  308250.0 1199400.0 309150.0 1200600.0 ;
      RECT  318450.0 1199400.0 319350.0 1200600.0 ;
      RECT  328650.0 1199400.0 329550.0 1200600.0 ;
      RECT  338850.0 1199400.0 339750.0 1200600.0 ;
      RECT  349050.0 1199400.0 349950.0 1200600.0 ;
      RECT  359250.0 1199400.0 360150.0 1200600.0 ;
      RECT  369450.0 1199400.0 370350.0 1200600.0 ;
      RECT  379650.0 1199400.0 380550.0 1200600.0 ;
      RECT  389850.0 1199400.0 390750.0 1200600.0 ;
      RECT  400050.0 1199400.0 400950.0 1200600.0 ;
      RECT  410250.0 1199400.0 411150.0 1200600.0 ;
      RECT  420450.0 1199400.0 421350.0 1200600.0 ;
      RECT  430650.0 1199400.0 431550.0 1200600.0 ;
      RECT  440850.0 1199400.0 441750.0 1200600.0 ;
      RECT  451050.0 1199400.0 451950.0 1200600.0 ;
      RECT  461250.0 1199400.0 462150.0 1200600.0 ;
      RECT  471450.0 1199400.0 472350.0 1200600.0 ;
      RECT  481650.0 1199400.0 482550.0 1200600.0 ;
      RECT  491850.0 1199400.0 492750.0 1200600.0 ;
      RECT  502050.0 1199400.0 502950.0 1200600.0 ;
      RECT  512250.0 1199400.0 513150.0 1200600.0 ;
      RECT  522450.0 1199400.0 523350.0 1200600.0 ;
      RECT  204750.0 79500.0 205650.0 80400.0 ;
      RECT  201600.0 79500.0 205200.0 80400.0 ;
      RECT  204750.0 79950.0 205650.0 81750.0 ;
      RECT  245550.0 79500.0 246450.0 80400.0 ;
      RECT  242400.0 79500.0 246000.0 80400.0 ;
      RECT  245550.0 79950.0 246450.0 81750.0 ;
      RECT  286350.0 79500.0 287250.0 80400.0 ;
      RECT  283200.0 79500.0 286800.0 80400.0 ;
      RECT  286350.0 79950.0 287250.0 81750.0 ;
      RECT  327150.0 79500.0 328050.0 80400.0 ;
      RECT  324000.0 79500.0 327600.0 80400.0 ;
      RECT  327150.0 79950.0 328050.0 81750.0 ;
      RECT  367950.0 79500.0 368850.0 80400.0 ;
      RECT  364800.0 79500.0 368400.0 80400.0 ;
      RECT  367950.0 79950.0 368850.0 81750.0 ;
      RECT  408750.0 79500.0 409650.0 80400.0 ;
      RECT  405600.0 79500.0 409200.0 80400.0 ;
      RECT  408750.0 79950.0 409650.0 81750.0 ;
      RECT  449550.0 79500.0 450450.0 80400.0 ;
      RECT  446400.0 79500.0 450000.0 80400.0 ;
      RECT  449550.0 79950.0 450450.0 81750.0 ;
      RECT  490350.0 79500.0 491250.0 80400.0 ;
      RECT  487200.0 79500.0 490800.0 80400.0 ;
      RECT  490350.0 79950.0 491250.0 81750.0 ;
      RECT  112200.0 1197000.0 113100.0 1199100.0 ;
      RECT  200100.0 313800.0 210300.0 327600.0 ;
      RECT  200100.0 341400.0 210300.0 327600.0 ;
      RECT  200100.0 341400.0 210300.0 355200.0 ;
      RECT  200100.0 369000.0 210300.0 355200.0 ;
      RECT  200100.0 369000.0 210300.0 382800.0 ;
      RECT  200100.0 396600.0 210300.0 382800.0 ;
      RECT  200100.0 396600.0 210300.0 410400.0 ;
      RECT  200100.0 424200.0 210300.0 410400.0 ;
      RECT  200100.0 424200.0 210300.0 438000.0 ;
      RECT  200100.0 451800.0 210300.0 438000.0 ;
      RECT  200100.0 451800.0 210300.0 465600.0 ;
      RECT  200100.0 479400.0 210300.0 465600.0 ;
      RECT  200100.0 479400.0 210300.0 493200.0 ;
      RECT  200100.0 507000.0 210300.0 493200.0 ;
      RECT  200100.0 507000.0 210300.0 520800.0 ;
      RECT  200100.0 534600.0 210300.0 520800.0 ;
      RECT  200100.0 534600.0 210300.0 548400.0 ;
      RECT  200100.0 562200.0 210300.0 548400.0 ;
      RECT  200100.0 562200.0 210300.0 576000.0 ;
      RECT  200100.0 589800.0 210300.0 576000.0 ;
      RECT  200100.0 589800.0 210300.0 603600.0 ;
      RECT  200100.0 617400.0 210300.0 603600.0 ;
      RECT  200100.0 617400.0 210300.0 631200.0 ;
      RECT  200100.0 645000.0 210300.0 631200.0 ;
      RECT  200100.0 645000.0 210300.0 658800.0 ;
      RECT  200100.0 672600.0 210300.0 658800.0 ;
      RECT  200100.0 672600.0 210300.0 686400.0 ;
      RECT  200100.0 700200.0 210300.0 686400.0 ;
      RECT  200100.0 700200.0 210300.0 714000.0 ;
      RECT  200100.0 727800.0 210300.0 714000.0 ;
      RECT  200100.0 727800.0 210300.0 741600.0 ;
      RECT  200100.0 755400.0 210300.0 741600.0 ;
      RECT  200100.0 755400.0 210300.0 769200.0 ;
      RECT  200100.0 783000.0 210300.0 769200.0 ;
      RECT  200100.0 783000.0 210300.0 796800.0 ;
      RECT  200100.0 810600.0 210300.0 796800.0 ;
      RECT  200100.0 810600.0 210300.0 824400.0 ;
      RECT  200100.0 838200.0 210300.0 824400.0 ;
      RECT  200100.0 838200.0 210300.0 852000.0 ;
      RECT  200100.0 865800.0 210300.0 852000.0 ;
      RECT  200100.0 865800.0 210300.0 879600.0 ;
      RECT  200100.0 893400.0 210300.0 879600.0 ;
      RECT  200100.0 893400.0 210300.0 907200.0 ;
      RECT  200100.0 921000.0 210300.0 907200.0 ;
      RECT  200100.0 921000.0 210300.0 934800.0 ;
      RECT  200100.0 948600.0 210300.0 934800.0 ;
      RECT  200100.0 948600.0 210300.0 962400.0 ;
      RECT  200100.0 976200.0 210300.0 962400.0 ;
      RECT  200100.0 976200.0 210300.0 990000.0 ;
      RECT  200100.0 1003800.0 210300.0 990000.0 ;
      RECT  200100.0 1003800.0 210300.0 1017600.0 ;
      RECT  200100.0 1031400.0 210300.0 1017600.0 ;
      RECT  200100.0 1031400.0 210300.0 1045200.0 ;
      RECT  200100.0 1059000.0 210300.0 1045200.0 ;
      RECT  200100.0 1059000.0 210300.0 1072800.0 ;
      RECT  200100.0 1086600.0 210300.0 1072800.0 ;
      RECT  200100.0 1086600.0 210300.0 1100400.0 ;
      RECT  200100.0 1114200.0 210300.0 1100400.0 ;
      RECT  200100.0 1114200.0 210300.0 1128000.0 ;
      RECT  200100.0 1141800.0 210300.0 1128000.0 ;
      RECT  200100.0 1141800.0 210300.0 1155600.0 ;
      RECT  200100.0 1169400.0 210300.0 1155600.0 ;
      RECT  200100.0 1169400.0 210300.0 1183200.0 ;
      RECT  200100.0 1197000.0 210300.0 1183200.0 ;
      RECT  210300.0 313800.0 220500.0 327600.0 ;
      RECT  210300.0 341400.0 220500.0 327600.0 ;
      RECT  210300.0 341400.0 220500.0 355200.0 ;
      RECT  210300.0 369000.0 220500.0 355200.0 ;
      RECT  210300.0 369000.0 220500.0 382800.0 ;
      RECT  210300.0 396600.0 220500.0 382800.0 ;
      RECT  210300.0 396600.0 220500.0 410400.0 ;
      RECT  210300.0 424200.0 220500.0 410400.0 ;
      RECT  210300.0 424200.0 220500.0 438000.0 ;
      RECT  210300.0 451800.0 220500.0 438000.0 ;
      RECT  210300.0 451800.0 220500.0 465600.0 ;
      RECT  210300.0 479400.0 220500.0 465600.0 ;
      RECT  210300.0 479400.0 220500.0 493200.0 ;
      RECT  210300.0 507000.0 220500.0 493200.0 ;
      RECT  210300.0 507000.0 220500.0 520800.0 ;
      RECT  210300.0 534600.0 220500.0 520800.0 ;
      RECT  210300.0 534600.0 220500.0 548400.0 ;
      RECT  210300.0 562200.0 220500.0 548400.0 ;
      RECT  210300.0 562200.0 220500.0 576000.0 ;
      RECT  210300.0 589800.0 220500.0 576000.0 ;
      RECT  210300.0 589800.0 220500.0 603600.0 ;
      RECT  210300.0 617400.0 220500.0 603600.0 ;
      RECT  210300.0 617400.0 220500.0 631200.0 ;
      RECT  210300.0 645000.0 220500.0 631200.0 ;
      RECT  210300.0 645000.0 220500.0 658800.0 ;
      RECT  210300.0 672600.0 220500.0 658800.0 ;
      RECT  210300.0 672600.0 220500.0 686400.0 ;
      RECT  210300.0 700200.0 220500.0 686400.0 ;
      RECT  210300.0 700200.0 220500.0 714000.0 ;
      RECT  210300.0 727800.0 220500.0 714000.0 ;
      RECT  210300.0 727800.0 220500.0 741600.0 ;
      RECT  210300.0 755400.0 220500.0 741600.0 ;
      RECT  210300.0 755400.0 220500.0 769200.0 ;
      RECT  210300.0 783000.0 220500.0 769200.0 ;
      RECT  210300.0 783000.0 220500.0 796800.0 ;
      RECT  210300.0 810600.0 220500.0 796800.0 ;
      RECT  210300.0 810600.0 220500.0 824400.0 ;
      RECT  210300.0 838200.0 220500.0 824400.0 ;
      RECT  210300.0 838200.0 220500.0 852000.0 ;
      RECT  210300.0 865800.0 220500.0 852000.0 ;
      RECT  210300.0 865800.0 220500.0 879600.0 ;
      RECT  210300.0 893400.0 220500.0 879600.0 ;
      RECT  210300.0 893400.0 220500.0 907200.0 ;
      RECT  210300.0 921000.0 220500.0 907200.0 ;
      RECT  210300.0 921000.0 220500.0 934800.0 ;
      RECT  210300.0 948600.0 220500.0 934800.0 ;
      RECT  210300.0 948600.0 220500.0 962400.0 ;
      RECT  210300.0 976200.0 220500.0 962400.0 ;
      RECT  210300.0 976200.0 220500.0 990000.0 ;
      RECT  210300.0 1003800.0 220500.0 990000.0 ;
      RECT  210300.0 1003800.0 220500.0 1017600.0 ;
      RECT  210300.0 1031400.0 220500.0 1017600.0 ;
      RECT  210300.0 1031400.0 220500.0 1045200.0 ;
      RECT  210300.0 1059000.0 220500.0 1045200.0 ;
      RECT  210300.0 1059000.0 220500.0 1072800.0 ;
      RECT  210300.0 1086600.0 220500.0 1072800.0 ;
      RECT  210300.0 1086600.0 220500.0 1100400.0 ;
      RECT  210300.0 1114200.0 220500.0 1100400.0 ;
      RECT  210300.0 1114200.0 220500.0 1128000.0 ;
      RECT  210300.0 1141800.0 220500.0 1128000.0 ;
      RECT  210300.0 1141800.0 220500.0 1155600.0 ;
      RECT  210300.0 1169400.0 220500.0 1155600.0 ;
      RECT  210300.0 1169400.0 220500.0 1183200.0 ;
      RECT  210300.0 1197000.0 220500.0 1183200.0 ;
      RECT  220500.0 313800.0 230700.0 327600.0 ;
      RECT  220500.0 341400.0 230700.0 327600.0 ;
      RECT  220500.0 341400.0 230700.0 355200.0 ;
      RECT  220500.0 369000.0 230700.0 355200.0 ;
      RECT  220500.0 369000.0 230700.0 382800.0 ;
      RECT  220500.0 396600.0 230700.0 382800.0 ;
      RECT  220500.0 396600.0 230700.0 410400.0 ;
      RECT  220500.0 424200.0 230700.0 410400.0 ;
      RECT  220500.0 424200.0 230700.0 438000.0 ;
      RECT  220500.0 451800.0 230700.0 438000.0 ;
      RECT  220500.0 451800.0 230700.0 465600.0 ;
      RECT  220500.0 479400.0 230700.0 465600.0 ;
      RECT  220500.0 479400.0 230700.0 493200.0 ;
      RECT  220500.0 507000.0 230700.0 493200.0 ;
      RECT  220500.0 507000.0 230700.0 520800.0 ;
      RECT  220500.0 534600.0 230700.0 520800.0 ;
      RECT  220500.0 534600.0 230700.0 548400.0 ;
      RECT  220500.0 562200.0 230700.0 548400.0 ;
      RECT  220500.0 562200.0 230700.0 576000.0 ;
      RECT  220500.0 589800.0 230700.0 576000.0 ;
      RECT  220500.0 589800.0 230700.0 603600.0 ;
      RECT  220500.0 617400.0 230700.0 603600.0 ;
      RECT  220500.0 617400.0 230700.0 631200.0 ;
      RECT  220500.0 645000.0 230700.0 631200.0 ;
      RECT  220500.0 645000.0 230700.0 658800.0 ;
      RECT  220500.0 672600.0 230700.0 658800.0 ;
      RECT  220500.0 672600.0 230700.0 686400.0 ;
      RECT  220500.0 700200.0 230700.0 686400.0 ;
      RECT  220500.0 700200.0 230700.0 714000.0 ;
      RECT  220500.0 727800.0 230700.0 714000.0 ;
      RECT  220500.0 727800.0 230700.0 741600.0 ;
      RECT  220500.0 755400.0 230700.0 741600.0 ;
      RECT  220500.0 755400.0 230700.0 769200.0 ;
      RECT  220500.0 783000.0 230700.0 769200.0 ;
      RECT  220500.0 783000.0 230700.0 796800.0 ;
      RECT  220500.0 810600.0 230700.0 796800.0 ;
      RECT  220500.0 810600.0 230700.0 824400.0 ;
      RECT  220500.0 838200.0 230700.0 824400.0 ;
      RECT  220500.0 838200.0 230700.0 852000.0 ;
      RECT  220500.0 865800.0 230700.0 852000.0 ;
      RECT  220500.0 865800.0 230700.0 879600.0 ;
      RECT  220500.0 893400.0 230700.0 879600.0 ;
      RECT  220500.0 893400.0 230700.0 907200.0 ;
      RECT  220500.0 921000.0 230700.0 907200.0 ;
      RECT  220500.0 921000.0 230700.0 934800.0 ;
      RECT  220500.0 948600.0 230700.0 934800.0 ;
      RECT  220500.0 948600.0 230700.0 962400.0 ;
      RECT  220500.0 976200.0 230700.0 962400.0 ;
      RECT  220500.0 976200.0 230700.0 990000.0 ;
      RECT  220500.0 1003800.0 230700.0 990000.0 ;
      RECT  220500.0 1003800.0 230700.0 1017600.0 ;
      RECT  220500.0 1031400.0 230700.0 1017600.0 ;
      RECT  220500.0 1031400.0 230700.0 1045200.0 ;
      RECT  220500.0 1059000.0 230700.0 1045200.0 ;
      RECT  220500.0 1059000.0 230700.0 1072800.0 ;
      RECT  220500.0 1086600.0 230700.0 1072800.0 ;
      RECT  220500.0 1086600.0 230700.0 1100400.0 ;
      RECT  220500.0 1114200.0 230700.0 1100400.0 ;
      RECT  220500.0 1114200.0 230700.0 1128000.0 ;
      RECT  220500.0 1141800.0 230700.0 1128000.0 ;
      RECT  220500.0 1141800.0 230700.0 1155600.0 ;
      RECT  220500.0 1169400.0 230700.0 1155600.0 ;
      RECT  220500.0 1169400.0 230700.0 1183200.0 ;
      RECT  220500.0 1197000.0 230700.0 1183200.0 ;
      RECT  230700.0 313800.0 240900.0 327600.0 ;
      RECT  230700.0 341400.0 240900.0 327600.0 ;
      RECT  230700.0 341400.0 240900.0 355200.0 ;
      RECT  230700.0 369000.0 240900.0 355200.0 ;
      RECT  230700.0 369000.0 240900.0 382800.0 ;
      RECT  230700.0 396600.0 240900.0 382800.0 ;
      RECT  230700.0 396600.0 240900.0 410400.0 ;
      RECT  230700.0 424200.0 240900.0 410400.0 ;
      RECT  230700.0 424200.0 240900.0 438000.0 ;
      RECT  230700.0 451800.0 240900.0 438000.0 ;
      RECT  230700.0 451800.0 240900.0 465600.0 ;
      RECT  230700.0 479400.0 240900.0 465600.0 ;
      RECT  230700.0 479400.0 240900.0 493200.0 ;
      RECT  230700.0 507000.0 240900.0 493200.0 ;
      RECT  230700.0 507000.0 240900.0 520800.0 ;
      RECT  230700.0 534600.0 240900.0 520800.0 ;
      RECT  230700.0 534600.0 240900.0 548400.0 ;
      RECT  230700.0 562200.0 240900.0 548400.0 ;
      RECT  230700.0 562200.0 240900.0 576000.0 ;
      RECT  230700.0 589800.0 240900.0 576000.0 ;
      RECT  230700.0 589800.0 240900.0 603600.0 ;
      RECT  230700.0 617400.0 240900.0 603600.0 ;
      RECT  230700.0 617400.0 240900.0 631200.0 ;
      RECT  230700.0 645000.0 240900.0 631200.0 ;
      RECT  230700.0 645000.0 240900.0 658800.0 ;
      RECT  230700.0 672600.0 240900.0 658800.0 ;
      RECT  230700.0 672600.0 240900.0 686400.0 ;
      RECT  230700.0 700200.0 240900.0 686400.0 ;
      RECT  230700.0 700200.0 240900.0 714000.0 ;
      RECT  230700.0 727800.0 240900.0 714000.0 ;
      RECT  230700.0 727800.0 240900.0 741600.0 ;
      RECT  230700.0 755400.0 240900.0 741600.0 ;
      RECT  230700.0 755400.0 240900.0 769200.0 ;
      RECT  230700.0 783000.0 240900.0 769200.0 ;
      RECT  230700.0 783000.0 240900.0 796800.0 ;
      RECT  230700.0 810600.0 240900.0 796800.0 ;
      RECT  230700.0 810600.0 240900.0 824400.0 ;
      RECT  230700.0 838200.0 240900.0 824400.0 ;
      RECT  230700.0 838200.0 240900.0 852000.0 ;
      RECT  230700.0 865800.0 240900.0 852000.0 ;
      RECT  230700.0 865800.0 240900.0 879600.0 ;
      RECT  230700.0 893400.0 240900.0 879600.0 ;
      RECT  230700.0 893400.0 240900.0 907200.0 ;
      RECT  230700.0 921000.0 240900.0 907200.0 ;
      RECT  230700.0 921000.0 240900.0 934800.0 ;
      RECT  230700.0 948600.0 240900.0 934800.0 ;
      RECT  230700.0 948600.0 240900.0 962400.0 ;
      RECT  230700.0 976200.0 240900.0 962400.0 ;
      RECT  230700.0 976200.0 240900.0 990000.0 ;
      RECT  230700.0 1003800.0 240900.0 990000.0 ;
      RECT  230700.0 1003800.0 240900.0 1017600.0 ;
      RECT  230700.0 1031400.0 240900.0 1017600.0 ;
      RECT  230700.0 1031400.0 240900.0 1045200.0 ;
      RECT  230700.0 1059000.0 240900.0 1045200.0 ;
      RECT  230700.0 1059000.0 240900.0 1072800.0 ;
      RECT  230700.0 1086600.0 240900.0 1072800.0 ;
      RECT  230700.0 1086600.0 240900.0 1100400.0 ;
      RECT  230700.0 1114200.0 240900.0 1100400.0 ;
      RECT  230700.0 1114200.0 240900.0 1128000.0 ;
      RECT  230700.0 1141800.0 240900.0 1128000.0 ;
      RECT  230700.0 1141800.0 240900.0 1155600.0 ;
      RECT  230700.0 1169400.0 240900.0 1155600.0 ;
      RECT  230700.0 1169400.0 240900.0 1183200.0 ;
      RECT  230700.0 1197000.0 240900.0 1183200.0 ;
      RECT  240900.0 313800.0 251100.0 327600.0 ;
      RECT  240900.0 341400.0 251100.0 327600.0 ;
      RECT  240900.0 341400.0 251100.0 355200.0 ;
      RECT  240900.0 369000.0 251100.0 355200.0 ;
      RECT  240900.0 369000.0 251100.0 382800.0 ;
      RECT  240900.0 396600.0 251100.0 382800.0 ;
      RECT  240900.0 396600.0 251100.0 410400.0 ;
      RECT  240900.0 424200.0 251100.0 410400.0 ;
      RECT  240900.0 424200.0 251100.0 438000.0 ;
      RECT  240900.0 451800.0 251100.0 438000.0 ;
      RECT  240900.0 451800.0 251100.0 465600.0 ;
      RECT  240900.0 479400.0 251100.0 465600.0 ;
      RECT  240900.0 479400.0 251100.0 493200.0 ;
      RECT  240900.0 507000.0 251100.0 493200.0 ;
      RECT  240900.0 507000.0 251100.0 520800.0 ;
      RECT  240900.0 534600.0 251100.0 520800.0 ;
      RECT  240900.0 534600.0 251100.0 548400.0 ;
      RECT  240900.0 562200.0 251100.0 548400.0 ;
      RECT  240900.0 562200.0 251100.0 576000.0 ;
      RECT  240900.0 589800.0 251100.0 576000.0 ;
      RECT  240900.0 589800.0 251100.0 603600.0 ;
      RECT  240900.0 617400.0 251100.0 603600.0 ;
      RECT  240900.0 617400.0 251100.0 631200.0 ;
      RECT  240900.0 645000.0 251100.0 631200.0 ;
      RECT  240900.0 645000.0 251100.0 658800.0 ;
      RECT  240900.0 672600.0 251100.0 658800.0 ;
      RECT  240900.0 672600.0 251100.0 686400.0 ;
      RECT  240900.0 700200.0 251100.0 686400.0 ;
      RECT  240900.0 700200.0 251100.0 714000.0 ;
      RECT  240900.0 727800.0 251100.0 714000.0 ;
      RECT  240900.0 727800.0 251100.0 741600.0 ;
      RECT  240900.0 755400.0 251100.0 741600.0 ;
      RECT  240900.0 755400.0 251100.0 769200.0 ;
      RECT  240900.0 783000.0 251100.0 769200.0 ;
      RECT  240900.0 783000.0 251100.0 796800.0 ;
      RECT  240900.0 810600.0 251100.0 796800.0 ;
      RECT  240900.0 810600.0 251100.0 824400.0 ;
      RECT  240900.0 838200.0 251100.0 824400.0 ;
      RECT  240900.0 838200.0 251100.0 852000.0 ;
      RECT  240900.0 865800.0 251100.0 852000.0 ;
      RECT  240900.0 865800.0 251100.0 879600.0 ;
      RECT  240900.0 893400.0 251100.0 879600.0 ;
      RECT  240900.0 893400.0 251100.0 907200.0 ;
      RECT  240900.0 921000.0 251100.0 907200.0 ;
      RECT  240900.0 921000.0 251100.0 934800.0 ;
      RECT  240900.0 948600.0 251100.0 934800.0 ;
      RECT  240900.0 948600.0 251100.0 962400.0 ;
      RECT  240900.0 976200.0 251100.0 962400.0 ;
      RECT  240900.0 976200.0 251100.0 990000.0 ;
      RECT  240900.0 1003800.0 251100.0 990000.0 ;
      RECT  240900.0 1003800.0 251100.0 1017600.0 ;
      RECT  240900.0 1031400.0 251100.0 1017600.0 ;
      RECT  240900.0 1031400.0 251100.0 1045200.0 ;
      RECT  240900.0 1059000.0 251100.0 1045200.0 ;
      RECT  240900.0 1059000.0 251100.0 1072800.0 ;
      RECT  240900.0 1086600.0 251100.0 1072800.0 ;
      RECT  240900.0 1086600.0 251100.0 1100400.0 ;
      RECT  240900.0 1114200.0 251100.0 1100400.0 ;
      RECT  240900.0 1114200.0 251100.0 1128000.0 ;
      RECT  240900.0 1141800.0 251100.0 1128000.0 ;
      RECT  240900.0 1141800.0 251100.0 1155600.0 ;
      RECT  240900.0 1169400.0 251100.0 1155600.0 ;
      RECT  240900.0 1169400.0 251100.0 1183200.0 ;
      RECT  240900.0 1197000.0 251100.0 1183200.0 ;
      RECT  251100.0 313800.0 261300.0 327600.0 ;
      RECT  251100.0 341400.0 261300.0 327600.0 ;
      RECT  251100.0 341400.0 261300.0 355200.0 ;
      RECT  251100.0 369000.0 261300.0 355200.0 ;
      RECT  251100.0 369000.0 261300.0 382800.0 ;
      RECT  251100.0 396600.0 261300.0 382800.0 ;
      RECT  251100.0 396600.0 261300.0 410400.0 ;
      RECT  251100.0 424200.0 261300.0 410400.0 ;
      RECT  251100.0 424200.0 261300.0 438000.0 ;
      RECT  251100.0 451800.0 261300.0 438000.0 ;
      RECT  251100.0 451800.0 261300.0 465600.0 ;
      RECT  251100.0 479400.0 261300.0 465600.0 ;
      RECT  251100.0 479400.0 261300.0 493200.0 ;
      RECT  251100.0 507000.0 261300.0 493200.0 ;
      RECT  251100.0 507000.0 261300.0 520800.0 ;
      RECT  251100.0 534600.0 261300.0 520800.0 ;
      RECT  251100.0 534600.0 261300.0 548400.0 ;
      RECT  251100.0 562200.0 261300.0 548400.0 ;
      RECT  251100.0 562200.0 261300.0 576000.0 ;
      RECT  251100.0 589800.0 261300.0 576000.0 ;
      RECT  251100.0 589800.0 261300.0 603600.0 ;
      RECT  251100.0 617400.0 261300.0 603600.0 ;
      RECT  251100.0 617400.0 261300.0 631200.0 ;
      RECT  251100.0 645000.0 261300.0 631200.0 ;
      RECT  251100.0 645000.0 261300.0 658800.0 ;
      RECT  251100.0 672600.0 261300.0 658800.0 ;
      RECT  251100.0 672600.0 261300.0 686400.0 ;
      RECT  251100.0 700200.0 261300.0 686400.0 ;
      RECT  251100.0 700200.0 261300.0 714000.0 ;
      RECT  251100.0 727800.0 261300.0 714000.0 ;
      RECT  251100.0 727800.0 261300.0 741600.0 ;
      RECT  251100.0 755400.0 261300.0 741600.0 ;
      RECT  251100.0 755400.0 261300.0 769200.0 ;
      RECT  251100.0 783000.0 261300.0 769200.0 ;
      RECT  251100.0 783000.0 261300.0 796800.0 ;
      RECT  251100.0 810600.0 261300.0 796800.0 ;
      RECT  251100.0 810600.0 261300.0 824400.0 ;
      RECT  251100.0 838200.0 261300.0 824400.0 ;
      RECT  251100.0 838200.0 261300.0 852000.0 ;
      RECT  251100.0 865800.0 261300.0 852000.0 ;
      RECT  251100.0 865800.0 261300.0 879600.0 ;
      RECT  251100.0 893400.0 261300.0 879600.0 ;
      RECT  251100.0 893400.0 261300.0 907200.0 ;
      RECT  251100.0 921000.0 261300.0 907200.0 ;
      RECT  251100.0 921000.0 261300.0 934800.0 ;
      RECT  251100.0 948600.0 261300.0 934800.0 ;
      RECT  251100.0 948600.0 261300.0 962400.0 ;
      RECT  251100.0 976200.0 261300.0 962400.0 ;
      RECT  251100.0 976200.0 261300.0 990000.0 ;
      RECT  251100.0 1003800.0 261300.0 990000.0 ;
      RECT  251100.0 1003800.0 261300.0 1017600.0 ;
      RECT  251100.0 1031400.0 261300.0 1017600.0 ;
      RECT  251100.0 1031400.0 261300.0 1045200.0 ;
      RECT  251100.0 1059000.0 261300.0 1045200.0 ;
      RECT  251100.0 1059000.0 261300.0 1072800.0 ;
      RECT  251100.0 1086600.0 261300.0 1072800.0 ;
      RECT  251100.0 1086600.0 261300.0 1100400.0 ;
      RECT  251100.0 1114200.0 261300.0 1100400.0 ;
      RECT  251100.0 1114200.0 261300.0 1128000.0 ;
      RECT  251100.0 1141800.0 261300.0 1128000.0 ;
      RECT  251100.0 1141800.0 261300.0 1155600.0 ;
      RECT  251100.0 1169400.0 261300.0 1155600.0 ;
      RECT  251100.0 1169400.0 261300.0 1183200.0 ;
      RECT  251100.0 1197000.0 261300.0 1183200.0 ;
      RECT  261300.0 313800.0 271500.0 327600.0 ;
      RECT  261300.0 341400.0 271500.0 327600.0 ;
      RECT  261300.0 341400.0 271500.0 355200.0 ;
      RECT  261300.0 369000.0 271500.0 355200.0 ;
      RECT  261300.0 369000.0 271500.0 382800.0 ;
      RECT  261300.0 396600.0 271500.0 382800.0 ;
      RECT  261300.0 396600.0 271500.0 410400.0 ;
      RECT  261300.0 424200.0 271500.0 410400.0 ;
      RECT  261300.0 424200.0 271500.0 438000.0 ;
      RECT  261300.0 451800.0 271500.0 438000.0 ;
      RECT  261300.0 451800.0 271500.0 465600.0 ;
      RECT  261300.0 479400.0 271500.0 465600.0 ;
      RECT  261300.0 479400.0 271500.0 493200.0 ;
      RECT  261300.0 507000.0 271500.0 493200.0 ;
      RECT  261300.0 507000.0 271500.0 520800.0 ;
      RECT  261300.0 534600.0 271500.0 520800.0 ;
      RECT  261300.0 534600.0 271500.0 548400.0 ;
      RECT  261300.0 562200.0 271500.0 548400.0 ;
      RECT  261300.0 562200.0 271500.0 576000.0 ;
      RECT  261300.0 589800.0 271500.0 576000.0 ;
      RECT  261300.0 589800.0 271500.0 603600.0 ;
      RECT  261300.0 617400.0 271500.0 603600.0 ;
      RECT  261300.0 617400.0 271500.0 631200.0 ;
      RECT  261300.0 645000.0 271500.0 631200.0 ;
      RECT  261300.0 645000.0 271500.0 658800.0 ;
      RECT  261300.0 672600.0 271500.0 658800.0 ;
      RECT  261300.0 672600.0 271500.0 686400.0 ;
      RECT  261300.0 700200.0 271500.0 686400.0 ;
      RECT  261300.0 700200.0 271500.0 714000.0 ;
      RECT  261300.0 727800.0 271500.0 714000.0 ;
      RECT  261300.0 727800.0 271500.0 741600.0 ;
      RECT  261300.0 755400.0 271500.0 741600.0 ;
      RECT  261300.0 755400.0 271500.0 769200.0 ;
      RECT  261300.0 783000.0 271500.0 769200.0 ;
      RECT  261300.0 783000.0 271500.0 796800.0 ;
      RECT  261300.0 810600.0 271500.0 796800.0 ;
      RECT  261300.0 810600.0 271500.0 824400.0 ;
      RECT  261300.0 838200.0 271500.0 824400.0 ;
      RECT  261300.0 838200.0 271500.0 852000.0 ;
      RECT  261300.0 865800.0 271500.0 852000.0 ;
      RECT  261300.0 865800.0 271500.0 879600.0 ;
      RECT  261300.0 893400.0 271500.0 879600.0 ;
      RECT  261300.0 893400.0 271500.0 907200.0 ;
      RECT  261300.0 921000.0 271500.0 907200.0 ;
      RECT  261300.0 921000.0 271500.0 934800.0 ;
      RECT  261300.0 948600.0 271500.0 934800.0 ;
      RECT  261300.0 948600.0 271500.0 962400.0 ;
      RECT  261300.0 976200.0 271500.0 962400.0 ;
      RECT  261300.0 976200.0 271500.0 990000.0 ;
      RECT  261300.0 1003800.0 271500.0 990000.0 ;
      RECT  261300.0 1003800.0 271500.0 1017600.0 ;
      RECT  261300.0 1031400.0 271500.0 1017600.0 ;
      RECT  261300.0 1031400.0 271500.0 1045200.0 ;
      RECT  261300.0 1059000.0 271500.0 1045200.0 ;
      RECT  261300.0 1059000.0 271500.0 1072800.0 ;
      RECT  261300.0 1086600.0 271500.0 1072800.0 ;
      RECT  261300.0 1086600.0 271500.0 1100400.0 ;
      RECT  261300.0 1114200.0 271500.0 1100400.0 ;
      RECT  261300.0 1114200.0 271500.0 1128000.0 ;
      RECT  261300.0 1141800.0 271500.0 1128000.0 ;
      RECT  261300.0 1141800.0 271500.0 1155600.0 ;
      RECT  261300.0 1169400.0 271500.0 1155600.0 ;
      RECT  261300.0 1169400.0 271500.0 1183200.0 ;
      RECT  261300.0 1197000.0 271500.0 1183200.0 ;
      RECT  271500.0 313800.0 281700.0 327600.0 ;
      RECT  271500.0 341400.0 281700.0 327600.0 ;
      RECT  271500.0 341400.0 281700.0 355200.0 ;
      RECT  271500.0 369000.0 281700.0 355200.0 ;
      RECT  271500.0 369000.0 281700.0 382800.0 ;
      RECT  271500.0 396600.0 281700.0 382800.0 ;
      RECT  271500.0 396600.0 281700.0 410400.0 ;
      RECT  271500.0 424200.0 281700.0 410400.0 ;
      RECT  271500.0 424200.0 281700.0 438000.0 ;
      RECT  271500.0 451800.0 281700.0 438000.0 ;
      RECT  271500.0 451800.0 281700.0 465600.0 ;
      RECT  271500.0 479400.0 281700.0 465600.0 ;
      RECT  271500.0 479400.0 281700.0 493200.0 ;
      RECT  271500.0 507000.0 281700.0 493200.0 ;
      RECT  271500.0 507000.0 281700.0 520800.0 ;
      RECT  271500.0 534600.0 281700.0 520800.0 ;
      RECT  271500.0 534600.0 281700.0 548400.0 ;
      RECT  271500.0 562200.0 281700.0 548400.0 ;
      RECT  271500.0 562200.0 281700.0 576000.0 ;
      RECT  271500.0 589800.0 281700.0 576000.0 ;
      RECT  271500.0 589800.0 281700.0 603600.0 ;
      RECT  271500.0 617400.0 281700.0 603600.0 ;
      RECT  271500.0 617400.0 281700.0 631200.0 ;
      RECT  271500.0 645000.0 281700.0 631200.0 ;
      RECT  271500.0 645000.0 281700.0 658800.0 ;
      RECT  271500.0 672600.0 281700.0 658800.0 ;
      RECT  271500.0 672600.0 281700.0 686400.0 ;
      RECT  271500.0 700200.0 281700.0 686400.0 ;
      RECT  271500.0 700200.0 281700.0 714000.0 ;
      RECT  271500.0 727800.0 281700.0 714000.0 ;
      RECT  271500.0 727800.0 281700.0 741600.0 ;
      RECT  271500.0 755400.0 281700.0 741600.0 ;
      RECT  271500.0 755400.0 281700.0 769200.0 ;
      RECT  271500.0 783000.0 281700.0 769200.0 ;
      RECT  271500.0 783000.0 281700.0 796800.0 ;
      RECT  271500.0 810600.0 281700.0 796800.0 ;
      RECT  271500.0 810600.0 281700.0 824400.0 ;
      RECT  271500.0 838200.0 281700.0 824400.0 ;
      RECT  271500.0 838200.0 281700.0 852000.0 ;
      RECT  271500.0 865800.0 281700.0 852000.0 ;
      RECT  271500.0 865800.0 281700.0 879600.0 ;
      RECT  271500.0 893400.0 281700.0 879600.0 ;
      RECT  271500.0 893400.0 281700.0 907200.0 ;
      RECT  271500.0 921000.0 281700.0 907200.0 ;
      RECT  271500.0 921000.0 281700.0 934800.0 ;
      RECT  271500.0 948600.0 281700.0 934800.0 ;
      RECT  271500.0 948600.0 281700.0 962400.0 ;
      RECT  271500.0 976200.0 281700.0 962400.0 ;
      RECT  271500.0 976200.0 281700.0 990000.0 ;
      RECT  271500.0 1003800.0 281700.0 990000.0 ;
      RECT  271500.0 1003800.0 281700.0 1017600.0 ;
      RECT  271500.0 1031400.0 281700.0 1017600.0 ;
      RECT  271500.0 1031400.0 281700.0 1045200.0 ;
      RECT  271500.0 1059000.0 281700.0 1045200.0 ;
      RECT  271500.0 1059000.0 281700.0 1072800.0 ;
      RECT  271500.0 1086600.0 281700.0 1072800.0 ;
      RECT  271500.0 1086600.0 281700.0 1100400.0 ;
      RECT  271500.0 1114200.0 281700.0 1100400.0 ;
      RECT  271500.0 1114200.0 281700.0 1128000.0 ;
      RECT  271500.0 1141800.0 281700.0 1128000.0 ;
      RECT  271500.0 1141800.0 281700.0 1155600.0 ;
      RECT  271500.0 1169400.0 281700.0 1155600.0 ;
      RECT  271500.0 1169400.0 281700.0 1183200.0 ;
      RECT  271500.0 1197000.0 281700.0 1183200.0 ;
      RECT  281700.0 313800.0 291900.0 327600.0 ;
      RECT  281700.0 341400.0 291900.0 327600.0 ;
      RECT  281700.0 341400.0 291900.0 355200.0 ;
      RECT  281700.0 369000.0 291900.0 355200.0 ;
      RECT  281700.0 369000.0 291900.0 382800.0 ;
      RECT  281700.0 396600.0 291900.0 382800.0 ;
      RECT  281700.0 396600.0 291900.0 410400.0 ;
      RECT  281700.0 424200.0 291900.0 410400.0 ;
      RECT  281700.0 424200.0 291900.0 438000.0 ;
      RECT  281700.0 451800.0 291900.0 438000.0 ;
      RECT  281700.0 451800.0 291900.0 465600.0 ;
      RECT  281700.0 479400.0 291900.0 465600.0 ;
      RECT  281700.0 479400.0 291900.0 493200.0 ;
      RECT  281700.0 507000.0 291900.0 493200.0 ;
      RECT  281700.0 507000.0 291900.0 520800.0 ;
      RECT  281700.0 534600.0 291900.0 520800.0 ;
      RECT  281700.0 534600.0 291900.0 548400.0 ;
      RECT  281700.0 562200.0 291900.0 548400.0 ;
      RECT  281700.0 562200.0 291900.0 576000.0 ;
      RECT  281700.0 589800.0 291900.0 576000.0 ;
      RECT  281700.0 589800.0 291900.0 603600.0 ;
      RECT  281700.0 617400.0 291900.0 603600.0 ;
      RECT  281700.0 617400.0 291900.0 631200.0 ;
      RECT  281700.0 645000.0 291900.0 631200.0 ;
      RECT  281700.0 645000.0 291900.0 658800.0 ;
      RECT  281700.0 672600.0 291900.0 658800.0 ;
      RECT  281700.0 672600.0 291900.0 686400.0 ;
      RECT  281700.0 700200.0 291900.0 686400.0 ;
      RECT  281700.0 700200.0 291900.0 714000.0 ;
      RECT  281700.0 727800.0 291900.0 714000.0 ;
      RECT  281700.0 727800.0 291900.0 741600.0 ;
      RECT  281700.0 755400.0 291900.0 741600.0 ;
      RECT  281700.0 755400.0 291900.0 769200.0 ;
      RECT  281700.0 783000.0 291900.0 769200.0 ;
      RECT  281700.0 783000.0 291900.0 796800.0 ;
      RECT  281700.0 810600.0 291900.0 796800.0 ;
      RECT  281700.0 810600.0 291900.0 824400.0 ;
      RECT  281700.0 838200.0 291900.0 824400.0 ;
      RECT  281700.0 838200.0 291900.0 852000.0 ;
      RECT  281700.0 865800.0 291900.0 852000.0 ;
      RECT  281700.0 865800.0 291900.0 879600.0 ;
      RECT  281700.0 893400.0 291900.0 879600.0 ;
      RECT  281700.0 893400.0 291900.0 907200.0 ;
      RECT  281700.0 921000.0 291900.0 907200.0 ;
      RECT  281700.0 921000.0 291900.0 934800.0 ;
      RECT  281700.0 948600.0 291900.0 934800.0 ;
      RECT  281700.0 948600.0 291900.0 962400.0 ;
      RECT  281700.0 976200.0 291900.0 962400.0 ;
      RECT  281700.0 976200.0 291900.0 990000.0 ;
      RECT  281700.0 1003800.0 291900.0 990000.0 ;
      RECT  281700.0 1003800.0 291900.0 1017600.0 ;
      RECT  281700.0 1031400.0 291900.0 1017600.0 ;
      RECT  281700.0 1031400.0 291900.0 1045200.0 ;
      RECT  281700.0 1059000.0 291900.0 1045200.0 ;
      RECT  281700.0 1059000.0 291900.0 1072800.0 ;
      RECT  281700.0 1086600.0 291900.0 1072800.0 ;
      RECT  281700.0 1086600.0 291900.0 1100400.0 ;
      RECT  281700.0 1114200.0 291900.0 1100400.0 ;
      RECT  281700.0 1114200.0 291900.0 1128000.0 ;
      RECT  281700.0 1141800.0 291900.0 1128000.0 ;
      RECT  281700.0 1141800.0 291900.0 1155600.0 ;
      RECT  281700.0 1169400.0 291900.0 1155600.0 ;
      RECT  281700.0 1169400.0 291900.0 1183200.0 ;
      RECT  281700.0 1197000.0 291900.0 1183200.0 ;
      RECT  291900.0 313800.0 302100.0 327600.0 ;
      RECT  291900.0 341400.0 302100.0 327600.0 ;
      RECT  291900.0 341400.0 302100.0 355200.0 ;
      RECT  291900.0 369000.0 302100.0 355200.0 ;
      RECT  291900.0 369000.0 302100.0 382800.0 ;
      RECT  291900.0 396600.0 302100.0 382800.0 ;
      RECT  291900.0 396600.0 302100.0 410400.0 ;
      RECT  291900.0 424200.0 302100.0 410400.0 ;
      RECT  291900.0 424200.0 302100.0 438000.0 ;
      RECT  291900.0 451800.0 302100.0 438000.0 ;
      RECT  291900.0 451800.0 302100.0 465600.0 ;
      RECT  291900.0 479400.0 302100.0 465600.0 ;
      RECT  291900.0 479400.0 302100.0 493200.0 ;
      RECT  291900.0 507000.0 302100.0 493200.0 ;
      RECT  291900.0 507000.0 302100.0 520800.0 ;
      RECT  291900.0 534600.0 302100.0 520800.0 ;
      RECT  291900.0 534600.0 302100.0 548400.0 ;
      RECT  291900.0 562200.0 302100.0 548400.0 ;
      RECT  291900.0 562200.0 302100.0 576000.0 ;
      RECT  291900.0 589800.0 302100.0 576000.0 ;
      RECT  291900.0 589800.0 302100.0 603600.0 ;
      RECT  291900.0 617400.0 302100.0 603600.0 ;
      RECT  291900.0 617400.0 302100.0 631200.0 ;
      RECT  291900.0 645000.0 302100.0 631200.0 ;
      RECT  291900.0 645000.0 302100.0 658800.0 ;
      RECT  291900.0 672600.0 302100.0 658800.0 ;
      RECT  291900.0 672600.0 302100.0 686400.0 ;
      RECT  291900.0 700200.0 302100.0 686400.0 ;
      RECT  291900.0 700200.0 302100.0 714000.0 ;
      RECT  291900.0 727800.0 302100.0 714000.0 ;
      RECT  291900.0 727800.0 302100.0 741600.0 ;
      RECT  291900.0 755400.0 302100.0 741600.0 ;
      RECT  291900.0 755400.0 302100.0 769200.0 ;
      RECT  291900.0 783000.0 302100.0 769200.0 ;
      RECT  291900.0 783000.0 302100.0 796800.0 ;
      RECT  291900.0 810600.0 302100.0 796800.0 ;
      RECT  291900.0 810600.0 302100.0 824400.0 ;
      RECT  291900.0 838200.0 302100.0 824400.0 ;
      RECT  291900.0 838200.0 302100.0 852000.0 ;
      RECT  291900.0 865800.0 302100.0 852000.0 ;
      RECT  291900.0 865800.0 302100.0 879600.0 ;
      RECT  291900.0 893400.0 302100.0 879600.0 ;
      RECT  291900.0 893400.0 302100.0 907200.0 ;
      RECT  291900.0 921000.0 302100.0 907200.0 ;
      RECT  291900.0 921000.0 302100.0 934800.0 ;
      RECT  291900.0 948600.0 302100.0 934800.0 ;
      RECT  291900.0 948600.0 302100.0 962400.0 ;
      RECT  291900.0 976200.0 302100.0 962400.0 ;
      RECT  291900.0 976200.0 302100.0 990000.0 ;
      RECT  291900.0 1003800.0 302100.0 990000.0 ;
      RECT  291900.0 1003800.0 302100.0 1017600.0 ;
      RECT  291900.0 1031400.0 302100.0 1017600.0 ;
      RECT  291900.0 1031400.0 302100.0 1045200.0 ;
      RECT  291900.0 1059000.0 302100.0 1045200.0 ;
      RECT  291900.0 1059000.0 302100.0 1072800.0 ;
      RECT  291900.0 1086600.0 302100.0 1072800.0 ;
      RECT  291900.0 1086600.0 302100.0 1100400.0 ;
      RECT  291900.0 1114200.0 302100.0 1100400.0 ;
      RECT  291900.0 1114200.0 302100.0 1128000.0 ;
      RECT  291900.0 1141800.0 302100.0 1128000.0 ;
      RECT  291900.0 1141800.0 302100.0 1155600.0 ;
      RECT  291900.0 1169400.0 302100.0 1155600.0 ;
      RECT  291900.0 1169400.0 302100.0 1183200.0 ;
      RECT  291900.0 1197000.0 302100.0 1183200.0 ;
      RECT  302100.0 313800.0 312300.0 327600.0 ;
      RECT  302100.0 341400.0 312300.0 327600.0 ;
      RECT  302100.0 341400.0 312300.0 355200.0 ;
      RECT  302100.0 369000.0 312300.0 355200.0 ;
      RECT  302100.0 369000.0 312300.0 382800.0 ;
      RECT  302100.0 396600.0 312300.0 382800.0 ;
      RECT  302100.0 396600.0 312300.0 410400.0 ;
      RECT  302100.0 424200.0 312300.0 410400.0 ;
      RECT  302100.0 424200.0 312300.0 438000.0 ;
      RECT  302100.0 451800.0 312300.0 438000.0 ;
      RECT  302100.0 451800.0 312300.0 465600.0 ;
      RECT  302100.0 479400.0 312300.0 465600.0 ;
      RECT  302100.0 479400.0 312300.0 493200.0 ;
      RECT  302100.0 507000.0 312300.0 493200.0 ;
      RECT  302100.0 507000.0 312300.0 520800.0 ;
      RECT  302100.0 534600.0 312300.0 520800.0 ;
      RECT  302100.0 534600.0 312300.0 548400.0 ;
      RECT  302100.0 562200.0 312300.0 548400.0 ;
      RECT  302100.0 562200.0 312300.0 576000.0 ;
      RECT  302100.0 589800.0 312300.0 576000.0 ;
      RECT  302100.0 589800.0 312300.0 603600.0 ;
      RECT  302100.0 617400.0 312300.0 603600.0 ;
      RECT  302100.0 617400.0 312300.0 631200.0 ;
      RECT  302100.0 645000.0 312300.0 631200.0 ;
      RECT  302100.0 645000.0 312300.0 658800.0 ;
      RECT  302100.0 672600.0 312300.0 658800.0 ;
      RECT  302100.0 672600.0 312300.0 686400.0 ;
      RECT  302100.0 700200.0 312300.0 686400.0 ;
      RECT  302100.0 700200.0 312300.0 714000.0 ;
      RECT  302100.0 727800.0 312300.0 714000.0 ;
      RECT  302100.0 727800.0 312300.0 741600.0 ;
      RECT  302100.0 755400.0 312300.0 741600.0 ;
      RECT  302100.0 755400.0 312300.0 769200.0 ;
      RECT  302100.0 783000.0 312300.0 769200.0 ;
      RECT  302100.0 783000.0 312300.0 796800.0 ;
      RECT  302100.0 810600.0 312300.0 796800.0 ;
      RECT  302100.0 810600.0 312300.0 824400.0 ;
      RECT  302100.0 838200.0 312300.0 824400.0 ;
      RECT  302100.0 838200.0 312300.0 852000.0 ;
      RECT  302100.0 865800.0 312300.0 852000.0 ;
      RECT  302100.0 865800.0 312300.0 879600.0 ;
      RECT  302100.0 893400.0 312300.0 879600.0 ;
      RECT  302100.0 893400.0 312300.0 907200.0 ;
      RECT  302100.0 921000.0 312300.0 907200.0 ;
      RECT  302100.0 921000.0 312300.0 934800.0 ;
      RECT  302100.0 948600.0 312300.0 934800.0 ;
      RECT  302100.0 948600.0 312300.0 962400.0 ;
      RECT  302100.0 976200.0 312300.0 962400.0 ;
      RECT  302100.0 976200.0 312300.0 990000.0 ;
      RECT  302100.0 1003800.0 312300.0 990000.0 ;
      RECT  302100.0 1003800.0 312300.0 1017600.0 ;
      RECT  302100.0 1031400.0 312300.0 1017600.0 ;
      RECT  302100.0 1031400.0 312300.0 1045200.0 ;
      RECT  302100.0 1059000.0 312300.0 1045200.0 ;
      RECT  302100.0 1059000.0 312300.0 1072800.0 ;
      RECT  302100.0 1086600.0 312300.0 1072800.0 ;
      RECT  302100.0 1086600.0 312300.0 1100400.0 ;
      RECT  302100.0 1114200.0 312300.0 1100400.0 ;
      RECT  302100.0 1114200.0 312300.0 1128000.0 ;
      RECT  302100.0 1141800.0 312300.0 1128000.0 ;
      RECT  302100.0 1141800.0 312300.0 1155600.0 ;
      RECT  302100.0 1169400.0 312300.0 1155600.0 ;
      RECT  302100.0 1169400.0 312300.0 1183200.0 ;
      RECT  302100.0 1197000.0 312300.0 1183200.0 ;
      RECT  312300.0 313800.0 322500.0 327600.0 ;
      RECT  312300.0 341400.0 322500.0 327600.0 ;
      RECT  312300.0 341400.0 322500.0 355200.0 ;
      RECT  312300.0 369000.0 322500.0 355200.0 ;
      RECT  312300.0 369000.0 322500.0 382800.0 ;
      RECT  312300.0 396600.0 322500.0 382800.0 ;
      RECT  312300.0 396600.0 322500.0 410400.0 ;
      RECT  312300.0 424200.0 322500.0 410400.0 ;
      RECT  312300.0 424200.0 322500.0 438000.0 ;
      RECT  312300.0 451800.0 322500.0 438000.0 ;
      RECT  312300.0 451800.0 322500.0 465600.0 ;
      RECT  312300.0 479400.0 322500.0 465600.0 ;
      RECT  312300.0 479400.0 322500.0 493200.0 ;
      RECT  312300.0 507000.0 322500.0 493200.0 ;
      RECT  312300.0 507000.0 322500.0 520800.0 ;
      RECT  312300.0 534600.0 322500.0 520800.0 ;
      RECT  312300.0 534600.0 322500.0 548400.0 ;
      RECT  312300.0 562200.0 322500.0 548400.0 ;
      RECT  312300.0 562200.0 322500.0 576000.0 ;
      RECT  312300.0 589800.0 322500.0 576000.0 ;
      RECT  312300.0 589800.0 322500.0 603600.0 ;
      RECT  312300.0 617400.0 322500.0 603600.0 ;
      RECT  312300.0 617400.0 322500.0 631200.0 ;
      RECT  312300.0 645000.0 322500.0 631200.0 ;
      RECT  312300.0 645000.0 322500.0 658800.0 ;
      RECT  312300.0 672600.0 322500.0 658800.0 ;
      RECT  312300.0 672600.0 322500.0 686400.0 ;
      RECT  312300.0 700200.0 322500.0 686400.0 ;
      RECT  312300.0 700200.0 322500.0 714000.0 ;
      RECT  312300.0 727800.0 322500.0 714000.0 ;
      RECT  312300.0 727800.0 322500.0 741600.0 ;
      RECT  312300.0 755400.0 322500.0 741600.0 ;
      RECT  312300.0 755400.0 322500.0 769200.0 ;
      RECT  312300.0 783000.0 322500.0 769200.0 ;
      RECT  312300.0 783000.0 322500.0 796800.0 ;
      RECT  312300.0 810600.0 322500.0 796800.0 ;
      RECT  312300.0 810600.0 322500.0 824400.0 ;
      RECT  312300.0 838200.0 322500.0 824400.0 ;
      RECT  312300.0 838200.0 322500.0 852000.0 ;
      RECT  312300.0 865800.0 322500.0 852000.0 ;
      RECT  312300.0 865800.0 322500.0 879600.0 ;
      RECT  312300.0 893400.0 322500.0 879600.0 ;
      RECT  312300.0 893400.0 322500.0 907200.0 ;
      RECT  312300.0 921000.0 322500.0 907200.0 ;
      RECT  312300.0 921000.0 322500.0 934800.0 ;
      RECT  312300.0 948600.0 322500.0 934800.0 ;
      RECT  312300.0 948600.0 322500.0 962400.0 ;
      RECT  312300.0 976200.0 322500.0 962400.0 ;
      RECT  312300.0 976200.0 322500.0 990000.0 ;
      RECT  312300.0 1003800.0 322500.0 990000.0 ;
      RECT  312300.0 1003800.0 322500.0 1017600.0 ;
      RECT  312300.0 1031400.0 322500.0 1017600.0 ;
      RECT  312300.0 1031400.0 322500.0 1045200.0 ;
      RECT  312300.0 1059000.0 322500.0 1045200.0 ;
      RECT  312300.0 1059000.0 322500.0 1072800.0 ;
      RECT  312300.0 1086600.0 322500.0 1072800.0 ;
      RECT  312300.0 1086600.0 322500.0 1100400.0 ;
      RECT  312300.0 1114200.0 322500.0 1100400.0 ;
      RECT  312300.0 1114200.0 322500.0 1128000.0 ;
      RECT  312300.0 1141800.0 322500.0 1128000.0 ;
      RECT  312300.0 1141800.0 322500.0 1155600.0 ;
      RECT  312300.0 1169400.0 322500.0 1155600.0 ;
      RECT  312300.0 1169400.0 322500.0 1183200.0 ;
      RECT  312300.0 1197000.0 322500.0 1183200.0 ;
      RECT  322500.0 313800.0 332700.0 327600.0 ;
      RECT  322500.0 341400.0 332700.0 327600.0 ;
      RECT  322500.0 341400.0 332700.0 355200.0 ;
      RECT  322500.0 369000.0 332700.0 355200.0 ;
      RECT  322500.0 369000.0 332700.0 382800.0 ;
      RECT  322500.0 396600.0 332700.0 382800.0 ;
      RECT  322500.0 396600.0 332700.0 410400.0 ;
      RECT  322500.0 424200.0 332700.0 410400.0 ;
      RECT  322500.0 424200.0 332700.0 438000.0 ;
      RECT  322500.0 451800.0 332700.0 438000.0 ;
      RECT  322500.0 451800.0 332700.0 465600.0 ;
      RECT  322500.0 479400.0 332700.0 465600.0 ;
      RECT  322500.0 479400.0 332700.0 493200.0 ;
      RECT  322500.0 507000.0 332700.0 493200.0 ;
      RECT  322500.0 507000.0 332700.0 520800.0 ;
      RECT  322500.0 534600.0 332700.0 520800.0 ;
      RECT  322500.0 534600.0 332700.0 548400.0 ;
      RECT  322500.0 562200.0 332700.0 548400.0 ;
      RECT  322500.0 562200.0 332700.0 576000.0 ;
      RECT  322500.0 589800.0 332700.0 576000.0 ;
      RECT  322500.0 589800.0 332700.0 603600.0 ;
      RECT  322500.0 617400.0 332700.0 603600.0 ;
      RECT  322500.0 617400.0 332700.0 631200.0 ;
      RECT  322500.0 645000.0 332700.0 631200.0 ;
      RECT  322500.0 645000.0 332700.0 658800.0 ;
      RECT  322500.0 672600.0 332700.0 658800.0 ;
      RECT  322500.0 672600.0 332700.0 686400.0 ;
      RECT  322500.0 700200.0 332700.0 686400.0 ;
      RECT  322500.0 700200.0 332700.0 714000.0 ;
      RECT  322500.0 727800.0 332700.0 714000.0 ;
      RECT  322500.0 727800.0 332700.0 741600.0 ;
      RECT  322500.0 755400.0 332700.0 741600.0 ;
      RECT  322500.0 755400.0 332700.0 769200.0 ;
      RECT  322500.0 783000.0 332700.0 769200.0 ;
      RECT  322500.0 783000.0 332700.0 796800.0 ;
      RECT  322500.0 810600.0 332700.0 796800.0 ;
      RECT  322500.0 810600.0 332700.0 824400.0 ;
      RECT  322500.0 838200.0 332700.0 824400.0 ;
      RECT  322500.0 838200.0 332700.0 852000.0 ;
      RECT  322500.0 865800.0 332700.0 852000.0 ;
      RECT  322500.0 865800.0 332700.0 879600.0 ;
      RECT  322500.0 893400.0 332700.0 879600.0 ;
      RECT  322500.0 893400.0 332700.0 907200.0 ;
      RECT  322500.0 921000.0 332700.0 907200.0 ;
      RECT  322500.0 921000.0 332700.0 934800.0 ;
      RECT  322500.0 948600.0 332700.0 934800.0 ;
      RECT  322500.0 948600.0 332700.0 962400.0 ;
      RECT  322500.0 976200.0 332700.0 962400.0 ;
      RECT  322500.0 976200.0 332700.0 990000.0 ;
      RECT  322500.0 1003800.0 332700.0 990000.0 ;
      RECT  322500.0 1003800.0 332700.0 1017600.0 ;
      RECT  322500.0 1031400.0 332700.0 1017600.0 ;
      RECT  322500.0 1031400.0 332700.0 1045200.0 ;
      RECT  322500.0 1059000.0 332700.0 1045200.0 ;
      RECT  322500.0 1059000.0 332700.0 1072800.0 ;
      RECT  322500.0 1086600.0 332700.0 1072800.0 ;
      RECT  322500.0 1086600.0 332700.0 1100400.0 ;
      RECT  322500.0 1114200.0 332700.0 1100400.0 ;
      RECT  322500.0 1114200.0 332700.0 1128000.0 ;
      RECT  322500.0 1141800.0 332700.0 1128000.0 ;
      RECT  322500.0 1141800.0 332700.0 1155600.0 ;
      RECT  322500.0 1169400.0 332700.0 1155600.0 ;
      RECT  322500.0 1169400.0 332700.0 1183200.0 ;
      RECT  322500.0 1197000.0 332700.0 1183200.0 ;
      RECT  332700.0 313800.0 342900.0 327600.0 ;
      RECT  332700.0 341400.0 342900.0 327600.0 ;
      RECT  332700.0 341400.0 342900.0 355200.0 ;
      RECT  332700.0 369000.0 342900.0 355200.0 ;
      RECT  332700.0 369000.0 342900.0 382800.0 ;
      RECT  332700.0 396600.0 342900.0 382800.0 ;
      RECT  332700.0 396600.0 342900.0 410400.0 ;
      RECT  332700.0 424200.0 342900.0 410400.0 ;
      RECT  332700.0 424200.0 342900.0 438000.0 ;
      RECT  332700.0 451800.0 342900.0 438000.0 ;
      RECT  332700.0 451800.0 342900.0 465600.0 ;
      RECT  332700.0 479400.0 342900.0 465600.0 ;
      RECT  332700.0 479400.0 342900.0 493200.0 ;
      RECT  332700.0 507000.0 342900.0 493200.0 ;
      RECT  332700.0 507000.0 342900.0 520800.0 ;
      RECT  332700.0 534600.0 342900.0 520800.0 ;
      RECT  332700.0 534600.0 342900.0 548400.0 ;
      RECT  332700.0 562200.0 342900.0 548400.0 ;
      RECT  332700.0 562200.0 342900.0 576000.0 ;
      RECT  332700.0 589800.0 342900.0 576000.0 ;
      RECT  332700.0 589800.0 342900.0 603600.0 ;
      RECT  332700.0 617400.0 342900.0 603600.0 ;
      RECT  332700.0 617400.0 342900.0 631200.0 ;
      RECT  332700.0 645000.0 342900.0 631200.0 ;
      RECT  332700.0 645000.0 342900.0 658800.0 ;
      RECT  332700.0 672600.0 342900.0 658800.0 ;
      RECT  332700.0 672600.0 342900.0 686400.0 ;
      RECT  332700.0 700200.0 342900.0 686400.0 ;
      RECT  332700.0 700200.0 342900.0 714000.0 ;
      RECT  332700.0 727800.0 342900.0 714000.0 ;
      RECT  332700.0 727800.0 342900.0 741600.0 ;
      RECT  332700.0 755400.0 342900.0 741600.0 ;
      RECT  332700.0 755400.0 342900.0 769200.0 ;
      RECT  332700.0 783000.0 342900.0 769200.0 ;
      RECT  332700.0 783000.0 342900.0 796800.0 ;
      RECT  332700.0 810600.0 342900.0 796800.0 ;
      RECT  332700.0 810600.0 342900.0 824400.0 ;
      RECT  332700.0 838200.0 342900.0 824400.0 ;
      RECT  332700.0 838200.0 342900.0 852000.0 ;
      RECT  332700.0 865800.0 342900.0 852000.0 ;
      RECT  332700.0 865800.0 342900.0 879600.0 ;
      RECT  332700.0 893400.0 342900.0 879600.0 ;
      RECT  332700.0 893400.0 342900.0 907200.0 ;
      RECT  332700.0 921000.0 342900.0 907200.0 ;
      RECT  332700.0 921000.0 342900.0 934800.0 ;
      RECT  332700.0 948600.0 342900.0 934800.0 ;
      RECT  332700.0 948600.0 342900.0 962400.0 ;
      RECT  332700.0 976200.0 342900.0 962400.0 ;
      RECT  332700.0 976200.0 342900.0 990000.0 ;
      RECT  332700.0 1003800.0 342900.0 990000.0 ;
      RECT  332700.0 1003800.0 342900.0 1017600.0 ;
      RECT  332700.0 1031400.0 342900.0 1017600.0 ;
      RECT  332700.0 1031400.0 342900.0 1045200.0 ;
      RECT  332700.0 1059000.0 342900.0 1045200.0 ;
      RECT  332700.0 1059000.0 342900.0 1072800.0 ;
      RECT  332700.0 1086600.0 342900.0 1072800.0 ;
      RECT  332700.0 1086600.0 342900.0 1100400.0 ;
      RECT  332700.0 1114200.0 342900.0 1100400.0 ;
      RECT  332700.0 1114200.0 342900.0 1128000.0 ;
      RECT  332700.0 1141800.0 342900.0 1128000.0 ;
      RECT  332700.0 1141800.0 342900.0 1155600.0 ;
      RECT  332700.0 1169400.0 342900.0 1155600.0 ;
      RECT  332700.0 1169400.0 342900.0 1183200.0 ;
      RECT  332700.0 1197000.0 342900.0 1183200.0 ;
      RECT  342900.0 313800.0 353100.0 327600.0 ;
      RECT  342900.0 341400.0 353100.0 327600.0 ;
      RECT  342900.0 341400.0 353100.0 355200.0 ;
      RECT  342900.0 369000.0 353100.0 355200.0 ;
      RECT  342900.0 369000.0 353100.0 382800.0 ;
      RECT  342900.0 396600.0 353100.0 382800.0 ;
      RECT  342900.0 396600.0 353100.0 410400.0 ;
      RECT  342900.0 424200.0 353100.0 410400.0 ;
      RECT  342900.0 424200.0 353100.0 438000.0 ;
      RECT  342900.0 451800.0 353100.0 438000.0 ;
      RECT  342900.0 451800.0 353100.0 465600.0 ;
      RECT  342900.0 479400.0 353100.0 465600.0 ;
      RECT  342900.0 479400.0 353100.0 493200.0 ;
      RECT  342900.0 507000.0 353100.0 493200.0 ;
      RECT  342900.0 507000.0 353100.0 520800.0 ;
      RECT  342900.0 534600.0 353100.0 520800.0 ;
      RECT  342900.0 534600.0 353100.0 548400.0 ;
      RECT  342900.0 562200.0 353100.0 548400.0 ;
      RECT  342900.0 562200.0 353100.0 576000.0 ;
      RECT  342900.0 589800.0 353100.0 576000.0 ;
      RECT  342900.0 589800.0 353100.0 603600.0 ;
      RECT  342900.0 617400.0 353100.0 603600.0 ;
      RECT  342900.0 617400.0 353100.0 631200.0 ;
      RECT  342900.0 645000.0 353100.0 631200.0 ;
      RECT  342900.0 645000.0 353100.0 658800.0 ;
      RECT  342900.0 672600.0 353100.0 658800.0 ;
      RECT  342900.0 672600.0 353100.0 686400.0 ;
      RECT  342900.0 700200.0 353100.0 686400.0 ;
      RECT  342900.0 700200.0 353100.0 714000.0 ;
      RECT  342900.0 727800.0 353100.0 714000.0 ;
      RECT  342900.0 727800.0 353100.0 741600.0 ;
      RECT  342900.0 755400.0 353100.0 741600.0 ;
      RECT  342900.0 755400.0 353100.0 769200.0 ;
      RECT  342900.0 783000.0 353100.0 769200.0 ;
      RECT  342900.0 783000.0 353100.0 796800.0 ;
      RECT  342900.0 810600.0 353100.0 796800.0 ;
      RECT  342900.0 810600.0 353100.0 824400.0 ;
      RECT  342900.0 838200.0 353100.0 824400.0 ;
      RECT  342900.0 838200.0 353100.0 852000.0 ;
      RECT  342900.0 865800.0 353100.0 852000.0 ;
      RECT  342900.0 865800.0 353100.0 879600.0 ;
      RECT  342900.0 893400.0 353100.0 879600.0 ;
      RECT  342900.0 893400.0 353100.0 907200.0 ;
      RECT  342900.0 921000.0 353100.0 907200.0 ;
      RECT  342900.0 921000.0 353100.0 934800.0 ;
      RECT  342900.0 948600.0 353100.0 934800.0 ;
      RECT  342900.0 948600.0 353100.0 962400.0 ;
      RECT  342900.0 976200.0 353100.0 962400.0 ;
      RECT  342900.0 976200.0 353100.0 990000.0 ;
      RECT  342900.0 1003800.0 353100.0 990000.0 ;
      RECT  342900.0 1003800.0 353100.0 1017600.0 ;
      RECT  342900.0 1031400.0 353100.0 1017600.0 ;
      RECT  342900.0 1031400.0 353100.0 1045200.0 ;
      RECT  342900.0 1059000.0 353100.0 1045200.0 ;
      RECT  342900.0 1059000.0 353100.0 1072800.0 ;
      RECT  342900.0 1086600.0 353100.0 1072800.0 ;
      RECT  342900.0 1086600.0 353100.0 1100400.0 ;
      RECT  342900.0 1114200.0 353100.0 1100400.0 ;
      RECT  342900.0 1114200.0 353100.0 1128000.0 ;
      RECT  342900.0 1141800.0 353100.0 1128000.0 ;
      RECT  342900.0 1141800.0 353100.0 1155600.0 ;
      RECT  342900.0 1169400.0 353100.0 1155600.0 ;
      RECT  342900.0 1169400.0 353100.0 1183200.0 ;
      RECT  342900.0 1197000.0 353100.0 1183200.0 ;
      RECT  353100.0 313800.0 363300.0 327600.0 ;
      RECT  353100.0 341400.0 363300.0 327600.0 ;
      RECT  353100.0 341400.0 363300.0 355200.0 ;
      RECT  353100.0 369000.0 363300.0 355200.0 ;
      RECT  353100.0 369000.0 363300.0 382800.0 ;
      RECT  353100.0 396600.0 363300.0 382800.0 ;
      RECT  353100.0 396600.0 363300.0 410400.0 ;
      RECT  353100.0 424200.0 363300.0 410400.0 ;
      RECT  353100.0 424200.0 363300.0 438000.0 ;
      RECT  353100.0 451800.0 363300.0 438000.0 ;
      RECT  353100.0 451800.0 363300.0 465600.0 ;
      RECT  353100.0 479400.0 363300.0 465600.0 ;
      RECT  353100.0 479400.0 363300.0 493200.0 ;
      RECT  353100.0 507000.0 363300.0 493200.0 ;
      RECT  353100.0 507000.0 363300.0 520800.0 ;
      RECT  353100.0 534600.0 363300.0 520800.0 ;
      RECT  353100.0 534600.0 363300.0 548400.0 ;
      RECT  353100.0 562200.0 363300.0 548400.0 ;
      RECT  353100.0 562200.0 363300.0 576000.0 ;
      RECT  353100.0 589800.0 363300.0 576000.0 ;
      RECT  353100.0 589800.0 363300.0 603600.0 ;
      RECT  353100.0 617400.0 363300.0 603600.0 ;
      RECT  353100.0 617400.0 363300.0 631200.0 ;
      RECT  353100.0 645000.0 363300.0 631200.0 ;
      RECT  353100.0 645000.0 363300.0 658800.0 ;
      RECT  353100.0 672600.0 363300.0 658800.0 ;
      RECT  353100.0 672600.0 363300.0 686400.0 ;
      RECT  353100.0 700200.0 363300.0 686400.0 ;
      RECT  353100.0 700200.0 363300.0 714000.0 ;
      RECT  353100.0 727800.0 363300.0 714000.0 ;
      RECT  353100.0 727800.0 363300.0 741600.0 ;
      RECT  353100.0 755400.0 363300.0 741600.0 ;
      RECT  353100.0 755400.0 363300.0 769200.0 ;
      RECT  353100.0 783000.0 363300.0 769200.0 ;
      RECT  353100.0 783000.0 363300.0 796800.0 ;
      RECT  353100.0 810600.0 363300.0 796800.0 ;
      RECT  353100.0 810600.0 363300.0 824400.0 ;
      RECT  353100.0 838200.0 363300.0 824400.0 ;
      RECT  353100.0 838200.0 363300.0 852000.0 ;
      RECT  353100.0 865800.0 363300.0 852000.0 ;
      RECT  353100.0 865800.0 363300.0 879600.0 ;
      RECT  353100.0 893400.0 363300.0 879600.0 ;
      RECT  353100.0 893400.0 363300.0 907200.0 ;
      RECT  353100.0 921000.0 363300.0 907200.0 ;
      RECT  353100.0 921000.0 363300.0 934800.0 ;
      RECT  353100.0 948600.0 363300.0 934800.0 ;
      RECT  353100.0 948600.0 363300.0 962400.0 ;
      RECT  353100.0 976200.0 363300.0 962400.0 ;
      RECT  353100.0 976200.0 363300.0 990000.0 ;
      RECT  353100.0 1003800.0 363300.0 990000.0 ;
      RECT  353100.0 1003800.0 363300.0 1017600.0 ;
      RECT  353100.0 1031400.0 363300.0 1017600.0 ;
      RECT  353100.0 1031400.0 363300.0 1045200.0 ;
      RECT  353100.0 1059000.0 363300.0 1045200.0 ;
      RECT  353100.0 1059000.0 363300.0 1072800.0 ;
      RECT  353100.0 1086600.0 363300.0 1072800.0 ;
      RECT  353100.0 1086600.0 363300.0 1100400.0 ;
      RECT  353100.0 1114200.0 363300.0 1100400.0 ;
      RECT  353100.0 1114200.0 363300.0 1128000.0 ;
      RECT  353100.0 1141800.0 363300.0 1128000.0 ;
      RECT  353100.0 1141800.0 363300.0 1155600.0 ;
      RECT  353100.0 1169400.0 363300.0 1155600.0 ;
      RECT  353100.0 1169400.0 363300.0 1183200.0 ;
      RECT  353100.0 1197000.0 363300.0 1183200.0 ;
      RECT  363300.0 313800.0 373500.0 327600.0 ;
      RECT  363300.0 341400.0 373500.0 327600.0 ;
      RECT  363300.0 341400.0 373500.0 355200.0 ;
      RECT  363300.0 369000.0 373500.0 355200.0 ;
      RECT  363300.0 369000.0 373500.0 382800.0 ;
      RECT  363300.0 396600.0 373500.0 382800.0 ;
      RECT  363300.0 396600.0 373500.0 410400.0 ;
      RECT  363300.0 424200.0 373500.0 410400.0 ;
      RECT  363300.0 424200.0 373500.0 438000.0 ;
      RECT  363300.0 451800.0 373500.0 438000.0 ;
      RECT  363300.0 451800.0 373500.0 465600.0 ;
      RECT  363300.0 479400.0 373500.0 465600.0 ;
      RECT  363300.0 479400.0 373500.0 493200.0 ;
      RECT  363300.0 507000.0 373500.0 493200.0 ;
      RECT  363300.0 507000.0 373500.0 520800.0 ;
      RECT  363300.0 534600.0 373500.0 520800.0 ;
      RECT  363300.0 534600.0 373500.0 548400.0 ;
      RECT  363300.0 562200.0 373500.0 548400.0 ;
      RECT  363300.0 562200.0 373500.0 576000.0 ;
      RECT  363300.0 589800.0 373500.0 576000.0 ;
      RECT  363300.0 589800.0 373500.0 603600.0 ;
      RECT  363300.0 617400.0 373500.0 603600.0 ;
      RECT  363300.0 617400.0 373500.0 631200.0 ;
      RECT  363300.0 645000.0 373500.0 631200.0 ;
      RECT  363300.0 645000.0 373500.0 658800.0 ;
      RECT  363300.0 672600.0 373500.0 658800.0 ;
      RECT  363300.0 672600.0 373500.0 686400.0 ;
      RECT  363300.0 700200.0 373500.0 686400.0 ;
      RECT  363300.0 700200.0 373500.0 714000.0 ;
      RECT  363300.0 727800.0 373500.0 714000.0 ;
      RECT  363300.0 727800.0 373500.0 741600.0 ;
      RECT  363300.0 755400.0 373500.0 741600.0 ;
      RECT  363300.0 755400.0 373500.0 769200.0 ;
      RECT  363300.0 783000.0 373500.0 769200.0 ;
      RECT  363300.0 783000.0 373500.0 796800.0 ;
      RECT  363300.0 810600.0 373500.0 796800.0 ;
      RECT  363300.0 810600.0 373500.0 824400.0 ;
      RECT  363300.0 838200.0 373500.0 824400.0 ;
      RECT  363300.0 838200.0 373500.0 852000.0 ;
      RECT  363300.0 865800.0 373500.0 852000.0 ;
      RECT  363300.0 865800.0 373500.0 879600.0 ;
      RECT  363300.0 893400.0 373500.0 879600.0 ;
      RECT  363300.0 893400.0 373500.0 907200.0 ;
      RECT  363300.0 921000.0 373500.0 907200.0 ;
      RECT  363300.0 921000.0 373500.0 934800.0 ;
      RECT  363300.0 948600.0 373500.0 934800.0 ;
      RECT  363300.0 948600.0 373500.0 962400.0 ;
      RECT  363300.0 976200.0 373500.0 962400.0 ;
      RECT  363300.0 976200.0 373500.0 990000.0 ;
      RECT  363300.0 1003800.0 373500.0 990000.0 ;
      RECT  363300.0 1003800.0 373500.0 1017600.0 ;
      RECT  363300.0 1031400.0 373500.0 1017600.0 ;
      RECT  363300.0 1031400.0 373500.0 1045200.0 ;
      RECT  363300.0 1059000.0 373500.0 1045200.0 ;
      RECT  363300.0 1059000.0 373500.0 1072800.0 ;
      RECT  363300.0 1086600.0 373500.0 1072800.0 ;
      RECT  363300.0 1086600.0 373500.0 1100400.0 ;
      RECT  363300.0 1114200.0 373500.0 1100400.0 ;
      RECT  363300.0 1114200.0 373500.0 1128000.0 ;
      RECT  363300.0 1141800.0 373500.0 1128000.0 ;
      RECT  363300.0 1141800.0 373500.0 1155600.0 ;
      RECT  363300.0 1169400.0 373500.0 1155600.0 ;
      RECT  363300.0 1169400.0 373500.0 1183200.0 ;
      RECT  363300.0 1197000.0 373500.0 1183200.0 ;
      RECT  373500.0 313800.0 383700.0 327600.0 ;
      RECT  373500.0 341400.0 383700.0 327600.0 ;
      RECT  373500.0 341400.0 383700.0 355200.0 ;
      RECT  373500.0 369000.0 383700.0 355200.0 ;
      RECT  373500.0 369000.0 383700.0 382800.0 ;
      RECT  373500.0 396600.0 383700.0 382800.0 ;
      RECT  373500.0 396600.0 383700.0 410400.0 ;
      RECT  373500.0 424200.0 383700.0 410400.0 ;
      RECT  373500.0 424200.0 383700.0 438000.0 ;
      RECT  373500.0 451800.0 383700.0 438000.0 ;
      RECT  373500.0 451800.0 383700.0 465600.0 ;
      RECT  373500.0 479400.0 383700.0 465600.0 ;
      RECT  373500.0 479400.0 383700.0 493200.0 ;
      RECT  373500.0 507000.0 383700.0 493200.0 ;
      RECT  373500.0 507000.0 383700.0 520800.0 ;
      RECT  373500.0 534600.0 383700.0 520800.0 ;
      RECT  373500.0 534600.0 383700.0 548400.0 ;
      RECT  373500.0 562200.0 383700.0 548400.0 ;
      RECT  373500.0 562200.0 383700.0 576000.0 ;
      RECT  373500.0 589800.0 383700.0 576000.0 ;
      RECT  373500.0 589800.0 383700.0 603600.0 ;
      RECT  373500.0 617400.0 383700.0 603600.0 ;
      RECT  373500.0 617400.0 383700.0 631200.0 ;
      RECT  373500.0 645000.0 383700.0 631200.0 ;
      RECT  373500.0 645000.0 383700.0 658800.0 ;
      RECT  373500.0 672600.0 383700.0 658800.0 ;
      RECT  373500.0 672600.0 383700.0 686400.0 ;
      RECT  373500.0 700200.0 383700.0 686400.0 ;
      RECT  373500.0 700200.0 383700.0 714000.0 ;
      RECT  373500.0 727800.0 383700.0 714000.0 ;
      RECT  373500.0 727800.0 383700.0 741600.0 ;
      RECT  373500.0 755400.0 383700.0 741600.0 ;
      RECT  373500.0 755400.0 383700.0 769200.0 ;
      RECT  373500.0 783000.0 383700.0 769200.0 ;
      RECT  373500.0 783000.0 383700.0 796800.0 ;
      RECT  373500.0 810600.0 383700.0 796800.0 ;
      RECT  373500.0 810600.0 383700.0 824400.0 ;
      RECT  373500.0 838200.0 383700.0 824400.0 ;
      RECT  373500.0 838200.0 383700.0 852000.0 ;
      RECT  373500.0 865800.0 383700.0 852000.0 ;
      RECT  373500.0 865800.0 383700.0 879600.0 ;
      RECT  373500.0 893400.0 383700.0 879600.0 ;
      RECT  373500.0 893400.0 383700.0 907200.0 ;
      RECT  373500.0 921000.0 383700.0 907200.0 ;
      RECT  373500.0 921000.0 383700.0 934800.0 ;
      RECT  373500.0 948600.0 383700.0 934800.0 ;
      RECT  373500.0 948600.0 383700.0 962400.0 ;
      RECT  373500.0 976200.0 383700.0 962400.0 ;
      RECT  373500.0 976200.0 383700.0 990000.0 ;
      RECT  373500.0 1003800.0 383700.0 990000.0 ;
      RECT  373500.0 1003800.0 383700.0 1017600.0 ;
      RECT  373500.0 1031400.0 383700.0 1017600.0 ;
      RECT  373500.0 1031400.0 383700.0 1045200.0 ;
      RECT  373500.0 1059000.0 383700.0 1045200.0 ;
      RECT  373500.0 1059000.0 383700.0 1072800.0 ;
      RECT  373500.0 1086600.0 383700.0 1072800.0 ;
      RECT  373500.0 1086600.0 383700.0 1100400.0 ;
      RECT  373500.0 1114200.0 383700.0 1100400.0 ;
      RECT  373500.0 1114200.0 383700.0 1128000.0 ;
      RECT  373500.0 1141800.0 383700.0 1128000.0 ;
      RECT  373500.0 1141800.0 383700.0 1155600.0 ;
      RECT  373500.0 1169400.0 383700.0 1155600.0 ;
      RECT  373500.0 1169400.0 383700.0 1183200.0 ;
      RECT  373500.0 1197000.0 383700.0 1183200.0 ;
      RECT  383700.0 313800.0 393900.0 327600.0 ;
      RECT  383700.0 341400.0 393900.0 327600.0 ;
      RECT  383700.0 341400.0 393900.0 355200.0 ;
      RECT  383700.0 369000.0 393900.0 355200.0 ;
      RECT  383700.0 369000.0 393900.0 382800.0 ;
      RECT  383700.0 396600.0 393900.0 382800.0 ;
      RECT  383700.0 396600.0 393900.0 410400.0 ;
      RECT  383700.0 424200.0 393900.0 410400.0 ;
      RECT  383700.0 424200.0 393900.0 438000.0 ;
      RECT  383700.0 451800.0 393900.0 438000.0 ;
      RECT  383700.0 451800.0 393900.0 465600.0 ;
      RECT  383700.0 479400.0 393900.0 465600.0 ;
      RECT  383700.0 479400.0 393900.0 493200.0 ;
      RECT  383700.0 507000.0 393900.0 493200.0 ;
      RECT  383700.0 507000.0 393900.0 520800.0 ;
      RECT  383700.0 534600.0 393900.0 520800.0 ;
      RECT  383700.0 534600.0 393900.0 548400.0 ;
      RECT  383700.0 562200.0 393900.0 548400.0 ;
      RECT  383700.0 562200.0 393900.0 576000.0 ;
      RECT  383700.0 589800.0 393900.0 576000.0 ;
      RECT  383700.0 589800.0 393900.0 603600.0 ;
      RECT  383700.0 617400.0 393900.0 603600.0 ;
      RECT  383700.0 617400.0 393900.0 631200.0 ;
      RECT  383700.0 645000.0 393900.0 631200.0 ;
      RECT  383700.0 645000.0 393900.0 658800.0 ;
      RECT  383700.0 672600.0 393900.0 658800.0 ;
      RECT  383700.0 672600.0 393900.0 686400.0 ;
      RECT  383700.0 700200.0 393900.0 686400.0 ;
      RECT  383700.0 700200.0 393900.0 714000.0 ;
      RECT  383700.0 727800.0 393900.0 714000.0 ;
      RECT  383700.0 727800.0 393900.0 741600.0 ;
      RECT  383700.0 755400.0 393900.0 741600.0 ;
      RECT  383700.0 755400.0 393900.0 769200.0 ;
      RECT  383700.0 783000.0 393900.0 769200.0 ;
      RECT  383700.0 783000.0 393900.0 796800.0 ;
      RECT  383700.0 810600.0 393900.0 796800.0 ;
      RECT  383700.0 810600.0 393900.0 824400.0 ;
      RECT  383700.0 838200.0 393900.0 824400.0 ;
      RECT  383700.0 838200.0 393900.0 852000.0 ;
      RECT  383700.0 865800.0 393900.0 852000.0 ;
      RECT  383700.0 865800.0 393900.0 879600.0 ;
      RECT  383700.0 893400.0 393900.0 879600.0 ;
      RECT  383700.0 893400.0 393900.0 907200.0 ;
      RECT  383700.0 921000.0 393900.0 907200.0 ;
      RECT  383700.0 921000.0 393900.0 934800.0 ;
      RECT  383700.0 948600.0 393900.0 934800.0 ;
      RECT  383700.0 948600.0 393900.0 962400.0 ;
      RECT  383700.0 976200.0 393900.0 962400.0 ;
      RECT  383700.0 976200.0 393900.0 990000.0 ;
      RECT  383700.0 1003800.0 393900.0 990000.0 ;
      RECT  383700.0 1003800.0 393900.0 1017600.0 ;
      RECT  383700.0 1031400.0 393900.0 1017600.0 ;
      RECT  383700.0 1031400.0 393900.0 1045200.0 ;
      RECT  383700.0 1059000.0 393900.0 1045200.0 ;
      RECT  383700.0 1059000.0 393900.0 1072800.0 ;
      RECT  383700.0 1086600.0 393900.0 1072800.0 ;
      RECT  383700.0 1086600.0 393900.0 1100400.0 ;
      RECT  383700.0 1114200.0 393900.0 1100400.0 ;
      RECT  383700.0 1114200.0 393900.0 1128000.0 ;
      RECT  383700.0 1141800.0 393900.0 1128000.0 ;
      RECT  383700.0 1141800.0 393900.0 1155600.0 ;
      RECT  383700.0 1169400.0 393900.0 1155600.0 ;
      RECT  383700.0 1169400.0 393900.0 1183200.0 ;
      RECT  383700.0 1197000.0 393900.0 1183200.0 ;
      RECT  393900.0 313800.0 404100.0 327600.0 ;
      RECT  393900.0 341400.0 404100.0 327600.0 ;
      RECT  393900.0 341400.0 404100.0 355200.0 ;
      RECT  393900.0 369000.0 404100.0 355200.0 ;
      RECT  393900.0 369000.0 404100.0 382800.0 ;
      RECT  393900.0 396600.0 404100.0 382800.0 ;
      RECT  393900.0 396600.0 404100.0 410400.0 ;
      RECT  393900.0 424200.0 404100.0 410400.0 ;
      RECT  393900.0 424200.0 404100.0 438000.0 ;
      RECT  393900.0 451800.0 404100.0 438000.0 ;
      RECT  393900.0 451800.0 404100.0 465600.0 ;
      RECT  393900.0 479400.0 404100.0 465600.0 ;
      RECT  393900.0 479400.0 404100.0 493200.0 ;
      RECT  393900.0 507000.0 404100.0 493200.0 ;
      RECT  393900.0 507000.0 404100.0 520800.0 ;
      RECT  393900.0 534600.0 404100.0 520800.0 ;
      RECT  393900.0 534600.0 404100.0 548400.0 ;
      RECT  393900.0 562200.0 404100.0 548400.0 ;
      RECT  393900.0 562200.0 404100.0 576000.0 ;
      RECT  393900.0 589800.0 404100.0 576000.0 ;
      RECT  393900.0 589800.0 404100.0 603600.0 ;
      RECT  393900.0 617400.0 404100.0 603600.0 ;
      RECT  393900.0 617400.0 404100.0 631200.0 ;
      RECT  393900.0 645000.0 404100.0 631200.0 ;
      RECT  393900.0 645000.0 404100.0 658800.0 ;
      RECT  393900.0 672600.0 404100.0 658800.0 ;
      RECT  393900.0 672600.0 404100.0 686400.0 ;
      RECT  393900.0 700200.0 404100.0 686400.0 ;
      RECT  393900.0 700200.0 404100.0 714000.0 ;
      RECT  393900.0 727800.0 404100.0 714000.0 ;
      RECT  393900.0 727800.0 404100.0 741600.0 ;
      RECT  393900.0 755400.0 404100.0 741600.0 ;
      RECT  393900.0 755400.0 404100.0 769200.0 ;
      RECT  393900.0 783000.0 404100.0 769200.0 ;
      RECT  393900.0 783000.0 404100.0 796800.0 ;
      RECT  393900.0 810600.0 404100.0 796800.0 ;
      RECT  393900.0 810600.0 404100.0 824400.0 ;
      RECT  393900.0 838200.0 404100.0 824400.0 ;
      RECT  393900.0 838200.0 404100.0 852000.0 ;
      RECT  393900.0 865800.0 404100.0 852000.0 ;
      RECT  393900.0 865800.0 404100.0 879600.0 ;
      RECT  393900.0 893400.0 404100.0 879600.0 ;
      RECT  393900.0 893400.0 404100.0 907200.0 ;
      RECT  393900.0 921000.0 404100.0 907200.0 ;
      RECT  393900.0 921000.0 404100.0 934800.0 ;
      RECT  393900.0 948600.0 404100.0 934800.0 ;
      RECT  393900.0 948600.0 404100.0 962400.0 ;
      RECT  393900.0 976200.0 404100.0 962400.0 ;
      RECT  393900.0 976200.0 404100.0 990000.0 ;
      RECT  393900.0 1003800.0 404100.0 990000.0 ;
      RECT  393900.0 1003800.0 404100.0 1017600.0 ;
      RECT  393900.0 1031400.0 404100.0 1017600.0 ;
      RECT  393900.0 1031400.0 404100.0 1045200.0 ;
      RECT  393900.0 1059000.0 404100.0 1045200.0 ;
      RECT  393900.0 1059000.0 404100.0 1072800.0 ;
      RECT  393900.0 1086600.0 404100.0 1072800.0 ;
      RECT  393900.0 1086600.0 404100.0 1100400.0 ;
      RECT  393900.0 1114200.0 404100.0 1100400.0 ;
      RECT  393900.0 1114200.0 404100.0 1128000.0 ;
      RECT  393900.0 1141800.0 404100.0 1128000.0 ;
      RECT  393900.0 1141800.0 404100.0 1155600.0 ;
      RECT  393900.0 1169400.0 404100.0 1155600.0 ;
      RECT  393900.0 1169400.0 404100.0 1183200.0 ;
      RECT  393900.0 1197000.0 404100.0 1183200.0 ;
      RECT  404100.0 313800.0 414300.0 327600.0 ;
      RECT  404100.0 341400.0 414300.0 327600.0 ;
      RECT  404100.0 341400.0 414300.0 355200.0 ;
      RECT  404100.0 369000.0 414300.0 355200.0 ;
      RECT  404100.0 369000.0 414300.0 382800.0 ;
      RECT  404100.0 396600.0 414300.0 382800.0 ;
      RECT  404100.0 396600.0 414300.0 410400.0 ;
      RECT  404100.0 424200.0 414300.0 410400.0 ;
      RECT  404100.0 424200.0 414300.0 438000.0 ;
      RECT  404100.0 451800.0 414300.0 438000.0 ;
      RECT  404100.0 451800.0 414300.0 465600.0 ;
      RECT  404100.0 479400.0 414300.0 465600.0 ;
      RECT  404100.0 479400.0 414300.0 493200.0 ;
      RECT  404100.0 507000.0 414300.0 493200.0 ;
      RECT  404100.0 507000.0 414300.0 520800.0 ;
      RECT  404100.0 534600.0 414300.0 520800.0 ;
      RECT  404100.0 534600.0 414300.0 548400.0 ;
      RECT  404100.0 562200.0 414300.0 548400.0 ;
      RECT  404100.0 562200.0 414300.0 576000.0 ;
      RECT  404100.0 589800.0 414300.0 576000.0 ;
      RECT  404100.0 589800.0 414300.0 603600.0 ;
      RECT  404100.0 617400.0 414300.0 603600.0 ;
      RECT  404100.0 617400.0 414300.0 631200.0 ;
      RECT  404100.0 645000.0 414300.0 631200.0 ;
      RECT  404100.0 645000.0 414300.0 658800.0 ;
      RECT  404100.0 672600.0 414300.0 658800.0 ;
      RECT  404100.0 672600.0 414300.0 686400.0 ;
      RECT  404100.0 700200.0 414300.0 686400.0 ;
      RECT  404100.0 700200.0 414300.0 714000.0 ;
      RECT  404100.0 727800.0 414300.0 714000.0 ;
      RECT  404100.0 727800.0 414300.0 741600.0 ;
      RECT  404100.0 755400.0 414300.0 741600.0 ;
      RECT  404100.0 755400.0 414300.0 769200.0 ;
      RECT  404100.0 783000.0 414300.0 769200.0 ;
      RECT  404100.0 783000.0 414300.0 796800.0 ;
      RECT  404100.0 810600.0 414300.0 796800.0 ;
      RECT  404100.0 810600.0 414300.0 824400.0 ;
      RECT  404100.0 838200.0 414300.0 824400.0 ;
      RECT  404100.0 838200.0 414300.0 852000.0 ;
      RECT  404100.0 865800.0 414300.0 852000.0 ;
      RECT  404100.0 865800.0 414300.0 879600.0 ;
      RECT  404100.0 893400.0 414300.0 879600.0 ;
      RECT  404100.0 893400.0 414300.0 907200.0 ;
      RECT  404100.0 921000.0 414300.0 907200.0 ;
      RECT  404100.0 921000.0 414300.0 934800.0 ;
      RECT  404100.0 948600.0 414300.0 934800.0 ;
      RECT  404100.0 948600.0 414300.0 962400.0 ;
      RECT  404100.0 976200.0 414300.0 962400.0 ;
      RECT  404100.0 976200.0 414300.0 990000.0 ;
      RECT  404100.0 1003800.0 414300.0 990000.0 ;
      RECT  404100.0 1003800.0 414300.0 1017600.0 ;
      RECT  404100.0 1031400.0 414300.0 1017600.0 ;
      RECT  404100.0 1031400.0 414300.0 1045200.0 ;
      RECT  404100.0 1059000.0 414300.0 1045200.0 ;
      RECT  404100.0 1059000.0 414300.0 1072800.0 ;
      RECT  404100.0 1086600.0 414300.0 1072800.0 ;
      RECT  404100.0 1086600.0 414300.0 1100400.0 ;
      RECT  404100.0 1114200.0 414300.0 1100400.0 ;
      RECT  404100.0 1114200.0 414300.0 1128000.0 ;
      RECT  404100.0 1141800.0 414300.0 1128000.0 ;
      RECT  404100.0 1141800.0 414300.0 1155600.0 ;
      RECT  404100.0 1169400.0 414300.0 1155600.0 ;
      RECT  404100.0 1169400.0 414300.0 1183200.0 ;
      RECT  404100.0 1197000.0 414300.0 1183200.0 ;
      RECT  414300.0 313800.0 424500.0 327600.0 ;
      RECT  414300.0 341400.0 424500.0 327600.0 ;
      RECT  414300.0 341400.0 424500.0 355200.0 ;
      RECT  414300.0 369000.0 424500.0 355200.0 ;
      RECT  414300.0 369000.0 424500.0 382800.0 ;
      RECT  414300.0 396600.0 424500.0 382800.0 ;
      RECT  414300.0 396600.0 424500.0 410400.0 ;
      RECT  414300.0 424200.0 424500.0 410400.0 ;
      RECT  414300.0 424200.0 424500.0 438000.0 ;
      RECT  414300.0 451800.0 424500.0 438000.0 ;
      RECT  414300.0 451800.0 424500.0 465600.0 ;
      RECT  414300.0 479400.0 424500.0 465600.0 ;
      RECT  414300.0 479400.0 424500.0 493200.0 ;
      RECT  414300.0 507000.0 424500.0 493200.0 ;
      RECT  414300.0 507000.0 424500.0 520800.0 ;
      RECT  414300.0 534600.0 424500.0 520800.0 ;
      RECT  414300.0 534600.0 424500.0 548400.0 ;
      RECT  414300.0 562200.0 424500.0 548400.0 ;
      RECT  414300.0 562200.0 424500.0 576000.0 ;
      RECT  414300.0 589800.0 424500.0 576000.0 ;
      RECT  414300.0 589800.0 424500.0 603600.0 ;
      RECT  414300.0 617400.0 424500.0 603600.0 ;
      RECT  414300.0 617400.0 424500.0 631200.0 ;
      RECT  414300.0 645000.0 424500.0 631200.0 ;
      RECT  414300.0 645000.0 424500.0 658800.0 ;
      RECT  414300.0 672600.0 424500.0 658800.0 ;
      RECT  414300.0 672600.0 424500.0 686400.0 ;
      RECT  414300.0 700200.0 424500.0 686400.0 ;
      RECT  414300.0 700200.0 424500.0 714000.0 ;
      RECT  414300.0 727800.0 424500.0 714000.0 ;
      RECT  414300.0 727800.0 424500.0 741600.0 ;
      RECT  414300.0 755400.0 424500.0 741600.0 ;
      RECT  414300.0 755400.0 424500.0 769200.0 ;
      RECT  414300.0 783000.0 424500.0 769200.0 ;
      RECT  414300.0 783000.0 424500.0 796800.0 ;
      RECT  414300.0 810600.0 424500.0 796800.0 ;
      RECT  414300.0 810600.0 424500.0 824400.0 ;
      RECT  414300.0 838200.0 424500.0 824400.0 ;
      RECT  414300.0 838200.0 424500.0 852000.0 ;
      RECT  414300.0 865800.0 424500.0 852000.0 ;
      RECT  414300.0 865800.0 424500.0 879600.0 ;
      RECT  414300.0 893400.0 424500.0 879600.0 ;
      RECT  414300.0 893400.0 424500.0 907200.0 ;
      RECT  414300.0 921000.0 424500.0 907200.0 ;
      RECT  414300.0 921000.0 424500.0 934800.0 ;
      RECT  414300.0 948600.0 424500.0 934800.0 ;
      RECT  414300.0 948600.0 424500.0 962400.0 ;
      RECT  414300.0 976200.0 424500.0 962400.0 ;
      RECT  414300.0 976200.0 424500.0 990000.0 ;
      RECT  414300.0 1003800.0 424500.0 990000.0 ;
      RECT  414300.0 1003800.0 424500.0 1017600.0 ;
      RECT  414300.0 1031400.0 424500.0 1017600.0 ;
      RECT  414300.0 1031400.0 424500.0 1045200.0 ;
      RECT  414300.0 1059000.0 424500.0 1045200.0 ;
      RECT  414300.0 1059000.0 424500.0 1072800.0 ;
      RECT  414300.0 1086600.0 424500.0 1072800.0 ;
      RECT  414300.0 1086600.0 424500.0 1100400.0 ;
      RECT  414300.0 1114200.0 424500.0 1100400.0 ;
      RECT  414300.0 1114200.0 424500.0 1128000.0 ;
      RECT  414300.0 1141800.0 424500.0 1128000.0 ;
      RECT  414300.0 1141800.0 424500.0 1155600.0 ;
      RECT  414300.0 1169400.0 424500.0 1155600.0 ;
      RECT  414300.0 1169400.0 424500.0 1183200.0 ;
      RECT  414300.0 1197000.0 424500.0 1183200.0 ;
      RECT  424500.0 313800.0 434700.0 327600.0 ;
      RECT  424500.0 341400.0 434700.0 327600.0 ;
      RECT  424500.0 341400.0 434700.0 355200.0 ;
      RECT  424500.0 369000.0 434700.0 355200.0 ;
      RECT  424500.0 369000.0 434700.0 382800.0 ;
      RECT  424500.0 396600.0 434700.0 382800.0 ;
      RECT  424500.0 396600.0 434700.0 410400.0 ;
      RECT  424500.0 424200.0 434700.0 410400.0 ;
      RECT  424500.0 424200.0 434700.0 438000.0 ;
      RECT  424500.0 451800.0 434700.0 438000.0 ;
      RECT  424500.0 451800.0 434700.0 465600.0 ;
      RECT  424500.0 479400.0 434700.0 465600.0 ;
      RECT  424500.0 479400.0 434700.0 493200.0 ;
      RECT  424500.0 507000.0 434700.0 493200.0 ;
      RECT  424500.0 507000.0 434700.0 520800.0 ;
      RECT  424500.0 534600.0 434700.0 520800.0 ;
      RECT  424500.0 534600.0 434700.0 548400.0 ;
      RECT  424500.0 562200.0 434700.0 548400.0 ;
      RECT  424500.0 562200.0 434700.0 576000.0 ;
      RECT  424500.0 589800.0 434700.0 576000.0 ;
      RECT  424500.0 589800.0 434700.0 603600.0 ;
      RECT  424500.0 617400.0 434700.0 603600.0 ;
      RECT  424500.0 617400.0 434700.0 631200.0 ;
      RECT  424500.0 645000.0 434700.0 631200.0 ;
      RECT  424500.0 645000.0 434700.0 658800.0 ;
      RECT  424500.0 672600.0 434700.0 658800.0 ;
      RECT  424500.0 672600.0 434700.0 686400.0 ;
      RECT  424500.0 700200.0 434700.0 686400.0 ;
      RECT  424500.0 700200.0 434700.0 714000.0 ;
      RECT  424500.0 727800.0 434700.0 714000.0 ;
      RECT  424500.0 727800.0 434700.0 741600.0 ;
      RECT  424500.0 755400.0 434700.0 741600.0 ;
      RECT  424500.0 755400.0 434700.0 769200.0 ;
      RECT  424500.0 783000.0 434700.0 769200.0 ;
      RECT  424500.0 783000.0 434700.0 796800.0 ;
      RECT  424500.0 810600.0 434700.0 796800.0 ;
      RECT  424500.0 810600.0 434700.0 824400.0 ;
      RECT  424500.0 838200.0 434700.0 824400.0 ;
      RECT  424500.0 838200.0 434700.0 852000.0 ;
      RECT  424500.0 865800.0 434700.0 852000.0 ;
      RECT  424500.0 865800.0 434700.0 879600.0 ;
      RECT  424500.0 893400.0 434700.0 879600.0 ;
      RECT  424500.0 893400.0 434700.0 907200.0 ;
      RECT  424500.0 921000.0 434700.0 907200.0 ;
      RECT  424500.0 921000.0 434700.0 934800.0 ;
      RECT  424500.0 948600.0 434700.0 934800.0 ;
      RECT  424500.0 948600.0 434700.0 962400.0 ;
      RECT  424500.0 976200.0 434700.0 962400.0 ;
      RECT  424500.0 976200.0 434700.0 990000.0 ;
      RECT  424500.0 1003800.0 434700.0 990000.0 ;
      RECT  424500.0 1003800.0 434700.0 1017600.0 ;
      RECT  424500.0 1031400.0 434700.0 1017600.0 ;
      RECT  424500.0 1031400.0 434700.0 1045200.0 ;
      RECT  424500.0 1059000.0 434700.0 1045200.0 ;
      RECT  424500.0 1059000.0 434700.0 1072800.0 ;
      RECT  424500.0 1086600.0 434700.0 1072800.0 ;
      RECT  424500.0 1086600.0 434700.0 1100400.0 ;
      RECT  424500.0 1114200.0 434700.0 1100400.0 ;
      RECT  424500.0 1114200.0 434700.0 1128000.0 ;
      RECT  424500.0 1141800.0 434700.0 1128000.0 ;
      RECT  424500.0 1141800.0 434700.0 1155600.0 ;
      RECT  424500.0 1169400.0 434700.0 1155600.0 ;
      RECT  424500.0 1169400.0 434700.0 1183200.0 ;
      RECT  424500.0 1197000.0 434700.0 1183200.0 ;
      RECT  434700.0 313800.0 444900.0 327600.0 ;
      RECT  434700.0 341400.0 444900.0 327600.0 ;
      RECT  434700.0 341400.0 444900.0 355200.0 ;
      RECT  434700.0 369000.0 444900.0 355200.0 ;
      RECT  434700.0 369000.0 444900.0 382800.0 ;
      RECT  434700.0 396600.0 444900.0 382800.0 ;
      RECT  434700.0 396600.0 444900.0 410400.0 ;
      RECT  434700.0 424200.0 444900.0 410400.0 ;
      RECT  434700.0 424200.0 444900.0 438000.0 ;
      RECT  434700.0 451800.0 444900.0 438000.0 ;
      RECT  434700.0 451800.0 444900.0 465600.0 ;
      RECT  434700.0 479400.0 444900.0 465600.0 ;
      RECT  434700.0 479400.0 444900.0 493200.0 ;
      RECT  434700.0 507000.0 444900.0 493200.0 ;
      RECT  434700.0 507000.0 444900.0 520800.0 ;
      RECT  434700.0 534600.0 444900.0 520800.0 ;
      RECT  434700.0 534600.0 444900.0 548400.0 ;
      RECT  434700.0 562200.0 444900.0 548400.0 ;
      RECT  434700.0 562200.0 444900.0 576000.0 ;
      RECT  434700.0 589800.0 444900.0 576000.0 ;
      RECT  434700.0 589800.0 444900.0 603600.0 ;
      RECT  434700.0 617400.0 444900.0 603600.0 ;
      RECT  434700.0 617400.0 444900.0 631200.0 ;
      RECT  434700.0 645000.0 444900.0 631200.0 ;
      RECT  434700.0 645000.0 444900.0 658800.0 ;
      RECT  434700.0 672600.0 444900.0 658800.0 ;
      RECT  434700.0 672600.0 444900.0 686400.0 ;
      RECT  434700.0 700200.0 444900.0 686400.0 ;
      RECT  434700.0 700200.0 444900.0 714000.0 ;
      RECT  434700.0 727800.0 444900.0 714000.0 ;
      RECT  434700.0 727800.0 444900.0 741600.0 ;
      RECT  434700.0 755400.0 444900.0 741600.0 ;
      RECT  434700.0 755400.0 444900.0 769200.0 ;
      RECT  434700.0 783000.0 444900.0 769200.0 ;
      RECT  434700.0 783000.0 444900.0 796800.0 ;
      RECT  434700.0 810600.0 444900.0 796800.0 ;
      RECT  434700.0 810600.0 444900.0 824400.0 ;
      RECT  434700.0 838200.0 444900.0 824400.0 ;
      RECT  434700.0 838200.0 444900.0 852000.0 ;
      RECT  434700.0 865800.0 444900.0 852000.0 ;
      RECT  434700.0 865800.0 444900.0 879600.0 ;
      RECT  434700.0 893400.0 444900.0 879600.0 ;
      RECT  434700.0 893400.0 444900.0 907200.0 ;
      RECT  434700.0 921000.0 444900.0 907200.0 ;
      RECT  434700.0 921000.0 444900.0 934800.0 ;
      RECT  434700.0 948600.0 444900.0 934800.0 ;
      RECT  434700.0 948600.0 444900.0 962400.0 ;
      RECT  434700.0 976200.0 444900.0 962400.0 ;
      RECT  434700.0 976200.0 444900.0 990000.0 ;
      RECT  434700.0 1003800.0 444900.0 990000.0 ;
      RECT  434700.0 1003800.0 444900.0 1017600.0 ;
      RECT  434700.0 1031400.0 444900.0 1017600.0 ;
      RECT  434700.0 1031400.0 444900.0 1045200.0 ;
      RECT  434700.0 1059000.0 444900.0 1045200.0 ;
      RECT  434700.0 1059000.0 444900.0 1072800.0 ;
      RECT  434700.0 1086600.0 444900.0 1072800.0 ;
      RECT  434700.0 1086600.0 444900.0 1100400.0 ;
      RECT  434700.0 1114200.0 444900.0 1100400.0 ;
      RECT  434700.0 1114200.0 444900.0 1128000.0 ;
      RECT  434700.0 1141800.0 444900.0 1128000.0 ;
      RECT  434700.0 1141800.0 444900.0 1155600.0 ;
      RECT  434700.0 1169400.0 444900.0 1155600.0 ;
      RECT  434700.0 1169400.0 444900.0 1183200.0 ;
      RECT  434700.0 1197000.0 444900.0 1183200.0 ;
      RECT  444900.0 313800.0 455100.0 327600.0 ;
      RECT  444900.0 341400.0 455100.0 327600.0 ;
      RECT  444900.0 341400.0 455100.0 355200.0 ;
      RECT  444900.0 369000.0 455100.0 355200.0 ;
      RECT  444900.0 369000.0 455100.0 382800.0 ;
      RECT  444900.0 396600.0 455100.0 382800.0 ;
      RECT  444900.0 396600.0 455100.0 410400.0 ;
      RECT  444900.0 424200.0 455100.0 410400.0 ;
      RECT  444900.0 424200.0 455100.0 438000.0 ;
      RECT  444900.0 451800.0 455100.0 438000.0 ;
      RECT  444900.0 451800.0 455100.0 465600.0 ;
      RECT  444900.0 479400.0 455100.0 465600.0 ;
      RECT  444900.0 479400.0 455100.0 493200.0 ;
      RECT  444900.0 507000.0 455100.0 493200.0 ;
      RECT  444900.0 507000.0 455100.0 520800.0 ;
      RECT  444900.0 534600.0 455100.0 520800.0 ;
      RECT  444900.0 534600.0 455100.0 548400.0 ;
      RECT  444900.0 562200.0 455100.0 548400.0 ;
      RECT  444900.0 562200.0 455100.0 576000.0 ;
      RECT  444900.0 589800.0 455100.0 576000.0 ;
      RECT  444900.0 589800.0 455100.0 603600.0 ;
      RECT  444900.0 617400.0 455100.0 603600.0 ;
      RECT  444900.0 617400.0 455100.0 631200.0 ;
      RECT  444900.0 645000.0 455100.0 631200.0 ;
      RECT  444900.0 645000.0 455100.0 658800.0 ;
      RECT  444900.0 672600.0 455100.0 658800.0 ;
      RECT  444900.0 672600.0 455100.0 686400.0 ;
      RECT  444900.0 700200.0 455100.0 686400.0 ;
      RECT  444900.0 700200.0 455100.0 714000.0 ;
      RECT  444900.0 727800.0 455100.0 714000.0 ;
      RECT  444900.0 727800.0 455100.0 741600.0 ;
      RECT  444900.0 755400.0 455100.0 741600.0 ;
      RECT  444900.0 755400.0 455100.0 769200.0 ;
      RECT  444900.0 783000.0 455100.0 769200.0 ;
      RECT  444900.0 783000.0 455100.0 796800.0 ;
      RECT  444900.0 810600.0 455100.0 796800.0 ;
      RECT  444900.0 810600.0 455100.0 824400.0 ;
      RECT  444900.0 838200.0 455100.0 824400.0 ;
      RECT  444900.0 838200.0 455100.0 852000.0 ;
      RECT  444900.0 865800.0 455100.0 852000.0 ;
      RECT  444900.0 865800.0 455100.0 879600.0 ;
      RECT  444900.0 893400.0 455100.0 879600.0 ;
      RECT  444900.0 893400.0 455100.0 907200.0 ;
      RECT  444900.0 921000.0 455100.0 907200.0 ;
      RECT  444900.0 921000.0 455100.0 934800.0 ;
      RECT  444900.0 948600.0 455100.0 934800.0 ;
      RECT  444900.0 948600.0 455100.0 962400.0 ;
      RECT  444900.0 976200.0 455100.0 962400.0 ;
      RECT  444900.0 976200.0 455100.0 990000.0 ;
      RECT  444900.0 1003800.0 455100.0 990000.0 ;
      RECT  444900.0 1003800.0 455100.0 1017600.0 ;
      RECT  444900.0 1031400.0 455100.0 1017600.0 ;
      RECT  444900.0 1031400.0 455100.0 1045200.0 ;
      RECT  444900.0 1059000.0 455100.0 1045200.0 ;
      RECT  444900.0 1059000.0 455100.0 1072800.0 ;
      RECT  444900.0 1086600.0 455100.0 1072800.0 ;
      RECT  444900.0 1086600.0 455100.0 1100400.0 ;
      RECT  444900.0 1114200.0 455100.0 1100400.0 ;
      RECT  444900.0 1114200.0 455100.0 1128000.0 ;
      RECT  444900.0 1141800.0 455100.0 1128000.0 ;
      RECT  444900.0 1141800.0 455100.0 1155600.0 ;
      RECT  444900.0 1169400.0 455100.0 1155600.0 ;
      RECT  444900.0 1169400.0 455100.0 1183200.0 ;
      RECT  444900.0 1197000.0 455100.0 1183200.0 ;
      RECT  455100.0 313800.0 465300.0 327600.0 ;
      RECT  455100.0 341400.0 465300.0 327600.0 ;
      RECT  455100.0 341400.0 465300.0 355200.0 ;
      RECT  455100.0 369000.0 465300.0 355200.0 ;
      RECT  455100.0 369000.0 465300.0 382800.0 ;
      RECT  455100.0 396600.0 465300.0 382800.0 ;
      RECT  455100.0 396600.0 465300.0 410400.0 ;
      RECT  455100.0 424200.0 465300.0 410400.0 ;
      RECT  455100.0 424200.0 465300.0 438000.0 ;
      RECT  455100.0 451800.0 465300.0 438000.0 ;
      RECT  455100.0 451800.0 465300.0 465600.0 ;
      RECT  455100.0 479400.0 465300.0 465600.0 ;
      RECT  455100.0 479400.0 465300.0 493200.0 ;
      RECT  455100.0 507000.0 465300.0 493200.0 ;
      RECT  455100.0 507000.0 465300.0 520800.0 ;
      RECT  455100.0 534600.0 465300.0 520800.0 ;
      RECT  455100.0 534600.0 465300.0 548400.0 ;
      RECT  455100.0 562200.0 465300.0 548400.0 ;
      RECT  455100.0 562200.0 465300.0 576000.0 ;
      RECT  455100.0 589800.0 465300.0 576000.0 ;
      RECT  455100.0 589800.0 465300.0 603600.0 ;
      RECT  455100.0 617400.0 465300.0 603600.0 ;
      RECT  455100.0 617400.0 465300.0 631200.0 ;
      RECT  455100.0 645000.0 465300.0 631200.0 ;
      RECT  455100.0 645000.0 465300.0 658800.0 ;
      RECT  455100.0 672600.0 465300.0 658800.0 ;
      RECT  455100.0 672600.0 465300.0 686400.0 ;
      RECT  455100.0 700200.0 465300.0 686400.0 ;
      RECT  455100.0 700200.0 465300.0 714000.0 ;
      RECT  455100.0 727800.0 465300.0 714000.0 ;
      RECT  455100.0 727800.0 465300.0 741600.0 ;
      RECT  455100.0 755400.0 465300.0 741600.0 ;
      RECT  455100.0 755400.0 465300.0 769200.0 ;
      RECT  455100.0 783000.0 465300.0 769200.0 ;
      RECT  455100.0 783000.0 465300.0 796800.0 ;
      RECT  455100.0 810600.0 465300.0 796800.0 ;
      RECT  455100.0 810600.0 465300.0 824400.0 ;
      RECT  455100.0 838200.0 465300.0 824400.0 ;
      RECT  455100.0 838200.0 465300.0 852000.0 ;
      RECT  455100.0 865800.0 465300.0 852000.0 ;
      RECT  455100.0 865800.0 465300.0 879600.0 ;
      RECT  455100.0 893400.0 465300.0 879600.0 ;
      RECT  455100.0 893400.0 465300.0 907200.0 ;
      RECT  455100.0 921000.0 465300.0 907200.0 ;
      RECT  455100.0 921000.0 465300.0 934800.0 ;
      RECT  455100.0 948600.0 465300.0 934800.0 ;
      RECT  455100.0 948600.0 465300.0 962400.0 ;
      RECT  455100.0 976200.0 465300.0 962400.0 ;
      RECT  455100.0 976200.0 465300.0 990000.0 ;
      RECT  455100.0 1003800.0 465300.0 990000.0 ;
      RECT  455100.0 1003800.0 465300.0 1017600.0 ;
      RECT  455100.0 1031400.0 465300.0 1017600.0 ;
      RECT  455100.0 1031400.0 465300.0 1045200.0 ;
      RECT  455100.0 1059000.0 465300.0 1045200.0 ;
      RECT  455100.0 1059000.0 465300.0 1072800.0 ;
      RECT  455100.0 1086600.0 465300.0 1072800.0 ;
      RECT  455100.0 1086600.0 465300.0 1100400.0 ;
      RECT  455100.0 1114200.0 465300.0 1100400.0 ;
      RECT  455100.0 1114200.0 465300.0 1128000.0 ;
      RECT  455100.0 1141800.0 465300.0 1128000.0 ;
      RECT  455100.0 1141800.0 465300.0 1155600.0 ;
      RECT  455100.0 1169400.0 465300.0 1155600.0 ;
      RECT  455100.0 1169400.0 465300.0 1183200.0 ;
      RECT  455100.0 1197000.0 465300.0 1183200.0 ;
      RECT  465300.0 313800.0 475500.0 327600.0 ;
      RECT  465300.0 341400.0 475500.0 327600.0 ;
      RECT  465300.0 341400.0 475500.0 355200.0 ;
      RECT  465300.0 369000.0 475500.0 355200.0 ;
      RECT  465300.0 369000.0 475500.0 382800.0 ;
      RECT  465300.0 396600.0 475500.0 382800.0 ;
      RECT  465300.0 396600.0 475500.0 410400.0 ;
      RECT  465300.0 424200.0 475500.0 410400.0 ;
      RECT  465300.0 424200.0 475500.0 438000.0 ;
      RECT  465300.0 451800.0 475500.0 438000.0 ;
      RECT  465300.0 451800.0 475500.0 465600.0 ;
      RECT  465300.0 479400.0 475500.0 465600.0 ;
      RECT  465300.0 479400.0 475500.0 493200.0 ;
      RECT  465300.0 507000.0 475500.0 493200.0 ;
      RECT  465300.0 507000.0 475500.0 520800.0 ;
      RECT  465300.0 534600.0 475500.0 520800.0 ;
      RECT  465300.0 534600.0 475500.0 548400.0 ;
      RECT  465300.0 562200.0 475500.0 548400.0 ;
      RECT  465300.0 562200.0 475500.0 576000.0 ;
      RECT  465300.0 589800.0 475500.0 576000.0 ;
      RECT  465300.0 589800.0 475500.0 603600.0 ;
      RECT  465300.0 617400.0 475500.0 603600.0 ;
      RECT  465300.0 617400.0 475500.0 631200.0 ;
      RECT  465300.0 645000.0 475500.0 631200.0 ;
      RECT  465300.0 645000.0 475500.0 658800.0 ;
      RECT  465300.0 672600.0 475500.0 658800.0 ;
      RECT  465300.0 672600.0 475500.0 686400.0 ;
      RECT  465300.0 700200.0 475500.0 686400.0 ;
      RECT  465300.0 700200.0 475500.0 714000.0 ;
      RECT  465300.0 727800.0 475500.0 714000.0 ;
      RECT  465300.0 727800.0 475500.0 741600.0 ;
      RECT  465300.0 755400.0 475500.0 741600.0 ;
      RECT  465300.0 755400.0 475500.0 769200.0 ;
      RECT  465300.0 783000.0 475500.0 769200.0 ;
      RECT  465300.0 783000.0 475500.0 796800.0 ;
      RECT  465300.0 810600.0 475500.0 796800.0 ;
      RECT  465300.0 810600.0 475500.0 824400.0 ;
      RECT  465300.0 838200.0 475500.0 824400.0 ;
      RECT  465300.0 838200.0 475500.0 852000.0 ;
      RECT  465300.0 865800.0 475500.0 852000.0 ;
      RECT  465300.0 865800.0 475500.0 879600.0 ;
      RECT  465300.0 893400.0 475500.0 879600.0 ;
      RECT  465300.0 893400.0 475500.0 907200.0 ;
      RECT  465300.0 921000.0 475500.0 907200.0 ;
      RECT  465300.0 921000.0 475500.0 934800.0 ;
      RECT  465300.0 948600.0 475500.0 934800.0 ;
      RECT  465300.0 948600.0 475500.0 962400.0 ;
      RECT  465300.0 976200.0 475500.0 962400.0 ;
      RECT  465300.0 976200.0 475500.0 990000.0 ;
      RECT  465300.0 1003800.0 475500.0 990000.0 ;
      RECT  465300.0 1003800.0 475500.0 1017600.0 ;
      RECT  465300.0 1031400.0 475500.0 1017600.0 ;
      RECT  465300.0 1031400.0 475500.0 1045200.0 ;
      RECT  465300.0 1059000.0 475500.0 1045200.0 ;
      RECT  465300.0 1059000.0 475500.0 1072800.0 ;
      RECT  465300.0 1086600.0 475500.0 1072800.0 ;
      RECT  465300.0 1086600.0 475500.0 1100400.0 ;
      RECT  465300.0 1114200.0 475500.0 1100400.0 ;
      RECT  465300.0 1114200.0 475500.0 1128000.0 ;
      RECT  465300.0 1141800.0 475500.0 1128000.0 ;
      RECT  465300.0 1141800.0 475500.0 1155600.0 ;
      RECT  465300.0 1169400.0 475500.0 1155600.0 ;
      RECT  465300.0 1169400.0 475500.0 1183200.0 ;
      RECT  465300.0 1197000.0 475500.0 1183200.0 ;
      RECT  475500.0 313800.0 485700.0 327600.0 ;
      RECT  475500.0 341400.0 485700.0 327600.0 ;
      RECT  475500.0 341400.0 485700.0 355200.0 ;
      RECT  475500.0 369000.0 485700.0 355200.0 ;
      RECT  475500.0 369000.0 485700.0 382800.0 ;
      RECT  475500.0 396600.0 485700.0 382800.0 ;
      RECT  475500.0 396600.0 485700.0 410400.0 ;
      RECT  475500.0 424200.0 485700.0 410400.0 ;
      RECT  475500.0 424200.0 485700.0 438000.0 ;
      RECT  475500.0 451800.0 485700.0 438000.0 ;
      RECT  475500.0 451800.0 485700.0 465600.0 ;
      RECT  475500.0 479400.0 485700.0 465600.0 ;
      RECT  475500.0 479400.0 485700.0 493200.0 ;
      RECT  475500.0 507000.0 485700.0 493200.0 ;
      RECT  475500.0 507000.0 485700.0 520800.0 ;
      RECT  475500.0 534600.0 485700.0 520800.0 ;
      RECT  475500.0 534600.0 485700.0 548400.0 ;
      RECT  475500.0 562200.0 485700.0 548400.0 ;
      RECT  475500.0 562200.0 485700.0 576000.0 ;
      RECT  475500.0 589800.0 485700.0 576000.0 ;
      RECT  475500.0 589800.0 485700.0 603600.0 ;
      RECT  475500.0 617400.0 485700.0 603600.0 ;
      RECT  475500.0 617400.0 485700.0 631200.0 ;
      RECT  475500.0 645000.0 485700.0 631200.0 ;
      RECT  475500.0 645000.0 485700.0 658800.0 ;
      RECT  475500.0 672600.0 485700.0 658800.0 ;
      RECT  475500.0 672600.0 485700.0 686400.0 ;
      RECT  475500.0 700200.0 485700.0 686400.0 ;
      RECT  475500.0 700200.0 485700.0 714000.0 ;
      RECT  475500.0 727800.0 485700.0 714000.0 ;
      RECT  475500.0 727800.0 485700.0 741600.0 ;
      RECT  475500.0 755400.0 485700.0 741600.0 ;
      RECT  475500.0 755400.0 485700.0 769200.0 ;
      RECT  475500.0 783000.0 485700.0 769200.0 ;
      RECT  475500.0 783000.0 485700.0 796800.0 ;
      RECT  475500.0 810600.0 485700.0 796800.0 ;
      RECT  475500.0 810600.0 485700.0 824400.0 ;
      RECT  475500.0 838200.0 485700.0 824400.0 ;
      RECT  475500.0 838200.0 485700.0 852000.0 ;
      RECT  475500.0 865800.0 485700.0 852000.0 ;
      RECT  475500.0 865800.0 485700.0 879600.0 ;
      RECT  475500.0 893400.0 485700.0 879600.0 ;
      RECT  475500.0 893400.0 485700.0 907200.0 ;
      RECT  475500.0 921000.0 485700.0 907200.0 ;
      RECT  475500.0 921000.0 485700.0 934800.0 ;
      RECT  475500.0 948600.0 485700.0 934800.0 ;
      RECT  475500.0 948600.0 485700.0 962400.0 ;
      RECT  475500.0 976200.0 485700.0 962400.0 ;
      RECT  475500.0 976200.0 485700.0 990000.0 ;
      RECT  475500.0 1003800.0 485700.0 990000.0 ;
      RECT  475500.0 1003800.0 485700.0 1017600.0 ;
      RECT  475500.0 1031400.0 485700.0 1017600.0 ;
      RECT  475500.0 1031400.0 485700.0 1045200.0 ;
      RECT  475500.0 1059000.0 485700.0 1045200.0 ;
      RECT  475500.0 1059000.0 485700.0 1072800.0 ;
      RECT  475500.0 1086600.0 485700.0 1072800.0 ;
      RECT  475500.0 1086600.0 485700.0 1100400.0 ;
      RECT  475500.0 1114200.0 485700.0 1100400.0 ;
      RECT  475500.0 1114200.0 485700.0 1128000.0 ;
      RECT  475500.0 1141800.0 485700.0 1128000.0 ;
      RECT  475500.0 1141800.0 485700.0 1155600.0 ;
      RECT  475500.0 1169400.0 485700.0 1155600.0 ;
      RECT  475500.0 1169400.0 485700.0 1183200.0 ;
      RECT  475500.0 1197000.0 485700.0 1183200.0 ;
      RECT  485700.0 313800.0 495900.0 327600.0 ;
      RECT  485700.0 341400.0 495900.0 327600.0 ;
      RECT  485700.0 341400.0 495900.0 355200.0 ;
      RECT  485700.0 369000.0 495900.0 355200.0 ;
      RECT  485700.0 369000.0 495900.0 382800.0 ;
      RECT  485700.0 396600.0 495900.0 382800.0 ;
      RECT  485700.0 396600.0 495900.0 410400.0 ;
      RECT  485700.0 424200.0 495900.0 410400.0 ;
      RECT  485700.0 424200.0 495900.0 438000.0 ;
      RECT  485700.0 451800.0 495900.0 438000.0 ;
      RECT  485700.0 451800.0 495900.0 465600.0 ;
      RECT  485700.0 479400.0 495900.0 465600.0 ;
      RECT  485700.0 479400.0 495900.0 493200.0 ;
      RECT  485700.0 507000.0 495900.0 493200.0 ;
      RECT  485700.0 507000.0 495900.0 520800.0 ;
      RECT  485700.0 534600.0 495900.0 520800.0 ;
      RECT  485700.0 534600.0 495900.0 548400.0 ;
      RECT  485700.0 562200.0 495900.0 548400.0 ;
      RECT  485700.0 562200.0 495900.0 576000.0 ;
      RECT  485700.0 589800.0 495900.0 576000.0 ;
      RECT  485700.0 589800.0 495900.0 603600.0 ;
      RECT  485700.0 617400.0 495900.0 603600.0 ;
      RECT  485700.0 617400.0 495900.0 631200.0 ;
      RECT  485700.0 645000.0 495900.0 631200.0 ;
      RECT  485700.0 645000.0 495900.0 658800.0 ;
      RECT  485700.0 672600.0 495900.0 658800.0 ;
      RECT  485700.0 672600.0 495900.0 686400.0 ;
      RECT  485700.0 700200.0 495900.0 686400.0 ;
      RECT  485700.0 700200.0 495900.0 714000.0 ;
      RECT  485700.0 727800.0 495900.0 714000.0 ;
      RECT  485700.0 727800.0 495900.0 741600.0 ;
      RECT  485700.0 755400.0 495900.0 741600.0 ;
      RECT  485700.0 755400.0 495900.0 769200.0 ;
      RECT  485700.0 783000.0 495900.0 769200.0 ;
      RECT  485700.0 783000.0 495900.0 796800.0 ;
      RECT  485700.0 810600.0 495900.0 796800.0 ;
      RECT  485700.0 810600.0 495900.0 824400.0 ;
      RECT  485700.0 838200.0 495900.0 824400.0 ;
      RECT  485700.0 838200.0 495900.0 852000.0 ;
      RECT  485700.0 865800.0 495900.0 852000.0 ;
      RECT  485700.0 865800.0 495900.0 879600.0 ;
      RECT  485700.0 893400.0 495900.0 879600.0 ;
      RECT  485700.0 893400.0 495900.0 907200.0 ;
      RECT  485700.0 921000.0 495900.0 907200.0 ;
      RECT  485700.0 921000.0 495900.0 934800.0 ;
      RECT  485700.0 948600.0 495900.0 934800.0 ;
      RECT  485700.0 948600.0 495900.0 962400.0 ;
      RECT  485700.0 976200.0 495900.0 962400.0 ;
      RECT  485700.0 976200.0 495900.0 990000.0 ;
      RECT  485700.0 1003800.0 495900.0 990000.0 ;
      RECT  485700.0 1003800.0 495900.0 1017600.0 ;
      RECT  485700.0 1031400.0 495900.0 1017600.0 ;
      RECT  485700.0 1031400.0 495900.0 1045200.0 ;
      RECT  485700.0 1059000.0 495900.0 1045200.0 ;
      RECT  485700.0 1059000.0 495900.0 1072800.0 ;
      RECT  485700.0 1086600.0 495900.0 1072800.0 ;
      RECT  485700.0 1086600.0 495900.0 1100400.0 ;
      RECT  485700.0 1114200.0 495900.0 1100400.0 ;
      RECT  485700.0 1114200.0 495900.0 1128000.0 ;
      RECT  485700.0 1141800.0 495900.0 1128000.0 ;
      RECT  485700.0 1141800.0 495900.0 1155600.0 ;
      RECT  485700.0 1169400.0 495900.0 1155600.0 ;
      RECT  485700.0 1169400.0 495900.0 1183200.0 ;
      RECT  485700.0 1197000.0 495900.0 1183200.0 ;
      RECT  495900.0 313800.0 506100.0 327600.0 ;
      RECT  495900.0 341400.0 506100.0 327600.0 ;
      RECT  495900.0 341400.0 506100.0 355200.0 ;
      RECT  495900.0 369000.0 506100.0 355200.0 ;
      RECT  495900.0 369000.0 506100.0 382800.0 ;
      RECT  495900.0 396600.0 506100.0 382800.0 ;
      RECT  495900.0 396600.0 506100.0 410400.0 ;
      RECT  495900.0 424200.0 506100.0 410400.0 ;
      RECT  495900.0 424200.0 506100.0 438000.0 ;
      RECT  495900.0 451800.0 506100.0 438000.0 ;
      RECT  495900.0 451800.0 506100.0 465600.0 ;
      RECT  495900.0 479400.0 506100.0 465600.0 ;
      RECT  495900.0 479400.0 506100.0 493200.0 ;
      RECT  495900.0 507000.0 506100.0 493200.0 ;
      RECT  495900.0 507000.0 506100.0 520800.0 ;
      RECT  495900.0 534600.0 506100.0 520800.0 ;
      RECT  495900.0 534600.0 506100.0 548400.0 ;
      RECT  495900.0 562200.0 506100.0 548400.0 ;
      RECT  495900.0 562200.0 506100.0 576000.0 ;
      RECT  495900.0 589800.0 506100.0 576000.0 ;
      RECT  495900.0 589800.0 506100.0 603600.0 ;
      RECT  495900.0 617400.0 506100.0 603600.0 ;
      RECT  495900.0 617400.0 506100.0 631200.0 ;
      RECT  495900.0 645000.0 506100.0 631200.0 ;
      RECT  495900.0 645000.0 506100.0 658800.0 ;
      RECT  495900.0 672600.0 506100.0 658800.0 ;
      RECT  495900.0 672600.0 506100.0 686400.0 ;
      RECT  495900.0 700200.0 506100.0 686400.0 ;
      RECT  495900.0 700200.0 506100.0 714000.0 ;
      RECT  495900.0 727800.0 506100.0 714000.0 ;
      RECT  495900.0 727800.0 506100.0 741600.0 ;
      RECT  495900.0 755400.0 506100.0 741600.0 ;
      RECT  495900.0 755400.0 506100.0 769200.0 ;
      RECT  495900.0 783000.0 506100.0 769200.0 ;
      RECT  495900.0 783000.0 506100.0 796800.0 ;
      RECT  495900.0 810600.0 506100.0 796800.0 ;
      RECT  495900.0 810600.0 506100.0 824400.0 ;
      RECT  495900.0 838200.0 506100.0 824400.0 ;
      RECT  495900.0 838200.0 506100.0 852000.0 ;
      RECT  495900.0 865800.0 506100.0 852000.0 ;
      RECT  495900.0 865800.0 506100.0 879600.0 ;
      RECT  495900.0 893400.0 506100.0 879600.0 ;
      RECT  495900.0 893400.0 506100.0 907200.0 ;
      RECT  495900.0 921000.0 506100.0 907200.0 ;
      RECT  495900.0 921000.0 506100.0 934800.0 ;
      RECT  495900.0 948600.0 506100.0 934800.0 ;
      RECT  495900.0 948600.0 506100.0 962400.0 ;
      RECT  495900.0 976200.0 506100.0 962400.0 ;
      RECT  495900.0 976200.0 506100.0 990000.0 ;
      RECT  495900.0 1003800.0 506100.0 990000.0 ;
      RECT  495900.0 1003800.0 506100.0 1017600.0 ;
      RECT  495900.0 1031400.0 506100.0 1017600.0 ;
      RECT  495900.0 1031400.0 506100.0 1045200.0 ;
      RECT  495900.0 1059000.0 506100.0 1045200.0 ;
      RECT  495900.0 1059000.0 506100.0 1072800.0 ;
      RECT  495900.0 1086600.0 506100.0 1072800.0 ;
      RECT  495900.0 1086600.0 506100.0 1100400.0 ;
      RECT  495900.0 1114200.0 506100.0 1100400.0 ;
      RECT  495900.0 1114200.0 506100.0 1128000.0 ;
      RECT  495900.0 1141800.0 506100.0 1128000.0 ;
      RECT  495900.0 1141800.0 506100.0 1155600.0 ;
      RECT  495900.0 1169400.0 506100.0 1155600.0 ;
      RECT  495900.0 1169400.0 506100.0 1183200.0 ;
      RECT  495900.0 1197000.0 506100.0 1183200.0 ;
      RECT  506100.0 313800.0 516300.0 327600.0 ;
      RECT  506100.0 341400.0 516300.0 327600.0 ;
      RECT  506100.0 341400.0 516300.0 355200.0 ;
      RECT  506100.0 369000.0 516300.0 355200.0 ;
      RECT  506100.0 369000.0 516300.0 382800.0 ;
      RECT  506100.0 396600.0 516300.0 382800.0 ;
      RECT  506100.0 396600.0 516300.0 410400.0 ;
      RECT  506100.0 424200.0 516300.0 410400.0 ;
      RECT  506100.0 424200.0 516300.0 438000.0 ;
      RECT  506100.0 451800.0 516300.0 438000.0 ;
      RECT  506100.0 451800.0 516300.0 465600.0 ;
      RECT  506100.0 479400.0 516300.0 465600.0 ;
      RECT  506100.0 479400.0 516300.0 493200.0 ;
      RECT  506100.0 507000.0 516300.0 493200.0 ;
      RECT  506100.0 507000.0 516300.0 520800.0 ;
      RECT  506100.0 534600.0 516300.0 520800.0 ;
      RECT  506100.0 534600.0 516300.0 548400.0 ;
      RECT  506100.0 562200.0 516300.0 548400.0 ;
      RECT  506100.0 562200.0 516300.0 576000.0 ;
      RECT  506100.0 589800.0 516300.0 576000.0 ;
      RECT  506100.0 589800.0 516300.0 603600.0 ;
      RECT  506100.0 617400.0 516300.0 603600.0 ;
      RECT  506100.0 617400.0 516300.0 631200.0 ;
      RECT  506100.0 645000.0 516300.0 631200.0 ;
      RECT  506100.0 645000.0 516300.0 658800.0 ;
      RECT  506100.0 672600.0 516300.0 658800.0 ;
      RECT  506100.0 672600.0 516300.0 686400.0 ;
      RECT  506100.0 700200.0 516300.0 686400.0 ;
      RECT  506100.0 700200.0 516300.0 714000.0 ;
      RECT  506100.0 727800.0 516300.0 714000.0 ;
      RECT  506100.0 727800.0 516300.0 741600.0 ;
      RECT  506100.0 755400.0 516300.0 741600.0 ;
      RECT  506100.0 755400.0 516300.0 769200.0 ;
      RECT  506100.0 783000.0 516300.0 769200.0 ;
      RECT  506100.0 783000.0 516300.0 796800.0 ;
      RECT  506100.0 810600.0 516300.0 796800.0 ;
      RECT  506100.0 810600.0 516300.0 824400.0 ;
      RECT  506100.0 838200.0 516300.0 824400.0 ;
      RECT  506100.0 838200.0 516300.0 852000.0 ;
      RECT  506100.0 865800.0 516300.0 852000.0 ;
      RECT  506100.0 865800.0 516300.0 879600.0 ;
      RECT  506100.0 893400.0 516300.0 879600.0 ;
      RECT  506100.0 893400.0 516300.0 907200.0 ;
      RECT  506100.0 921000.0 516300.0 907200.0 ;
      RECT  506100.0 921000.0 516300.0 934800.0 ;
      RECT  506100.0 948600.0 516300.0 934800.0 ;
      RECT  506100.0 948600.0 516300.0 962400.0 ;
      RECT  506100.0 976200.0 516300.0 962400.0 ;
      RECT  506100.0 976200.0 516300.0 990000.0 ;
      RECT  506100.0 1003800.0 516300.0 990000.0 ;
      RECT  506100.0 1003800.0 516300.0 1017600.0 ;
      RECT  506100.0 1031400.0 516300.0 1017600.0 ;
      RECT  506100.0 1031400.0 516300.0 1045200.0 ;
      RECT  506100.0 1059000.0 516300.0 1045200.0 ;
      RECT  506100.0 1059000.0 516300.0 1072800.0 ;
      RECT  506100.0 1086600.0 516300.0 1072800.0 ;
      RECT  506100.0 1086600.0 516300.0 1100400.0 ;
      RECT  506100.0 1114200.0 516300.0 1100400.0 ;
      RECT  506100.0 1114200.0 516300.0 1128000.0 ;
      RECT  506100.0 1141800.0 516300.0 1128000.0 ;
      RECT  506100.0 1141800.0 516300.0 1155600.0 ;
      RECT  506100.0 1169400.0 516300.0 1155600.0 ;
      RECT  506100.0 1169400.0 516300.0 1183200.0 ;
      RECT  506100.0 1197000.0 516300.0 1183200.0 ;
      RECT  516300.0 313800.0 526500.0 327600.0 ;
      RECT  516300.0 341400.0 526500.0 327600.0 ;
      RECT  516300.0 341400.0 526500.0 355200.0 ;
      RECT  516300.0 369000.0 526500.0 355200.0 ;
      RECT  516300.0 369000.0 526500.0 382800.0 ;
      RECT  516300.0 396600.0 526500.0 382800.0 ;
      RECT  516300.0 396600.0 526500.0 410400.0 ;
      RECT  516300.0 424200.0 526500.0 410400.0 ;
      RECT  516300.0 424200.0 526500.0 438000.0 ;
      RECT  516300.0 451800.0 526500.0 438000.0 ;
      RECT  516300.0 451800.0 526500.0 465600.0 ;
      RECT  516300.0 479400.0 526500.0 465600.0 ;
      RECT  516300.0 479400.0 526500.0 493200.0 ;
      RECT  516300.0 507000.0 526500.0 493200.0 ;
      RECT  516300.0 507000.0 526500.0 520800.0 ;
      RECT  516300.0 534600.0 526500.0 520800.0 ;
      RECT  516300.0 534600.0 526500.0 548400.0 ;
      RECT  516300.0 562200.0 526500.0 548400.0 ;
      RECT  516300.0 562200.0 526500.0 576000.0 ;
      RECT  516300.0 589800.0 526500.0 576000.0 ;
      RECT  516300.0 589800.0 526500.0 603600.0 ;
      RECT  516300.0 617400.0 526500.0 603600.0 ;
      RECT  516300.0 617400.0 526500.0 631200.0 ;
      RECT  516300.0 645000.0 526500.0 631200.0 ;
      RECT  516300.0 645000.0 526500.0 658800.0 ;
      RECT  516300.0 672600.0 526500.0 658800.0 ;
      RECT  516300.0 672600.0 526500.0 686400.0 ;
      RECT  516300.0 700200.0 526500.0 686400.0 ;
      RECT  516300.0 700200.0 526500.0 714000.0 ;
      RECT  516300.0 727800.0 526500.0 714000.0 ;
      RECT  516300.0 727800.0 526500.0 741600.0 ;
      RECT  516300.0 755400.0 526500.0 741600.0 ;
      RECT  516300.0 755400.0 526500.0 769200.0 ;
      RECT  516300.0 783000.0 526500.0 769200.0 ;
      RECT  516300.0 783000.0 526500.0 796800.0 ;
      RECT  516300.0 810600.0 526500.0 796800.0 ;
      RECT  516300.0 810600.0 526500.0 824400.0 ;
      RECT  516300.0 838200.0 526500.0 824400.0 ;
      RECT  516300.0 838200.0 526500.0 852000.0 ;
      RECT  516300.0 865800.0 526500.0 852000.0 ;
      RECT  516300.0 865800.0 526500.0 879600.0 ;
      RECT  516300.0 893400.0 526500.0 879600.0 ;
      RECT  516300.0 893400.0 526500.0 907200.0 ;
      RECT  516300.0 921000.0 526500.0 907200.0 ;
      RECT  516300.0 921000.0 526500.0 934800.0 ;
      RECT  516300.0 948600.0 526500.0 934800.0 ;
      RECT  516300.0 948600.0 526500.0 962400.0 ;
      RECT  516300.0 976200.0 526500.0 962400.0 ;
      RECT  516300.0 976200.0 526500.0 990000.0 ;
      RECT  516300.0 1003800.0 526500.0 990000.0 ;
      RECT  516300.0 1003800.0 526500.0 1017600.0 ;
      RECT  516300.0 1031400.0 526500.0 1017600.0 ;
      RECT  516300.0 1031400.0 526500.0 1045200.0 ;
      RECT  516300.0 1059000.0 526500.0 1045200.0 ;
      RECT  516300.0 1059000.0 526500.0 1072800.0 ;
      RECT  516300.0 1086600.0 526500.0 1072800.0 ;
      RECT  516300.0 1086600.0 526500.0 1100400.0 ;
      RECT  516300.0 1114200.0 526500.0 1100400.0 ;
      RECT  516300.0 1114200.0 526500.0 1128000.0 ;
      RECT  516300.0 1141800.0 526500.0 1128000.0 ;
      RECT  516300.0 1141800.0 526500.0 1155600.0 ;
      RECT  516300.0 1169400.0 526500.0 1155600.0 ;
      RECT  516300.0 1169400.0 526500.0 1183200.0 ;
      RECT  516300.0 1197000.0 526500.0 1183200.0 ;
      RECT  203100.0 314400.0 204300.0 1200600.0 ;
      RECT  206100.0 313200.0 207300.0 1199400.0 ;
      RECT  213300.0 314400.0 214500.0 1200600.0 ;
      RECT  216300.0 313200.0 217500.0 1199400.0 ;
      RECT  223500.0 314400.0 224700.0 1200600.0 ;
      RECT  226500.0 313200.0 227700.0 1199400.0 ;
      RECT  233700.0 314400.0 234900.0 1200600.0 ;
      RECT  236700.0 313200.0 237900.0 1199400.0 ;
      RECT  243900.0 314400.0 245100.0 1200600.0 ;
      RECT  246900.0 313200.0 248100.0 1199400.0 ;
      RECT  254100.0 314400.0 255300.0 1200600.0 ;
      RECT  257100.0 313200.0 258300.0 1199400.0 ;
      RECT  264300.0 314400.0 265500.0 1200600.0 ;
      RECT  267300.0 313200.0 268500.0 1199400.0 ;
      RECT  274500.0 314400.0 275700.0 1200600.0 ;
      RECT  277500.0 313200.0 278700.0 1199400.0 ;
      RECT  284700.0 314400.0 285900.0 1200600.0 ;
      RECT  287700.0 313200.0 288900.0 1199400.0 ;
      RECT  294900.0 314400.0 296100.0 1200600.0 ;
      RECT  297900.0 313200.0 299100.0 1199400.0 ;
      RECT  305100.0 314400.0 306300.0 1200600.0 ;
      RECT  308100.0 313200.0 309300.0 1199400.0 ;
      RECT  315300.0 314400.0 316500.0 1200600.0 ;
      RECT  318300.0 313200.0 319500.0 1199400.0 ;
      RECT  325500.0 314400.0 326700.0 1200600.0 ;
      RECT  328500.0 313200.0 329700.0 1199400.0 ;
      RECT  335700.0 314400.0 336900.0 1200600.0 ;
      RECT  338700.0 313200.0 339900.0 1199400.0 ;
      RECT  345900.0 314400.0 347100.0 1200600.0 ;
      RECT  348900.0 313200.0 350100.0 1199400.0 ;
      RECT  356100.0 314400.0 357300.0 1200600.0 ;
      RECT  359100.0 313200.0 360300.0 1199400.0 ;
      RECT  366300.0 314400.0 367500.0 1200600.0 ;
      RECT  369300.0 313200.0 370500.0 1199400.0 ;
      RECT  376500.0 314400.0 377700.0 1200600.0 ;
      RECT  379500.0 313200.0 380700.0 1199400.0 ;
      RECT  386700.0 314400.0 387900.0 1200600.0 ;
      RECT  389700.0 313200.0 390900.0 1199400.0 ;
      RECT  396900.0 314400.0 398100.0 1200600.0 ;
      RECT  399900.0 313200.0 401100.0 1199400.0 ;
      RECT  407100.0 314400.0 408300.0 1200600.0 ;
      RECT  410100.0 313200.0 411300.0 1199400.0 ;
      RECT  417300.0 314400.0 418500.0 1200600.0 ;
      RECT  420300.0 313200.0 421500.0 1199400.0 ;
      RECT  427500.0 314400.0 428700.0 1200600.0 ;
      RECT  430500.0 313200.0 431700.0 1199400.0 ;
      RECT  437700.0 314400.0 438900.0 1200600.0 ;
      RECT  440700.0 313200.0 441900.0 1199400.0 ;
      RECT  447900.0 314400.0 449100.0 1200600.0 ;
      RECT  450900.0 313200.0 452100.0 1199400.0 ;
      RECT  458100.0 314400.0 459300.0 1200600.0 ;
      RECT  461100.0 313200.0 462300.0 1199400.0 ;
      RECT  468300.0 314400.0 469500.0 1200600.0 ;
      RECT  471300.0 313200.0 472500.0 1199400.0 ;
      RECT  478500.0 314400.0 479700.0 1200600.0 ;
      RECT  481500.0 313200.0 482700.0 1199400.0 ;
      RECT  488700.0 314400.0 489900.0 1200600.0 ;
      RECT  491700.0 313200.0 492900.0 1199400.0 ;
      RECT  498900.0 314400.0 500100.0 1200600.0 ;
      RECT  501900.0 313200.0 503100.0 1199400.0 ;
      RECT  509100.0 314400.0 510300.0 1200600.0 ;
      RECT  512100.0 313200.0 513300.0 1199400.0 ;
      RECT  519300.0 314400.0 520500.0 1200600.0 ;
      RECT  522300.0 313200.0 523500.0 1199400.0 ;
      RECT  199500.0 313200.0 200700.0 1199400.0 ;
      RECT  209700.0 313200.0 210900.0 1199400.0 ;
      RECT  219900.0 313200.0 221100.0 1199400.0 ;
      RECT  230100.0 313200.0 231300.0 1199400.0 ;
      RECT  240300.0 313200.0 241500.0 1199400.0 ;
      RECT  250500.0 313200.0 251700.0 1199400.0 ;
      RECT  260700.0 313200.0 261900.0 1199400.0 ;
      RECT  270900.0 313200.0 272100.0 1199400.0 ;
      RECT  281100.0 313200.0 282300.0 1199400.0 ;
      RECT  291300.0 313200.0 292500.0 1199400.0 ;
      RECT  301500.0 313200.0 302700.0 1199400.0 ;
      RECT  311700.0 313200.0 312900.0 1199400.0 ;
      RECT  321900.0 313200.0 323100.0 1199400.0 ;
      RECT  332100.0 313200.0 333300.0 1199400.0 ;
      RECT  342300.0 313200.0 343500.0 1199400.0 ;
      RECT  352500.0 313200.0 353700.0 1199400.0 ;
      RECT  362700.0 313200.0 363900.0 1199400.0 ;
      RECT  372900.0 313200.0 374100.0 1199400.0 ;
      RECT  383100.0 313200.0 384300.0 1199400.0 ;
      RECT  393300.0 313200.0 394500.0 1199400.0 ;
      RECT  403500.0 313200.0 404700.0 1199400.0 ;
      RECT  413700.0 313200.0 414900.0 1199400.0 ;
      RECT  423900.0 313200.0 425100.0 1199400.0 ;
      RECT  434100.0 313200.0 435300.0 1199400.0 ;
      RECT  444300.0 313200.0 445500.0 1199400.0 ;
      RECT  454500.0 313200.0 455700.0 1199400.0 ;
      RECT  464700.0 313200.0 465900.0 1199400.0 ;
      RECT  474900.0 313200.0 476100.0 1199400.0 ;
      RECT  485100.0 313200.0 486300.0 1199400.0 ;
      RECT  495300.0 313200.0 496500.0 1199400.0 ;
      RECT  505500.0 313200.0 506700.0 1199400.0 ;
      RECT  515700.0 313200.0 516900.0 1199400.0 ;
      RECT  525900.0 313200.0 527100.0 1199400.0 ;
      RECT  203100.0 1203000.0 204300.0 1204200.0 ;
      RECT  205500.0 1203000.0 207150.0 1204200.0 ;
      RECT  203100.0 1210200.0 204300.0 1211400.0 ;
      RECT  206250.0 1210200.0 209100.0 1211400.0 ;
      RECT  203100.0 1203000.0 204300.0 1204200.0 ;
      RECT  205500.0 1203000.0 206700.0 1204200.0 ;
      RECT  203100.0 1210200.0 204300.0 1211400.0 ;
      RECT  207900.0 1210200.0 209100.0 1211400.0 ;
      RECT  203250.0 1200600.0 204150.0 1217400.0 ;
      RECT  206250.0 1200600.0 207150.0 1217400.0 ;
      RECT  213300.0 1203000.0 214500.0 1204200.0 ;
      RECT  215700.0 1203000.0 217350.0 1204200.0 ;
      RECT  213300.0 1210200.0 214500.0 1211400.0 ;
      RECT  216450.0 1210200.0 219300.0 1211400.0 ;
      RECT  213300.0 1203000.0 214500.0 1204200.0 ;
      RECT  215700.0 1203000.0 216900.0 1204200.0 ;
      RECT  213300.0 1210200.0 214500.0 1211400.0 ;
      RECT  218100.0 1210200.0 219300.0 1211400.0 ;
      RECT  213450.0 1200600.0 214350.0 1217400.0 ;
      RECT  216450.0 1200600.0 217350.0 1217400.0 ;
      RECT  223500.0 1203000.0 224700.0 1204200.0 ;
      RECT  225900.0 1203000.0 227550.0 1204200.0 ;
      RECT  223500.0 1210200.0 224700.0 1211400.0 ;
      RECT  226650.0 1210200.0 229500.0 1211400.0 ;
      RECT  223500.0 1203000.0 224700.0 1204200.0 ;
      RECT  225900.0 1203000.0 227100.0 1204200.0 ;
      RECT  223500.0 1210200.0 224700.0 1211400.0 ;
      RECT  228300.0 1210200.0 229500.0 1211400.0 ;
      RECT  223650.0 1200600.0 224550.0 1217400.0 ;
      RECT  226650.0 1200600.0 227550.0 1217400.0 ;
      RECT  233700.0 1203000.0 234900.0 1204200.0 ;
      RECT  236100.0 1203000.0 237750.0 1204200.0 ;
      RECT  233700.0 1210200.0 234900.0 1211400.0 ;
      RECT  236850.0 1210200.0 239700.0 1211400.0 ;
      RECT  233700.0 1203000.0 234900.0 1204200.0 ;
      RECT  236100.0 1203000.0 237300.0 1204200.0 ;
      RECT  233700.0 1210200.0 234900.0 1211400.0 ;
      RECT  238500.0 1210200.0 239700.0 1211400.0 ;
      RECT  233850.0 1200600.0 234750.0 1217400.0 ;
      RECT  236850.0 1200600.0 237750.0 1217400.0 ;
      RECT  243900.0 1203000.0 245100.0 1204200.0 ;
      RECT  246300.0 1203000.0 247950.0 1204200.0 ;
      RECT  243900.0 1210200.0 245100.0 1211400.0 ;
      RECT  247050.0 1210200.0 249900.0 1211400.0 ;
      RECT  243900.0 1203000.0 245100.0 1204200.0 ;
      RECT  246300.0 1203000.0 247500.0 1204200.0 ;
      RECT  243900.0 1210200.0 245100.0 1211400.0 ;
      RECT  248700.0 1210200.0 249900.0 1211400.0 ;
      RECT  244050.0 1200600.0 244950.0 1217400.0 ;
      RECT  247050.0 1200600.0 247950.0 1217400.0 ;
      RECT  254100.0 1203000.0 255300.0 1204200.0 ;
      RECT  256500.0 1203000.0 258150.0 1204200.0 ;
      RECT  254100.0 1210200.0 255300.0 1211400.0 ;
      RECT  257250.0 1210200.0 260100.0 1211400.0 ;
      RECT  254100.0 1203000.0 255300.0 1204200.0 ;
      RECT  256500.0 1203000.0 257700.0 1204200.0 ;
      RECT  254100.0 1210200.0 255300.0 1211400.0 ;
      RECT  258900.0 1210200.0 260100.0 1211400.0 ;
      RECT  254250.0 1200600.0 255150.0 1217400.0 ;
      RECT  257250.0 1200600.0 258150.0 1217400.0 ;
      RECT  264300.0 1203000.0 265500.0 1204200.0 ;
      RECT  266700.0 1203000.0 268350.0 1204200.0 ;
      RECT  264300.0 1210200.0 265500.0 1211400.0 ;
      RECT  267450.0 1210200.0 270300.0 1211400.0 ;
      RECT  264300.0 1203000.0 265500.0 1204200.0 ;
      RECT  266700.0 1203000.0 267900.0 1204200.0 ;
      RECT  264300.0 1210200.0 265500.0 1211400.0 ;
      RECT  269100.0 1210200.0 270300.0 1211400.0 ;
      RECT  264450.0 1200600.0 265350.0 1217400.0 ;
      RECT  267450.0 1200600.0 268350.0 1217400.0 ;
      RECT  274500.0 1203000.0 275700.0 1204200.0 ;
      RECT  276900.0 1203000.0 278550.0 1204200.0 ;
      RECT  274500.0 1210200.0 275700.0 1211400.0 ;
      RECT  277650.0 1210200.0 280500.0 1211400.0 ;
      RECT  274500.0 1203000.0 275700.0 1204200.0 ;
      RECT  276900.0 1203000.0 278100.0 1204200.0 ;
      RECT  274500.0 1210200.0 275700.0 1211400.0 ;
      RECT  279300.0 1210200.0 280500.0 1211400.0 ;
      RECT  274650.0 1200600.0 275550.0 1217400.0 ;
      RECT  277650.0 1200600.0 278550.0 1217400.0 ;
      RECT  284700.0 1203000.0 285900.0 1204200.0 ;
      RECT  287100.0 1203000.0 288750.0 1204200.0 ;
      RECT  284700.0 1210200.0 285900.0 1211400.0 ;
      RECT  287850.0 1210200.0 290700.0 1211400.0 ;
      RECT  284700.0 1203000.0 285900.0 1204200.0 ;
      RECT  287100.0 1203000.0 288300.0 1204200.0 ;
      RECT  284700.0 1210200.0 285900.0 1211400.0 ;
      RECT  289500.0 1210200.0 290700.0 1211400.0 ;
      RECT  284850.0 1200600.0 285750.0 1217400.0 ;
      RECT  287850.0 1200600.0 288750.0 1217400.0 ;
      RECT  294900.0 1203000.0 296100.0 1204200.0 ;
      RECT  297300.0 1203000.0 298950.0 1204200.0 ;
      RECT  294900.0 1210200.0 296100.0 1211400.0 ;
      RECT  298050.0 1210200.0 300900.0 1211400.0 ;
      RECT  294900.0 1203000.0 296100.0 1204200.0 ;
      RECT  297300.0 1203000.0 298500.0 1204200.0 ;
      RECT  294900.0 1210200.0 296100.0 1211400.0 ;
      RECT  299700.0 1210200.0 300900.0 1211400.0 ;
      RECT  295050.0 1200600.0 295950.0 1217400.0 ;
      RECT  298050.0 1200600.0 298950.0 1217400.0 ;
      RECT  305100.0 1203000.0 306300.0 1204200.0 ;
      RECT  307500.0 1203000.0 309150.0 1204200.0 ;
      RECT  305100.0 1210200.0 306300.0 1211400.0 ;
      RECT  308250.0 1210200.0 311100.0 1211400.0 ;
      RECT  305100.0 1203000.0 306300.0 1204200.0 ;
      RECT  307500.0 1203000.0 308700.0 1204200.0 ;
      RECT  305100.0 1210200.0 306300.0 1211400.0 ;
      RECT  309900.0 1210200.0 311100.0 1211400.0 ;
      RECT  305250.0 1200600.0 306150.0 1217400.0 ;
      RECT  308250.0 1200600.0 309150.0 1217400.0 ;
      RECT  315300.0 1203000.0 316500.0 1204200.0 ;
      RECT  317700.0 1203000.0 319350.0 1204200.0 ;
      RECT  315300.0 1210200.0 316500.0 1211400.0 ;
      RECT  318450.0 1210200.0 321300.0 1211400.0 ;
      RECT  315300.0 1203000.0 316500.0 1204200.0 ;
      RECT  317700.0 1203000.0 318900.0 1204200.0 ;
      RECT  315300.0 1210200.0 316500.0 1211400.0 ;
      RECT  320100.0 1210200.0 321300.0 1211400.0 ;
      RECT  315450.0 1200600.0 316350.0 1217400.0 ;
      RECT  318450.0 1200600.0 319350.0 1217400.0 ;
      RECT  325500.0 1203000.0 326700.0 1204200.0 ;
      RECT  327900.0 1203000.0 329550.0 1204200.0 ;
      RECT  325500.0 1210200.0 326700.0 1211400.0 ;
      RECT  328650.0 1210200.0 331500.0 1211400.0 ;
      RECT  325500.0 1203000.0 326700.0 1204200.0 ;
      RECT  327900.0 1203000.0 329100.0 1204200.0 ;
      RECT  325500.0 1210200.0 326700.0 1211400.0 ;
      RECT  330300.0 1210200.0 331500.0 1211400.0 ;
      RECT  325650.0 1200600.0 326550.0 1217400.0 ;
      RECT  328650.0 1200600.0 329550.0 1217400.0 ;
      RECT  335700.0 1203000.0 336900.0 1204200.0 ;
      RECT  338100.0 1203000.0 339750.0 1204200.0 ;
      RECT  335700.0 1210200.0 336900.0 1211400.0 ;
      RECT  338850.0 1210200.0 341700.0 1211400.0 ;
      RECT  335700.0 1203000.0 336900.0 1204200.0 ;
      RECT  338100.0 1203000.0 339300.0 1204200.0 ;
      RECT  335700.0 1210200.0 336900.0 1211400.0 ;
      RECT  340500.0 1210200.0 341700.0 1211400.0 ;
      RECT  335850.0 1200600.0 336750.0 1217400.0 ;
      RECT  338850.0 1200600.0 339750.0 1217400.0 ;
      RECT  345900.0 1203000.0 347100.0 1204200.0 ;
      RECT  348300.0 1203000.0 349950.0 1204200.0 ;
      RECT  345900.0 1210200.0 347100.0 1211400.0 ;
      RECT  349050.0 1210200.0 351900.0 1211400.0 ;
      RECT  345900.0 1203000.0 347100.0 1204200.0 ;
      RECT  348300.0 1203000.0 349500.0 1204200.0 ;
      RECT  345900.0 1210200.0 347100.0 1211400.0 ;
      RECT  350700.0 1210200.0 351900.0 1211400.0 ;
      RECT  346050.0 1200600.0 346950.0 1217400.0 ;
      RECT  349050.0 1200600.0 349950.0 1217400.0 ;
      RECT  356100.0 1203000.0 357300.0 1204200.0 ;
      RECT  358500.0 1203000.0 360150.0 1204200.0 ;
      RECT  356100.0 1210200.0 357300.0 1211400.0 ;
      RECT  359250.0 1210200.0 362100.0 1211400.0 ;
      RECT  356100.0 1203000.0 357300.0 1204200.0 ;
      RECT  358500.0 1203000.0 359700.0 1204200.0 ;
      RECT  356100.0 1210200.0 357300.0 1211400.0 ;
      RECT  360900.0 1210200.0 362100.0 1211400.0 ;
      RECT  356250.0 1200600.0 357150.0 1217400.0 ;
      RECT  359250.0 1200600.0 360150.0 1217400.0 ;
      RECT  366300.0 1203000.0 367500.0 1204200.0 ;
      RECT  368700.0 1203000.0 370350.0 1204200.0 ;
      RECT  366300.0 1210200.0 367500.0 1211400.0 ;
      RECT  369450.0 1210200.0 372300.0 1211400.0 ;
      RECT  366300.0 1203000.0 367500.0 1204200.0 ;
      RECT  368700.0 1203000.0 369900.0 1204200.0 ;
      RECT  366300.0 1210200.0 367500.0 1211400.0 ;
      RECT  371100.0 1210200.0 372300.0 1211400.0 ;
      RECT  366450.0 1200600.0 367350.0 1217400.0 ;
      RECT  369450.0 1200600.0 370350.0 1217400.0 ;
      RECT  376500.0 1203000.0 377700.0 1204200.0 ;
      RECT  378900.0 1203000.0 380550.0 1204200.0 ;
      RECT  376500.0 1210200.0 377700.0 1211400.0 ;
      RECT  379650.0 1210200.0 382500.0 1211400.0 ;
      RECT  376500.0 1203000.0 377700.0 1204200.0 ;
      RECT  378900.0 1203000.0 380100.0 1204200.0 ;
      RECT  376500.0 1210200.0 377700.0 1211400.0 ;
      RECT  381300.0 1210200.0 382500.0 1211400.0 ;
      RECT  376650.0 1200600.0 377550.0 1217400.0 ;
      RECT  379650.0 1200600.0 380550.0 1217400.0 ;
      RECT  386700.0 1203000.0 387900.0 1204200.0 ;
      RECT  389100.0 1203000.0 390750.0 1204200.0 ;
      RECT  386700.0 1210200.0 387900.0 1211400.0 ;
      RECT  389850.0 1210200.0 392700.0 1211400.0 ;
      RECT  386700.0 1203000.0 387900.0 1204200.0 ;
      RECT  389100.0 1203000.0 390300.0 1204200.0 ;
      RECT  386700.0 1210200.0 387900.0 1211400.0 ;
      RECT  391500.0 1210200.0 392700.0 1211400.0 ;
      RECT  386850.0 1200600.0 387750.0 1217400.0 ;
      RECT  389850.0 1200600.0 390750.0 1217400.0 ;
      RECT  396900.0 1203000.0 398100.0 1204200.0 ;
      RECT  399300.0 1203000.0 400950.0 1204200.0 ;
      RECT  396900.0 1210200.0 398100.0 1211400.0 ;
      RECT  400050.0 1210200.0 402900.0 1211400.0 ;
      RECT  396900.0 1203000.0 398100.0 1204200.0 ;
      RECT  399300.0 1203000.0 400500.0 1204200.0 ;
      RECT  396900.0 1210200.0 398100.0 1211400.0 ;
      RECT  401700.0 1210200.0 402900.0 1211400.0 ;
      RECT  397050.0 1200600.0 397950.0 1217400.0 ;
      RECT  400050.0 1200600.0 400950.0 1217400.0 ;
      RECT  407100.0 1203000.0 408300.0 1204200.0 ;
      RECT  409500.0 1203000.0 411150.0 1204200.0 ;
      RECT  407100.0 1210200.0 408300.0 1211400.0 ;
      RECT  410250.0 1210200.0 413100.0 1211400.0 ;
      RECT  407100.0 1203000.0 408300.0 1204200.0 ;
      RECT  409500.0 1203000.0 410700.0 1204200.0 ;
      RECT  407100.0 1210200.0 408300.0 1211400.0 ;
      RECT  411900.0 1210200.0 413100.0 1211400.0 ;
      RECT  407250.0 1200600.0 408150.0 1217400.0 ;
      RECT  410250.0 1200600.0 411150.0 1217400.0 ;
      RECT  417300.0 1203000.0 418500.0 1204200.0 ;
      RECT  419700.0 1203000.0 421350.0 1204200.0 ;
      RECT  417300.0 1210200.0 418500.0 1211400.0 ;
      RECT  420450.0 1210200.0 423300.0 1211400.0 ;
      RECT  417300.0 1203000.0 418500.0 1204200.0 ;
      RECT  419700.0 1203000.0 420900.0 1204200.0 ;
      RECT  417300.0 1210200.0 418500.0 1211400.0 ;
      RECT  422100.0 1210200.0 423300.0 1211400.0 ;
      RECT  417450.0 1200600.0 418350.0 1217400.0 ;
      RECT  420450.0 1200600.0 421350.0 1217400.0 ;
      RECT  427500.0 1203000.0 428700.0 1204200.0 ;
      RECT  429900.0 1203000.0 431550.0 1204200.0 ;
      RECT  427500.0 1210200.0 428700.0 1211400.0 ;
      RECT  430650.0 1210200.0 433500.0 1211400.0 ;
      RECT  427500.0 1203000.0 428700.0 1204200.0 ;
      RECT  429900.0 1203000.0 431100.0 1204200.0 ;
      RECT  427500.0 1210200.0 428700.0 1211400.0 ;
      RECT  432300.0 1210200.0 433500.0 1211400.0 ;
      RECT  427650.0 1200600.0 428550.0 1217400.0 ;
      RECT  430650.0 1200600.0 431550.0 1217400.0 ;
      RECT  437700.0 1203000.0 438900.0 1204200.0 ;
      RECT  440100.0 1203000.0 441750.0 1204200.0 ;
      RECT  437700.0 1210200.0 438900.0 1211400.0 ;
      RECT  440850.0 1210200.0 443700.0 1211400.0 ;
      RECT  437700.0 1203000.0 438900.0 1204200.0 ;
      RECT  440100.0 1203000.0 441300.0 1204200.0 ;
      RECT  437700.0 1210200.0 438900.0 1211400.0 ;
      RECT  442500.0 1210200.0 443700.0 1211400.0 ;
      RECT  437850.0 1200600.0 438750.0 1217400.0 ;
      RECT  440850.0 1200600.0 441750.0 1217400.0 ;
      RECT  447900.0 1203000.0 449100.0 1204200.0 ;
      RECT  450300.0 1203000.0 451950.0 1204200.0 ;
      RECT  447900.0 1210200.0 449100.0 1211400.0 ;
      RECT  451050.0 1210200.0 453900.0 1211400.0 ;
      RECT  447900.0 1203000.0 449100.0 1204200.0 ;
      RECT  450300.0 1203000.0 451500.0 1204200.0 ;
      RECT  447900.0 1210200.0 449100.0 1211400.0 ;
      RECT  452700.0 1210200.0 453900.0 1211400.0 ;
      RECT  448050.0 1200600.0 448950.0 1217400.0 ;
      RECT  451050.0 1200600.0 451950.0 1217400.0 ;
      RECT  458100.0 1203000.0 459300.0 1204200.0 ;
      RECT  460500.0 1203000.0 462150.0 1204200.0 ;
      RECT  458100.0 1210200.0 459300.0 1211400.0 ;
      RECT  461250.0 1210200.0 464100.0 1211400.0 ;
      RECT  458100.0 1203000.0 459300.0 1204200.0 ;
      RECT  460500.0 1203000.0 461700.0 1204200.0 ;
      RECT  458100.0 1210200.0 459300.0 1211400.0 ;
      RECT  462900.0 1210200.0 464100.0 1211400.0 ;
      RECT  458250.0 1200600.0 459150.0 1217400.0 ;
      RECT  461250.0 1200600.0 462150.0 1217400.0 ;
      RECT  468300.0 1203000.0 469500.0 1204200.0 ;
      RECT  470700.0 1203000.0 472350.0 1204200.0 ;
      RECT  468300.0 1210200.0 469500.0 1211400.0 ;
      RECT  471450.0 1210200.0 474300.0 1211400.0 ;
      RECT  468300.0 1203000.0 469500.0 1204200.0 ;
      RECT  470700.0 1203000.0 471900.0 1204200.0 ;
      RECT  468300.0 1210200.0 469500.0 1211400.0 ;
      RECT  473100.0 1210200.0 474300.0 1211400.0 ;
      RECT  468450.0 1200600.0 469350.0 1217400.0 ;
      RECT  471450.0 1200600.0 472350.0 1217400.0 ;
      RECT  478500.0 1203000.0 479700.0 1204200.0 ;
      RECT  480900.0 1203000.0 482550.0 1204200.0 ;
      RECT  478500.0 1210200.0 479700.0 1211400.0 ;
      RECT  481650.0 1210200.0 484500.0 1211400.0 ;
      RECT  478500.0 1203000.0 479700.0 1204200.0 ;
      RECT  480900.0 1203000.0 482100.0 1204200.0 ;
      RECT  478500.0 1210200.0 479700.0 1211400.0 ;
      RECT  483300.0 1210200.0 484500.0 1211400.0 ;
      RECT  478650.0 1200600.0 479550.0 1217400.0 ;
      RECT  481650.0 1200600.0 482550.0 1217400.0 ;
      RECT  488700.0 1203000.0 489900.0 1204200.0 ;
      RECT  491100.0 1203000.0 492750.0 1204200.0 ;
      RECT  488700.0 1210200.0 489900.0 1211400.0 ;
      RECT  491850.0 1210200.0 494700.0 1211400.0 ;
      RECT  488700.0 1203000.0 489900.0 1204200.0 ;
      RECT  491100.0 1203000.0 492300.0 1204200.0 ;
      RECT  488700.0 1210200.0 489900.0 1211400.0 ;
      RECT  493500.0 1210200.0 494700.0 1211400.0 ;
      RECT  488850.0 1200600.0 489750.0 1217400.0 ;
      RECT  491850.0 1200600.0 492750.0 1217400.0 ;
      RECT  498900.0 1203000.0 500100.0 1204200.0 ;
      RECT  501300.0 1203000.0 502950.0 1204200.0 ;
      RECT  498900.0 1210200.0 500100.0 1211400.0 ;
      RECT  502050.0 1210200.0 504900.0 1211400.0 ;
      RECT  498900.0 1203000.0 500100.0 1204200.0 ;
      RECT  501300.0 1203000.0 502500.0 1204200.0 ;
      RECT  498900.0 1210200.0 500100.0 1211400.0 ;
      RECT  503700.0 1210200.0 504900.0 1211400.0 ;
      RECT  499050.0 1200600.0 499950.0 1217400.0 ;
      RECT  502050.0 1200600.0 502950.0 1217400.0 ;
      RECT  509100.0 1203000.0 510300.0 1204200.0 ;
      RECT  511500.0 1203000.0 513150.0 1204200.0 ;
      RECT  509100.0 1210200.0 510300.0 1211400.0 ;
      RECT  512250.0 1210200.0 515100.0 1211400.0 ;
      RECT  509100.0 1203000.0 510300.0 1204200.0 ;
      RECT  511500.0 1203000.0 512700.0 1204200.0 ;
      RECT  509100.0 1210200.0 510300.0 1211400.0 ;
      RECT  513900.0 1210200.0 515100.0 1211400.0 ;
      RECT  509250.0 1200600.0 510150.0 1217400.0 ;
      RECT  512250.0 1200600.0 513150.0 1217400.0 ;
      RECT  519300.0 1203000.0 520500.0 1204200.0 ;
      RECT  521700.0 1203000.0 523350.0 1204200.0 ;
      RECT  519300.0 1210200.0 520500.0 1211400.0 ;
      RECT  522450.0 1210200.0 525300.0 1211400.0 ;
      RECT  519300.0 1203000.0 520500.0 1204200.0 ;
      RECT  521700.0 1203000.0 522900.0 1204200.0 ;
      RECT  519300.0 1210200.0 520500.0 1211400.0 ;
      RECT  524100.0 1210200.0 525300.0 1211400.0 ;
      RECT  519450.0 1200600.0 520350.0 1217400.0 ;
      RECT  522450.0 1200600.0 523350.0 1217400.0 ;
      RECT  203250.0 1200600.0 204150.0 1217400.0 ;
      RECT  206250.0 1200600.0 207150.0 1217400.0 ;
      RECT  213450.0 1200600.0 214350.0 1217400.0 ;
      RECT  216450.0 1200600.0 217350.0 1217400.0 ;
      RECT  223650.0 1200600.0 224550.0 1217400.0 ;
      RECT  226650.0 1200600.0 227550.0 1217400.0 ;
      RECT  233850.0 1200600.0 234750.0 1217400.0 ;
      RECT  236850.0 1200600.0 237750.0 1217400.0 ;
      RECT  244050.0 1200600.0 244950.0 1217400.0 ;
      RECT  247050.0 1200600.0 247950.0 1217400.0 ;
      RECT  254250.0 1200600.0 255150.0 1217400.0 ;
      RECT  257250.0 1200600.0 258150.0 1217400.0 ;
      RECT  264450.0 1200600.0 265350.0 1217400.0 ;
      RECT  267450.0 1200600.0 268350.0 1217400.0 ;
      RECT  274650.0 1200600.0 275550.0 1217400.0 ;
      RECT  277650.0 1200600.0 278550.0 1217400.0 ;
      RECT  284850.0 1200600.0 285750.0 1217400.0 ;
      RECT  287850.0 1200600.0 288750.0 1217400.0 ;
      RECT  295050.0 1200600.0 295950.0 1217400.0 ;
      RECT  298050.0 1200600.0 298950.0 1217400.0 ;
      RECT  305250.0 1200600.0 306150.0 1217400.0 ;
      RECT  308250.0 1200600.0 309150.0 1217400.0 ;
      RECT  315450.0 1200600.0 316350.0 1217400.0 ;
      RECT  318450.0 1200600.0 319350.0 1217400.0 ;
      RECT  325650.0 1200600.0 326550.0 1217400.0 ;
      RECT  328650.0 1200600.0 329550.0 1217400.0 ;
      RECT  335850.0 1200600.0 336750.0 1217400.0 ;
      RECT  338850.0 1200600.0 339750.0 1217400.0 ;
      RECT  346050.0 1200600.0 346950.0 1217400.0 ;
      RECT  349050.0 1200600.0 349950.0 1217400.0 ;
      RECT  356250.0 1200600.0 357150.0 1217400.0 ;
      RECT  359250.0 1200600.0 360150.0 1217400.0 ;
      RECT  366450.0 1200600.0 367350.0 1217400.0 ;
      RECT  369450.0 1200600.0 370350.0 1217400.0 ;
      RECT  376650.0 1200600.0 377550.0 1217400.0 ;
      RECT  379650.0 1200600.0 380550.0 1217400.0 ;
      RECT  386850.0 1200600.0 387750.0 1217400.0 ;
      RECT  389850.0 1200600.0 390750.0 1217400.0 ;
      RECT  397050.0 1200600.0 397950.0 1217400.0 ;
      RECT  400050.0 1200600.0 400950.0 1217400.0 ;
      RECT  407250.0 1200600.0 408150.0 1217400.0 ;
      RECT  410250.0 1200600.0 411150.0 1217400.0 ;
      RECT  417450.0 1200600.0 418350.0 1217400.0 ;
      RECT  420450.0 1200600.0 421350.0 1217400.0 ;
      RECT  427650.0 1200600.0 428550.0 1217400.0 ;
      RECT  430650.0 1200600.0 431550.0 1217400.0 ;
      RECT  437850.0 1200600.0 438750.0 1217400.0 ;
      RECT  440850.0 1200600.0 441750.0 1217400.0 ;
      RECT  448050.0 1200600.0 448950.0 1217400.0 ;
      RECT  451050.0 1200600.0 451950.0 1217400.0 ;
      RECT  458250.0 1200600.0 459150.0 1217400.0 ;
      RECT  461250.0 1200600.0 462150.0 1217400.0 ;
      RECT  468450.0 1200600.0 469350.0 1217400.0 ;
      RECT  471450.0 1200600.0 472350.0 1217400.0 ;
      RECT  478650.0 1200600.0 479550.0 1217400.0 ;
      RECT  481650.0 1200600.0 482550.0 1217400.0 ;
      RECT  488850.0 1200600.0 489750.0 1217400.0 ;
      RECT  491850.0 1200600.0 492750.0 1217400.0 ;
      RECT  499050.0 1200600.0 499950.0 1217400.0 ;
      RECT  502050.0 1200600.0 502950.0 1217400.0 ;
      RECT  509250.0 1200600.0 510150.0 1217400.0 ;
      RECT  512250.0 1200600.0 513150.0 1217400.0 ;
      RECT  519450.0 1200600.0 520350.0 1217400.0 ;
      RECT  522450.0 1200600.0 523350.0 1217400.0 ;
      RECT  213300.0 277350.0 214200.0 287850.0 ;
      RECT  216300.0 275250.0 217200.0 287850.0 ;
      RECT  223500.0 277350.0 224400.0 287850.0 ;
      RECT  226500.0 275250.0 227400.0 287850.0 ;
      RECT  233700.0 277350.0 234600.0 287850.0 ;
      RECT  236700.0 275250.0 237600.0 287850.0 ;
      RECT  254100.0 277350.0 255000.0 287850.0 ;
      RECT  257100.0 275250.0 258000.0 287850.0 ;
      RECT  264300.0 277350.0 265200.0 287850.0 ;
      RECT  267300.0 275250.0 268200.0 287850.0 ;
      RECT  274500.0 277350.0 275400.0 287850.0 ;
      RECT  277500.0 275250.0 278400.0 287850.0 ;
      RECT  294900.0 277350.0 295800.0 287850.0 ;
      RECT  297900.0 275250.0 298800.0 287850.0 ;
      RECT  305100.0 277350.0 306000.0 287850.0 ;
      RECT  308100.0 275250.0 309000.0 287850.0 ;
      RECT  315300.0 277350.0 316200.0 287850.0 ;
      RECT  318300.0 275250.0 319200.0 287850.0 ;
      RECT  335700.0 277350.0 336600.0 287850.0 ;
      RECT  338700.0 275250.0 339600.0 287850.0 ;
      RECT  345900.0 277350.0 346800.0 287850.0 ;
      RECT  348900.0 275250.0 349800.0 287850.0 ;
      RECT  356100.0 277350.0 357000.0 287850.0 ;
      RECT  359100.0 275250.0 360000.0 287850.0 ;
      RECT  376500.0 277350.0 377400.0 287850.0 ;
      RECT  379500.0 275250.0 380400.0 287850.0 ;
      RECT  386700.0 277350.0 387600.0 287850.0 ;
      RECT  389700.0 275250.0 390600.0 287850.0 ;
      RECT  396900.0 277350.0 397800.0 287850.0 ;
      RECT  399900.0 275250.0 400800.0 287850.0 ;
      RECT  417300.0 277350.0 418200.0 287850.0 ;
      RECT  420300.0 275250.0 421200.0 287850.0 ;
      RECT  427500.0 277350.0 428400.0 287850.0 ;
      RECT  430500.0 275250.0 431400.0 287850.0 ;
      RECT  437700.0 277350.0 438600.0 287850.0 ;
      RECT  440700.0 275250.0 441600.0 287850.0 ;
      RECT  458100.0 277350.0 459000.0 287850.0 ;
      RECT  461100.0 275250.0 462000.0 287850.0 ;
      RECT  468300.0 277350.0 469200.0 287850.0 ;
      RECT  471300.0 275250.0 472200.0 287850.0 ;
      RECT  478500.0 277350.0 479400.0 287850.0 ;
      RECT  481500.0 275250.0 482400.0 287850.0 ;
      RECT  498900.0 277350.0 499800.0 287850.0 ;
      RECT  501900.0 275250.0 502800.0 287850.0 ;
      RECT  509100.0 277350.0 510000.0 287850.0 ;
      RECT  512100.0 275250.0 513000.0 287850.0 ;
      RECT  519300.0 277350.0 520200.0 287850.0 ;
      RECT  522300.0 275250.0 523200.0 287850.0 ;
      RECT  203100.0 296550.0 204000.0 297450.0 ;
      RECT  203550.0 296550.0 204450.0 297450.0 ;
      RECT  203100.0 289650.0 204000.0 297000.0 ;
      RECT  203550.0 296550.0 204000.0 297450.0 ;
      RECT  203550.0 297000.0 204450.0 304350.0 ;
      RECT  206100.0 302850.0 207000.0 303750.0 ;
      RECT  205950.0 302850.0 206850.0 303750.0 ;
      RECT  206100.0 303300.0 207000.0 311550.0 ;
      RECT  206400.0 302850.0 206550.0 303750.0 ;
      RECT  205950.0 295050.0 206850.0 303300.0 ;
      RECT  202950.0 310950.0 204150.0 312150.0 ;
      RECT  205950.0 289050.0 207150.0 290250.0 ;
      RECT  203400.0 304350.0 204600.0 305550.0 ;
      RECT  205800.0 293850.0 207000.0 295050.0 ;
      RECT  209700.0 292050.0 210900.0 293250.0 ;
      RECT  203100.0 311550.0 204000.0 313350.0 ;
      RECT  206100.0 311550.0 207000.0 313350.0 ;
      RECT  203100.0 287850.0 204000.0 289650.0 ;
      RECT  206100.0 287850.0 207000.0 289650.0 ;
      RECT  199500.0 287850.0 200400.0 313350.0 ;
      RECT  209700.0 287850.0 210600.0 313350.0 ;
      RECT  213300.0 296550.0 214200.0 297450.0 ;
      RECT  213750.0 296550.0 214650.0 297450.0 ;
      RECT  213300.0 289650.0 214200.0 297000.0 ;
      RECT  213750.0 296550.0 214200.0 297450.0 ;
      RECT  213750.0 297000.0 214650.0 304350.0 ;
      RECT  216300.0 302850.0 217200.0 303750.0 ;
      RECT  216150.0 302850.0 217050.0 303750.0 ;
      RECT  216300.0 303300.0 217200.0 311550.0 ;
      RECT  216600.0 302850.0 216750.0 303750.0 ;
      RECT  216150.0 295050.0 217050.0 303300.0 ;
      RECT  213150.0 310950.0 214350.0 312150.0 ;
      RECT  216150.0 289050.0 217350.0 290250.0 ;
      RECT  213600.0 304350.0 214800.0 305550.0 ;
      RECT  216000.0 293850.0 217200.0 295050.0 ;
      RECT  219900.0 292050.0 221100.0 293250.0 ;
      RECT  213300.0 311550.0 214200.0 313350.0 ;
      RECT  216300.0 311550.0 217200.0 313350.0 ;
      RECT  213300.0 287850.0 214200.0 289650.0 ;
      RECT  216300.0 287850.0 217200.0 289650.0 ;
      RECT  209700.0 287850.0 210600.0 313350.0 ;
      RECT  219900.0 287850.0 220800.0 313350.0 ;
      RECT  223500.0 296550.0 224400.0 297450.0 ;
      RECT  223950.0 296550.0 224850.0 297450.0 ;
      RECT  223500.0 289650.0 224400.0 297000.0 ;
      RECT  223950.0 296550.0 224400.0 297450.0 ;
      RECT  223950.0 297000.0 224850.0 304350.0 ;
      RECT  226500.0 302850.0 227400.0 303750.0 ;
      RECT  226350.0 302850.0 227250.0 303750.0 ;
      RECT  226500.0 303300.0 227400.0 311550.0 ;
      RECT  226800.0 302850.0 226950.0 303750.0 ;
      RECT  226350.0 295050.0 227250.0 303300.0 ;
      RECT  223350.0 310950.0 224550.0 312150.0 ;
      RECT  226350.0 289050.0 227550.0 290250.0 ;
      RECT  223800.0 304350.0 225000.0 305550.0 ;
      RECT  226200.0 293850.0 227400.0 295050.0 ;
      RECT  230100.0 292050.0 231300.0 293250.0 ;
      RECT  223500.0 311550.0 224400.0 313350.0 ;
      RECT  226500.0 311550.0 227400.0 313350.0 ;
      RECT  223500.0 287850.0 224400.0 289650.0 ;
      RECT  226500.0 287850.0 227400.0 289650.0 ;
      RECT  219900.0 287850.0 220800.0 313350.0 ;
      RECT  230100.0 287850.0 231000.0 313350.0 ;
      RECT  233700.0 296550.0 234600.0 297450.0 ;
      RECT  234150.0 296550.0 235050.0 297450.0 ;
      RECT  233700.0 289650.0 234600.0 297000.0 ;
      RECT  234150.0 296550.0 234600.0 297450.0 ;
      RECT  234150.0 297000.0 235050.0 304350.0 ;
      RECT  236700.0 302850.0 237600.0 303750.0 ;
      RECT  236550.0 302850.0 237450.0 303750.0 ;
      RECT  236700.0 303300.0 237600.0 311550.0 ;
      RECT  237000.0 302850.0 237150.0 303750.0 ;
      RECT  236550.0 295050.0 237450.0 303300.0 ;
      RECT  233550.0 310950.0 234750.0 312150.0 ;
      RECT  236550.0 289050.0 237750.0 290250.0 ;
      RECT  234000.0 304350.0 235200.0 305550.0 ;
      RECT  236400.0 293850.0 237600.0 295050.0 ;
      RECT  240300.0 292050.0 241500.0 293250.0 ;
      RECT  233700.0 311550.0 234600.0 313350.0 ;
      RECT  236700.0 311550.0 237600.0 313350.0 ;
      RECT  233700.0 287850.0 234600.0 289650.0 ;
      RECT  236700.0 287850.0 237600.0 289650.0 ;
      RECT  230100.0 287850.0 231000.0 313350.0 ;
      RECT  240300.0 287850.0 241200.0 313350.0 ;
      RECT  243900.0 296550.0 244800.0 297450.0 ;
      RECT  244350.0 296550.0 245250.0 297450.0 ;
      RECT  243900.0 289650.0 244800.0 297000.0 ;
      RECT  244350.0 296550.0 244800.0 297450.0 ;
      RECT  244350.0 297000.0 245250.0 304350.0 ;
      RECT  246900.0 302850.0 247800.0 303750.0 ;
      RECT  246750.0 302850.0 247650.0 303750.0 ;
      RECT  246900.0 303300.0 247800.0 311550.0 ;
      RECT  247200.0 302850.0 247350.0 303750.0 ;
      RECT  246750.0 295050.0 247650.0 303300.0 ;
      RECT  243750.0 310950.0 244950.0 312150.0 ;
      RECT  246750.0 289050.0 247950.0 290250.0 ;
      RECT  244200.0 304350.0 245400.0 305550.0 ;
      RECT  246600.0 293850.0 247800.0 295050.0 ;
      RECT  250500.0 292050.0 251700.0 293250.0 ;
      RECT  243900.0 311550.0 244800.0 313350.0 ;
      RECT  246900.0 311550.0 247800.0 313350.0 ;
      RECT  243900.0 287850.0 244800.0 289650.0 ;
      RECT  246900.0 287850.0 247800.0 289650.0 ;
      RECT  240300.0 287850.0 241200.0 313350.0 ;
      RECT  250500.0 287850.0 251400.0 313350.0 ;
      RECT  254100.0 296550.0 255000.0 297450.0 ;
      RECT  254550.0 296550.0 255450.0 297450.0 ;
      RECT  254100.0 289650.0 255000.0 297000.0 ;
      RECT  254550.0 296550.0 255000.0 297450.0 ;
      RECT  254550.0 297000.0 255450.0 304350.0 ;
      RECT  257100.0 302850.0 258000.0 303750.0 ;
      RECT  256950.0 302850.0 257850.0 303750.0 ;
      RECT  257100.0 303300.0 258000.0 311550.0 ;
      RECT  257400.0 302850.0 257550.0 303750.0 ;
      RECT  256950.0 295050.0 257850.0 303300.0 ;
      RECT  253950.0 310950.0 255150.0 312150.0 ;
      RECT  256950.0 289050.0 258150.0 290250.0 ;
      RECT  254400.0 304350.0 255600.0 305550.0 ;
      RECT  256800.0 293850.0 258000.0 295050.0 ;
      RECT  260700.0 292050.0 261900.0 293250.0 ;
      RECT  254100.0 311550.0 255000.0 313350.0 ;
      RECT  257100.0 311550.0 258000.0 313350.0 ;
      RECT  254100.0 287850.0 255000.0 289650.0 ;
      RECT  257100.0 287850.0 258000.0 289650.0 ;
      RECT  250500.0 287850.0 251400.0 313350.0 ;
      RECT  260700.0 287850.0 261600.0 313350.0 ;
      RECT  264300.0 296550.0 265200.0 297450.0 ;
      RECT  264750.0 296550.0 265650.0 297450.0 ;
      RECT  264300.0 289650.0 265200.0 297000.0 ;
      RECT  264750.0 296550.0 265200.0 297450.0 ;
      RECT  264750.0 297000.0 265650.0 304350.0 ;
      RECT  267300.0 302850.0 268200.0 303750.0 ;
      RECT  267150.0 302850.0 268050.0 303750.0 ;
      RECT  267300.0 303300.0 268200.0 311550.0 ;
      RECT  267600.0 302850.0 267750.0 303750.0 ;
      RECT  267150.0 295050.0 268050.0 303300.0 ;
      RECT  264150.0 310950.0 265350.0 312150.0 ;
      RECT  267150.0 289050.0 268350.0 290250.0 ;
      RECT  264600.0 304350.0 265800.0 305550.0 ;
      RECT  267000.0 293850.0 268200.0 295050.0 ;
      RECT  270900.0 292050.0 272100.0 293250.0 ;
      RECT  264300.0 311550.0 265200.0 313350.0 ;
      RECT  267300.0 311550.0 268200.0 313350.0 ;
      RECT  264300.0 287850.0 265200.0 289650.0 ;
      RECT  267300.0 287850.0 268200.0 289650.0 ;
      RECT  260700.0 287850.0 261600.0 313350.0 ;
      RECT  270900.0 287850.0 271800.0 313350.0 ;
      RECT  274500.0 296550.0 275400.0 297450.0 ;
      RECT  274950.0 296550.0 275850.0 297450.0 ;
      RECT  274500.0 289650.0 275400.0 297000.0 ;
      RECT  274950.0 296550.0 275400.0 297450.0 ;
      RECT  274950.0 297000.0 275850.0 304350.0 ;
      RECT  277500.0 302850.0 278400.0 303750.0 ;
      RECT  277350.0 302850.0 278250.0 303750.0 ;
      RECT  277500.0 303300.0 278400.0 311550.0 ;
      RECT  277800.0 302850.0 277950.0 303750.0 ;
      RECT  277350.0 295050.0 278250.0 303300.0 ;
      RECT  274350.0 310950.0 275550.0 312150.0 ;
      RECT  277350.0 289050.0 278550.0 290250.0 ;
      RECT  274800.0 304350.0 276000.0 305550.0 ;
      RECT  277200.0 293850.0 278400.0 295050.0 ;
      RECT  281100.0 292050.0 282300.0 293250.0 ;
      RECT  274500.0 311550.0 275400.0 313350.0 ;
      RECT  277500.0 311550.0 278400.0 313350.0 ;
      RECT  274500.0 287850.0 275400.0 289650.0 ;
      RECT  277500.0 287850.0 278400.0 289650.0 ;
      RECT  270900.0 287850.0 271800.0 313350.0 ;
      RECT  281100.0 287850.0 282000.0 313350.0 ;
      RECT  284700.0 296550.0 285600.0 297450.0 ;
      RECT  285150.0 296550.0 286050.0 297450.0 ;
      RECT  284700.0 289650.0 285600.0 297000.0 ;
      RECT  285150.0 296550.0 285600.0 297450.0 ;
      RECT  285150.0 297000.0 286050.0 304350.0 ;
      RECT  287700.0 302850.0 288600.0 303750.0 ;
      RECT  287550.0 302850.0 288450.0 303750.0 ;
      RECT  287700.0 303300.0 288600.0 311550.0 ;
      RECT  288000.0 302850.0 288150.0 303750.0 ;
      RECT  287550.0 295050.0 288450.0 303300.0 ;
      RECT  284550.0 310950.0 285750.0 312150.0 ;
      RECT  287550.0 289050.0 288750.0 290250.0 ;
      RECT  285000.0 304350.0 286200.0 305550.0 ;
      RECT  287400.0 293850.0 288600.0 295050.0 ;
      RECT  291300.0 292050.0 292500.0 293250.0 ;
      RECT  284700.0 311550.0 285600.0 313350.0 ;
      RECT  287700.0 311550.0 288600.0 313350.0 ;
      RECT  284700.0 287850.0 285600.0 289650.0 ;
      RECT  287700.0 287850.0 288600.0 289650.0 ;
      RECT  281100.0 287850.0 282000.0 313350.0 ;
      RECT  291300.0 287850.0 292200.0 313350.0 ;
      RECT  294900.0 296550.0 295800.0 297450.0 ;
      RECT  295350.0 296550.0 296250.0 297450.0 ;
      RECT  294900.0 289650.0 295800.0 297000.0 ;
      RECT  295350.0 296550.0 295800.0 297450.0 ;
      RECT  295350.0 297000.0 296250.0 304350.0 ;
      RECT  297900.0 302850.0 298800.0 303750.0 ;
      RECT  297750.0 302850.0 298650.0 303750.0 ;
      RECT  297900.0 303300.0 298800.0 311550.0 ;
      RECT  298200.0 302850.0 298350.0 303750.0 ;
      RECT  297750.0 295050.0 298650.0 303300.0 ;
      RECT  294750.0 310950.0 295950.0 312150.0 ;
      RECT  297750.0 289050.0 298950.0 290250.0 ;
      RECT  295200.0 304350.0 296400.0 305550.0 ;
      RECT  297600.0 293850.0 298800.0 295050.0 ;
      RECT  301500.0 292050.0 302700.0 293250.0 ;
      RECT  294900.0 311550.0 295800.0 313350.0 ;
      RECT  297900.0 311550.0 298800.0 313350.0 ;
      RECT  294900.0 287850.0 295800.0 289650.0 ;
      RECT  297900.0 287850.0 298800.0 289650.0 ;
      RECT  291300.0 287850.0 292200.0 313350.0 ;
      RECT  301500.0 287850.0 302400.0 313350.0 ;
      RECT  305100.0 296550.0 306000.0 297450.0 ;
      RECT  305550.0 296550.0 306450.0 297450.0 ;
      RECT  305100.0 289650.0 306000.0 297000.0 ;
      RECT  305550.0 296550.0 306000.0 297450.0 ;
      RECT  305550.0 297000.0 306450.0 304350.0 ;
      RECT  308100.0 302850.0 309000.0 303750.0 ;
      RECT  307950.0 302850.0 308850.0 303750.0 ;
      RECT  308100.0 303300.0 309000.0 311550.0 ;
      RECT  308400.0 302850.0 308550.0 303750.0 ;
      RECT  307950.0 295050.0 308850.0 303300.0 ;
      RECT  304950.0 310950.0 306150.0 312150.0 ;
      RECT  307950.0 289050.0 309150.0 290250.0 ;
      RECT  305400.0 304350.0 306600.0 305550.0 ;
      RECT  307800.0 293850.0 309000.0 295050.0 ;
      RECT  311700.0 292050.0 312900.0 293250.0 ;
      RECT  305100.0 311550.0 306000.0 313350.0 ;
      RECT  308100.0 311550.0 309000.0 313350.0 ;
      RECT  305100.0 287850.0 306000.0 289650.0 ;
      RECT  308100.0 287850.0 309000.0 289650.0 ;
      RECT  301500.0 287850.0 302400.0 313350.0 ;
      RECT  311700.0 287850.0 312600.0 313350.0 ;
      RECT  315300.0 296550.0 316200.0 297450.0 ;
      RECT  315750.0 296550.0 316650.0 297450.0 ;
      RECT  315300.0 289650.0 316200.0 297000.0 ;
      RECT  315750.0 296550.0 316200.0 297450.0 ;
      RECT  315750.0 297000.0 316650.0 304350.0 ;
      RECT  318300.0 302850.0 319200.0 303750.0 ;
      RECT  318150.0 302850.0 319050.0 303750.0 ;
      RECT  318300.0 303300.0 319200.0 311550.0 ;
      RECT  318600.0 302850.0 318750.0 303750.0 ;
      RECT  318150.0 295050.0 319050.0 303300.0 ;
      RECT  315150.0 310950.0 316350.0 312150.0 ;
      RECT  318150.0 289050.0 319350.0 290250.0 ;
      RECT  315600.0 304350.0 316800.0 305550.0 ;
      RECT  318000.0 293850.0 319200.0 295050.0 ;
      RECT  321900.0 292050.0 323100.0 293250.0 ;
      RECT  315300.0 311550.0 316200.0 313350.0 ;
      RECT  318300.0 311550.0 319200.0 313350.0 ;
      RECT  315300.0 287850.0 316200.0 289650.0 ;
      RECT  318300.0 287850.0 319200.0 289650.0 ;
      RECT  311700.0 287850.0 312600.0 313350.0 ;
      RECT  321900.0 287850.0 322800.0 313350.0 ;
      RECT  325500.0 296550.0 326400.0 297450.0 ;
      RECT  325950.0 296550.0 326850.0 297450.0 ;
      RECT  325500.0 289650.0 326400.0 297000.0 ;
      RECT  325950.0 296550.0 326400.0 297450.0 ;
      RECT  325950.0 297000.0 326850.0 304350.0 ;
      RECT  328500.0 302850.0 329400.0 303750.0 ;
      RECT  328350.0 302850.0 329250.0 303750.0 ;
      RECT  328500.0 303300.0 329400.0 311550.0 ;
      RECT  328800.0 302850.0 328950.0 303750.0 ;
      RECT  328350.0 295050.0 329250.0 303300.0 ;
      RECT  325350.0 310950.0 326550.0 312150.0 ;
      RECT  328350.0 289050.0 329550.0 290250.0 ;
      RECT  325800.0 304350.0 327000.0 305550.0 ;
      RECT  328200.0 293850.0 329400.0 295050.0 ;
      RECT  332100.0 292050.0 333300.0 293250.0 ;
      RECT  325500.0 311550.0 326400.0 313350.0 ;
      RECT  328500.0 311550.0 329400.0 313350.0 ;
      RECT  325500.0 287850.0 326400.0 289650.0 ;
      RECT  328500.0 287850.0 329400.0 289650.0 ;
      RECT  321900.0 287850.0 322800.0 313350.0 ;
      RECT  332100.0 287850.0 333000.0 313350.0 ;
      RECT  335700.0 296550.0 336600.0 297450.0 ;
      RECT  336150.0 296550.0 337050.0 297450.0 ;
      RECT  335700.0 289650.0 336600.0 297000.0 ;
      RECT  336150.0 296550.0 336600.0 297450.0 ;
      RECT  336150.0 297000.0 337050.0 304350.0 ;
      RECT  338700.0 302850.0 339600.0 303750.0 ;
      RECT  338550.0 302850.0 339450.0 303750.0 ;
      RECT  338700.0 303300.0 339600.0 311550.0 ;
      RECT  339000.0 302850.0 339150.0 303750.0 ;
      RECT  338550.0 295050.0 339450.0 303300.0 ;
      RECT  335550.0 310950.0 336750.0 312150.0 ;
      RECT  338550.0 289050.0 339750.0 290250.0 ;
      RECT  336000.0 304350.0 337200.0 305550.0 ;
      RECT  338400.0 293850.0 339600.0 295050.0 ;
      RECT  342300.0 292050.0 343500.0 293250.0 ;
      RECT  335700.0 311550.0 336600.0 313350.0 ;
      RECT  338700.0 311550.0 339600.0 313350.0 ;
      RECT  335700.0 287850.0 336600.0 289650.0 ;
      RECT  338700.0 287850.0 339600.0 289650.0 ;
      RECT  332100.0 287850.0 333000.0 313350.0 ;
      RECT  342300.0 287850.0 343200.0 313350.0 ;
      RECT  345900.0 296550.0 346800.0 297450.0 ;
      RECT  346350.0 296550.0 347250.0 297450.0 ;
      RECT  345900.0 289650.0 346800.0 297000.0 ;
      RECT  346350.0 296550.0 346800.0 297450.0 ;
      RECT  346350.0 297000.0 347250.0 304350.0 ;
      RECT  348900.0 302850.0 349800.0 303750.0 ;
      RECT  348750.0 302850.0 349650.0 303750.0 ;
      RECT  348900.0 303300.0 349800.0 311550.0 ;
      RECT  349200.0 302850.0 349350.0 303750.0 ;
      RECT  348750.0 295050.0 349650.0 303300.0 ;
      RECT  345750.0 310950.0 346950.0 312150.0 ;
      RECT  348750.0 289050.0 349950.0 290250.0 ;
      RECT  346200.0 304350.0 347400.0 305550.0 ;
      RECT  348600.0 293850.0 349800.0 295050.0 ;
      RECT  352500.0 292050.0 353700.0 293250.0 ;
      RECT  345900.0 311550.0 346800.0 313350.0 ;
      RECT  348900.0 311550.0 349800.0 313350.0 ;
      RECT  345900.0 287850.0 346800.0 289650.0 ;
      RECT  348900.0 287850.0 349800.0 289650.0 ;
      RECT  342300.0 287850.0 343200.0 313350.0 ;
      RECT  352500.0 287850.0 353400.0 313350.0 ;
      RECT  356100.0 296550.0 357000.0 297450.0 ;
      RECT  356550.0 296550.0 357450.0 297450.0 ;
      RECT  356100.0 289650.0 357000.0 297000.0 ;
      RECT  356550.0 296550.0 357000.0 297450.0 ;
      RECT  356550.0 297000.0 357450.0 304350.0 ;
      RECT  359100.0 302850.0 360000.0 303750.0 ;
      RECT  358950.0 302850.0 359850.0 303750.0 ;
      RECT  359100.0 303300.0 360000.0 311550.0 ;
      RECT  359400.0 302850.0 359550.0 303750.0 ;
      RECT  358950.0 295050.0 359850.0 303300.0 ;
      RECT  355950.0 310950.0 357150.0 312150.0 ;
      RECT  358950.0 289050.0 360150.0 290250.0 ;
      RECT  356400.0 304350.0 357600.0 305550.0 ;
      RECT  358800.0 293850.0 360000.0 295050.0 ;
      RECT  362700.0 292050.0 363900.0 293250.0 ;
      RECT  356100.0 311550.0 357000.0 313350.0 ;
      RECT  359100.0 311550.0 360000.0 313350.0 ;
      RECT  356100.0 287850.0 357000.0 289650.0 ;
      RECT  359100.0 287850.0 360000.0 289650.0 ;
      RECT  352500.0 287850.0 353400.0 313350.0 ;
      RECT  362700.0 287850.0 363600.0 313350.0 ;
      RECT  366300.0 296550.0 367200.0 297450.0 ;
      RECT  366750.0 296550.0 367650.0 297450.0 ;
      RECT  366300.0 289650.0 367200.0 297000.0 ;
      RECT  366750.0 296550.0 367200.0 297450.0 ;
      RECT  366750.0 297000.0 367650.0 304350.0 ;
      RECT  369300.0 302850.0 370200.0 303750.0 ;
      RECT  369150.0 302850.0 370050.0 303750.0 ;
      RECT  369300.0 303300.0 370200.0 311550.0 ;
      RECT  369600.0 302850.0 369750.0 303750.0 ;
      RECT  369150.0 295050.0 370050.0 303300.0 ;
      RECT  366150.0 310950.0 367350.0 312150.0 ;
      RECT  369150.0 289050.0 370350.0 290250.0 ;
      RECT  366600.0 304350.0 367800.0 305550.0 ;
      RECT  369000.0 293850.0 370200.0 295050.0 ;
      RECT  372900.0 292050.0 374100.0 293250.0 ;
      RECT  366300.0 311550.0 367200.0 313350.0 ;
      RECT  369300.0 311550.0 370200.0 313350.0 ;
      RECT  366300.0 287850.0 367200.0 289650.0 ;
      RECT  369300.0 287850.0 370200.0 289650.0 ;
      RECT  362700.0 287850.0 363600.0 313350.0 ;
      RECT  372900.0 287850.0 373800.0 313350.0 ;
      RECT  376500.0 296550.0 377400.0 297450.0 ;
      RECT  376950.0 296550.0 377850.0 297450.0 ;
      RECT  376500.0 289650.0 377400.0 297000.0 ;
      RECT  376950.0 296550.0 377400.0 297450.0 ;
      RECT  376950.0 297000.0 377850.0 304350.0 ;
      RECT  379500.0 302850.0 380400.0 303750.0 ;
      RECT  379350.0 302850.0 380250.0 303750.0 ;
      RECT  379500.0 303300.0 380400.0 311550.0 ;
      RECT  379800.0 302850.0 379950.0 303750.0 ;
      RECT  379350.0 295050.0 380250.0 303300.0 ;
      RECT  376350.0 310950.0 377550.0 312150.0 ;
      RECT  379350.0 289050.0 380550.0 290250.0 ;
      RECT  376800.0 304350.0 378000.0 305550.0 ;
      RECT  379200.0 293850.0 380400.0 295050.0 ;
      RECT  383100.0 292050.0 384300.0 293250.0 ;
      RECT  376500.0 311550.0 377400.0 313350.0 ;
      RECT  379500.0 311550.0 380400.0 313350.0 ;
      RECT  376500.0 287850.0 377400.0 289650.0 ;
      RECT  379500.0 287850.0 380400.0 289650.0 ;
      RECT  372900.0 287850.0 373800.0 313350.0 ;
      RECT  383100.0 287850.0 384000.0 313350.0 ;
      RECT  386700.0 296550.0 387600.0 297450.0 ;
      RECT  387150.0 296550.0 388050.0 297450.0 ;
      RECT  386700.0 289650.0 387600.0 297000.0 ;
      RECT  387150.0 296550.0 387600.0 297450.0 ;
      RECT  387150.0 297000.0 388050.0 304350.0 ;
      RECT  389700.0 302850.0 390600.0 303750.0 ;
      RECT  389550.0 302850.0 390450.0 303750.0 ;
      RECT  389700.0 303300.0 390600.0 311550.0 ;
      RECT  390000.0 302850.0 390150.0 303750.0 ;
      RECT  389550.0 295050.0 390450.0 303300.0 ;
      RECT  386550.0 310950.0 387750.0 312150.0 ;
      RECT  389550.0 289050.0 390750.0 290250.0 ;
      RECT  387000.0 304350.0 388200.0 305550.0 ;
      RECT  389400.0 293850.0 390600.0 295050.0 ;
      RECT  393300.0 292050.0 394500.0 293250.0 ;
      RECT  386700.0 311550.0 387600.0 313350.0 ;
      RECT  389700.0 311550.0 390600.0 313350.0 ;
      RECT  386700.0 287850.0 387600.0 289650.0 ;
      RECT  389700.0 287850.0 390600.0 289650.0 ;
      RECT  383100.0 287850.0 384000.0 313350.0 ;
      RECT  393300.0 287850.0 394200.0 313350.0 ;
      RECT  396900.0 296550.0 397800.0 297450.0 ;
      RECT  397350.0 296550.0 398250.0 297450.0 ;
      RECT  396900.0 289650.0 397800.0 297000.0 ;
      RECT  397350.0 296550.0 397800.0 297450.0 ;
      RECT  397350.0 297000.0 398250.0 304350.0 ;
      RECT  399900.0 302850.0 400800.0 303750.0 ;
      RECT  399750.0 302850.0 400650.0 303750.0 ;
      RECT  399900.0 303300.0 400800.0 311550.0 ;
      RECT  400200.0 302850.0 400350.0 303750.0 ;
      RECT  399750.0 295050.0 400650.0 303300.0 ;
      RECT  396750.0 310950.0 397950.0 312150.0 ;
      RECT  399750.0 289050.0 400950.0 290250.0 ;
      RECT  397200.0 304350.0 398400.0 305550.0 ;
      RECT  399600.0 293850.0 400800.0 295050.0 ;
      RECT  403500.0 292050.0 404700.0 293250.0 ;
      RECT  396900.0 311550.0 397800.0 313350.0 ;
      RECT  399900.0 311550.0 400800.0 313350.0 ;
      RECT  396900.0 287850.0 397800.0 289650.0 ;
      RECT  399900.0 287850.0 400800.0 289650.0 ;
      RECT  393300.0 287850.0 394200.0 313350.0 ;
      RECT  403500.0 287850.0 404400.0 313350.0 ;
      RECT  407100.0 296550.0 408000.0 297450.0 ;
      RECT  407550.0 296550.0 408450.0 297450.0 ;
      RECT  407100.0 289650.0 408000.0 297000.0 ;
      RECT  407550.0 296550.0 408000.0 297450.0 ;
      RECT  407550.0 297000.0 408450.0 304350.0 ;
      RECT  410100.0 302850.0 411000.0 303750.0 ;
      RECT  409950.0 302850.0 410850.0 303750.0 ;
      RECT  410100.0 303300.0 411000.0 311550.0 ;
      RECT  410400.0 302850.0 410550.0 303750.0 ;
      RECT  409950.0 295050.0 410850.0 303300.0 ;
      RECT  406950.0 310950.0 408150.0 312150.0 ;
      RECT  409950.0 289050.0 411150.0 290250.0 ;
      RECT  407400.0 304350.0 408600.0 305550.0 ;
      RECT  409800.0 293850.0 411000.0 295050.0 ;
      RECT  413700.0 292050.0 414900.0 293250.0 ;
      RECT  407100.0 311550.0 408000.0 313350.0 ;
      RECT  410100.0 311550.0 411000.0 313350.0 ;
      RECT  407100.0 287850.0 408000.0 289650.0 ;
      RECT  410100.0 287850.0 411000.0 289650.0 ;
      RECT  403500.0 287850.0 404400.0 313350.0 ;
      RECT  413700.0 287850.0 414600.0 313350.0 ;
      RECT  417300.0 296550.0 418200.0 297450.0 ;
      RECT  417750.0 296550.0 418650.0 297450.0 ;
      RECT  417300.0 289650.0 418200.0 297000.0 ;
      RECT  417750.0 296550.0 418200.0 297450.0 ;
      RECT  417750.0 297000.0 418650.0 304350.0 ;
      RECT  420300.0 302850.0 421200.0 303750.0 ;
      RECT  420150.0 302850.0 421050.0 303750.0 ;
      RECT  420300.0 303300.0 421200.0 311550.0 ;
      RECT  420600.0 302850.0 420750.0 303750.0 ;
      RECT  420150.0 295050.0 421050.0 303300.0 ;
      RECT  417150.0 310950.0 418350.0 312150.0 ;
      RECT  420150.0 289050.0 421350.0 290250.0 ;
      RECT  417600.0 304350.0 418800.0 305550.0 ;
      RECT  420000.0 293850.0 421200.0 295050.0 ;
      RECT  423900.0 292050.0 425100.0 293250.0 ;
      RECT  417300.0 311550.0 418200.0 313350.0 ;
      RECT  420300.0 311550.0 421200.0 313350.0 ;
      RECT  417300.0 287850.0 418200.0 289650.0 ;
      RECT  420300.0 287850.0 421200.0 289650.0 ;
      RECT  413700.0 287850.0 414600.0 313350.0 ;
      RECT  423900.0 287850.0 424800.0 313350.0 ;
      RECT  427500.0 296550.0 428400.0 297450.0 ;
      RECT  427950.0 296550.0 428850.0 297450.0 ;
      RECT  427500.0 289650.0 428400.0 297000.0 ;
      RECT  427950.0 296550.0 428400.0 297450.0 ;
      RECT  427950.0 297000.0 428850.0 304350.0 ;
      RECT  430500.0 302850.0 431400.0 303750.0 ;
      RECT  430350.0 302850.0 431250.0 303750.0 ;
      RECT  430500.0 303300.0 431400.0 311550.0 ;
      RECT  430800.0 302850.0 430950.0 303750.0 ;
      RECT  430350.0 295050.0 431250.0 303300.0 ;
      RECT  427350.0 310950.0 428550.0 312150.0 ;
      RECT  430350.0 289050.0 431550.0 290250.0 ;
      RECT  427800.0 304350.0 429000.0 305550.0 ;
      RECT  430200.0 293850.0 431400.0 295050.0 ;
      RECT  434100.0 292050.0 435300.0 293250.0 ;
      RECT  427500.0 311550.0 428400.0 313350.0 ;
      RECT  430500.0 311550.0 431400.0 313350.0 ;
      RECT  427500.0 287850.0 428400.0 289650.0 ;
      RECT  430500.0 287850.0 431400.0 289650.0 ;
      RECT  423900.0 287850.0 424800.0 313350.0 ;
      RECT  434100.0 287850.0 435000.0 313350.0 ;
      RECT  437700.0 296550.0 438600.0 297450.0 ;
      RECT  438150.0 296550.0 439050.0 297450.0 ;
      RECT  437700.0 289650.0 438600.0 297000.0 ;
      RECT  438150.0 296550.0 438600.0 297450.0 ;
      RECT  438150.0 297000.0 439050.0 304350.0 ;
      RECT  440700.0 302850.0 441600.0 303750.0 ;
      RECT  440550.0 302850.0 441450.0 303750.0 ;
      RECT  440700.0 303300.0 441600.0 311550.0 ;
      RECT  441000.0 302850.0 441150.0 303750.0 ;
      RECT  440550.0 295050.0 441450.0 303300.0 ;
      RECT  437550.0 310950.0 438750.0 312150.0 ;
      RECT  440550.0 289050.0 441750.0 290250.0 ;
      RECT  438000.0 304350.0 439200.0 305550.0 ;
      RECT  440400.0 293850.0 441600.0 295050.0 ;
      RECT  444300.0 292050.0 445500.0 293250.0 ;
      RECT  437700.0 311550.0 438600.0 313350.0 ;
      RECT  440700.0 311550.0 441600.0 313350.0 ;
      RECT  437700.0 287850.0 438600.0 289650.0 ;
      RECT  440700.0 287850.0 441600.0 289650.0 ;
      RECT  434100.0 287850.0 435000.0 313350.0 ;
      RECT  444300.0 287850.0 445200.0 313350.0 ;
      RECT  447900.0 296550.0 448800.0 297450.0 ;
      RECT  448350.0 296550.0 449250.0 297450.0 ;
      RECT  447900.0 289650.0 448800.0 297000.0 ;
      RECT  448350.0 296550.0 448800.0 297450.0 ;
      RECT  448350.0 297000.0 449250.0 304350.0 ;
      RECT  450900.0 302850.0 451800.0 303750.0 ;
      RECT  450750.0 302850.0 451650.0 303750.0 ;
      RECT  450900.0 303300.0 451800.0 311550.0 ;
      RECT  451200.0 302850.0 451350.0 303750.0 ;
      RECT  450750.0 295050.0 451650.0 303300.0 ;
      RECT  447750.0 310950.0 448950.0 312150.0 ;
      RECT  450750.0 289050.0 451950.0 290250.0 ;
      RECT  448200.0 304350.0 449400.0 305550.0 ;
      RECT  450600.0 293850.0 451800.0 295050.0 ;
      RECT  454500.0 292050.0 455700.0 293250.0 ;
      RECT  447900.0 311550.0 448800.0 313350.0 ;
      RECT  450900.0 311550.0 451800.0 313350.0 ;
      RECT  447900.0 287850.0 448800.0 289650.0 ;
      RECT  450900.0 287850.0 451800.0 289650.0 ;
      RECT  444300.0 287850.0 445200.0 313350.0 ;
      RECT  454500.0 287850.0 455400.0 313350.0 ;
      RECT  458100.0 296550.0 459000.0 297450.0 ;
      RECT  458550.0 296550.0 459450.0 297450.0 ;
      RECT  458100.0 289650.0 459000.0 297000.0 ;
      RECT  458550.0 296550.0 459000.0 297450.0 ;
      RECT  458550.0 297000.0 459450.0 304350.0 ;
      RECT  461100.0 302850.0 462000.0 303750.0 ;
      RECT  460950.0 302850.0 461850.0 303750.0 ;
      RECT  461100.0 303300.0 462000.0 311550.0 ;
      RECT  461400.0 302850.0 461550.0 303750.0 ;
      RECT  460950.0 295050.0 461850.0 303300.0 ;
      RECT  457950.0 310950.0 459150.0 312150.0 ;
      RECT  460950.0 289050.0 462150.0 290250.0 ;
      RECT  458400.0 304350.0 459600.0 305550.0 ;
      RECT  460800.0 293850.0 462000.0 295050.0 ;
      RECT  464700.0 292050.0 465900.0 293250.0 ;
      RECT  458100.0 311550.0 459000.0 313350.0 ;
      RECT  461100.0 311550.0 462000.0 313350.0 ;
      RECT  458100.0 287850.0 459000.0 289650.0 ;
      RECT  461100.0 287850.0 462000.0 289650.0 ;
      RECT  454500.0 287850.0 455400.0 313350.0 ;
      RECT  464700.0 287850.0 465600.0 313350.0 ;
      RECT  468300.0 296550.0 469200.0 297450.0 ;
      RECT  468750.0 296550.0 469650.0 297450.0 ;
      RECT  468300.0 289650.0 469200.0 297000.0 ;
      RECT  468750.0 296550.0 469200.0 297450.0 ;
      RECT  468750.0 297000.0 469650.0 304350.0 ;
      RECT  471300.0 302850.0 472200.0 303750.0 ;
      RECT  471150.0 302850.0 472050.0 303750.0 ;
      RECT  471300.0 303300.0 472200.0 311550.0 ;
      RECT  471600.0 302850.0 471750.0 303750.0 ;
      RECT  471150.0 295050.0 472050.0 303300.0 ;
      RECT  468150.0 310950.0 469350.0 312150.0 ;
      RECT  471150.0 289050.0 472350.0 290250.0 ;
      RECT  468600.0 304350.0 469800.0 305550.0 ;
      RECT  471000.0 293850.0 472200.0 295050.0 ;
      RECT  474900.0 292050.0 476100.0 293250.0 ;
      RECT  468300.0 311550.0 469200.0 313350.0 ;
      RECT  471300.0 311550.0 472200.0 313350.0 ;
      RECT  468300.0 287850.0 469200.0 289650.0 ;
      RECT  471300.0 287850.0 472200.0 289650.0 ;
      RECT  464700.0 287850.0 465600.0 313350.0 ;
      RECT  474900.0 287850.0 475800.0 313350.0 ;
      RECT  478500.0 296550.0 479400.0 297450.0 ;
      RECT  478950.0 296550.0 479850.0 297450.0 ;
      RECT  478500.0 289650.0 479400.0 297000.0 ;
      RECT  478950.0 296550.0 479400.0 297450.0 ;
      RECT  478950.0 297000.0 479850.0 304350.0 ;
      RECT  481500.0 302850.0 482400.0 303750.0 ;
      RECT  481350.0 302850.0 482250.0 303750.0 ;
      RECT  481500.0 303300.0 482400.0 311550.0 ;
      RECT  481800.0 302850.0 481950.0 303750.0 ;
      RECT  481350.0 295050.0 482250.0 303300.0 ;
      RECT  478350.0 310950.0 479550.0 312150.0 ;
      RECT  481350.0 289050.0 482550.0 290250.0 ;
      RECT  478800.0 304350.0 480000.0 305550.0 ;
      RECT  481200.0 293850.0 482400.0 295050.0 ;
      RECT  485100.0 292050.0 486300.0 293250.0 ;
      RECT  478500.0 311550.0 479400.0 313350.0 ;
      RECT  481500.0 311550.0 482400.0 313350.0 ;
      RECT  478500.0 287850.0 479400.0 289650.0 ;
      RECT  481500.0 287850.0 482400.0 289650.0 ;
      RECT  474900.0 287850.0 475800.0 313350.0 ;
      RECT  485100.0 287850.0 486000.0 313350.0 ;
      RECT  488700.0 296550.0 489600.0 297450.0 ;
      RECT  489150.0 296550.0 490050.0 297450.0 ;
      RECT  488700.0 289650.0 489600.0 297000.0 ;
      RECT  489150.0 296550.0 489600.0 297450.0 ;
      RECT  489150.0 297000.0 490050.0 304350.0 ;
      RECT  491700.0 302850.0 492600.0 303750.0 ;
      RECT  491550.0 302850.0 492450.0 303750.0 ;
      RECT  491700.0 303300.0 492600.0 311550.0 ;
      RECT  492000.0 302850.0 492150.0 303750.0 ;
      RECT  491550.0 295050.0 492450.0 303300.0 ;
      RECT  488550.0 310950.0 489750.0 312150.0 ;
      RECT  491550.0 289050.0 492750.0 290250.0 ;
      RECT  489000.0 304350.0 490200.0 305550.0 ;
      RECT  491400.0 293850.0 492600.0 295050.0 ;
      RECT  495300.0 292050.0 496500.0 293250.0 ;
      RECT  488700.0 311550.0 489600.0 313350.0 ;
      RECT  491700.0 311550.0 492600.0 313350.0 ;
      RECT  488700.0 287850.0 489600.0 289650.0 ;
      RECT  491700.0 287850.0 492600.0 289650.0 ;
      RECT  485100.0 287850.0 486000.0 313350.0 ;
      RECT  495300.0 287850.0 496200.0 313350.0 ;
      RECT  498900.0 296550.0 499800.0 297450.0 ;
      RECT  499350.0 296550.0 500250.0 297450.0 ;
      RECT  498900.0 289650.0 499800.0 297000.0 ;
      RECT  499350.0 296550.0 499800.0 297450.0 ;
      RECT  499350.0 297000.0 500250.0 304350.0 ;
      RECT  501900.0 302850.0 502800.0 303750.0 ;
      RECT  501750.0 302850.0 502650.0 303750.0 ;
      RECT  501900.0 303300.0 502800.0 311550.0 ;
      RECT  502200.0 302850.0 502350.0 303750.0 ;
      RECT  501750.0 295050.0 502650.0 303300.0 ;
      RECT  498750.0 310950.0 499950.0 312150.0 ;
      RECT  501750.0 289050.0 502950.0 290250.0 ;
      RECT  499200.0 304350.0 500400.0 305550.0 ;
      RECT  501600.0 293850.0 502800.0 295050.0 ;
      RECT  505500.0 292050.0 506700.0 293250.0 ;
      RECT  498900.0 311550.0 499800.0 313350.0 ;
      RECT  501900.0 311550.0 502800.0 313350.0 ;
      RECT  498900.0 287850.0 499800.0 289650.0 ;
      RECT  501900.0 287850.0 502800.0 289650.0 ;
      RECT  495300.0 287850.0 496200.0 313350.0 ;
      RECT  505500.0 287850.0 506400.0 313350.0 ;
      RECT  509100.0 296550.0 510000.0 297450.0 ;
      RECT  509550.0 296550.0 510450.0 297450.0 ;
      RECT  509100.0 289650.0 510000.0 297000.0 ;
      RECT  509550.0 296550.0 510000.0 297450.0 ;
      RECT  509550.0 297000.0 510450.0 304350.0 ;
      RECT  512100.0 302850.0 513000.0 303750.0 ;
      RECT  511950.0 302850.0 512850.0 303750.0 ;
      RECT  512100.0 303300.0 513000.0 311550.0 ;
      RECT  512400.0 302850.0 512550.0 303750.0 ;
      RECT  511950.0 295050.0 512850.0 303300.0 ;
      RECT  508950.0 310950.0 510150.0 312150.0 ;
      RECT  511950.0 289050.0 513150.0 290250.0 ;
      RECT  509400.0 304350.0 510600.0 305550.0 ;
      RECT  511800.0 293850.0 513000.0 295050.0 ;
      RECT  515700.0 292050.0 516900.0 293250.0 ;
      RECT  509100.0 311550.0 510000.0 313350.0 ;
      RECT  512100.0 311550.0 513000.0 313350.0 ;
      RECT  509100.0 287850.0 510000.0 289650.0 ;
      RECT  512100.0 287850.0 513000.0 289650.0 ;
      RECT  505500.0 287850.0 506400.0 313350.0 ;
      RECT  515700.0 287850.0 516600.0 313350.0 ;
      RECT  519300.0 296550.0 520200.0 297450.0 ;
      RECT  519750.0 296550.0 520650.0 297450.0 ;
      RECT  519300.0 289650.0 520200.0 297000.0 ;
      RECT  519750.0 296550.0 520200.0 297450.0 ;
      RECT  519750.0 297000.0 520650.0 304350.0 ;
      RECT  522300.0 302850.0 523200.0 303750.0 ;
      RECT  522150.0 302850.0 523050.0 303750.0 ;
      RECT  522300.0 303300.0 523200.0 311550.0 ;
      RECT  522600.0 302850.0 522750.0 303750.0 ;
      RECT  522150.0 295050.0 523050.0 303300.0 ;
      RECT  519150.0 310950.0 520350.0 312150.0 ;
      RECT  522150.0 289050.0 523350.0 290250.0 ;
      RECT  519600.0 304350.0 520800.0 305550.0 ;
      RECT  522000.0 293850.0 523200.0 295050.0 ;
      RECT  525900.0 292050.0 527100.0 293250.0 ;
      RECT  519300.0 311550.0 520200.0 313350.0 ;
      RECT  522300.0 311550.0 523200.0 313350.0 ;
      RECT  519300.0 287850.0 520200.0 289650.0 ;
      RECT  522300.0 287850.0 523200.0 289650.0 ;
      RECT  515700.0 287850.0 516600.0 313350.0 ;
      RECT  525900.0 287850.0 526800.0 313350.0 ;
      RECT  204300.0 277350.0 203100.0 278550.0 ;
      RECT  206100.0 275250.0 204900.0 276450.0 ;
      RECT  214500.0 277350.0 213300.0 278550.0 ;
      RECT  216300.0 275250.0 215100.0 276450.0 ;
      RECT  224700.0 277350.0 223500.0 278550.0 ;
      RECT  226500.0 275250.0 225300.0 276450.0 ;
      RECT  234900.0 277350.0 233700.0 278550.0 ;
      RECT  236700.0 275250.0 235500.0 276450.0 ;
      RECT  245100.0 277350.0 243900.0 278550.0 ;
      RECT  246900.0 275250.0 245700.0 276450.0 ;
      RECT  255300.0 277350.0 254100.0 278550.0 ;
      RECT  257100.0 275250.0 255900.0 276450.0 ;
      RECT  265500.0 277350.0 264300.0 278550.0 ;
      RECT  267300.0 275250.0 266100.0 276450.0 ;
      RECT  275700.0 277350.0 274500.0 278550.0 ;
      RECT  277500.0 275250.0 276300.0 276450.0 ;
      RECT  285900.0 277350.0 284700.0 278550.0 ;
      RECT  287700.0 275250.0 286500.0 276450.0 ;
      RECT  296100.0 277350.0 294900.0 278550.0 ;
      RECT  297900.0 275250.0 296700.0 276450.0 ;
      RECT  306300.0 277350.0 305100.0 278550.0 ;
      RECT  308100.0 275250.0 306900.0 276450.0 ;
      RECT  316500.0 277350.0 315300.0 278550.0 ;
      RECT  318300.0 275250.0 317100.0 276450.0 ;
      RECT  326700.0 277350.0 325500.0 278550.0 ;
      RECT  328500.0 275250.0 327300.0 276450.0 ;
      RECT  336900.0 277350.0 335700.0 278550.0 ;
      RECT  338700.0 275250.0 337500.0 276450.0 ;
      RECT  347100.0 277350.0 345900.0 278550.0 ;
      RECT  348900.0 275250.0 347700.0 276450.0 ;
      RECT  357300.0 277350.0 356100.0 278550.0 ;
      RECT  359100.0 275250.0 357900.0 276450.0 ;
      RECT  367500.0 277350.0 366300.0 278550.0 ;
      RECT  369300.0 275250.0 368100.0 276450.0 ;
      RECT  377700.0 277350.0 376500.0 278550.0 ;
      RECT  379500.0 275250.0 378300.0 276450.0 ;
      RECT  387900.0 277350.0 386700.0 278550.0 ;
      RECT  389700.0 275250.0 388500.0 276450.0 ;
      RECT  398100.0 277350.0 396900.0 278550.0 ;
      RECT  399900.0 275250.0 398700.0 276450.0 ;
      RECT  408300.0 277350.0 407100.0 278550.0 ;
      RECT  410100.0 275250.0 408900.0 276450.0 ;
      RECT  418500.0 277350.0 417300.0 278550.0 ;
      RECT  420300.0 275250.0 419100.0 276450.0 ;
      RECT  428700.0 277350.0 427500.0 278550.0 ;
      RECT  430500.0 275250.0 429300.0 276450.0 ;
      RECT  438900.0 277350.0 437700.0 278550.0 ;
      RECT  440700.0 275250.0 439500.0 276450.0 ;
      RECT  449100.0 277350.0 447900.0 278550.0 ;
      RECT  450900.0 275250.0 449700.0 276450.0 ;
      RECT  459300.0 277350.0 458100.0 278550.0 ;
      RECT  461100.0 275250.0 459900.0 276450.0 ;
      RECT  469500.0 277350.0 468300.0 278550.0 ;
      RECT  471300.0 275250.0 470100.0 276450.0 ;
      RECT  479700.0 277350.0 478500.0 278550.0 ;
      RECT  481500.0 275250.0 480300.0 276450.0 ;
      RECT  489900.0 277350.0 488700.0 278550.0 ;
      RECT  491700.0 275250.0 490500.0 276450.0 ;
      RECT  500100.0 277350.0 498900.0 278550.0 ;
      RECT  501900.0 275250.0 500700.0 276450.0 ;
      RECT  510300.0 277350.0 509100.0 278550.0 ;
      RECT  512100.0 275250.0 510900.0 276450.0 ;
      RECT  520500.0 277350.0 519300.0 278550.0 ;
      RECT  522300.0 275250.0 521100.0 276450.0 ;
      RECT  203100.0 311550.0 204000.0 313350.0 ;
      RECT  206100.0 311550.0 207000.0 313350.0 ;
      RECT  213300.0 311550.0 214200.0 313350.0 ;
      RECT  216300.0 311550.0 217200.0 313350.0 ;
      RECT  223500.0 311550.0 224400.0 313350.0 ;
      RECT  226500.0 311550.0 227400.0 313350.0 ;
      RECT  233700.0 311550.0 234600.0 313350.0 ;
      RECT  236700.0 311550.0 237600.0 313350.0 ;
      RECT  243900.0 311550.0 244800.0 313350.0 ;
      RECT  246900.0 311550.0 247800.0 313350.0 ;
      RECT  254100.0 311550.0 255000.0 313350.0 ;
      RECT  257100.0 311550.0 258000.0 313350.0 ;
      RECT  264300.0 311550.0 265200.0 313350.0 ;
      RECT  267300.0 311550.0 268200.0 313350.0 ;
      RECT  274500.0 311550.0 275400.0 313350.0 ;
      RECT  277500.0 311550.0 278400.0 313350.0 ;
      RECT  284700.0 311550.0 285600.0 313350.0 ;
      RECT  287700.0 311550.0 288600.0 313350.0 ;
      RECT  294900.0 311550.0 295800.0 313350.0 ;
      RECT  297900.0 311550.0 298800.0 313350.0 ;
      RECT  305100.0 311550.0 306000.0 313350.0 ;
      RECT  308100.0 311550.0 309000.0 313350.0 ;
      RECT  315300.0 311550.0 316200.0 313350.0 ;
      RECT  318300.0 311550.0 319200.0 313350.0 ;
      RECT  325500.0 311550.0 326400.0 313350.0 ;
      RECT  328500.0 311550.0 329400.0 313350.0 ;
      RECT  335700.0 311550.0 336600.0 313350.0 ;
      RECT  338700.0 311550.0 339600.0 313350.0 ;
      RECT  345900.0 311550.0 346800.0 313350.0 ;
      RECT  348900.0 311550.0 349800.0 313350.0 ;
      RECT  356100.0 311550.0 357000.0 313350.0 ;
      RECT  359100.0 311550.0 360000.0 313350.0 ;
      RECT  366300.0 311550.0 367200.0 313350.0 ;
      RECT  369300.0 311550.0 370200.0 313350.0 ;
      RECT  376500.0 311550.0 377400.0 313350.0 ;
      RECT  379500.0 311550.0 380400.0 313350.0 ;
      RECT  386700.0 311550.0 387600.0 313350.0 ;
      RECT  389700.0 311550.0 390600.0 313350.0 ;
      RECT  396900.0 311550.0 397800.0 313350.0 ;
      RECT  399900.0 311550.0 400800.0 313350.0 ;
      RECT  407100.0 311550.0 408000.0 313350.0 ;
      RECT  410100.0 311550.0 411000.0 313350.0 ;
      RECT  417300.0 311550.0 418200.0 313350.0 ;
      RECT  420300.0 311550.0 421200.0 313350.0 ;
      RECT  427500.0 311550.0 428400.0 313350.0 ;
      RECT  430500.0 311550.0 431400.0 313350.0 ;
      RECT  437700.0 311550.0 438600.0 313350.0 ;
      RECT  440700.0 311550.0 441600.0 313350.0 ;
      RECT  447900.0 311550.0 448800.0 313350.0 ;
      RECT  450900.0 311550.0 451800.0 313350.0 ;
      RECT  458100.0 311550.0 459000.0 313350.0 ;
      RECT  461100.0 311550.0 462000.0 313350.0 ;
      RECT  468300.0 311550.0 469200.0 313350.0 ;
      RECT  471300.0 311550.0 472200.0 313350.0 ;
      RECT  478500.0 311550.0 479400.0 313350.0 ;
      RECT  481500.0 311550.0 482400.0 313350.0 ;
      RECT  488700.0 311550.0 489600.0 313350.0 ;
      RECT  491700.0 311550.0 492600.0 313350.0 ;
      RECT  498900.0 311550.0 499800.0 313350.0 ;
      RECT  501900.0 311550.0 502800.0 313350.0 ;
      RECT  509100.0 311550.0 510000.0 313350.0 ;
      RECT  512100.0 311550.0 513000.0 313350.0 ;
      RECT  519300.0 311550.0 520200.0 313350.0 ;
      RECT  522300.0 311550.0 523200.0 313350.0 ;
      RECT  203100.0 273150.0 204000.0 287850.0 ;
      RECT  206100.0 273150.0 207000.0 287850.0 ;
      RECT  243900.0 273150.0 244800.0 287850.0 ;
      RECT  246900.0 273150.0 247800.0 287850.0 ;
      RECT  284700.0 273150.0 285600.0 287850.0 ;
      RECT  287700.0 273150.0 288600.0 287850.0 ;
      RECT  325500.0 273150.0 326400.0 287850.0 ;
      RECT  328500.0 273150.0 329400.0 287850.0 ;
      RECT  366300.0 273150.0 367200.0 287850.0 ;
      RECT  369300.0 273150.0 370200.0 287850.0 ;
      RECT  407100.0 273150.0 408000.0 287850.0 ;
      RECT  410100.0 273150.0 411000.0 287850.0 ;
      RECT  447900.0 273150.0 448800.0 287850.0 ;
      RECT  450900.0 273150.0 451800.0 287850.0 ;
      RECT  488700.0 273150.0 489600.0 287850.0 ;
      RECT  491700.0 273150.0 492600.0 287850.0 ;
      RECT  199500.0 273150.0 200400.0 313350.0 ;
      RECT  209700.0 273150.0 210600.0 313350.0 ;
      RECT  219900.0 273150.0 220800.0 313350.0 ;
      RECT  230100.0 273150.0 231000.0 313350.0 ;
      RECT  240300.0 273150.0 241200.0 313350.0 ;
      RECT  250500.0 273150.0 251400.0 313350.0 ;
      RECT  260700.0 273150.0 261600.0 313350.0 ;
      RECT  270900.0 273150.0 271800.0 313350.0 ;
      RECT  281100.0 273150.0 282000.0 313350.0 ;
      RECT  291300.0 273150.0 292200.0 313350.0 ;
      RECT  301500.0 273150.0 302400.0 313350.0 ;
      RECT  311700.0 273150.0 312600.0 313350.0 ;
      RECT  321900.0 273150.0 322800.0 313350.0 ;
      RECT  332100.0 273150.0 333000.0 313350.0 ;
      RECT  342300.0 273150.0 343200.0 313350.0 ;
      RECT  352500.0 273150.0 353400.0 313350.0 ;
      RECT  362700.0 273150.0 363600.0 313350.0 ;
      RECT  372900.0 273150.0 373800.0 313350.0 ;
      RECT  383100.0 273150.0 384000.0 313350.0 ;
      RECT  393300.0 273150.0 394200.0 313350.0 ;
      RECT  403500.0 273150.0 404400.0 313350.0 ;
      RECT  413700.0 273150.0 414600.0 313350.0 ;
      RECT  423900.0 273150.0 424800.0 313350.0 ;
      RECT  434100.0 273150.0 435000.0 313350.0 ;
      RECT  444300.0 273150.0 445200.0 313350.0 ;
      RECT  454500.0 273150.0 455400.0 313350.0 ;
      RECT  464700.0 273150.0 465600.0 313350.0 ;
      RECT  474900.0 273150.0 475800.0 313350.0 ;
      RECT  485100.0 273150.0 486000.0 313350.0 ;
      RECT  495300.0 273150.0 496200.0 313350.0 ;
      RECT  505500.0 273150.0 506400.0 313350.0 ;
      RECT  515700.0 273150.0 516600.0 313350.0 ;
      RECT  103500.0 600.0 104400.0 54000.0 ;
      RECT  106500.0 600.0 107400.0 54000.0 ;
      RECT  97500.0 600.0 98400.0 54000.0 ;
      RECT  100500.0 600.0 101400.0 54000.0 ;
      RECT  113850.0 7950.0 114750.0 8850.0 ;
      RECT  116250.0 7950.0 117150.0 8850.0 ;
      RECT  113850.0 8400.0 114750.0 11250.0 ;
      RECT  114300.0 7950.0 116700.0 8850.0 ;
      RECT  116250.0 3750.0 117150.0 8400.0 ;
      RECT  113700.0 11250.0 114900.0 12450.0 ;
      RECT  116100.0 2550.0 117300.0 3750.0 ;
      RECT  117300.0 7800.0 116100.0 9000.0 ;
      RECT  113850.0 20850.0 114750.0 19950.0 ;
      RECT  116250.0 20850.0 117150.0 19950.0 ;
      RECT  113850.0 20400.0 114750.0 17550.0 ;
      RECT  114300.0 20850.0 116700.0 19950.0 ;
      RECT  116250.0 25050.0 117150.0 20400.0 ;
      RECT  113700.0 17550.0 114900.0 16350.0 ;
      RECT  116100.0 26250.0 117300.0 25050.0 ;
      RECT  117300.0 21000.0 116100.0 19800.0 ;
      RECT  113850.0 35550.0 114750.0 36450.0 ;
      RECT  116250.0 35550.0 117150.0 36450.0 ;
      RECT  113850.0 36000.0 114750.0 38850.0 ;
      RECT  114300.0 35550.0 116700.0 36450.0 ;
      RECT  116250.0 31350.0 117150.0 36000.0 ;
      RECT  113700.0 38850.0 114900.0 40050.0 ;
      RECT  116100.0 30150.0 117300.0 31350.0 ;
      RECT  117300.0 35400.0 116100.0 36600.0 ;
      RECT  113850.0 48450.0 114750.0 47550.0 ;
      RECT  116250.0 48450.0 117150.0 47550.0 ;
      RECT  113850.0 48000.0 114750.0 45150.0 ;
      RECT  114300.0 48450.0 116700.0 47550.0 ;
      RECT  116250.0 52650.0 117150.0 48000.0 ;
      RECT  113700.0 45150.0 114900.0 43950.0 ;
      RECT  116100.0 53850.0 117300.0 52650.0 ;
      RECT  117300.0 48600.0 116100.0 47400.0 ;
      RECT  98550.0 11100.0 97350.0 12300.0 ;
      RECT  79950.0 6600.0 78750.0 7800.0 ;
      RECT  101550.0 24900.0 100350.0 26100.0 ;
      RECT  82950.0 21000.0 81750.0 22200.0 ;
      RECT  79950.0 29700.0 78750.0 30900.0 ;
      RECT  104550.0 29700.0 103350.0 30900.0 ;
      RECT  82950.0 43500.0 81750.0 44700.0 ;
      RECT  107550.0 43500.0 106350.0 44700.0 ;
      RECT  98550.0 7800.0 97350.0 9000.0 ;
      RECT  101550.0 5100.0 100350.0 6300.0 ;
      RECT  104550.0 19800.0 103350.0 21000.0 ;
      RECT  101550.0 22500.0 100350.0 23700.0 ;
      RECT  98550.0 35400.0 97350.0 36600.0 ;
      RECT  107550.0 32700.0 106350.0 33900.0 ;
      RECT  104550.0 47400.0 103350.0 48600.0 ;
      RECT  107550.0 50100.0 106350.0 51300.0 ;
      RECT  78900.0 600.0 79800.0 54000.0 ;
      RECT  81900.0 600.0 82800.0 54000.0 ;
      RECT  200100.0 224250.0 210300.0 273150.0 ;
      RECT  240900.0 224250.0 251100.0 273150.0 ;
      RECT  281700.0 224250.0 291900.0 273150.0 ;
      RECT  322500.0 224250.0 332700.0 273150.0 ;
      RECT  363300.0 224250.0 373500.0 273150.0 ;
      RECT  404100.0 224250.0 414300.0 273150.0 ;
      RECT  444900.0 224250.0 455100.0 273150.0 ;
      RECT  485700.0 224250.0 495900.0 273150.0 ;
      RECT  203100.0 224250.0 204300.0 237450.0 ;
      RECT  206100.0 224250.0 207300.0 237450.0 ;
      RECT  243900.0 224250.0 245100.0 237450.0 ;
      RECT  246900.0 224250.0 248100.0 237450.0 ;
      RECT  284700.0 224250.0 285900.0 237450.0 ;
      RECT  287700.0 224250.0 288900.0 237450.0 ;
      RECT  325500.0 224250.0 326700.0 237450.0 ;
      RECT  328500.0 224250.0 329700.0 237450.0 ;
      RECT  366300.0 224250.0 367500.0 237450.0 ;
      RECT  369300.0 224250.0 370500.0 237450.0 ;
      RECT  407100.0 224250.0 408300.0 237450.0 ;
      RECT  410100.0 224250.0 411300.0 237450.0 ;
      RECT  447900.0 224250.0 449100.0 237450.0 ;
      RECT  450900.0 224250.0 452100.0 237450.0 ;
      RECT  488700.0 224250.0 489900.0 237450.0 ;
      RECT  491700.0 224250.0 492900.0 237450.0 ;
      RECT  200100.0 163650.0 210300.0 224250.0 ;
      RECT  240900.0 163650.0 251100.0 224250.0 ;
      RECT  281700.0 163650.0 291900.0 224250.0 ;
      RECT  322500.0 163650.0 332700.0 224250.0 ;
      RECT  363300.0 163650.0 373500.0 224250.0 ;
      RECT  404100.0 163650.0 414300.0 224250.0 ;
      RECT  444900.0 163650.0 455100.0 224250.0 ;
      RECT  485700.0 163650.0 495900.0 224250.0 ;
      RECT  204600.0 163650.0 205800.0 166650.0 ;
      RECT  245400.0 163650.0 246600.0 166650.0 ;
      RECT  286200.0 163650.0 287400.0 166650.0 ;
      RECT  327000.0 163650.0 328200.0 166650.0 ;
      RECT  367800.0 163650.0 369000.0 166650.0 ;
      RECT  408600.0 163650.0 409800.0 166650.0 ;
      RECT  449400.0 163650.0 450600.0 166650.0 ;
      RECT  490200.0 163650.0 491400.0 166650.0 ;
      RECT  203100.0 222150.0 204300.0 224250.0 ;
      RECT  206100.0 216750.0 207300.0 224250.0 ;
      RECT  243900.0 222150.0 245100.0 224250.0 ;
      RECT  246900.0 216750.0 248100.0 224250.0 ;
      RECT  284700.0 222150.0 285900.0 224250.0 ;
      RECT  287700.0 216750.0 288900.0 224250.0 ;
      RECT  325500.0 222150.0 326700.0 224250.0 ;
      RECT  328500.0 216750.0 329700.0 224250.0 ;
      RECT  366300.0 222150.0 367500.0 224250.0 ;
      RECT  369300.0 216750.0 370500.0 224250.0 ;
      RECT  407100.0 222150.0 408300.0 224250.0 ;
      RECT  410100.0 216750.0 411300.0 224250.0 ;
      RECT  447900.0 222150.0 449100.0 224250.0 ;
      RECT  450900.0 216750.0 452100.0 224250.0 ;
      RECT  488700.0 222150.0 489900.0 224250.0 ;
      RECT  491700.0 216750.0 492900.0 224250.0 ;
      RECT  200100.0 103650.0 210300.0 163650.0 ;
      RECT  240900.0 103650.0 251100.0 163650.0 ;
      RECT  281700.0 103650.0 291900.0 163650.0 ;
      RECT  322500.0 103650.0 332700.0 163650.0 ;
      RECT  363300.0 103650.0 373500.0 163650.0 ;
      RECT  404100.0 103650.0 414300.0 163650.0 ;
      RECT  444900.0 103650.0 455100.0 163650.0 ;
      RECT  485700.0 103650.0 495900.0 163650.0 ;
      RECT  204600.0 161250.0 207300.0 162450.0 ;
      RECT  201900.0 159150.0 203100.0 163650.0 ;
      RECT  245400.0 161250.0 248100.0 162450.0 ;
      RECT  242700.0 159150.0 243900.0 163650.0 ;
      RECT  286200.0 161250.0 288900.0 162450.0 ;
      RECT  283500.0 159150.0 284700.0 163650.0 ;
      RECT  327000.0 161250.0 329700.0 162450.0 ;
      RECT  324300.0 159150.0 325500.0 163650.0 ;
      RECT  367800.0 161250.0 370500.0 162450.0 ;
      RECT  365100.0 159150.0 366300.0 163650.0 ;
      RECT  408600.0 161250.0 411300.0 162450.0 ;
      RECT  405900.0 159150.0 407100.0 163650.0 ;
      RECT  449400.0 161250.0 452100.0 162450.0 ;
      RECT  446700.0 159150.0 447900.0 163650.0 ;
      RECT  490200.0 161250.0 492900.0 162450.0 ;
      RECT  487500.0 159150.0 488700.0 163650.0 ;
      RECT  209700.0 103650.0 210900.0 163650.0 ;
      RECT  250500.0 103650.0 251700.0 163650.0 ;
      RECT  291300.0 103650.0 292500.0 163650.0 ;
      RECT  332100.0 103650.0 333300.0 163650.0 ;
      RECT  372900.0 103650.0 374100.0 163650.0 ;
      RECT  413700.0 103650.0 414900.0 163650.0 ;
      RECT  454500.0 103650.0 455700.0 163650.0 ;
      RECT  495300.0 103650.0 496500.0 163650.0 ;
      RECT  200100.0 103650.0 210300.0 81750.0 ;
      RECT  240900.0 103650.0 251100.0 81750.0 ;
      RECT  281700.0 103650.0 291900.0 81750.0 ;
      RECT  322500.0 103650.0 332700.0 81750.0 ;
      RECT  363300.0 103650.0 373500.0 81750.0 ;
      RECT  404100.0 103650.0 414300.0 81750.0 ;
      RECT  444900.0 103650.0 455100.0 81750.0 ;
      RECT  485700.0 103650.0 495900.0 81750.0 ;
      RECT  204600.0 88650.0 205800.0 81750.0 ;
      RECT  245400.0 88650.0 246600.0 81750.0 ;
      RECT  286200.0 88650.0 287400.0 81750.0 ;
      RECT  327000.0 88650.0 328200.0 81750.0 ;
      RECT  367800.0 88650.0 369000.0 81750.0 ;
      RECT  408600.0 88650.0 409800.0 81750.0 ;
      RECT  449400.0 88650.0 450600.0 81750.0 ;
      RECT  490200.0 88650.0 491400.0 81750.0 ;
      RECT  204600.0 103650.0 205800.0 102150.0 ;
      RECT  245400.0 103650.0 246600.0 102150.0 ;
      RECT  286200.0 103650.0 287400.0 102150.0 ;
      RECT  327000.0 103650.0 328200.0 102150.0 ;
      RECT  367800.0 103650.0 369000.0 102150.0 ;
      RECT  408600.0 103650.0 409800.0 102150.0 ;
      RECT  449400.0 103650.0 450600.0 102150.0 ;
      RECT  490200.0 103650.0 491400.0 102150.0 ;
      RECT  59100.0 148200.0 60000.0 1197000.0 ;
      RECT  61200.0 148200.0 62100.0 1197000.0 ;
      RECT  63300.0 148200.0 64200.0 1197000.0 ;
      RECT  65400.0 148200.0 66300.0 1197000.0 ;
      RECT  67500.0 148200.0 68400.0 1197000.0 ;
      RECT  69600.0 148200.0 70500.0 1197000.0 ;
      RECT  71700.0 148200.0 72600.0 1197000.0 ;
      RECT  73800.0 148200.0 74700.0 1197000.0 ;
      RECT  75900.0 148200.0 76800.0 1197000.0 ;
      RECT  78000.0 148200.0 78900.0 1197000.0 ;
      RECT  80100.0 148200.0 81000.0 1197000.0 ;
      RECT  82200.0 148200.0 83100.0 1197000.0 ;
      RECT  114300.0 148200.0 113400.0 201600.0 ;
      RECT  111300.0 148200.0 110400.0 201600.0 ;
      RECT  120300.0 148200.0 119400.0 201600.0 ;
      RECT  117300.0 148200.0 116400.0 201600.0 ;
      RECT  103950.0 155550.0 103050.0 156450.0 ;
      RECT  101550.0 155550.0 100650.0 156450.0 ;
      RECT  103950.0 156000.0 103050.0 158850.0 ;
      RECT  103500.0 155550.0 101100.0 156450.0 ;
      RECT  101550.0 151350.0 100650.0 156000.0 ;
      RECT  104100.0 158850.0 102900.0 160050.0 ;
      RECT  101700.0 150150.0 100500.0 151350.0 ;
      RECT  100500.0 155400.0 101700.0 156600.0 ;
      RECT  103950.0 168450.0 103050.0 167550.0 ;
      RECT  101550.0 168450.0 100650.0 167550.0 ;
      RECT  103950.0 168000.0 103050.0 165150.0 ;
      RECT  103500.0 168450.0 101100.0 167550.0 ;
      RECT  101550.0 172650.0 100650.0 168000.0 ;
      RECT  104100.0 165150.0 102900.0 163950.0 ;
      RECT  101700.0 173850.0 100500.0 172650.0 ;
      RECT  100500.0 168600.0 101700.0 167400.0 ;
      RECT  103950.0 183150.0 103050.0 184050.0 ;
      RECT  101550.0 183150.0 100650.0 184050.0 ;
      RECT  103950.0 183600.0 103050.0 186450.0 ;
      RECT  103500.0 183150.0 101100.0 184050.0 ;
      RECT  101550.0 178950.0 100650.0 183600.0 ;
      RECT  104100.0 186450.0 102900.0 187650.0 ;
      RECT  101700.0 177750.0 100500.0 178950.0 ;
      RECT  100500.0 183000.0 101700.0 184200.0 ;
      RECT  103950.0 196050.0 103050.0 195150.0 ;
      RECT  101550.0 196050.0 100650.0 195150.0 ;
      RECT  103950.0 195600.0 103050.0 192750.0 ;
      RECT  103500.0 196050.0 101100.0 195150.0 ;
      RECT  101550.0 200250.0 100650.0 195600.0 ;
      RECT  104100.0 192750.0 102900.0 191550.0 ;
      RECT  101700.0 201450.0 100500.0 200250.0 ;
      RECT  100500.0 196200.0 101700.0 195000.0 ;
      RECT  119250.0 158700.0 120450.0 159900.0 ;
      RECT  137850.0 154200.0 139050.0 155400.0 ;
      RECT  116250.0 172500.0 117450.0 173700.0 ;
      RECT  134850.0 168600.0 136050.0 169800.0 ;
      RECT  137850.0 177300.0 139050.0 178500.0 ;
      RECT  113250.0 177300.0 114450.0 178500.0 ;
      RECT  134850.0 191100.0 136050.0 192300.0 ;
      RECT  110250.0 191100.0 111450.0 192300.0 ;
      RECT  119250.0 155400.0 120450.0 156600.0 ;
      RECT  116250.0 152700.0 117450.0 153900.0 ;
      RECT  113250.0 167400.0 114450.0 168600.0 ;
      RECT  116250.0 170100.0 117450.0 171300.0 ;
      RECT  119250.0 183000.0 120450.0 184200.0 ;
      RECT  110250.0 180300.0 111450.0 181500.0 ;
      RECT  113250.0 195000.0 114450.0 196200.0 ;
      RECT  110250.0 197700.0 111450.0 198900.0 ;
      RECT  138900.0 148200.0 138000.0 201600.0 ;
      RECT  135900.0 148200.0 135000.0 201600.0 ;
      RECT  114300.0 203400.0 113400.0 256800.0 ;
      RECT  111300.0 203400.0 110400.0 256800.0 ;
      RECT  120300.0 203400.0 119400.0 256800.0 ;
      RECT  117300.0 203400.0 116400.0 256800.0 ;
      RECT  103950.0 210750.0 103050.0 211650.0 ;
      RECT  101550.0 210750.0 100650.0 211650.0 ;
      RECT  103950.0 211200.0 103050.0 214050.0 ;
      RECT  103500.0 210750.0 101100.0 211650.0 ;
      RECT  101550.0 206550.0 100650.0 211200.0 ;
      RECT  104100.0 214050.0 102900.0 215250.0 ;
      RECT  101700.0 205350.0 100500.0 206550.0 ;
      RECT  100500.0 210600.0 101700.0 211800.0 ;
      RECT  103950.0 223650.0 103050.0 222750.0 ;
      RECT  101550.0 223650.0 100650.0 222750.0 ;
      RECT  103950.0 223200.0 103050.0 220350.0 ;
      RECT  103500.0 223650.0 101100.0 222750.0 ;
      RECT  101550.0 227850.0 100650.0 223200.0 ;
      RECT  104100.0 220350.0 102900.0 219150.0 ;
      RECT  101700.0 229050.0 100500.0 227850.0 ;
      RECT  100500.0 223800.0 101700.0 222600.0 ;
      RECT  103950.0 238350.0 103050.0 239250.0 ;
      RECT  101550.0 238350.0 100650.0 239250.0 ;
      RECT  103950.0 238800.0 103050.0 241650.0 ;
      RECT  103500.0 238350.0 101100.0 239250.0 ;
      RECT  101550.0 234150.0 100650.0 238800.0 ;
      RECT  104100.0 241650.0 102900.0 242850.0 ;
      RECT  101700.0 232950.0 100500.0 234150.0 ;
      RECT  100500.0 238200.0 101700.0 239400.0 ;
      RECT  103950.0 251250.0 103050.0 250350.0 ;
      RECT  101550.0 251250.0 100650.0 250350.0 ;
      RECT  103950.0 250800.0 103050.0 247950.0 ;
      RECT  103500.0 251250.0 101100.0 250350.0 ;
      RECT  101550.0 255450.0 100650.0 250800.0 ;
      RECT  104100.0 247950.0 102900.0 246750.0 ;
      RECT  101700.0 256650.0 100500.0 255450.0 ;
      RECT  100500.0 251400.0 101700.0 250200.0 ;
      RECT  119250.0 213900.0 120450.0 215100.0 ;
      RECT  137850.0 209400.0 139050.0 210600.0 ;
      RECT  116250.0 227700.0 117450.0 228900.0 ;
      RECT  134850.0 223800.0 136050.0 225000.0 ;
      RECT  137850.0 232500.0 139050.0 233700.0 ;
      RECT  113250.0 232500.0 114450.0 233700.0 ;
      RECT  134850.0 246300.0 136050.0 247500.0 ;
      RECT  110250.0 246300.0 111450.0 247500.0 ;
      RECT  119250.0 210600.0 120450.0 211800.0 ;
      RECT  116250.0 207900.0 117450.0 209100.0 ;
      RECT  113250.0 222600.0 114450.0 223800.0 ;
      RECT  116250.0 225300.0 117450.0 226500.0 ;
      RECT  119250.0 238200.0 120450.0 239400.0 ;
      RECT  110250.0 235500.0 111450.0 236700.0 ;
      RECT  113250.0 250200.0 114450.0 251400.0 ;
      RECT  110250.0 252900.0 111450.0 254100.0 ;
      RECT  138900.0 203400.0 138000.0 256800.0 ;
      RECT  135900.0 203400.0 135000.0 256800.0 ;
      RECT  114300.0 258600.0 113400.0 312000.0 ;
      RECT  111300.0 258600.0 110400.0 312000.0 ;
      RECT  120300.0 258600.0 119400.0 312000.0 ;
      RECT  117300.0 258600.0 116400.0 312000.0 ;
      RECT  103950.0 265950.0 103050.0 266850.0 ;
      RECT  101550.0 265950.0 100650.0 266850.0 ;
      RECT  103950.0 266400.0 103050.0 269250.0 ;
      RECT  103500.0 265950.0 101100.0 266850.0 ;
      RECT  101550.0 261750.0 100650.0 266400.0 ;
      RECT  104100.0 269250.0 102900.0 270450.0 ;
      RECT  101700.0 260550.0 100500.0 261750.0 ;
      RECT  100500.0 265800.0 101700.0 267000.0 ;
      RECT  103950.0 278850.0 103050.0 277950.0 ;
      RECT  101550.0 278850.0 100650.0 277950.0 ;
      RECT  103950.0 278400.0 103050.0 275550.0 ;
      RECT  103500.0 278850.0 101100.0 277950.0 ;
      RECT  101550.0 283050.0 100650.0 278400.0 ;
      RECT  104100.0 275550.0 102900.0 274350.0 ;
      RECT  101700.0 284250.0 100500.0 283050.0 ;
      RECT  100500.0 279000.0 101700.0 277800.0 ;
      RECT  103950.0 293550.0 103050.0 294450.0 ;
      RECT  101550.0 293550.0 100650.0 294450.0 ;
      RECT  103950.0 294000.0 103050.0 296850.0 ;
      RECT  103500.0 293550.0 101100.0 294450.0 ;
      RECT  101550.0 289350.0 100650.0 294000.0 ;
      RECT  104100.0 296850.0 102900.0 298050.0 ;
      RECT  101700.0 288150.0 100500.0 289350.0 ;
      RECT  100500.0 293400.0 101700.0 294600.0 ;
      RECT  103950.0 306450.0 103050.0 305550.0 ;
      RECT  101550.0 306450.0 100650.0 305550.0 ;
      RECT  103950.0 306000.0 103050.0 303150.0 ;
      RECT  103500.0 306450.0 101100.0 305550.0 ;
      RECT  101550.0 310650.0 100650.0 306000.0 ;
      RECT  104100.0 303150.0 102900.0 301950.0 ;
      RECT  101700.0 311850.0 100500.0 310650.0 ;
      RECT  100500.0 306600.0 101700.0 305400.0 ;
      RECT  119250.0 269100.0 120450.0 270300.0 ;
      RECT  137850.0 264600.0 139050.0 265800.0 ;
      RECT  116250.0 282900.0 117450.0 284100.0 ;
      RECT  134850.0 279000.0 136050.0 280200.0 ;
      RECT  137850.0 287700.0 139050.0 288900.0 ;
      RECT  113250.0 287700.0 114450.0 288900.0 ;
      RECT  134850.0 301500.0 136050.0 302700.0 ;
      RECT  110250.0 301500.0 111450.0 302700.0 ;
      RECT  119250.0 265800.0 120450.0 267000.0 ;
      RECT  116250.0 263100.0 117450.0 264300.0 ;
      RECT  113250.0 277800.0 114450.0 279000.0 ;
      RECT  116250.0 280500.0 117450.0 281700.0 ;
      RECT  119250.0 293400.0 120450.0 294600.0 ;
      RECT  110250.0 290700.0 111450.0 291900.0 ;
      RECT  113250.0 305400.0 114450.0 306600.0 ;
      RECT  110250.0 308100.0 111450.0 309300.0 ;
      RECT  138900.0 258600.0 138000.0 312000.0 ;
      RECT  135900.0 258600.0 135000.0 312000.0 ;
      RECT  93450.0 316950.0 94350.0 324450.0 ;
      RECT  88650.0 321900.0 89550.0 322800.0 ;
      RECT  93450.0 321900.0 94350.0 322800.0 ;
      RECT  88650.0 322350.0 89550.0 324450.0 ;
      RECT  89100.0 321900.0 93900.0 322800.0 ;
      RECT  93450.0 316950.0 94350.0 322350.0 ;
      RECT  88500.0 324450.0 89700.0 325650.0 ;
      RECT  93300.0 324450.0 94500.0 325650.0 ;
      RECT  93300.0 315750.0 94500.0 316950.0 ;
      RECT  93300.0 321750.0 94500.0 322950.0 ;
      RECT  93450.0 338250.0 94350.0 330750.0 ;
      RECT  88650.0 333300.0 89550.0 332400.0 ;
      RECT  93450.0 333300.0 94350.0 332400.0 ;
      RECT  88650.0 332850.0 89550.0 330750.0 ;
      RECT  89100.0 333300.0 93900.0 332400.0 ;
      RECT  93450.0 338250.0 94350.0 332850.0 ;
      RECT  88500.0 330750.0 89700.0 329550.0 ;
      RECT  93300.0 330750.0 94500.0 329550.0 ;
      RECT  93300.0 339450.0 94500.0 338250.0 ;
      RECT  93300.0 333450.0 94500.0 332250.0 ;
      RECT  93450.0 344550.0 94350.0 352050.0 ;
      RECT  88650.0 349500.0 89550.0 350400.0 ;
      RECT  93450.0 349500.0 94350.0 350400.0 ;
      RECT  88650.0 349950.0 89550.0 352050.0 ;
      RECT  89100.0 349500.0 93900.0 350400.0 ;
      RECT  93450.0 344550.0 94350.0 349950.0 ;
      RECT  88500.0 352050.0 89700.0 353250.0 ;
      RECT  93300.0 352050.0 94500.0 353250.0 ;
      RECT  93300.0 343350.0 94500.0 344550.0 ;
      RECT  93300.0 349350.0 94500.0 350550.0 ;
      RECT  93450.0 365850.0 94350.0 358350.0 ;
      RECT  88650.0 360900.0 89550.0 360000.0 ;
      RECT  93450.0 360900.0 94350.0 360000.0 ;
      RECT  88650.0 360450.0 89550.0 358350.0 ;
      RECT  89100.0 360900.0 93900.0 360000.0 ;
      RECT  93450.0 365850.0 94350.0 360450.0 ;
      RECT  88500.0 358350.0 89700.0 357150.0 ;
      RECT  93300.0 358350.0 94500.0 357150.0 ;
      RECT  93300.0 367050.0 94500.0 365850.0 ;
      RECT  93300.0 361050.0 94500.0 359850.0 ;
      RECT  93450.0 372150.0 94350.0 379650.0 ;
      RECT  88650.0 377100.0 89550.0 378000.0 ;
      RECT  93450.0 377100.0 94350.0 378000.0 ;
      RECT  88650.0 377550.0 89550.0 379650.0 ;
      RECT  89100.0 377100.0 93900.0 378000.0 ;
      RECT  93450.0 372150.0 94350.0 377550.0 ;
      RECT  88500.0 379650.0 89700.0 380850.0 ;
      RECT  93300.0 379650.0 94500.0 380850.0 ;
      RECT  93300.0 370950.0 94500.0 372150.0 ;
      RECT  93300.0 376950.0 94500.0 378150.0 ;
      RECT  93450.0 393450.0 94350.0 385950.0 ;
      RECT  88650.0 388500.0 89550.0 387600.0 ;
      RECT  93450.0 388500.0 94350.0 387600.0 ;
      RECT  88650.0 388050.0 89550.0 385950.0 ;
      RECT  89100.0 388500.0 93900.0 387600.0 ;
      RECT  93450.0 393450.0 94350.0 388050.0 ;
      RECT  88500.0 385950.0 89700.0 384750.0 ;
      RECT  93300.0 385950.0 94500.0 384750.0 ;
      RECT  93300.0 394650.0 94500.0 393450.0 ;
      RECT  93300.0 388650.0 94500.0 387450.0 ;
      RECT  93450.0 399750.0 94350.0 407250.0 ;
      RECT  88650.0 404700.0 89550.0 405600.0 ;
      RECT  93450.0 404700.0 94350.0 405600.0 ;
      RECT  88650.0 405150.0 89550.0 407250.0 ;
      RECT  89100.0 404700.0 93900.0 405600.0 ;
      RECT  93450.0 399750.0 94350.0 405150.0 ;
      RECT  88500.0 407250.0 89700.0 408450.0 ;
      RECT  93300.0 407250.0 94500.0 408450.0 ;
      RECT  93300.0 398550.0 94500.0 399750.0 ;
      RECT  93300.0 404550.0 94500.0 405750.0 ;
      RECT  93450.0 421050.0 94350.0 413550.0 ;
      RECT  88650.0 416100.0 89550.0 415200.0 ;
      RECT  93450.0 416100.0 94350.0 415200.0 ;
      RECT  88650.0 415650.0 89550.0 413550.0 ;
      RECT  89100.0 416100.0 93900.0 415200.0 ;
      RECT  93450.0 421050.0 94350.0 415650.0 ;
      RECT  88500.0 413550.0 89700.0 412350.0 ;
      RECT  93300.0 413550.0 94500.0 412350.0 ;
      RECT  93300.0 422250.0 94500.0 421050.0 ;
      RECT  93300.0 416250.0 94500.0 415050.0 ;
      RECT  93450.0 427350.0 94350.0 434850.0 ;
      RECT  88650.0 432300.0 89550.0 433200.0 ;
      RECT  93450.0 432300.0 94350.0 433200.0 ;
      RECT  88650.0 432750.0 89550.0 434850.0 ;
      RECT  89100.0 432300.0 93900.0 433200.0 ;
      RECT  93450.0 427350.0 94350.0 432750.0 ;
      RECT  88500.0 434850.0 89700.0 436050.0 ;
      RECT  93300.0 434850.0 94500.0 436050.0 ;
      RECT  93300.0 426150.0 94500.0 427350.0 ;
      RECT  93300.0 432150.0 94500.0 433350.0 ;
      RECT  93450.0 448650.0 94350.0 441150.0 ;
      RECT  88650.0 443700.0 89550.0 442800.0 ;
      RECT  93450.0 443700.0 94350.0 442800.0 ;
      RECT  88650.0 443250.0 89550.0 441150.0 ;
      RECT  89100.0 443700.0 93900.0 442800.0 ;
      RECT  93450.0 448650.0 94350.0 443250.0 ;
      RECT  88500.0 441150.0 89700.0 439950.0 ;
      RECT  93300.0 441150.0 94500.0 439950.0 ;
      RECT  93300.0 449850.0 94500.0 448650.0 ;
      RECT  93300.0 443850.0 94500.0 442650.0 ;
      RECT  93450.0 454950.0 94350.0 462450.0 ;
      RECT  88650.0 459900.0 89550.0 460800.0 ;
      RECT  93450.0 459900.0 94350.0 460800.0 ;
      RECT  88650.0 460350.0 89550.0 462450.0 ;
      RECT  89100.0 459900.0 93900.0 460800.0 ;
      RECT  93450.0 454950.0 94350.0 460350.0 ;
      RECT  88500.0 462450.0 89700.0 463650.0 ;
      RECT  93300.0 462450.0 94500.0 463650.0 ;
      RECT  93300.0 453750.0 94500.0 454950.0 ;
      RECT  93300.0 459750.0 94500.0 460950.0 ;
      RECT  93450.0 476250.0 94350.0 468750.0 ;
      RECT  88650.0 471300.0 89550.0 470400.0 ;
      RECT  93450.0 471300.0 94350.0 470400.0 ;
      RECT  88650.0 470850.0 89550.0 468750.0 ;
      RECT  89100.0 471300.0 93900.0 470400.0 ;
      RECT  93450.0 476250.0 94350.0 470850.0 ;
      RECT  88500.0 468750.0 89700.0 467550.0 ;
      RECT  93300.0 468750.0 94500.0 467550.0 ;
      RECT  93300.0 477450.0 94500.0 476250.0 ;
      RECT  93300.0 471450.0 94500.0 470250.0 ;
      RECT  93450.0 482550.0 94350.0 490050.0 ;
      RECT  88650.0 487500.0 89550.0 488400.0 ;
      RECT  93450.0 487500.0 94350.0 488400.0 ;
      RECT  88650.0 487950.0 89550.0 490050.0 ;
      RECT  89100.0 487500.0 93900.0 488400.0 ;
      RECT  93450.0 482550.0 94350.0 487950.0 ;
      RECT  88500.0 490050.0 89700.0 491250.0 ;
      RECT  93300.0 490050.0 94500.0 491250.0 ;
      RECT  93300.0 481350.0 94500.0 482550.0 ;
      RECT  93300.0 487350.0 94500.0 488550.0 ;
      RECT  93450.0 503850.0 94350.0 496350.0 ;
      RECT  88650.0 498900.0 89550.0 498000.0 ;
      RECT  93450.0 498900.0 94350.0 498000.0 ;
      RECT  88650.0 498450.0 89550.0 496350.0 ;
      RECT  89100.0 498900.0 93900.0 498000.0 ;
      RECT  93450.0 503850.0 94350.0 498450.0 ;
      RECT  88500.0 496350.0 89700.0 495150.0 ;
      RECT  93300.0 496350.0 94500.0 495150.0 ;
      RECT  93300.0 505050.0 94500.0 503850.0 ;
      RECT  93300.0 499050.0 94500.0 497850.0 ;
      RECT  93450.0 510150.0 94350.0 517650.0 ;
      RECT  88650.0 515100.0 89550.0 516000.0 ;
      RECT  93450.0 515100.0 94350.0 516000.0 ;
      RECT  88650.0 515550.0 89550.0 517650.0 ;
      RECT  89100.0 515100.0 93900.0 516000.0 ;
      RECT  93450.0 510150.0 94350.0 515550.0 ;
      RECT  88500.0 517650.0 89700.0 518850.0 ;
      RECT  93300.0 517650.0 94500.0 518850.0 ;
      RECT  93300.0 508950.0 94500.0 510150.0 ;
      RECT  93300.0 514950.0 94500.0 516150.0 ;
      RECT  93450.0 531450.0 94350.0 523950.0 ;
      RECT  88650.0 526500.0 89550.0 525600.0 ;
      RECT  93450.0 526500.0 94350.0 525600.0 ;
      RECT  88650.0 526050.0 89550.0 523950.0 ;
      RECT  89100.0 526500.0 93900.0 525600.0 ;
      RECT  93450.0 531450.0 94350.0 526050.0 ;
      RECT  88500.0 523950.0 89700.0 522750.0 ;
      RECT  93300.0 523950.0 94500.0 522750.0 ;
      RECT  93300.0 532650.0 94500.0 531450.0 ;
      RECT  93300.0 526650.0 94500.0 525450.0 ;
      RECT  93450.0 537750.0 94350.0 545250.0 ;
      RECT  88650.0 542700.0 89550.0 543600.0 ;
      RECT  93450.0 542700.0 94350.0 543600.0 ;
      RECT  88650.0 543150.0 89550.0 545250.0 ;
      RECT  89100.0 542700.0 93900.0 543600.0 ;
      RECT  93450.0 537750.0 94350.0 543150.0 ;
      RECT  88500.0 545250.0 89700.0 546450.0 ;
      RECT  93300.0 545250.0 94500.0 546450.0 ;
      RECT  93300.0 536550.0 94500.0 537750.0 ;
      RECT  93300.0 542550.0 94500.0 543750.0 ;
      RECT  93450.0 559050.0 94350.0 551550.0 ;
      RECT  88650.0 554100.0 89550.0 553200.0 ;
      RECT  93450.0 554100.0 94350.0 553200.0 ;
      RECT  88650.0 553650.0 89550.0 551550.0 ;
      RECT  89100.0 554100.0 93900.0 553200.0 ;
      RECT  93450.0 559050.0 94350.0 553650.0 ;
      RECT  88500.0 551550.0 89700.0 550350.0 ;
      RECT  93300.0 551550.0 94500.0 550350.0 ;
      RECT  93300.0 560250.0 94500.0 559050.0 ;
      RECT  93300.0 554250.0 94500.0 553050.0 ;
      RECT  93450.0 565350.0 94350.0 572850.0 ;
      RECT  88650.0 570300.0 89550.0 571200.0 ;
      RECT  93450.0 570300.0 94350.0 571200.0 ;
      RECT  88650.0 570750.0 89550.0 572850.0 ;
      RECT  89100.0 570300.0 93900.0 571200.0 ;
      RECT  93450.0 565350.0 94350.0 570750.0 ;
      RECT  88500.0 572850.0 89700.0 574050.0 ;
      RECT  93300.0 572850.0 94500.0 574050.0 ;
      RECT  93300.0 564150.0 94500.0 565350.0 ;
      RECT  93300.0 570150.0 94500.0 571350.0 ;
      RECT  93450.0 586650.0 94350.0 579150.0 ;
      RECT  88650.0 581700.0 89550.0 580800.0 ;
      RECT  93450.0 581700.0 94350.0 580800.0 ;
      RECT  88650.0 581250.0 89550.0 579150.0 ;
      RECT  89100.0 581700.0 93900.0 580800.0 ;
      RECT  93450.0 586650.0 94350.0 581250.0 ;
      RECT  88500.0 579150.0 89700.0 577950.0 ;
      RECT  93300.0 579150.0 94500.0 577950.0 ;
      RECT  93300.0 587850.0 94500.0 586650.0 ;
      RECT  93300.0 581850.0 94500.0 580650.0 ;
      RECT  93450.0 592950.0 94350.0 600450.0 ;
      RECT  88650.0 597900.0 89550.0 598800.0 ;
      RECT  93450.0 597900.0 94350.0 598800.0 ;
      RECT  88650.0 598350.0 89550.0 600450.0 ;
      RECT  89100.0 597900.0 93900.0 598800.0 ;
      RECT  93450.0 592950.0 94350.0 598350.0 ;
      RECT  88500.0 600450.0 89700.0 601650.0 ;
      RECT  93300.0 600450.0 94500.0 601650.0 ;
      RECT  93300.0 591750.0 94500.0 592950.0 ;
      RECT  93300.0 597750.0 94500.0 598950.0 ;
      RECT  93450.0 614250.0 94350.0 606750.0 ;
      RECT  88650.0 609300.0 89550.0 608400.0 ;
      RECT  93450.0 609300.0 94350.0 608400.0 ;
      RECT  88650.0 608850.0 89550.0 606750.0 ;
      RECT  89100.0 609300.0 93900.0 608400.0 ;
      RECT  93450.0 614250.0 94350.0 608850.0 ;
      RECT  88500.0 606750.0 89700.0 605550.0 ;
      RECT  93300.0 606750.0 94500.0 605550.0 ;
      RECT  93300.0 615450.0 94500.0 614250.0 ;
      RECT  93300.0 609450.0 94500.0 608250.0 ;
      RECT  93450.0 620550.0 94350.0 628050.0 ;
      RECT  88650.0 625500.0 89550.0 626400.0 ;
      RECT  93450.0 625500.0 94350.0 626400.0 ;
      RECT  88650.0 625950.0 89550.0 628050.0 ;
      RECT  89100.0 625500.0 93900.0 626400.0 ;
      RECT  93450.0 620550.0 94350.0 625950.0 ;
      RECT  88500.0 628050.0 89700.0 629250.0 ;
      RECT  93300.0 628050.0 94500.0 629250.0 ;
      RECT  93300.0 619350.0 94500.0 620550.0 ;
      RECT  93300.0 625350.0 94500.0 626550.0 ;
      RECT  93450.0 641850.0 94350.0 634350.0 ;
      RECT  88650.0 636900.0 89550.0 636000.0 ;
      RECT  93450.0 636900.0 94350.0 636000.0 ;
      RECT  88650.0 636450.0 89550.0 634350.0 ;
      RECT  89100.0 636900.0 93900.0 636000.0 ;
      RECT  93450.0 641850.0 94350.0 636450.0 ;
      RECT  88500.0 634350.0 89700.0 633150.0 ;
      RECT  93300.0 634350.0 94500.0 633150.0 ;
      RECT  93300.0 643050.0 94500.0 641850.0 ;
      RECT  93300.0 637050.0 94500.0 635850.0 ;
      RECT  93450.0 648150.0 94350.0 655650.0 ;
      RECT  88650.0 653100.0 89550.0 654000.0 ;
      RECT  93450.0 653100.0 94350.0 654000.0 ;
      RECT  88650.0 653550.0 89550.0 655650.0 ;
      RECT  89100.0 653100.0 93900.0 654000.0 ;
      RECT  93450.0 648150.0 94350.0 653550.0 ;
      RECT  88500.0 655650.0 89700.0 656850.0 ;
      RECT  93300.0 655650.0 94500.0 656850.0 ;
      RECT  93300.0 646950.0 94500.0 648150.0 ;
      RECT  93300.0 652950.0 94500.0 654150.0 ;
      RECT  93450.0 669450.0 94350.0 661950.0 ;
      RECT  88650.0 664500.0 89550.0 663600.0 ;
      RECT  93450.0 664500.0 94350.0 663600.0 ;
      RECT  88650.0 664050.0 89550.0 661950.0 ;
      RECT  89100.0 664500.0 93900.0 663600.0 ;
      RECT  93450.0 669450.0 94350.0 664050.0 ;
      RECT  88500.0 661950.0 89700.0 660750.0 ;
      RECT  93300.0 661950.0 94500.0 660750.0 ;
      RECT  93300.0 670650.0 94500.0 669450.0 ;
      RECT  93300.0 664650.0 94500.0 663450.0 ;
      RECT  93450.0 675750.0 94350.0 683250.0 ;
      RECT  88650.0 680700.0 89550.0 681600.0 ;
      RECT  93450.0 680700.0 94350.0 681600.0 ;
      RECT  88650.0 681150.0 89550.0 683250.0 ;
      RECT  89100.0 680700.0 93900.0 681600.0 ;
      RECT  93450.0 675750.0 94350.0 681150.0 ;
      RECT  88500.0 683250.0 89700.0 684450.0 ;
      RECT  93300.0 683250.0 94500.0 684450.0 ;
      RECT  93300.0 674550.0 94500.0 675750.0 ;
      RECT  93300.0 680550.0 94500.0 681750.0 ;
      RECT  93450.0 697050.0 94350.0 689550.0 ;
      RECT  88650.0 692100.0 89550.0 691200.0 ;
      RECT  93450.0 692100.0 94350.0 691200.0 ;
      RECT  88650.0 691650.0 89550.0 689550.0 ;
      RECT  89100.0 692100.0 93900.0 691200.0 ;
      RECT  93450.0 697050.0 94350.0 691650.0 ;
      RECT  88500.0 689550.0 89700.0 688350.0 ;
      RECT  93300.0 689550.0 94500.0 688350.0 ;
      RECT  93300.0 698250.0 94500.0 697050.0 ;
      RECT  93300.0 692250.0 94500.0 691050.0 ;
      RECT  93450.0 703350.0 94350.0 710850.0 ;
      RECT  88650.0 708300.0 89550.0 709200.0 ;
      RECT  93450.0 708300.0 94350.0 709200.0 ;
      RECT  88650.0 708750.0 89550.0 710850.0 ;
      RECT  89100.0 708300.0 93900.0 709200.0 ;
      RECT  93450.0 703350.0 94350.0 708750.0 ;
      RECT  88500.0 710850.0 89700.0 712050.0 ;
      RECT  93300.0 710850.0 94500.0 712050.0 ;
      RECT  93300.0 702150.0 94500.0 703350.0 ;
      RECT  93300.0 708150.0 94500.0 709350.0 ;
      RECT  93450.0 724650.0 94350.0 717150.0 ;
      RECT  88650.0 719700.0 89550.0 718800.0 ;
      RECT  93450.0 719700.0 94350.0 718800.0 ;
      RECT  88650.0 719250.0 89550.0 717150.0 ;
      RECT  89100.0 719700.0 93900.0 718800.0 ;
      RECT  93450.0 724650.0 94350.0 719250.0 ;
      RECT  88500.0 717150.0 89700.0 715950.0 ;
      RECT  93300.0 717150.0 94500.0 715950.0 ;
      RECT  93300.0 725850.0 94500.0 724650.0 ;
      RECT  93300.0 719850.0 94500.0 718650.0 ;
      RECT  93450.0 730950.0 94350.0 738450.0 ;
      RECT  88650.0 735900.0 89550.0 736800.0 ;
      RECT  93450.0 735900.0 94350.0 736800.0 ;
      RECT  88650.0 736350.0 89550.0 738450.0 ;
      RECT  89100.0 735900.0 93900.0 736800.0 ;
      RECT  93450.0 730950.0 94350.0 736350.0 ;
      RECT  88500.0 738450.0 89700.0 739650.0 ;
      RECT  93300.0 738450.0 94500.0 739650.0 ;
      RECT  93300.0 729750.0 94500.0 730950.0 ;
      RECT  93300.0 735750.0 94500.0 736950.0 ;
      RECT  93450.0 752250.0 94350.0 744750.0 ;
      RECT  88650.0 747300.0 89550.0 746400.0 ;
      RECT  93450.0 747300.0 94350.0 746400.0 ;
      RECT  88650.0 746850.0 89550.0 744750.0 ;
      RECT  89100.0 747300.0 93900.0 746400.0 ;
      RECT  93450.0 752250.0 94350.0 746850.0 ;
      RECT  88500.0 744750.0 89700.0 743550.0 ;
      RECT  93300.0 744750.0 94500.0 743550.0 ;
      RECT  93300.0 753450.0 94500.0 752250.0 ;
      RECT  93300.0 747450.0 94500.0 746250.0 ;
      RECT  93450.0 758550.0 94350.0 766050.0 ;
      RECT  88650.0 763500.0 89550.0 764400.0 ;
      RECT  93450.0 763500.0 94350.0 764400.0 ;
      RECT  88650.0 763950.0 89550.0 766050.0 ;
      RECT  89100.0 763500.0 93900.0 764400.0 ;
      RECT  93450.0 758550.0 94350.0 763950.0 ;
      RECT  88500.0 766050.0 89700.0 767250.0 ;
      RECT  93300.0 766050.0 94500.0 767250.0 ;
      RECT  93300.0 757350.0 94500.0 758550.0 ;
      RECT  93300.0 763350.0 94500.0 764550.0 ;
      RECT  93450.0 779850.0 94350.0 772350.0 ;
      RECT  88650.0 774900.0 89550.0 774000.0 ;
      RECT  93450.0 774900.0 94350.0 774000.0 ;
      RECT  88650.0 774450.0 89550.0 772350.0 ;
      RECT  89100.0 774900.0 93900.0 774000.0 ;
      RECT  93450.0 779850.0 94350.0 774450.0 ;
      RECT  88500.0 772350.0 89700.0 771150.0 ;
      RECT  93300.0 772350.0 94500.0 771150.0 ;
      RECT  93300.0 781050.0 94500.0 779850.0 ;
      RECT  93300.0 775050.0 94500.0 773850.0 ;
      RECT  93450.0 786150.0 94350.0 793650.0 ;
      RECT  88650.0 791100.0 89550.0 792000.0 ;
      RECT  93450.0 791100.0 94350.0 792000.0 ;
      RECT  88650.0 791550.0 89550.0 793650.0 ;
      RECT  89100.0 791100.0 93900.0 792000.0 ;
      RECT  93450.0 786150.0 94350.0 791550.0 ;
      RECT  88500.0 793650.0 89700.0 794850.0 ;
      RECT  93300.0 793650.0 94500.0 794850.0 ;
      RECT  93300.0 784950.0 94500.0 786150.0 ;
      RECT  93300.0 790950.0 94500.0 792150.0 ;
      RECT  93450.0 807450.0 94350.0 799950.0 ;
      RECT  88650.0 802500.0 89550.0 801600.0 ;
      RECT  93450.0 802500.0 94350.0 801600.0 ;
      RECT  88650.0 802050.0 89550.0 799950.0 ;
      RECT  89100.0 802500.0 93900.0 801600.0 ;
      RECT  93450.0 807450.0 94350.0 802050.0 ;
      RECT  88500.0 799950.0 89700.0 798750.0 ;
      RECT  93300.0 799950.0 94500.0 798750.0 ;
      RECT  93300.0 808650.0 94500.0 807450.0 ;
      RECT  93300.0 802650.0 94500.0 801450.0 ;
      RECT  93450.0 813750.0 94350.0 821250.0 ;
      RECT  88650.0 818700.0 89550.0 819600.0 ;
      RECT  93450.0 818700.0 94350.0 819600.0 ;
      RECT  88650.0 819150.0 89550.0 821250.0 ;
      RECT  89100.0 818700.0 93900.0 819600.0 ;
      RECT  93450.0 813750.0 94350.0 819150.0 ;
      RECT  88500.0 821250.0 89700.0 822450.0 ;
      RECT  93300.0 821250.0 94500.0 822450.0 ;
      RECT  93300.0 812550.0 94500.0 813750.0 ;
      RECT  93300.0 818550.0 94500.0 819750.0 ;
      RECT  93450.0 835050.0 94350.0 827550.0 ;
      RECT  88650.0 830100.0 89550.0 829200.0 ;
      RECT  93450.0 830100.0 94350.0 829200.0 ;
      RECT  88650.0 829650.0 89550.0 827550.0 ;
      RECT  89100.0 830100.0 93900.0 829200.0 ;
      RECT  93450.0 835050.0 94350.0 829650.0 ;
      RECT  88500.0 827550.0 89700.0 826350.0 ;
      RECT  93300.0 827550.0 94500.0 826350.0 ;
      RECT  93300.0 836250.0 94500.0 835050.0 ;
      RECT  93300.0 830250.0 94500.0 829050.0 ;
      RECT  93450.0 841350.0 94350.0 848850.0 ;
      RECT  88650.0 846300.0 89550.0 847200.0 ;
      RECT  93450.0 846300.0 94350.0 847200.0 ;
      RECT  88650.0 846750.0 89550.0 848850.0 ;
      RECT  89100.0 846300.0 93900.0 847200.0 ;
      RECT  93450.0 841350.0 94350.0 846750.0 ;
      RECT  88500.0 848850.0 89700.0 850050.0 ;
      RECT  93300.0 848850.0 94500.0 850050.0 ;
      RECT  93300.0 840150.0 94500.0 841350.0 ;
      RECT  93300.0 846150.0 94500.0 847350.0 ;
      RECT  93450.0 862650.0 94350.0 855150.0 ;
      RECT  88650.0 857700.0 89550.0 856800.0 ;
      RECT  93450.0 857700.0 94350.0 856800.0 ;
      RECT  88650.0 857250.0 89550.0 855150.0 ;
      RECT  89100.0 857700.0 93900.0 856800.0 ;
      RECT  93450.0 862650.0 94350.0 857250.0 ;
      RECT  88500.0 855150.0 89700.0 853950.0 ;
      RECT  93300.0 855150.0 94500.0 853950.0 ;
      RECT  93300.0 863850.0 94500.0 862650.0 ;
      RECT  93300.0 857850.0 94500.0 856650.0 ;
      RECT  93450.0 868950.0 94350.0 876450.0 ;
      RECT  88650.0 873900.0 89550.0 874800.0 ;
      RECT  93450.0 873900.0 94350.0 874800.0 ;
      RECT  88650.0 874350.0 89550.0 876450.0 ;
      RECT  89100.0 873900.0 93900.0 874800.0 ;
      RECT  93450.0 868950.0 94350.0 874350.0 ;
      RECT  88500.0 876450.0 89700.0 877650.0 ;
      RECT  93300.0 876450.0 94500.0 877650.0 ;
      RECT  93300.0 867750.0 94500.0 868950.0 ;
      RECT  93300.0 873750.0 94500.0 874950.0 ;
      RECT  93450.0 890250.0 94350.0 882750.0 ;
      RECT  88650.0 885300.0 89550.0 884400.0 ;
      RECT  93450.0 885300.0 94350.0 884400.0 ;
      RECT  88650.0 884850.0 89550.0 882750.0 ;
      RECT  89100.0 885300.0 93900.0 884400.0 ;
      RECT  93450.0 890250.0 94350.0 884850.0 ;
      RECT  88500.0 882750.0 89700.0 881550.0 ;
      RECT  93300.0 882750.0 94500.0 881550.0 ;
      RECT  93300.0 891450.0 94500.0 890250.0 ;
      RECT  93300.0 885450.0 94500.0 884250.0 ;
      RECT  93450.0 896550.0 94350.0 904050.0 ;
      RECT  88650.0 901500.0 89550.0 902400.0 ;
      RECT  93450.0 901500.0 94350.0 902400.0 ;
      RECT  88650.0 901950.0 89550.0 904050.0 ;
      RECT  89100.0 901500.0 93900.0 902400.0 ;
      RECT  93450.0 896550.0 94350.0 901950.0 ;
      RECT  88500.0 904050.0 89700.0 905250.0 ;
      RECT  93300.0 904050.0 94500.0 905250.0 ;
      RECT  93300.0 895350.0 94500.0 896550.0 ;
      RECT  93300.0 901350.0 94500.0 902550.0 ;
      RECT  93450.0 917850.0 94350.0 910350.0 ;
      RECT  88650.0 912900.0 89550.0 912000.0 ;
      RECT  93450.0 912900.0 94350.0 912000.0 ;
      RECT  88650.0 912450.0 89550.0 910350.0 ;
      RECT  89100.0 912900.0 93900.0 912000.0 ;
      RECT  93450.0 917850.0 94350.0 912450.0 ;
      RECT  88500.0 910350.0 89700.0 909150.0 ;
      RECT  93300.0 910350.0 94500.0 909150.0 ;
      RECT  93300.0 919050.0 94500.0 917850.0 ;
      RECT  93300.0 913050.0 94500.0 911850.0 ;
      RECT  93450.0 924150.0 94350.0 931650.0 ;
      RECT  88650.0 929100.0 89550.0 930000.0 ;
      RECT  93450.0 929100.0 94350.0 930000.0 ;
      RECT  88650.0 929550.0 89550.0 931650.0 ;
      RECT  89100.0 929100.0 93900.0 930000.0 ;
      RECT  93450.0 924150.0 94350.0 929550.0 ;
      RECT  88500.0 931650.0 89700.0 932850.0 ;
      RECT  93300.0 931650.0 94500.0 932850.0 ;
      RECT  93300.0 922950.0 94500.0 924150.0 ;
      RECT  93300.0 928950.0 94500.0 930150.0 ;
      RECT  93450.0 945450.0 94350.0 937950.0 ;
      RECT  88650.0 940500.0 89550.0 939600.0 ;
      RECT  93450.0 940500.0 94350.0 939600.0 ;
      RECT  88650.0 940050.0 89550.0 937950.0 ;
      RECT  89100.0 940500.0 93900.0 939600.0 ;
      RECT  93450.0 945450.0 94350.0 940050.0 ;
      RECT  88500.0 937950.0 89700.0 936750.0 ;
      RECT  93300.0 937950.0 94500.0 936750.0 ;
      RECT  93300.0 946650.0 94500.0 945450.0 ;
      RECT  93300.0 940650.0 94500.0 939450.0 ;
      RECT  93450.0 951750.0 94350.0 959250.0 ;
      RECT  88650.0 956700.0 89550.0 957600.0 ;
      RECT  93450.0 956700.0 94350.0 957600.0 ;
      RECT  88650.0 957150.0 89550.0 959250.0 ;
      RECT  89100.0 956700.0 93900.0 957600.0 ;
      RECT  93450.0 951750.0 94350.0 957150.0 ;
      RECT  88500.0 959250.0 89700.0 960450.0 ;
      RECT  93300.0 959250.0 94500.0 960450.0 ;
      RECT  93300.0 950550.0 94500.0 951750.0 ;
      RECT  93300.0 956550.0 94500.0 957750.0 ;
      RECT  93450.0 973050.0 94350.0 965550.0 ;
      RECT  88650.0 968100.0 89550.0 967200.0 ;
      RECT  93450.0 968100.0 94350.0 967200.0 ;
      RECT  88650.0 967650.0 89550.0 965550.0 ;
      RECT  89100.0 968100.0 93900.0 967200.0 ;
      RECT  93450.0 973050.0 94350.0 967650.0 ;
      RECT  88500.0 965550.0 89700.0 964350.0 ;
      RECT  93300.0 965550.0 94500.0 964350.0 ;
      RECT  93300.0 974250.0 94500.0 973050.0 ;
      RECT  93300.0 968250.0 94500.0 967050.0 ;
      RECT  93450.0 979350.0 94350.0 986850.0 ;
      RECT  88650.0 984300.0 89550.0 985200.0 ;
      RECT  93450.0 984300.0 94350.0 985200.0 ;
      RECT  88650.0 984750.0 89550.0 986850.0 ;
      RECT  89100.0 984300.0 93900.0 985200.0 ;
      RECT  93450.0 979350.0 94350.0 984750.0 ;
      RECT  88500.0 986850.0 89700.0 988050.0 ;
      RECT  93300.0 986850.0 94500.0 988050.0 ;
      RECT  93300.0 978150.0 94500.0 979350.0 ;
      RECT  93300.0 984150.0 94500.0 985350.0 ;
      RECT  93450.0 1000650.0 94350.0 993150.0 ;
      RECT  88650.0 995700.0 89550.0 994800.0 ;
      RECT  93450.0 995700.0 94350.0 994800.0 ;
      RECT  88650.0 995250.0 89550.0 993150.0 ;
      RECT  89100.0 995700.0 93900.0 994800.0 ;
      RECT  93450.0 1000650.0 94350.0 995250.0 ;
      RECT  88500.0 993150.0 89700.0 991950.0 ;
      RECT  93300.0 993150.0 94500.0 991950.0 ;
      RECT  93300.0 1001850.0 94500.0 1000650.0 ;
      RECT  93300.0 995850.0 94500.0 994650.0 ;
      RECT  93450.0 1006950.0 94350.0 1014450.0 ;
      RECT  88650.0 1011900.0 89550.0 1012800.0 ;
      RECT  93450.0 1011900.0 94350.0 1012800.0 ;
      RECT  88650.0 1012350.0 89550.0 1014450.0 ;
      RECT  89100.0 1011900.0 93900.0 1012800.0 ;
      RECT  93450.0 1006950.0 94350.0 1012350.0 ;
      RECT  88500.0 1014450.0 89700.0 1015650.0 ;
      RECT  93300.0 1014450.0 94500.0 1015650.0 ;
      RECT  93300.0 1005750.0 94500.0 1006950.0 ;
      RECT  93300.0 1011750.0 94500.0 1012950.0 ;
      RECT  93450.0 1028250.0 94350.0 1020750.0 ;
      RECT  88650.0 1023300.0 89550.0 1022400.0 ;
      RECT  93450.0 1023300.0 94350.0 1022400.0 ;
      RECT  88650.0 1022850.0 89550.0 1020750.0 ;
      RECT  89100.0 1023300.0 93900.0 1022400.0 ;
      RECT  93450.0 1028250.0 94350.0 1022850.0 ;
      RECT  88500.0 1020750.0 89700.0 1019550.0 ;
      RECT  93300.0 1020750.0 94500.0 1019550.0 ;
      RECT  93300.0 1029450.0 94500.0 1028250.0 ;
      RECT  93300.0 1023450.0 94500.0 1022250.0 ;
      RECT  93450.0 1034550.0 94350.0 1042050.0 ;
      RECT  88650.0 1039500.0 89550.0 1040400.0 ;
      RECT  93450.0 1039500.0 94350.0 1040400.0 ;
      RECT  88650.0 1039950.0 89550.0 1042050.0 ;
      RECT  89100.0 1039500.0 93900.0 1040400.0 ;
      RECT  93450.0 1034550.0 94350.0 1039950.0 ;
      RECT  88500.0 1042050.0 89700.0 1043250.0 ;
      RECT  93300.0 1042050.0 94500.0 1043250.0 ;
      RECT  93300.0 1033350.0 94500.0 1034550.0 ;
      RECT  93300.0 1039350.0 94500.0 1040550.0 ;
      RECT  93450.0 1055850.0 94350.0 1048350.0 ;
      RECT  88650.0 1050900.0 89550.0 1050000.0 ;
      RECT  93450.0 1050900.0 94350.0 1050000.0 ;
      RECT  88650.0 1050450.0 89550.0 1048350.0 ;
      RECT  89100.0 1050900.0 93900.0 1050000.0 ;
      RECT  93450.0 1055850.0 94350.0 1050450.0 ;
      RECT  88500.0 1048350.0 89700.0 1047150.0 ;
      RECT  93300.0 1048350.0 94500.0 1047150.0 ;
      RECT  93300.0 1057050.0 94500.0 1055850.0 ;
      RECT  93300.0 1051050.0 94500.0 1049850.0 ;
      RECT  93450.0 1062150.0 94350.0 1069650.0 ;
      RECT  88650.0 1067100.0 89550.0 1068000.0 ;
      RECT  93450.0 1067100.0 94350.0 1068000.0 ;
      RECT  88650.0 1067550.0 89550.0 1069650.0 ;
      RECT  89100.0 1067100.0 93900.0 1068000.0 ;
      RECT  93450.0 1062150.0 94350.0 1067550.0 ;
      RECT  88500.0 1069650.0 89700.0 1070850.0 ;
      RECT  93300.0 1069650.0 94500.0 1070850.0 ;
      RECT  93300.0 1060950.0 94500.0 1062150.0 ;
      RECT  93300.0 1066950.0 94500.0 1068150.0 ;
      RECT  93450.0 1083450.0 94350.0 1075950.0 ;
      RECT  88650.0 1078500.0 89550.0 1077600.0 ;
      RECT  93450.0 1078500.0 94350.0 1077600.0 ;
      RECT  88650.0 1078050.0 89550.0 1075950.0 ;
      RECT  89100.0 1078500.0 93900.0 1077600.0 ;
      RECT  93450.0 1083450.0 94350.0 1078050.0 ;
      RECT  88500.0 1075950.0 89700.0 1074750.0 ;
      RECT  93300.0 1075950.0 94500.0 1074750.0 ;
      RECT  93300.0 1084650.0 94500.0 1083450.0 ;
      RECT  93300.0 1078650.0 94500.0 1077450.0 ;
      RECT  93450.0 1089750.0 94350.0 1097250.0 ;
      RECT  88650.0 1094700.0 89550.0 1095600.0 ;
      RECT  93450.0 1094700.0 94350.0 1095600.0 ;
      RECT  88650.0 1095150.0 89550.0 1097250.0 ;
      RECT  89100.0 1094700.0 93900.0 1095600.0 ;
      RECT  93450.0 1089750.0 94350.0 1095150.0 ;
      RECT  88500.0 1097250.0 89700.0 1098450.0 ;
      RECT  93300.0 1097250.0 94500.0 1098450.0 ;
      RECT  93300.0 1088550.0 94500.0 1089750.0 ;
      RECT  93300.0 1094550.0 94500.0 1095750.0 ;
      RECT  93450.0 1111050.0 94350.0 1103550.0 ;
      RECT  88650.0 1106100.0 89550.0 1105200.0 ;
      RECT  93450.0 1106100.0 94350.0 1105200.0 ;
      RECT  88650.0 1105650.0 89550.0 1103550.0 ;
      RECT  89100.0 1106100.0 93900.0 1105200.0 ;
      RECT  93450.0 1111050.0 94350.0 1105650.0 ;
      RECT  88500.0 1103550.0 89700.0 1102350.0 ;
      RECT  93300.0 1103550.0 94500.0 1102350.0 ;
      RECT  93300.0 1112250.0 94500.0 1111050.0 ;
      RECT  93300.0 1106250.0 94500.0 1105050.0 ;
      RECT  93450.0 1117350.0 94350.0 1124850.0 ;
      RECT  88650.0 1122300.0 89550.0 1123200.0 ;
      RECT  93450.0 1122300.0 94350.0 1123200.0 ;
      RECT  88650.0 1122750.0 89550.0 1124850.0 ;
      RECT  89100.0 1122300.0 93900.0 1123200.0 ;
      RECT  93450.0 1117350.0 94350.0 1122750.0 ;
      RECT  88500.0 1124850.0 89700.0 1126050.0 ;
      RECT  93300.0 1124850.0 94500.0 1126050.0 ;
      RECT  93300.0 1116150.0 94500.0 1117350.0 ;
      RECT  93300.0 1122150.0 94500.0 1123350.0 ;
      RECT  93450.0 1138650.0 94350.0 1131150.0 ;
      RECT  88650.0 1133700.0 89550.0 1132800.0 ;
      RECT  93450.0 1133700.0 94350.0 1132800.0 ;
      RECT  88650.0 1133250.0 89550.0 1131150.0 ;
      RECT  89100.0 1133700.0 93900.0 1132800.0 ;
      RECT  93450.0 1138650.0 94350.0 1133250.0 ;
      RECT  88500.0 1131150.0 89700.0 1129950.0 ;
      RECT  93300.0 1131150.0 94500.0 1129950.0 ;
      RECT  93300.0 1139850.0 94500.0 1138650.0 ;
      RECT  93300.0 1133850.0 94500.0 1132650.0 ;
      RECT  93450.0 1144950.0 94350.0 1152450.0 ;
      RECT  88650.0 1149900.0 89550.0 1150800.0 ;
      RECT  93450.0 1149900.0 94350.0 1150800.0 ;
      RECT  88650.0 1150350.0 89550.0 1152450.0 ;
      RECT  89100.0 1149900.0 93900.0 1150800.0 ;
      RECT  93450.0 1144950.0 94350.0 1150350.0 ;
      RECT  88500.0 1152450.0 89700.0 1153650.0 ;
      RECT  93300.0 1152450.0 94500.0 1153650.0 ;
      RECT  93300.0 1143750.0 94500.0 1144950.0 ;
      RECT  93300.0 1149750.0 94500.0 1150950.0 ;
      RECT  93450.0 1166250.0 94350.0 1158750.0 ;
      RECT  88650.0 1161300.0 89550.0 1160400.0 ;
      RECT  93450.0 1161300.0 94350.0 1160400.0 ;
      RECT  88650.0 1160850.0 89550.0 1158750.0 ;
      RECT  89100.0 1161300.0 93900.0 1160400.0 ;
      RECT  93450.0 1166250.0 94350.0 1160850.0 ;
      RECT  88500.0 1158750.0 89700.0 1157550.0 ;
      RECT  93300.0 1158750.0 94500.0 1157550.0 ;
      RECT  93300.0 1167450.0 94500.0 1166250.0 ;
      RECT  93300.0 1161450.0 94500.0 1160250.0 ;
      RECT  93450.0 1172550.0 94350.0 1180050.0 ;
      RECT  88650.0 1177500.0 89550.0 1178400.0 ;
      RECT  93450.0 1177500.0 94350.0 1178400.0 ;
      RECT  88650.0 1177950.0 89550.0 1180050.0 ;
      RECT  89100.0 1177500.0 93900.0 1178400.0 ;
      RECT  93450.0 1172550.0 94350.0 1177950.0 ;
      RECT  88500.0 1180050.0 89700.0 1181250.0 ;
      RECT  93300.0 1180050.0 94500.0 1181250.0 ;
      RECT  93300.0 1171350.0 94500.0 1172550.0 ;
      RECT  93300.0 1177350.0 94500.0 1178550.0 ;
      RECT  93450.0 1193850.0 94350.0 1186350.0 ;
      RECT  88650.0 1188900.0 89550.0 1188000.0 ;
      RECT  93450.0 1188900.0 94350.0 1188000.0 ;
      RECT  88650.0 1188450.0 89550.0 1186350.0 ;
      RECT  89100.0 1188900.0 93900.0 1188000.0 ;
      RECT  93450.0 1193850.0 94350.0 1188450.0 ;
      RECT  88500.0 1186350.0 89700.0 1185150.0 ;
      RECT  93300.0 1186350.0 94500.0 1185150.0 ;
      RECT  93300.0 1195050.0 94500.0 1193850.0 ;
      RECT  93300.0 1189050.0 94500.0 1187850.0 ;
      RECT  60150.0 154200.0 58950.0 155400.0 ;
      RECT  62250.0 168600.0 61050.0 169800.0 ;
      RECT  64350.0 181800.0 63150.0 183000.0 ;
      RECT  66450.0 196200.0 65250.0 197400.0 ;
      RECT  68550.0 209400.0 67350.0 210600.0 ;
      RECT  70650.0 223800.0 69450.0 225000.0 ;
      RECT  72750.0 237000.0 71550.0 238200.0 ;
      RECT  74850.0 251400.0 73650.0 252600.0 ;
      RECT  76950.0 264600.0 75750.0 265800.0 ;
      RECT  79050.0 279000.0 77850.0 280200.0 ;
      RECT  81150.0 292200.0 79950.0 293400.0 ;
      RECT  83250.0 306600.0 82050.0 307800.0 ;
      RECT  60150.0 321750.0 58950.0 322950.0 ;
      RECT  68550.0 319800.0 67350.0 321000.0 ;
      RECT  76950.0 317850.0 75750.0 319050.0 ;
      RECT  60150.0 332250.0 58950.0 333450.0 ;
      RECT  68550.0 334200.0 67350.0 335400.0 ;
      RECT  79050.0 336150.0 77850.0 337350.0 ;
      RECT  60150.0 349350.0 58950.0 350550.0 ;
      RECT  68550.0 347400.0 67350.0 348600.0 ;
      RECT  81150.0 345450.0 79950.0 346650.0 ;
      RECT  60150.0 359850.0 58950.0 361050.0 ;
      RECT  68550.0 361800.0 67350.0 363000.0 ;
      RECT  83250.0 363750.0 82050.0 364950.0 ;
      RECT  60150.0 376950.0 58950.0 378150.0 ;
      RECT  70650.0 375000.0 69450.0 376200.0 ;
      RECT  76950.0 373050.0 75750.0 374250.0 ;
      RECT  60150.0 387450.0 58950.0 388650.0 ;
      RECT  70650.0 389400.0 69450.0 390600.0 ;
      RECT  79050.0 391350.0 77850.0 392550.0 ;
      RECT  60150.0 404550.0 58950.0 405750.0 ;
      RECT  70650.0 402600.0 69450.0 403800.0 ;
      RECT  81150.0 400650.0 79950.0 401850.0 ;
      RECT  60150.0 415050.0 58950.0 416250.0 ;
      RECT  70650.0 417000.0 69450.0 418200.0 ;
      RECT  83250.0 418950.0 82050.0 420150.0 ;
      RECT  60150.0 432150.0 58950.0 433350.0 ;
      RECT  72750.0 430200.0 71550.0 431400.0 ;
      RECT  76950.0 428250.0 75750.0 429450.0 ;
      RECT  60150.0 442650.0 58950.0 443850.0 ;
      RECT  72750.0 444600.0 71550.0 445800.0 ;
      RECT  79050.0 446550.0 77850.0 447750.0 ;
      RECT  60150.0 459750.0 58950.0 460950.0 ;
      RECT  72750.0 457800.0 71550.0 459000.0 ;
      RECT  81150.0 455850.0 79950.0 457050.0 ;
      RECT  60150.0 470250.0 58950.0 471450.0 ;
      RECT  72750.0 472200.0 71550.0 473400.0 ;
      RECT  83250.0 474150.0 82050.0 475350.0 ;
      RECT  60150.0 487350.0 58950.0 488550.0 ;
      RECT  74850.0 485400.0 73650.0 486600.0 ;
      RECT  76950.0 483450.0 75750.0 484650.0 ;
      RECT  60150.0 497850.0 58950.0 499050.0 ;
      RECT  74850.0 499800.0 73650.0 501000.0 ;
      RECT  79050.0 501750.0 77850.0 502950.0 ;
      RECT  60150.0 514950.0 58950.0 516150.0 ;
      RECT  74850.0 513000.0 73650.0 514200.0 ;
      RECT  81150.0 511050.0 79950.0 512250.0 ;
      RECT  60150.0 525450.0 58950.0 526650.0 ;
      RECT  74850.0 527400.0 73650.0 528600.0 ;
      RECT  83250.0 529350.0 82050.0 530550.0 ;
      RECT  62250.0 542550.0 61050.0 543750.0 ;
      RECT  68550.0 540600.0 67350.0 541800.0 ;
      RECT  76950.0 538650.0 75750.0 539850.0 ;
      RECT  62250.0 553050.0 61050.0 554250.0 ;
      RECT  68550.0 555000.0 67350.0 556200.0 ;
      RECT  79050.0 556950.0 77850.0 558150.0 ;
      RECT  62250.0 570150.0 61050.0 571350.0 ;
      RECT  68550.0 568200.0 67350.0 569400.0 ;
      RECT  81150.0 566250.0 79950.0 567450.0 ;
      RECT  62250.0 580650.0 61050.0 581850.0 ;
      RECT  68550.0 582600.0 67350.0 583800.0 ;
      RECT  83250.0 584550.0 82050.0 585750.0 ;
      RECT  62250.0 597750.0 61050.0 598950.0 ;
      RECT  70650.0 595800.0 69450.0 597000.0 ;
      RECT  76950.0 593850.0 75750.0 595050.0 ;
      RECT  62250.0 608250.0 61050.0 609450.0 ;
      RECT  70650.0 610200.0 69450.0 611400.0 ;
      RECT  79050.0 612150.0 77850.0 613350.0 ;
      RECT  62250.0 625350.0 61050.0 626550.0 ;
      RECT  70650.0 623400.0 69450.0 624600.0 ;
      RECT  81150.0 621450.0 79950.0 622650.0 ;
      RECT  62250.0 635850.0 61050.0 637050.0 ;
      RECT  70650.0 637800.0 69450.0 639000.0 ;
      RECT  83250.0 639750.0 82050.0 640950.0 ;
      RECT  62250.0 652950.0 61050.0 654150.0 ;
      RECT  72750.0 651000.0 71550.0 652200.0 ;
      RECT  76950.0 649050.0 75750.0 650250.0 ;
      RECT  62250.0 663450.0 61050.0 664650.0 ;
      RECT  72750.0 665400.0 71550.0 666600.0 ;
      RECT  79050.0 667350.0 77850.0 668550.0 ;
      RECT  62250.0 680550.0 61050.0 681750.0 ;
      RECT  72750.0 678600.0 71550.0 679800.0 ;
      RECT  81150.0 676650.0 79950.0 677850.0 ;
      RECT  62250.0 691050.0 61050.0 692250.0 ;
      RECT  72750.0 693000.0 71550.0 694200.0 ;
      RECT  83250.0 694950.0 82050.0 696150.0 ;
      RECT  62250.0 708150.0 61050.0 709350.0 ;
      RECT  74850.0 706200.0 73650.0 707400.0 ;
      RECT  76950.0 704250.0 75750.0 705450.0 ;
      RECT  62250.0 718650.0 61050.0 719850.0 ;
      RECT  74850.0 720600.0 73650.0 721800.0 ;
      RECT  79050.0 722550.0 77850.0 723750.0 ;
      RECT  62250.0 735750.0 61050.0 736950.0 ;
      RECT  74850.0 733800.0 73650.0 735000.0 ;
      RECT  81150.0 731850.0 79950.0 733050.0 ;
      RECT  62250.0 746250.0 61050.0 747450.0 ;
      RECT  74850.0 748200.0 73650.0 749400.0 ;
      RECT  83250.0 750150.0 82050.0 751350.0 ;
      RECT  64350.0 763350.0 63150.0 764550.0 ;
      RECT  68550.0 761400.0 67350.0 762600.0 ;
      RECT  76950.0 759450.0 75750.0 760650.0 ;
      RECT  64350.0 773850.0 63150.0 775050.0 ;
      RECT  68550.0 775800.0 67350.0 777000.0 ;
      RECT  79050.0 777750.0 77850.0 778950.0 ;
      RECT  64350.0 790950.0 63150.0 792150.0 ;
      RECT  68550.0 789000.0 67350.0 790200.0 ;
      RECT  81150.0 787050.0 79950.0 788250.0 ;
      RECT  64350.0 801450.0 63150.0 802650.0 ;
      RECT  68550.0 803400.0 67350.0 804600.0 ;
      RECT  83250.0 805350.0 82050.0 806550.0 ;
      RECT  64350.0 818550.0 63150.0 819750.0 ;
      RECT  70650.0 816600.0 69450.0 817800.0 ;
      RECT  76950.0 814650.0 75750.0 815850.0 ;
      RECT  64350.0 829050.0 63150.0 830250.0 ;
      RECT  70650.0 831000.0 69450.0 832200.0 ;
      RECT  79050.0 832950.0 77850.0 834150.0 ;
      RECT  64350.0 846150.0 63150.0 847350.0 ;
      RECT  70650.0 844200.0 69450.0 845400.0 ;
      RECT  81150.0 842250.0 79950.0 843450.0 ;
      RECT  64350.0 856650.0 63150.0 857850.0 ;
      RECT  70650.0 858600.0 69450.0 859800.0 ;
      RECT  83250.0 860550.0 82050.0 861750.0 ;
      RECT  64350.0 873750.0 63150.0 874950.0 ;
      RECT  72750.0 871800.0 71550.0 873000.0 ;
      RECT  76950.0 869850.0 75750.0 871050.0 ;
      RECT  64350.0 884250.0 63150.0 885450.0 ;
      RECT  72750.0 886200.0 71550.0 887400.0 ;
      RECT  79050.0 888150.0 77850.0 889350.0 ;
      RECT  64350.0 901350.0 63150.0 902550.0 ;
      RECT  72750.0 899400.0 71550.0 900600.0 ;
      RECT  81150.0 897450.0 79950.0 898650.0 ;
      RECT  64350.0 911850.0 63150.0 913050.0 ;
      RECT  72750.0 913800.0 71550.0 915000.0 ;
      RECT  83250.0 915750.0 82050.0 916950.0 ;
      RECT  64350.0 928950.0 63150.0 930150.0 ;
      RECT  74850.0 927000.0 73650.0 928200.0 ;
      RECT  76950.0 925050.0 75750.0 926250.0 ;
      RECT  64350.0 939450.0 63150.0 940650.0 ;
      RECT  74850.0 941400.0 73650.0 942600.0 ;
      RECT  79050.0 943350.0 77850.0 944550.0 ;
      RECT  64350.0 956550.0 63150.0 957750.0 ;
      RECT  74850.0 954600.0 73650.0 955800.0 ;
      RECT  81150.0 952650.0 79950.0 953850.0 ;
      RECT  64350.0 967050.0 63150.0 968250.0 ;
      RECT  74850.0 969000.0 73650.0 970200.0 ;
      RECT  83250.0 970950.0 82050.0 972150.0 ;
      RECT  66450.0 984150.0 65250.0 985350.0 ;
      RECT  68550.0 982200.0 67350.0 983400.0 ;
      RECT  76950.0 980250.0 75750.0 981450.0 ;
      RECT  66450.0 994650.0 65250.0 995850.0 ;
      RECT  68550.0 996600.0 67350.0 997800.0 ;
      RECT  79050.0 998550.0 77850.0 999750.0 ;
      RECT  66450.0 1011750.0 65250.0 1012950.0 ;
      RECT  68550.0 1009800.0 67350.0 1011000.0 ;
      RECT  81150.0 1007850.0 79950.0 1009050.0 ;
      RECT  66450.0 1022250.0 65250.0 1023450.0 ;
      RECT  68550.0 1024200.0 67350.0 1025400.0 ;
      RECT  83250.0 1026150.0 82050.0 1027350.0 ;
      RECT  66450.0 1039350.0 65250.0 1040550.0 ;
      RECT  70650.0 1037400.0 69450.0 1038600.0 ;
      RECT  76950.0 1035450.0 75750.0 1036650.0 ;
      RECT  66450.0 1049850.0 65250.0 1051050.0 ;
      RECT  70650.0 1051800.0 69450.0 1053000.0 ;
      RECT  79050.0 1053750.0 77850.0 1054950.0 ;
      RECT  66450.0 1066950.0 65250.0 1068150.0 ;
      RECT  70650.0 1065000.0 69450.0 1066200.0 ;
      RECT  81150.0 1063050.0 79950.0 1064250.0 ;
      RECT  66450.0 1077450.0 65250.0 1078650.0 ;
      RECT  70650.0 1079400.0 69450.0 1080600.0 ;
      RECT  83250.0 1081350.0 82050.0 1082550.0 ;
      RECT  66450.0 1094550.0 65250.0 1095750.0 ;
      RECT  72750.0 1092600.0 71550.0 1093800.0 ;
      RECT  76950.0 1090650.0 75750.0 1091850.0 ;
      RECT  66450.0 1105050.0 65250.0 1106250.0 ;
      RECT  72750.0 1107000.0 71550.0 1108200.0 ;
      RECT  79050.0 1108950.0 77850.0 1110150.0 ;
      RECT  66450.0 1122150.0 65250.0 1123350.0 ;
      RECT  72750.0 1120200.0 71550.0 1121400.0 ;
      RECT  81150.0 1118250.0 79950.0 1119450.0 ;
      RECT  66450.0 1132650.0 65250.0 1133850.0 ;
      RECT  72750.0 1134600.0 71550.0 1135800.0 ;
      RECT  83250.0 1136550.0 82050.0 1137750.0 ;
      RECT  66450.0 1149750.0 65250.0 1150950.0 ;
      RECT  74850.0 1147800.0 73650.0 1149000.0 ;
      RECT  76950.0 1145850.0 75750.0 1147050.0 ;
      RECT  66450.0 1160250.0 65250.0 1161450.0 ;
      RECT  74850.0 1162200.0 73650.0 1163400.0 ;
      RECT  79050.0 1164150.0 77850.0 1165350.0 ;
      RECT  66450.0 1177350.0 65250.0 1178550.0 ;
      RECT  74850.0 1175400.0 73650.0 1176600.0 ;
      RECT  81150.0 1173450.0 79950.0 1174650.0 ;
      RECT  66450.0 1187850.0 65250.0 1189050.0 ;
      RECT  74850.0 1189800.0 73650.0 1191000.0 ;
      RECT  83250.0 1191750.0 82050.0 1192950.0 ;
      RECT  138000.0 148200.0 138900.0 201600.0 ;
      RECT  135000.0 148200.0 135900.0 201600.0 ;
      RECT  138000.0 203400.0 138900.0 256800.0 ;
      RECT  135000.0 203400.0 135900.0 256800.0 ;
      RECT  138000.0 258600.0 138900.0 312000.0 ;
      RECT  135000.0 258600.0 135900.0 312000.0 ;
      RECT  114150.0 318450.0 115050.0 319350.0 ;
      RECT  114150.0 318000.0 115050.0 318900.0 ;
      RECT  114600.0 318450.0 130800.0 319350.0 ;
      RECT  114150.0 335850.0 115050.0 336750.0 ;
      RECT  114150.0 336300.0 115050.0 337200.0 ;
      RECT  114600.0 335850.0 130800.0 336750.0 ;
      RECT  114150.0 346050.0 115050.0 346950.0 ;
      RECT  114150.0 345600.0 115050.0 346500.0 ;
      RECT  114600.0 346050.0 130800.0 346950.0 ;
      RECT  114150.0 363450.0 115050.0 364350.0 ;
      RECT  114150.0 363900.0 115050.0 364800.0 ;
      RECT  114600.0 363450.0 130800.0 364350.0 ;
      RECT  114150.0 373650.0 115050.0 374550.0 ;
      RECT  114150.0 373200.0 115050.0 374100.0 ;
      RECT  114600.0 373650.0 130800.0 374550.0 ;
      RECT  114150.0 391050.0 115050.0 391950.0 ;
      RECT  114150.0 391500.0 115050.0 392400.0 ;
      RECT  114600.0 391050.0 130800.0 391950.0 ;
      RECT  114150.0 401250.0 115050.0 402150.0 ;
      RECT  114150.0 400800.0 115050.0 401700.0 ;
      RECT  114600.0 401250.0 130800.0 402150.0 ;
      RECT  114150.0 418650.0 115050.0 419550.0 ;
      RECT  114150.0 419100.0 115050.0 420000.0 ;
      RECT  114600.0 418650.0 130800.0 419550.0 ;
      RECT  114150.0 428850.0 115050.0 429750.0 ;
      RECT  114150.0 428400.0 115050.0 429300.0 ;
      RECT  114600.0 428850.0 130800.0 429750.0 ;
      RECT  114150.0 446250.0 115050.0 447150.0 ;
      RECT  114150.0 446700.0 115050.0 447600.0 ;
      RECT  114600.0 446250.0 130800.0 447150.0 ;
      RECT  114150.0 456450.0 115050.0 457350.0 ;
      RECT  114150.0 456000.0 115050.0 456900.0 ;
      RECT  114600.0 456450.0 130800.0 457350.0 ;
      RECT  114150.0 473850.0 115050.0 474750.0 ;
      RECT  114150.0 474300.0 115050.0 475200.0 ;
      RECT  114600.0 473850.0 130800.0 474750.0 ;
      RECT  114150.0 484050.0 115050.0 484950.0 ;
      RECT  114150.0 483600.0 115050.0 484500.0 ;
      RECT  114600.0 484050.0 130800.0 484950.0 ;
      RECT  114150.0 501450.0 115050.0 502350.0 ;
      RECT  114150.0 501900.0 115050.0 502800.0 ;
      RECT  114600.0 501450.0 130800.0 502350.0 ;
      RECT  114150.0 511650.0 115050.0 512550.0 ;
      RECT  114150.0 511200.0 115050.0 512100.0 ;
      RECT  114600.0 511650.0 130800.0 512550.0 ;
      RECT  114150.0 529050.0 115050.0 529950.0 ;
      RECT  114150.0 529500.0 115050.0 530400.0 ;
      RECT  114600.0 529050.0 130800.0 529950.0 ;
      RECT  114150.0 539250.0 115050.0 540150.0 ;
      RECT  114150.0 538800.0 115050.0 539700.0 ;
      RECT  114600.0 539250.0 130800.0 540150.0 ;
      RECT  114150.0 556650.0 115050.0 557550.0 ;
      RECT  114150.0 557100.0 115050.0 558000.0 ;
      RECT  114600.0 556650.0 130800.0 557550.0 ;
      RECT  114150.0 566850.0 115050.0 567750.0 ;
      RECT  114150.0 566400.0 115050.0 567300.0 ;
      RECT  114600.0 566850.0 130800.0 567750.0 ;
      RECT  114150.0 584250.0 115050.0 585150.0 ;
      RECT  114150.0 584700.0 115050.0 585600.0 ;
      RECT  114600.0 584250.0 130800.0 585150.0 ;
      RECT  114150.0 594450.0 115050.0 595350.0 ;
      RECT  114150.0 594000.0 115050.0 594900.0 ;
      RECT  114600.0 594450.0 130800.0 595350.0 ;
      RECT  114150.0 611850.0 115050.0 612750.0 ;
      RECT  114150.0 612300.0 115050.0 613200.0 ;
      RECT  114600.0 611850.0 130800.0 612750.0 ;
      RECT  114150.0 622050.0 115050.0 622950.0 ;
      RECT  114150.0 621600.0 115050.0 622500.0 ;
      RECT  114600.0 622050.0 130800.0 622950.0 ;
      RECT  114150.0 639450.0 115050.0 640350.0 ;
      RECT  114150.0 639900.0 115050.0 640800.0 ;
      RECT  114600.0 639450.0 130800.0 640350.0 ;
      RECT  114150.0 649650.0 115050.0 650550.0 ;
      RECT  114150.0 649200.0 115050.0 650100.0 ;
      RECT  114600.0 649650.0 130800.0 650550.0 ;
      RECT  114150.0 667050.0 115050.0 667950.0 ;
      RECT  114150.0 667500.0 115050.0 668400.0 ;
      RECT  114600.0 667050.0 130800.0 667950.0 ;
      RECT  114150.0 677250.0 115050.0 678150.0 ;
      RECT  114150.0 676800.0 115050.0 677700.0 ;
      RECT  114600.0 677250.0 130800.0 678150.0 ;
      RECT  114150.0 694650.0 115050.0 695550.0 ;
      RECT  114150.0 695100.0 115050.0 696000.0 ;
      RECT  114600.0 694650.0 130800.0 695550.0 ;
      RECT  114150.0 704850.0 115050.0 705750.0 ;
      RECT  114150.0 704400.0 115050.0 705300.0 ;
      RECT  114600.0 704850.0 130800.0 705750.0 ;
      RECT  114150.0 722250.0 115050.0 723150.0 ;
      RECT  114150.0 722700.0 115050.0 723600.0 ;
      RECT  114600.0 722250.0 130800.0 723150.0 ;
      RECT  114150.0 732450.0 115050.0 733350.0 ;
      RECT  114150.0 732000.0 115050.0 732900.0 ;
      RECT  114600.0 732450.0 130800.0 733350.0 ;
      RECT  114150.0 749850.0 115050.0 750750.0 ;
      RECT  114150.0 750300.0 115050.0 751200.0 ;
      RECT  114600.0 749850.0 130800.0 750750.0 ;
      RECT  114150.0 760050.0 115050.0 760950.0 ;
      RECT  114150.0 759600.0 115050.0 760500.0 ;
      RECT  114600.0 760050.0 130800.0 760950.0 ;
      RECT  114150.0 777450.0 115050.0 778350.0 ;
      RECT  114150.0 777900.0 115050.0 778800.0 ;
      RECT  114600.0 777450.0 130800.0 778350.0 ;
      RECT  114150.0 787650.0 115050.0 788550.0 ;
      RECT  114150.0 787200.0 115050.0 788100.0 ;
      RECT  114600.0 787650.0 130800.0 788550.0 ;
      RECT  114150.0 805050.0 115050.0 805950.0 ;
      RECT  114150.0 805500.0 115050.0 806400.0 ;
      RECT  114600.0 805050.0 130800.0 805950.0 ;
      RECT  114150.0 815250.0 115050.0 816150.0 ;
      RECT  114150.0 814800.0 115050.0 815700.0 ;
      RECT  114600.0 815250.0 130800.0 816150.0 ;
      RECT  114150.0 832650.0 115050.0 833550.0 ;
      RECT  114150.0 833100.0 115050.0 834000.0 ;
      RECT  114600.0 832650.0 130800.0 833550.0 ;
      RECT  114150.0 842850.0 115050.0 843750.0 ;
      RECT  114150.0 842400.0 115050.0 843300.0 ;
      RECT  114600.0 842850.0 130800.0 843750.0 ;
      RECT  114150.0 860250.0 115050.0 861150.0 ;
      RECT  114150.0 860700.0 115050.0 861600.0 ;
      RECT  114600.0 860250.0 130800.0 861150.0 ;
      RECT  114150.0 870450.0 115050.0 871350.0 ;
      RECT  114150.0 870000.0 115050.0 870900.0 ;
      RECT  114600.0 870450.0 130800.0 871350.0 ;
      RECT  114150.0 887850.0 115050.0 888750.0 ;
      RECT  114150.0 888300.0 115050.0 889200.0 ;
      RECT  114600.0 887850.0 130800.0 888750.0 ;
      RECT  114150.0 898050.0 115050.0 898950.0 ;
      RECT  114150.0 897600.0 115050.0 898500.0 ;
      RECT  114600.0 898050.0 130800.0 898950.0 ;
      RECT  114150.0 915450.0 115050.0 916350.0 ;
      RECT  114150.0 915900.0 115050.0 916800.0 ;
      RECT  114600.0 915450.0 130800.0 916350.0 ;
      RECT  114150.0 925650.0 115050.0 926550.0 ;
      RECT  114150.0 925200.0 115050.0 926100.0 ;
      RECT  114600.0 925650.0 130800.0 926550.0 ;
      RECT  114150.0 943050.0 115050.0 943950.0 ;
      RECT  114150.0 943500.0 115050.0 944400.0 ;
      RECT  114600.0 943050.0 130800.0 943950.0 ;
      RECT  114150.0 953250.0 115050.0 954150.0 ;
      RECT  114150.0 952800.0 115050.0 953700.0 ;
      RECT  114600.0 953250.0 130800.0 954150.0 ;
      RECT  114150.0 970650.0 115050.0 971550.0 ;
      RECT  114150.0 971100.0 115050.0 972000.0 ;
      RECT  114600.0 970650.0 130800.0 971550.0 ;
      RECT  114150.0 980850.0 115050.0 981750.0 ;
      RECT  114150.0 980400.0 115050.0 981300.0 ;
      RECT  114600.0 980850.0 130800.0 981750.0 ;
      RECT  114150.0 998250.0 115050.0 999150.0 ;
      RECT  114150.0 998700.0 115050.0 999600.0 ;
      RECT  114600.0 998250.0 130800.0 999150.0 ;
      RECT  114150.0 1008450.0 115050.0 1009350.0 ;
      RECT  114150.0 1008000.0 115050.0 1008900.0 ;
      RECT  114600.0 1008450.0 130800.0 1009350.0 ;
      RECT  114150.0 1025850.0 115050.0 1026750.0 ;
      RECT  114150.0 1026300.0 115050.0 1027200.0 ;
      RECT  114600.0 1025850.0 130800.0 1026750.0 ;
      RECT  114150.0 1036050.0 115050.0 1036950.0 ;
      RECT  114150.0 1035600.0 115050.0 1036500.0 ;
      RECT  114600.0 1036050.0 130800.0 1036950.0 ;
      RECT  114150.0 1053450.0 115050.0 1054350.0 ;
      RECT  114150.0 1053900.0 115050.0 1054800.0 ;
      RECT  114600.0 1053450.0 130800.0 1054350.0 ;
      RECT  114150.0 1063650.0 115050.0 1064550.0 ;
      RECT  114150.0 1063200.0 115050.0 1064100.0 ;
      RECT  114600.0 1063650.0 130800.0 1064550.0 ;
      RECT  114150.0 1081050.0 115050.0 1081950.0 ;
      RECT  114150.0 1081500.0 115050.0 1082400.0 ;
      RECT  114600.0 1081050.0 130800.0 1081950.0 ;
      RECT  114150.0 1091250.0 115050.0 1092150.0 ;
      RECT  114150.0 1090800.0 115050.0 1091700.0 ;
      RECT  114600.0 1091250.0 130800.0 1092150.0 ;
      RECT  114150.0 1108650.0 115050.0 1109550.0 ;
      RECT  114150.0 1109100.0 115050.0 1110000.0 ;
      RECT  114600.0 1108650.0 130800.0 1109550.0 ;
      RECT  114150.0 1118850.0 115050.0 1119750.0 ;
      RECT  114150.0 1118400.0 115050.0 1119300.0 ;
      RECT  114600.0 1118850.0 130800.0 1119750.0 ;
      RECT  114150.0 1136250.0 115050.0 1137150.0 ;
      RECT  114150.0 1136700.0 115050.0 1137600.0 ;
      RECT  114600.0 1136250.0 130800.0 1137150.0 ;
      RECT  114150.0 1146450.0 115050.0 1147350.0 ;
      RECT  114150.0 1146000.0 115050.0 1146900.0 ;
      RECT  114600.0 1146450.0 130800.0 1147350.0 ;
      RECT  114150.0 1163850.0 115050.0 1164750.0 ;
      RECT  114150.0 1164300.0 115050.0 1165200.0 ;
      RECT  114600.0 1163850.0 130800.0 1164750.0 ;
      RECT  114150.0 1174050.0 115050.0 1174950.0 ;
      RECT  114150.0 1173600.0 115050.0 1174500.0 ;
      RECT  114600.0 1174050.0 130800.0 1174950.0 ;
      RECT  114150.0 1191450.0 115050.0 1192350.0 ;
      RECT  114150.0 1191900.0 115050.0 1192800.0 ;
      RECT  114600.0 1191450.0 130800.0 1192350.0 ;
      RECT  129750.0 321150.0 130650.0 322050.0 ;
      RECT  132150.0 321150.0 133050.0 322050.0 ;
      RECT  129750.0 321600.0 130650.0 324450.0 ;
      RECT  130200.0 321150.0 132600.0 322050.0 ;
      RECT  132150.0 316950.0 133050.0 321600.0 ;
      RECT  129600.0 324450.0 130800.0 325650.0 ;
      RECT  132000.0 315750.0 133200.0 316950.0 ;
      RECT  133200.0 321000.0 132000.0 322200.0 ;
      RECT  112050.0 319800.0 113250.0 321000.0 ;
      RECT  114000.0 317400.0 115200.0 318600.0 ;
      RECT  130800.0 318300.0 129600.0 319500.0 ;
      RECT  129750.0 334050.0 130650.0 333150.0 ;
      RECT  132150.0 334050.0 133050.0 333150.0 ;
      RECT  129750.0 333600.0 130650.0 330750.0 ;
      RECT  130200.0 334050.0 132600.0 333150.0 ;
      RECT  132150.0 338250.0 133050.0 333600.0 ;
      RECT  129600.0 330750.0 130800.0 329550.0 ;
      RECT  132000.0 339450.0 133200.0 338250.0 ;
      RECT  133200.0 334200.0 132000.0 333000.0 ;
      RECT  112050.0 334200.0 113250.0 335400.0 ;
      RECT  114000.0 336600.0 115200.0 337800.0 ;
      RECT  130800.0 335700.0 129600.0 336900.0 ;
      RECT  129750.0 348750.0 130650.0 349650.0 ;
      RECT  132150.0 348750.0 133050.0 349650.0 ;
      RECT  129750.0 349200.0 130650.0 352050.0 ;
      RECT  130200.0 348750.0 132600.0 349650.0 ;
      RECT  132150.0 344550.0 133050.0 349200.0 ;
      RECT  129600.0 352050.0 130800.0 353250.0 ;
      RECT  132000.0 343350.0 133200.0 344550.0 ;
      RECT  133200.0 348600.0 132000.0 349800.0 ;
      RECT  112050.0 347400.0 113250.0 348600.0 ;
      RECT  114000.0 345000.0 115200.0 346200.0 ;
      RECT  130800.0 345900.0 129600.0 347100.0 ;
      RECT  129750.0 361650.0 130650.0 360750.0 ;
      RECT  132150.0 361650.0 133050.0 360750.0 ;
      RECT  129750.0 361200.0 130650.0 358350.0 ;
      RECT  130200.0 361650.0 132600.0 360750.0 ;
      RECT  132150.0 365850.0 133050.0 361200.0 ;
      RECT  129600.0 358350.0 130800.0 357150.0 ;
      RECT  132000.0 367050.0 133200.0 365850.0 ;
      RECT  133200.0 361800.0 132000.0 360600.0 ;
      RECT  112050.0 361800.0 113250.0 363000.0 ;
      RECT  114000.0 364200.0 115200.0 365400.0 ;
      RECT  130800.0 363300.0 129600.0 364500.0 ;
      RECT  129750.0 376350.0 130650.0 377250.0 ;
      RECT  132150.0 376350.0 133050.0 377250.0 ;
      RECT  129750.0 376800.0 130650.0 379650.0 ;
      RECT  130200.0 376350.0 132600.0 377250.0 ;
      RECT  132150.0 372150.0 133050.0 376800.0 ;
      RECT  129600.0 379650.0 130800.0 380850.0 ;
      RECT  132000.0 370950.0 133200.0 372150.0 ;
      RECT  133200.0 376200.0 132000.0 377400.0 ;
      RECT  112050.0 375000.0 113250.0 376200.0 ;
      RECT  114000.0 372600.0 115200.0 373800.0 ;
      RECT  130800.0 373500.0 129600.0 374700.0 ;
      RECT  129750.0 389250.0 130650.0 388350.0 ;
      RECT  132150.0 389250.0 133050.0 388350.0 ;
      RECT  129750.0 388800.0 130650.0 385950.0 ;
      RECT  130200.0 389250.0 132600.0 388350.0 ;
      RECT  132150.0 393450.0 133050.0 388800.0 ;
      RECT  129600.0 385950.0 130800.0 384750.0 ;
      RECT  132000.0 394650.0 133200.0 393450.0 ;
      RECT  133200.0 389400.0 132000.0 388200.0 ;
      RECT  112050.0 389400.0 113250.0 390600.0 ;
      RECT  114000.0 391800.0 115200.0 393000.0 ;
      RECT  130800.0 390900.0 129600.0 392100.0 ;
      RECT  129750.0 403950.0 130650.0 404850.0 ;
      RECT  132150.0 403950.0 133050.0 404850.0 ;
      RECT  129750.0 404400.0 130650.0 407250.0 ;
      RECT  130200.0 403950.0 132600.0 404850.0 ;
      RECT  132150.0 399750.0 133050.0 404400.0 ;
      RECT  129600.0 407250.0 130800.0 408450.0 ;
      RECT  132000.0 398550.0 133200.0 399750.0 ;
      RECT  133200.0 403800.0 132000.0 405000.0 ;
      RECT  112050.0 402600.0 113250.0 403800.0 ;
      RECT  114000.0 400200.0 115200.0 401400.0 ;
      RECT  130800.0 401100.0 129600.0 402300.0 ;
      RECT  129750.0 416850.0 130650.0 415950.0 ;
      RECT  132150.0 416850.0 133050.0 415950.0 ;
      RECT  129750.0 416400.0 130650.0 413550.0 ;
      RECT  130200.0 416850.0 132600.0 415950.0 ;
      RECT  132150.0 421050.0 133050.0 416400.0 ;
      RECT  129600.0 413550.0 130800.0 412350.0 ;
      RECT  132000.0 422250.0 133200.0 421050.0 ;
      RECT  133200.0 417000.0 132000.0 415800.0 ;
      RECT  112050.0 417000.0 113250.0 418200.0 ;
      RECT  114000.0 419400.0 115200.0 420600.0 ;
      RECT  130800.0 418500.0 129600.0 419700.0 ;
      RECT  129750.0 431550.0 130650.0 432450.0 ;
      RECT  132150.0 431550.0 133050.0 432450.0 ;
      RECT  129750.0 432000.0 130650.0 434850.0 ;
      RECT  130200.0 431550.0 132600.0 432450.0 ;
      RECT  132150.0 427350.0 133050.0 432000.0 ;
      RECT  129600.0 434850.0 130800.0 436050.0 ;
      RECT  132000.0 426150.0 133200.0 427350.0 ;
      RECT  133200.0 431400.0 132000.0 432600.0 ;
      RECT  112050.0 430200.0 113250.0 431400.0 ;
      RECT  114000.0 427800.0 115200.0 429000.0 ;
      RECT  130800.0 428700.0 129600.0 429900.0 ;
      RECT  129750.0 444450.0 130650.0 443550.0 ;
      RECT  132150.0 444450.0 133050.0 443550.0 ;
      RECT  129750.0 444000.0 130650.0 441150.0 ;
      RECT  130200.0 444450.0 132600.0 443550.0 ;
      RECT  132150.0 448650.0 133050.0 444000.0 ;
      RECT  129600.0 441150.0 130800.0 439950.0 ;
      RECT  132000.0 449850.0 133200.0 448650.0 ;
      RECT  133200.0 444600.0 132000.0 443400.0 ;
      RECT  112050.0 444600.0 113250.0 445800.0 ;
      RECT  114000.0 447000.0 115200.0 448200.0 ;
      RECT  130800.0 446100.0 129600.0 447300.0 ;
      RECT  129750.0 459150.0 130650.0 460050.0 ;
      RECT  132150.0 459150.0 133050.0 460050.0 ;
      RECT  129750.0 459600.0 130650.0 462450.0 ;
      RECT  130200.0 459150.0 132600.0 460050.0 ;
      RECT  132150.0 454950.0 133050.0 459600.0 ;
      RECT  129600.0 462450.0 130800.0 463650.0 ;
      RECT  132000.0 453750.0 133200.0 454950.0 ;
      RECT  133200.0 459000.0 132000.0 460200.0 ;
      RECT  112050.0 457800.0 113250.0 459000.0 ;
      RECT  114000.0 455400.0 115200.0 456600.0 ;
      RECT  130800.0 456300.0 129600.0 457500.0 ;
      RECT  129750.0 472050.0 130650.0 471150.0 ;
      RECT  132150.0 472050.0 133050.0 471150.0 ;
      RECT  129750.0 471600.0 130650.0 468750.0 ;
      RECT  130200.0 472050.0 132600.0 471150.0 ;
      RECT  132150.0 476250.0 133050.0 471600.0 ;
      RECT  129600.0 468750.0 130800.0 467550.0 ;
      RECT  132000.0 477450.0 133200.0 476250.0 ;
      RECT  133200.0 472200.0 132000.0 471000.0 ;
      RECT  112050.0 472200.0 113250.0 473400.0 ;
      RECT  114000.0 474600.0 115200.0 475800.0 ;
      RECT  130800.0 473700.0 129600.0 474900.0 ;
      RECT  129750.0 486750.0 130650.0 487650.0 ;
      RECT  132150.0 486750.0 133050.0 487650.0 ;
      RECT  129750.0 487200.0 130650.0 490050.0 ;
      RECT  130200.0 486750.0 132600.0 487650.0 ;
      RECT  132150.0 482550.0 133050.0 487200.0 ;
      RECT  129600.0 490050.0 130800.0 491250.0 ;
      RECT  132000.0 481350.0 133200.0 482550.0 ;
      RECT  133200.0 486600.0 132000.0 487800.0 ;
      RECT  112050.0 485400.0 113250.0 486600.0 ;
      RECT  114000.0 483000.0 115200.0 484200.0 ;
      RECT  130800.0 483900.0 129600.0 485100.0 ;
      RECT  129750.0 499650.0 130650.0 498750.0 ;
      RECT  132150.0 499650.0 133050.0 498750.0 ;
      RECT  129750.0 499200.0 130650.0 496350.0 ;
      RECT  130200.0 499650.0 132600.0 498750.0 ;
      RECT  132150.0 503850.0 133050.0 499200.0 ;
      RECT  129600.0 496350.0 130800.0 495150.0 ;
      RECT  132000.0 505050.0 133200.0 503850.0 ;
      RECT  133200.0 499800.0 132000.0 498600.0 ;
      RECT  112050.0 499800.0 113250.0 501000.0 ;
      RECT  114000.0 502200.0 115200.0 503400.0 ;
      RECT  130800.0 501300.0 129600.0 502500.0 ;
      RECT  129750.0 514350.0 130650.0 515250.0 ;
      RECT  132150.0 514350.0 133050.0 515250.0 ;
      RECT  129750.0 514800.0 130650.0 517650.0 ;
      RECT  130200.0 514350.0 132600.0 515250.0 ;
      RECT  132150.0 510150.0 133050.0 514800.0 ;
      RECT  129600.0 517650.0 130800.0 518850.0 ;
      RECT  132000.0 508950.0 133200.0 510150.0 ;
      RECT  133200.0 514200.0 132000.0 515400.0 ;
      RECT  112050.0 513000.0 113250.0 514200.0 ;
      RECT  114000.0 510600.0 115200.0 511800.0 ;
      RECT  130800.0 511500.0 129600.0 512700.0 ;
      RECT  129750.0 527250.0 130650.0 526350.0 ;
      RECT  132150.0 527250.0 133050.0 526350.0 ;
      RECT  129750.0 526800.0 130650.0 523950.0 ;
      RECT  130200.0 527250.0 132600.0 526350.0 ;
      RECT  132150.0 531450.0 133050.0 526800.0 ;
      RECT  129600.0 523950.0 130800.0 522750.0 ;
      RECT  132000.0 532650.0 133200.0 531450.0 ;
      RECT  133200.0 527400.0 132000.0 526200.0 ;
      RECT  112050.0 527400.0 113250.0 528600.0 ;
      RECT  114000.0 529800.0 115200.0 531000.0 ;
      RECT  130800.0 528900.0 129600.0 530100.0 ;
      RECT  129750.0 541950.0 130650.0 542850.0 ;
      RECT  132150.0 541950.0 133050.0 542850.0 ;
      RECT  129750.0 542400.0 130650.0 545250.0 ;
      RECT  130200.0 541950.0 132600.0 542850.0 ;
      RECT  132150.0 537750.0 133050.0 542400.0 ;
      RECT  129600.0 545250.0 130800.0 546450.0 ;
      RECT  132000.0 536550.0 133200.0 537750.0 ;
      RECT  133200.0 541800.0 132000.0 543000.0 ;
      RECT  112050.0 540600.0 113250.0 541800.0 ;
      RECT  114000.0 538200.0 115200.0 539400.0 ;
      RECT  130800.0 539100.0 129600.0 540300.0 ;
      RECT  129750.0 554850.0 130650.0 553950.0 ;
      RECT  132150.0 554850.0 133050.0 553950.0 ;
      RECT  129750.0 554400.0 130650.0 551550.0 ;
      RECT  130200.0 554850.0 132600.0 553950.0 ;
      RECT  132150.0 559050.0 133050.0 554400.0 ;
      RECT  129600.0 551550.0 130800.0 550350.0 ;
      RECT  132000.0 560250.0 133200.0 559050.0 ;
      RECT  133200.0 555000.0 132000.0 553800.0 ;
      RECT  112050.0 555000.0 113250.0 556200.0 ;
      RECT  114000.0 557400.0 115200.0 558600.0 ;
      RECT  130800.0 556500.0 129600.0 557700.0 ;
      RECT  129750.0 569550.0 130650.0 570450.0 ;
      RECT  132150.0 569550.0 133050.0 570450.0 ;
      RECT  129750.0 570000.0 130650.0 572850.0 ;
      RECT  130200.0 569550.0 132600.0 570450.0 ;
      RECT  132150.0 565350.0 133050.0 570000.0 ;
      RECT  129600.0 572850.0 130800.0 574050.0 ;
      RECT  132000.0 564150.0 133200.0 565350.0 ;
      RECT  133200.0 569400.0 132000.0 570600.0 ;
      RECT  112050.0 568200.0 113250.0 569400.0 ;
      RECT  114000.0 565800.0 115200.0 567000.0 ;
      RECT  130800.0 566700.0 129600.0 567900.0 ;
      RECT  129750.0 582450.0 130650.0 581550.0 ;
      RECT  132150.0 582450.0 133050.0 581550.0 ;
      RECT  129750.0 582000.0 130650.0 579150.0 ;
      RECT  130200.0 582450.0 132600.0 581550.0 ;
      RECT  132150.0 586650.0 133050.0 582000.0 ;
      RECT  129600.0 579150.0 130800.0 577950.0 ;
      RECT  132000.0 587850.0 133200.0 586650.0 ;
      RECT  133200.0 582600.0 132000.0 581400.0 ;
      RECT  112050.0 582600.0 113250.0 583800.0 ;
      RECT  114000.0 585000.0 115200.0 586200.0 ;
      RECT  130800.0 584100.0 129600.0 585300.0 ;
      RECT  129750.0 597150.0 130650.0 598050.0 ;
      RECT  132150.0 597150.0 133050.0 598050.0 ;
      RECT  129750.0 597600.0 130650.0 600450.0 ;
      RECT  130200.0 597150.0 132600.0 598050.0 ;
      RECT  132150.0 592950.0 133050.0 597600.0 ;
      RECT  129600.0 600450.0 130800.0 601650.0 ;
      RECT  132000.0 591750.0 133200.0 592950.0 ;
      RECT  133200.0 597000.0 132000.0 598200.0 ;
      RECT  112050.0 595800.0 113250.0 597000.0 ;
      RECT  114000.0 593400.0 115200.0 594600.0 ;
      RECT  130800.0 594300.0 129600.0 595500.0 ;
      RECT  129750.0 610050.0 130650.0 609150.0 ;
      RECT  132150.0 610050.0 133050.0 609150.0 ;
      RECT  129750.0 609600.0 130650.0 606750.0 ;
      RECT  130200.0 610050.0 132600.0 609150.0 ;
      RECT  132150.0 614250.0 133050.0 609600.0 ;
      RECT  129600.0 606750.0 130800.0 605550.0 ;
      RECT  132000.0 615450.0 133200.0 614250.0 ;
      RECT  133200.0 610200.0 132000.0 609000.0 ;
      RECT  112050.0 610200.0 113250.0 611400.0 ;
      RECT  114000.0 612600.0 115200.0 613800.0 ;
      RECT  130800.0 611700.0 129600.0 612900.0 ;
      RECT  129750.0 624750.0 130650.0 625650.0 ;
      RECT  132150.0 624750.0 133050.0 625650.0 ;
      RECT  129750.0 625200.0 130650.0 628050.0 ;
      RECT  130200.0 624750.0 132600.0 625650.0 ;
      RECT  132150.0 620550.0 133050.0 625200.0 ;
      RECT  129600.0 628050.0 130800.0 629250.0 ;
      RECT  132000.0 619350.0 133200.0 620550.0 ;
      RECT  133200.0 624600.0 132000.0 625800.0 ;
      RECT  112050.0 623400.0 113250.0 624600.0 ;
      RECT  114000.0 621000.0 115200.0 622200.0 ;
      RECT  130800.0 621900.0 129600.0 623100.0 ;
      RECT  129750.0 637650.0 130650.0 636750.0 ;
      RECT  132150.0 637650.0 133050.0 636750.0 ;
      RECT  129750.0 637200.0 130650.0 634350.0 ;
      RECT  130200.0 637650.0 132600.0 636750.0 ;
      RECT  132150.0 641850.0 133050.0 637200.0 ;
      RECT  129600.0 634350.0 130800.0 633150.0 ;
      RECT  132000.0 643050.0 133200.0 641850.0 ;
      RECT  133200.0 637800.0 132000.0 636600.0 ;
      RECT  112050.0 637800.0 113250.0 639000.0 ;
      RECT  114000.0 640200.0 115200.0 641400.0 ;
      RECT  130800.0 639300.0 129600.0 640500.0 ;
      RECT  129750.0 652350.0 130650.0 653250.0 ;
      RECT  132150.0 652350.0 133050.0 653250.0 ;
      RECT  129750.0 652800.0 130650.0 655650.0 ;
      RECT  130200.0 652350.0 132600.0 653250.0 ;
      RECT  132150.0 648150.0 133050.0 652800.0 ;
      RECT  129600.0 655650.0 130800.0 656850.0 ;
      RECT  132000.0 646950.0 133200.0 648150.0 ;
      RECT  133200.0 652200.0 132000.0 653400.0 ;
      RECT  112050.0 651000.0 113250.0 652200.0 ;
      RECT  114000.0 648600.0 115200.0 649800.0 ;
      RECT  130800.0 649500.0 129600.0 650700.0 ;
      RECT  129750.0 665250.0 130650.0 664350.0 ;
      RECT  132150.0 665250.0 133050.0 664350.0 ;
      RECT  129750.0 664800.0 130650.0 661950.0 ;
      RECT  130200.0 665250.0 132600.0 664350.0 ;
      RECT  132150.0 669450.0 133050.0 664800.0 ;
      RECT  129600.0 661950.0 130800.0 660750.0 ;
      RECT  132000.0 670650.0 133200.0 669450.0 ;
      RECT  133200.0 665400.0 132000.0 664200.0 ;
      RECT  112050.0 665400.0 113250.0 666600.0 ;
      RECT  114000.0 667800.0 115200.0 669000.0 ;
      RECT  130800.0 666900.0 129600.0 668100.0 ;
      RECT  129750.0 679950.0 130650.0 680850.0 ;
      RECT  132150.0 679950.0 133050.0 680850.0 ;
      RECT  129750.0 680400.0 130650.0 683250.0 ;
      RECT  130200.0 679950.0 132600.0 680850.0 ;
      RECT  132150.0 675750.0 133050.0 680400.0 ;
      RECT  129600.0 683250.0 130800.0 684450.0 ;
      RECT  132000.0 674550.0 133200.0 675750.0 ;
      RECT  133200.0 679800.0 132000.0 681000.0 ;
      RECT  112050.0 678600.0 113250.0 679800.0 ;
      RECT  114000.0 676200.0 115200.0 677400.0 ;
      RECT  130800.0 677100.0 129600.0 678300.0 ;
      RECT  129750.0 692850.0 130650.0 691950.0 ;
      RECT  132150.0 692850.0 133050.0 691950.0 ;
      RECT  129750.0 692400.0 130650.0 689550.0 ;
      RECT  130200.0 692850.0 132600.0 691950.0 ;
      RECT  132150.0 697050.0 133050.0 692400.0 ;
      RECT  129600.0 689550.0 130800.0 688350.0 ;
      RECT  132000.0 698250.0 133200.0 697050.0 ;
      RECT  133200.0 693000.0 132000.0 691800.0 ;
      RECT  112050.0 693000.0 113250.0 694200.0 ;
      RECT  114000.0 695400.0 115200.0 696600.0 ;
      RECT  130800.0 694500.0 129600.0 695700.0 ;
      RECT  129750.0 707550.0 130650.0 708450.0 ;
      RECT  132150.0 707550.0 133050.0 708450.0 ;
      RECT  129750.0 708000.0 130650.0 710850.0 ;
      RECT  130200.0 707550.0 132600.0 708450.0 ;
      RECT  132150.0 703350.0 133050.0 708000.0 ;
      RECT  129600.0 710850.0 130800.0 712050.0 ;
      RECT  132000.0 702150.0 133200.0 703350.0 ;
      RECT  133200.0 707400.0 132000.0 708600.0 ;
      RECT  112050.0 706200.0 113250.0 707400.0 ;
      RECT  114000.0 703800.0 115200.0 705000.0 ;
      RECT  130800.0 704700.0 129600.0 705900.0 ;
      RECT  129750.0 720450.0 130650.0 719550.0 ;
      RECT  132150.0 720450.0 133050.0 719550.0 ;
      RECT  129750.0 720000.0 130650.0 717150.0 ;
      RECT  130200.0 720450.0 132600.0 719550.0 ;
      RECT  132150.0 724650.0 133050.0 720000.0 ;
      RECT  129600.0 717150.0 130800.0 715950.0 ;
      RECT  132000.0 725850.0 133200.0 724650.0 ;
      RECT  133200.0 720600.0 132000.0 719400.0 ;
      RECT  112050.0 720600.0 113250.0 721800.0 ;
      RECT  114000.0 723000.0 115200.0 724200.0 ;
      RECT  130800.0 722100.0 129600.0 723300.0 ;
      RECT  129750.0 735150.0 130650.0 736050.0 ;
      RECT  132150.0 735150.0 133050.0 736050.0 ;
      RECT  129750.0 735600.0 130650.0 738450.0 ;
      RECT  130200.0 735150.0 132600.0 736050.0 ;
      RECT  132150.0 730950.0 133050.0 735600.0 ;
      RECT  129600.0 738450.0 130800.0 739650.0 ;
      RECT  132000.0 729750.0 133200.0 730950.0 ;
      RECT  133200.0 735000.0 132000.0 736200.0 ;
      RECT  112050.0 733800.0 113250.0 735000.0 ;
      RECT  114000.0 731400.0 115200.0 732600.0 ;
      RECT  130800.0 732300.0 129600.0 733500.0 ;
      RECT  129750.0 748050.0 130650.0 747150.0 ;
      RECT  132150.0 748050.0 133050.0 747150.0 ;
      RECT  129750.0 747600.0 130650.0 744750.0 ;
      RECT  130200.0 748050.0 132600.0 747150.0 ;
      RECT  132150.0 752250.0 133050.0 747600.0 ;
      RECT  129600.0 744750.0 130800.0 743550.0 ;
      RECT  132000.0 753450.0 133200.0 752250.0 ;
      RECT  133200.0 748200.0 132000.0 747000.0 ;
      RECT  112050.0 748200.0 113250.0 749400.0 ;
      RECT  114000.0 750600.0 115200.0 751800.0 ;
      RECT  130800.0 749700.0 129600.0 750900.0 ;
      RECT  129750.0 762750.0 130650.0 763650.0 ;
      RECT  132150.0 762750.0 133050.0 763650.0 ;
      RECT  129750.0 763200.0 130650.0 766050.0 ;
      RECT  130200.0 762750.0 132600.0 763650.0 ;
      RECT  132150.0 758550.0 133050.0 763200.0 ;
      RECT  129600.0 766050.0 130800.0 767250.0 ;
      RECT  132000.0 757350.0 133200.0 758550.0 ;
      RECT  133200.0 762600.0 132000.0 763800.0 ;
      RECT  112050.0 761400.0 113250.0 762600.0 ;
      RECT  114000.0 759000.0 115200.0 760200.0 ;
      RECT  130800.0 759900.0 129600.0 761100.0 ;
      RECT  129750.0 775650.0 130650.0 774750.0 ;
      RECT  132150.0 775650.0 133050.0 774750.0 ;
      RECT  129750.0 775200.0 130650.0 772350.0 ;
      RECT  130200.0 775650.0 132600.0 774750.0 ;
      RECT  132150.0 779850.0 133050.0 775200.0 ;
      RECT  129600.0 772350.0 130800.0 771150.0 ;
      RECT  132000.0 781050.0 133200.0 779850.0 ;
      RECT  133200.0 775800.0 132000.0 774600.0 ;
      RECT  112050.0 775800.0 113250.0 777000.0 ;
      RECT  114000.0 778200.0 115200.0 779400.0 ;
      RECT  130800.0 777300.0 129600.0 778500.0 ;
      RECT  129750.0 790350.0 130650.0 791250.0 ;
      RECT  132150.0 790350.0 133050.0 791250.0 ;
      RECT  129750.0 790800.0 130650.0 793650.0 ;
      RECT  130200.0 790350.0 132600.0 791250.0 ;
      RECT  132150.0 786150.0 133050.0 790800.0 ;
      RECT  129600.0 793650.0 130800.0 794850.0 ;
      RECT  132000.0 784950.0 133200.0 786150.0 ;
      RECT  133200.0 790200.0 132000.0 791400.0 ;
      RECT  112050.0 789000.0 113250.0 790200.0 ;
      RECT  114000.0 786600.0 115200.0 787800.0 ;
      RECT  130800.0 787500.0 129600.0 788700.0 ;
      RECT  129750.0 803250.0 130650.0 802350.0 ;
      RECT  132150.0 803250.0 133050.0 802350.0 ;
      RECT  129750.0 802800.0 130650.0 799950.0 ;
      RECT  130200.0 803250.0 132600.0 802350.0 ;
      RECT  132150.0 807450.0 133050.0 802800.0 ;
      RECT  129600.0 799950.0 130800.0 798750.0 ;
      RECT  132000.0 808650.0 133200.0 807450.0 ;
      RECT  133200.0 803400.0 132000.0 802200.0 ;
      RECT  112050.0 803400.0 113250.0 804600.0 ;
      RECT  114000.0 805800.0 115200.0 807000.0 ;
      RECT  130800.0 804900.0 129600.0 806100.0 ;
      RECT  129750.0 817950.0 130650.0 818850.0 ;
      RECT  132150.0 817950.0 133050.0 818850.0 ;
      RECT  129750.0 818400.0 130650.0 821250.0 ;
      RECT  130200.0 817950.0 132600.0 818850.0 ;
      RECT  132150.0 813750.0 133050.0 818400.0 ;
      RECT  129600.0 821250.0 130800.0 822450.0 ;
      RECT  132000.0 812550.0 133200.0 813750.0 ;
      RECT  133200.0 817800.0 132000.0 819000.0 ;
      RECT  112050.0 816600.0 113250.0 817800.0 ;
      RECT  114000.0 814200.0 115200.0 815400.0 ;
      RECT  130800.0 815100.0 129600.0 816300.0 ;
      RECT  129750.0 830850.0 130650.0 829950.0 ;
      RECT  132150.0 830850.0 133050.0 829950.0 ;
      RECT  129750.0 830400.0 130650.0 827550.0 ;
      RECT  130200.0 830850.0 132600.0 829950.0 ;
      RECT  132150.0 835050.0 133050.0 830400.0 ;
      RECT  129600.0 827550.0 130800.0 826350.0 ;
      RECT  132000.0 836250.0 133200.0 835050.0 ;
      RECT  133200.0 831000.0 132000.0 829800.0 ;
      RECT  112050.0 831000.0 113250.0 832200.0 ;
      RECT  114000.0 833400.0 115200.0 834600.0 ;
      RECT  130800.0 832500.0 129600.0 833700.0 ;
      RECT  129750.0 845550.0 130650.0 846450.0 ;
      RECT  132150.0 845550.0 133050.0 846450.0 ;
      RECT  129750.0 846000.0 130650.0 848850.0 ;
      RECT  130200.0 845550.0 132600.0 846450.0 ;
      RECT  132150.0 841350.0 133050.0 846000.0 ;
      RECT  129600.0 848850.0 130800.0 850050.0 ;
      RECT  132000.0 840150.0 133200.0 841350.0 ;
      RECT  133200.0 845400.0 132000.0 846600.0 ;
      RECT  112050.0 844200.0 113250.0 845400.0 ;
      RECT  114000.0 841800.0 115200.0 843000.0 ;
      RECT  130800.0 842700.0 129600.0 843900.0 ;
      RECT  129750.0 858450.0 130650.0 857550.0 ;
      RECT  132150.0 858450.0 133050.0 857550.0 ;
      RECT  129750.0 858000.0 130650.0 855150.0 ;
      RECT  130200.0 858450.0 132600.0 857550.0 ;
      RECT  132150.0 862650.0 133050.0 858000.0 ;
      RECT  129600.0 855150.0 130800.0 853950.0 ;
      RECT  132000.0 863850.0 133200.0 862650.0 ;
      RECT  133200.0 858600.0 132000.0 857400.0 ;
      RECT  112050.0 858600.0 113250.0 859800.0 ;
      RECT  114000.0 861000.0 115200.0 862200.0 ;
      RECT  130800.0 860100.0 129600.0 861300.0 ;
      RECT  129750.0 873150.0 130650.0 874050.0 ;
      RECT  132150.0 873150.0 133050.0 874050.0 ;
      RECT  129750.0 873600.0 130650.0 876450.0 ;
      RECT  130200.0 873150.0 132600.0 874050.0 ;
      RECT  132150.0 868950.0 133050.0 873600.0 ;
      RECT  129600.0 876450.0 130800.0 877650.0 ;
      RECT  132000.0 867750.0 133200.0 868950.0 ;
      RECT  133200.0 873000.0 132000.0 874200.0 ;
      RECT  112050.0 871800.0 113250.0 873000.0 ;
      RECT  114000.0 869400.0 115200.0 870600.0 ;
      RECT  130800.0 870300.0 129600.0 871500.0 ;
      RECT  129750.0 886050.0 130650.0 885150.0 ;
      RECT  132150.0 886050.0 133050.0 885150.0 ;
      RECT  129750.0 885600.0 130650.0 882750.0 ;
      RECT  130200.0 886050.0 132600.0 885150.0 ;
      RECT  132150.0 890250.0 133050.0 885600.0 ;
      RECT  129600.0 882750.0 130800.0 881550.0 ;
      RECT  132000.0 891450.0 133200.0 890250.0 ;
      RECT  133200.0 886200.0 132000.0 885000.0 ;
      RECT  112050.0 886200.0 113250.0 887400.0 ;
      RECT  114000.0 888600.0 115200.0 889800.0 ;
      RECT  130800.0 887700.0 129600.0 888900.0 ;
      RECT  129750.0 900750.0 130650.0 901650.0 ;
      RECT  132150.0 900750.0 133050.0 901650.0 ;
      RECT  129750.0 901200.0 130650.0 904050.0 ;
      RECT  130200.0 900750.0 132600.0 901650.0 ;
      RECT  132150.0 896550.0 133050.0 901200.0 ;
      RECT  129600.0 904050.0 130800.0 905250.0 ;
      RECT  132000.0 895350.0 133200.0 896550.0 ;
      RECT  133200.0 900600.0 132000.0 901800.0 ;
      RECT  112050.0 899400.0 113250.0 900600.0 ;
      RECT  114000.0 897000.0 115200.0 898200.0 ;
      RECT  130800.0 897900.0 129600.0 899100.0 ;
      RECT  129750.0 913650.0 130650.0 912750.0 ;
      RECT  132150.0 913650.0 133050.0 912750.0 ;
      RECT  129750.0 913200.0 130650.0 910350.0 ;
      RECT  130200.0 913650.0 132600.0 912750.0 ;
      RECT  132150.0 917850.0 133050.0 913200.0 ;
      RECT  129600.0 910350.0 130800.0 909150.0 ;
      RECT  132000.0 919050.0 133200.0 917850.0 ;
      RECT  133200.0 913800.0 132000.0 912600.0 ;
      RECT  112050.0 913800.0 113250.0 915000.0 ;
      RECT  114000.0 916200.0 115200.0 917400.0 ;
      RECT  130800.0 915300.0 129600.0 916500.0 ;
      RECT  129750.0 928350.0 130650.0 929250.0 ;
      RECT  132150.0 928350.0 133050.0 929250.0 ;
      RECT  129750.0 928800.0 130650.0 931650.0 ;
      RECT  130200.0 928350.0 132600.0 929250.0 ;
      RECT  132150.0 924150.0 133050.0 928800.0 ;
      RECT  129600.0 931650.0 130800.0 932850.0 ;
      RECT  132000.0 922950.0 133200.0 924150.0 ;
      RECT  133200.0 928200.0 132000.0 929400.0 ;
      RECT  112050.0 927000.0 113250.0 928200.0 ;
      RECT  114000.0 924600.0 115200.0 925800.0 ;
      RECT  130800.0 925500.0 129600.0 926700.0 ;
      RECT  129750.0 941250.0 130650.0 940350.0 ;
      RECT  132150.0 941250.0 133050.0 940350.0 ;
      RECT  129750.0 940800.0 130650.0 937950.0 ;
      RECT  130200.0 941250.0 132600.0 940350.0 ;
      RECT  132150.0 945450.0 133050.0 940800.0 ;
      RECT  129600.0 937950.0 130800.0 936750.0 ;
      RECT  132000.0 946650.0 133200.0 945450.0 ;
      RECT  133200.0 941400.0 132000.0 940200.0 ;
      RECT  112050.0 941400.0 113250.0 942600.0 ;
      RECT  114000.0 943800.0 115200.0 945000.0 ;
      RECT  130800.0 942900.0 129600.0 944100.0 ;
      RECT  129750.0 955950.0 130650.0 956850.0 ;
      RECT  132150.0 955950.0 133050.0 956850.0 ;
      RECT  129750.0 956400.0 130650.0 959250.0 ;
      RECT  130200.0 955950.0 132600.0 956850.0 ;
      RECT  132150.0 951750.0 133050.0 956400.0 ;
      RECT  129600.0 959250.0 130800.0 960450.0 ;
      RECT  132000.0 950550.0 133200.0 951750.0 ;
      RECT  133200.0 955800.0 132000.0 957000.0 ;
      RECT  112050.0 954600.0 113250.0 955800.0 ;
      RECT  114000.0 952200.0 115200.0 953400.0 ;
      RECT  130800.0 953100.0 129600.0 954300.0 ;
      RECT  129750.0 968850.0 130650.0 967950.0 ;
      RECT  132150.0 968850.0 133050.0 967950.0 ;
      RECT  129750.0 968400.0 130650.0 965550.0 ;
      RECT  130200.0 968850.0 132600.0 967950.0 ;
      RECT  132150.0 973050.0 133050.0 968400.0 ;
      RECT  129600.0 965550.0 130800.0 964350.0 ;
      RECT  132000.0 974250.0 133200.0 973050.0 ;
      RECT  133200.0 969000.0 132000.0 967800.0 ;
      RECT  112050.0 969000.0 113250.0 970200.0 ;
      RECT  114000.0 971400.0 115200.0 972600.0 ;
      RECT  130800.0 970500.0 129600.0 971700.0 ;
      RECT  129750.0 983550.0 130650.0 984450.0 ;
      RECT  132150.0 983550.0 133050.0 984450.0 ;
      RECT  129750.0 984000.0 130650.0 986850.0 ;
      RECT  130200.0 983550.0 132600.0 984450.0 ;
      RECT  132150.0 979350.0 133050.0 984000.0 ;
      RECT  129600.0 986850.0 130800.0 988050.0 ;
      RECT  132000.0 978150.0 133200.0 979350.0 ;
      RECT  133200.0 983400.0 132000.0 984600.0 ;
      RECT  112050.0 982200.0 113250.0 983400.0 ;
      RECT  114000.0 979800.0 115200.0 981000.0 ;
      RECT  130800.0 980700.0 129600.0 981900.0 ;
      RECT  129750.0 996450.0 130650.0 995550.0 ;
      RECT  132150.0 996450.0 133050.0 995550.0 ;
      RECT  129750.0 996000.0 130650.0 993150.0 ;
      RECT  130200.0 996450.0 132600.0 995550.0 ;
      RECT  132150.0 1000650.0 133050.0 996000.0 ;
      RECT  129600.0 993150.0 130800.0 991950.0 ;
      RECT  132000.0 1001850.0 133200.0 1000650.0 ;
      RECT  133200.0 996600.0 132000.0 995400.0 ;
      RECT  112050.0 996600.0 113250.0 997800.0 ;
      RECT  114000.0 999000.0 115200.0 1000200.0 ;
      RECT  130800.0 998100.0 129600.0 999300.0 ;
      RECT  129750.0 1011150.0 130650.0 1012050.0 ;
      RECT  132150.0 1011150.0 133050.0 1012050.0 ;
      RECT  129750.0 1011600.0 130650.0 1014450.0 ;
      RECT  130200.0 1011150.0 132600.0 1012050.0 ;
      RECT  132150.0 1006950.0 133050.0 1011600.0 ;
      RECT  129600.0 1014450.0 130800.0 1015650.0 ;
      RECT  132000.0 1005750.0 133200.0 1006950.0 ;
      RECT  133200.0 1011000.0 132000.0 1012200.0 ;
      RECT  112050.0 1009800.0 113250.0 1011000.0 ;
      RECT  114000.0 1007400.0 115200.0 1008600.0 ;
      RECT  130800.0 1008300.0 129600.0 1009500.0 ;
      RECT  129750.0 1024050.0 130650.0 1023150.0 ;
      RECT  132150.0 1024050.0 133050.0 1023150.0 ;
      RECT  129750.0 1023600.0 130650.0 1020750.0 ;
      RECT  130200.0 1024050.0 132600.0 1023150.0 ;
      RECT  132150.0 1028250.0 133050.0 1023600.0 ;
      RECT  129600.0 1020750.0 130800.0 1019550.0 ;
      RECT  132000.0 1029450.0 133200.0 1028250.0 ;
      RECT  133200.0 1024200.0 132000.0 1023000.0 ;
      RECT  112050.0 1024200.0 113250.0 1025400.0 ;
      RECT  114000.0 1026600.0 115200.0 1027800.0 ;
      RECT  130800.0 1025700.0 129600.0 1026900.0 ;
      RECT  129750.0 1038750.0 130650.0 1039650.0 ;
      RECT  132150.0 1038750.0 133050.0 1039650.0 ;
      RECT  129750.0 1039200.0 130650.0 1042050.0 ;
      RECT  130200.0 1038750.0 132600.0 1039650.0 ;
      RECT  132150.0 1034550.0 133050.0 1039200.0 ;
      RECT  129600.0 1042050.0 130800.0 1043250.0 ;
      RECT  132000.0 1033350.0 133200.0 1034550.0 ;
      RECT  133200.0 1038600.0 132000.0 1039800.0 ;
      RECT  112050.0 1037400.0 113250.0 1038600.0 ;
      RECT  114000.0 1035000.0 115200.0 1036200.0 ;
      RECT  130800.0 1035900.0 129600.0 1037100.0 ;
      RECT  129750.0 1051650.0 130650.0 1050750.0 ;
      RECT  132150.0 1051650.0 133050.0 1050750.0 ;
      RECT  129750.0 1051200.0 130650.0 1048350.0 ;
      RECT  130200.0 1051650.0 132600.0 1050750.0 ;
      RECT  132150.0 1055850.0 133050.0 1051200.0 ;
      RECT  129600.0 1048350.0 130800.0 1047150.0 ;
      RECT  132000.0 1057050.0 133200.0 1055850.0 ;
      RECT  133200.0 1051800.0 132000.0 1050600.0 ;
      RECT  112050.0 1051800.0 113250.0 1053000.0 ;
      RECT  114000.0 1054200.0 115200.0 1055400.0 ;
      RECT  130800.0 1053300.0 129600.0 1054500.0 ;
      RECT  129750.0 1066350.0 130650.0 1067250.0 ;
      RECT  132150.0 1066350.0 133050.0 1067250.0 ;
      RECT  129750.0 1066800.0 130650.0 1069650.0 ;
      RECT  130200.0 1066350.0 132600.0 1067250.0 ;
      RECT  132150.0 1062150.0 133050.0 1066800.0 ;
      RECT  129600.0 1069650.0 130800.0 1070850.0 ;
      RECT  132000.0 1060950.0 133200.0 1062150.0 ;
      RECT  133200.0 1066200.0 132000.0 1067400.0 ;
      RECT  112050.0 1065000.0 113250.0 1066200.0 ;
      RECT  114000.0 1062600.0 115200.0 1063800.0 ;
      RECT  130800.0 1063500.0 129600.0 1064700.0 ;
      RECT  129750.0 1079250.0 130650.0 1078350.0 ;
      RECT  132150.0 1079250.0 133050.0 1078350.0 ;
      RECT  129750.0 1078800.0 130650.0 1075950.0 ;
      RECT  130200.0 1079250.0 132600.0 1078350.0 ;
      RECT  132150.0 1083450.0 133050.0 1078800.0 ;
      RECT  129600.0 1075950.0 130800.0 1074750.0 ;
      RECT  132000.0 1084650.0 133200.0 1083450.0 ;
      RECT  133200.0 1079400.0 132000.0 1078200.0 ;
      RECT  112050.0 1079400.0 113250.0 1080600.0 ;
      RECT  114000.0 1081800.0 115200.0 1083000.0 ;
      RECT  130800.0 1080900.0 129600.0 1082100.0 ;
      RECT  129750.0 1093950.0 130650.0 1094850.0 ;
      RECT  132150.0 1093950.0 133050.0 1094850.0 ;
      RECT  129750.0 1094400.0 130650.0 1097250.0 ;
      RECT  130200.0 1093950.0 132600.0 1094850.0 ;
      RECT  132150.0 1089750.0 133050.0 1094400.0 ;
      RECT  129600.0 1097250.0 130800.0 1098450.0 ;
      RECT  132000.0 1088550.0 133200.0 1089750.0 ;
      RECT  133200.0 1093800.0 132000.0 1095000.0 ;
      RECT  112050.0 1092600.0 113250.0 1093800.0 ;
      RECT  114000.0 1090200.0 115200.0 1091400.0 ;
      RECT  130800.0 1091100.0 129600.0 1092300.0 ;
      RECT  129750.0 1106850.0 130650.0 1105950.0 ;
      RECT  132150.0 1106850.0 133050.0 1105950.0 ;
      RECT  129750.0 1106400.0 130650.0 1103550.0 ;
      RECT  130200.0 1106850.0 132600.0 1105950.0 ;
      RECT  132150.0 1111050.0 133050.0 1106400.0 ;
      RECT  129600.0 1103550.0 130800.0 1102350.0 ;
      RECT  132000.0 1112250.0 133200.0 1111050.0 ;
      RECT  133200.0 1107000.0 132000.0 1105800.0 ;
      RECT  112050.0 1107000.0 113250.0 1108200.0 ;
      RECT  114000.0 1109400.0 115200.0 1110600.0 ;
      RECT  130800.0 1108500.0 129600.0 1109700.0 ;
      RECT  129750.0 1121550.0 130650.0 1122450.0 ;
      RECT  132150.0 1121550.0 133050.0 1122450.0 ;
      RECT  129750.0 1122000.0 130650.0 1124850.0 ;
      RECT  130200.0 1121550.0 132600.0 1122450.0 ;
      RECT  132150.0 1117350.0 133050.0 1122000.0 ;
      RECT  129600.0 1124850.0 130800.0 1126050.0 ;
      RECT  132000.0 1116150.0 133200.0 1117350.0 ;
      RECT  133200.0 1121400.0 132000.0 1122600.0 ;
      RECT  112050.0 1120200.0 113250.0 1121400.0 ;
      RECT  114000.0 1117800.0 115200.0 1119000.0 ;
      RECT  130800.0 1118700.0 129600.0 1119900.0 ;
      RECT  129750.0 1134450.0 130650.0 1133550.0 ;
      RECT  132150.0 1134450.0 133050.0 1133550.0 ;
      RECT  129750.0 1134000.0 130650.0 1131150.0 ;
      RECT  130200.0 1134450.0 132600.0 1133550.0 ;
      RECT  132150.0 1138650.0 133050.0 1134000.0 ;
      RECT  129600.0 1131150.0 130800.0 1129950.0 ;
      RECT  132000.0 1139850.0 133200.0 1138650.0 ;
      RECT  133200.0 1134600.0 132000.0 1133400.0 ;
      RECT  112050.0 1134600.0 113250.0 1135800.0 ;
      RECT  114000.0 1137000.0 115200.0 1138200.0 ;
      RECT  130800.0 1136100.0 129600.0 1137300.0 ;
      RECT  129750.0 1149150.0 130650.0 1150050.0 ;
      RECT  132150.0 1149150.0 133050.0 1150050.0 ;
      RECT  129750.0 1149600.0 130650.0 1152450.0 ;
      RECT  130200.0 1149150.0 132600.0 1150050.0 ;
      RECT  132150.0 1144950.0 133050.0 1149600.0 ;
      RECT  129600.0 1152450.0 130800.0 1153650.0 ;
      RECT  132000.0 1143750.0 133200.0 1144950.0 ;
      RECT  133200.0 1149000.0 132000.0 1150200.0 ;
      RECT  112050.0 1147800.0 113250.0 1149000.0 ;
      RECT  114000.0 1145400.0 115200.0 1146600.0 ;
      RECT  130800.0 1146300.0 129600.0 1147500.0 ;
      RECT  129750.0 1162050.0 130650.0 1161150.0 ;
      RECT  132150.0 1162050.0 133050.0 1161150.0 ;
      RECT  129750.0 1161600.0 130650.0 1158750.0 ;
      RECT  130200.0 1162050.0 132600.0 1161150.0 ;
      RECT  132150.0 1166250.0 133050.0 1161600.0 ;
      RECT  129600.0 1158750.0 130800.0 1157550.0 ;
      RECT  132000.0 1167450.0 133200.0 1166250.0 ;
      RECT  133200.0 1162200.0 132000.0 1161000.0 ;
      RECT  112050.0 1162200.0 113250.0 1163400.0 ;
      RECT  114000.0 1164600.0 115200.0 1165800.0 ;
      RECT  130800.0 1163700.0 129600.0 1164900.0 ;
      RECT  129750.0 1176750.0 130650.0 1177650.0 ;
      RECT  132150.0 1176750.0 133050.0 1177650.0 ;
      RECT  129750.0 1177200.0 130650.0 1180050.0 ;
      RECT  130200.0 1176750.0 132600.0 1177650.0 ;
      RECT  132150.0 1172550.0 133050.0 1177200.0 ;
      RECT  129600.0 1180050.0 130800.0 1181250.0 ;
      RECT  132000.0 1171350.0 133200.0 1172550.0 ;
      RECT  133200.0 1176600.0 132000.0 1177800.0 ;
      RECT  112050.0 1175400.0 113250.0 1176600.0 ;
      RECT  114000.0 1173000.0 115200.0 1174200.0 ;
      RECT  130800.0 1173900.0 129600.0 1175100.0 ;
      RECT  129750.0 1189650.0 130650.0 1188750.0 ;
      RECT  132150.0 1189650.0 133050.0 1188750.0 ;
      RECT  129750.0 1189200.0 130650.0 1186350.0 ;
      RECT  130200.0 1189650.0 132600.0 1188750.0 ;
      RECT  132150.0 1193850.0 133050.0 1189200.0 ;
      RECT  129600.0 1186350.0 130800.0 1185150.0 ;
      RECT  132000.0 1195050.0 133200.0 1193850.0 ;
      RECT  133200.0 1189800.0 132000.0 1188600.0 ;
      RECT  112050.0 1189800.0 113250.0 1191000.0 ;
      RECT  114000.0 1192200.0 115200.0 1193400.0 ;
      RECT  130800.0 1191300.0 129600.0 1192500.0 ;
      RECT  112200.0 313800.0 113100.0 1197000.0 ;
      RECT  59100.0 142800.0 119100.0 132600.0 ;
      RECT  59100.0 122400.0 119100.0 132600.0 ;
      RECT  59100.0 122400.0 119100.0 112200.0 ;
      RECT  59100.0 102000.0 119100.0 112200.0 ;
      RECT  59100.0 102000.0 119100.0 91800.0 ;
      RECT  59100.0 81600.0 119100.0 91800.0 ;
      RECT  59100.0 81600.0 119100.0 71400.0 ;
      RECT  59100.0 61200.0 119100.0 71400.0 ;
      RECT  116700.0 138300.0 117900.0 135600.0 ;
      RECT  114600.0 141000.0 119100.0 139800.0 ;
      RECT  116700.0 129600.0 117900.0 126900.0 ;
      RECT  114600.0 125400.0 119100.0 124200.0 ;
      RECT  116700.0 117900.0 117900.0 115200.0 ;
      RECT  114600.0 120600.0 119100.0 119400.0 ;
      RECT  116700.0 109200.0 117900.0 106500.0 ;
      RECT  114600.0 105000.0 119100.0 103800.0 ;
      RECT  116700.0 97500.0 117900.0 94800.0 ;
      RECT  114600.0 100200.0 119100.0 99000.0 ;
      RECT  116700.0 88800.0 117900.0 86100.0 ;
      RECT  114600.0 84600.0 119100.0 83400.0 ;
      RECT  116700.0 77100.0 117900.0 74400.0 ;
      RECT  114600.0 79800.0 119100.0 78600.0 ;
      RECT  116700.0 68400.0 117900.0 65700.0 ;
      RECT  114600.0 64200.0 119100.0 63000.0 ;
      RECT  59100.0 133200.0 119100.0 132000.0 ;
      RECT  59100.0 112800.0 119100.0 111600.0 ;
      RECT  59100.0 92400.0 119100.0 91200.0 ;
      RECT  59100.0 72000.0 119100.0 70800.0 ;
      RECT  201150.0 79500.0 202350.0 80700.0 ;
      RECT  241950.0 79500.0 243150.0 80700.0 ;
      RECT  282750.0 79500.0 283950.0 80700.0 ;
      RECT  323550.0 79500.0 324750.0 80700.0 ;
      RECT  364350.0 79500.0 365550.0 80700.0 ;
      RECT  405150.0 79500.0 406350.0 80700.0 ;
      RECT  445950.0 79500.0 447150.0 80700.0 ;
      RECT  486750.0 79500.0 487950.0 80700.0 ;
      RECT  204900.0 900.0 206100.0 2100.0 ;
      RECT  245700.0 900.0 246900.0 2100.0 ;
      RECT  286500.0 900.0 287700.0 2100.0 ;
      RECT  327300.0 900.0 328500.0 2100.0 ;
      RECT  368100.0 900.0 369300.0 2100.0 ;
      RECT  408900.0 900.0 410100.0 2100.0 ;
      RECT  449700.0 900.0 450900.0 2100.0 ;
      RECT  490500.0 900.0 491700.0 2100.0 ;
      RECT  172650.0 314400.0 173850.0 313200.0 ;
      RECT  172650.0 342000.0 173850.0 340800.0 ;
      RECT  172650.0 369600.0 173850.0 368400.0 ;
      RECT  172650.0 397200.0 173850.0 396000.0 ;
      RECT  172650.0 424800.0 173850.0 423600.0 ;
      RECT  172650.0 452400.0 173850.0 451200.0 ;
      RECT  172650.0 480000.0 173850.0 478800.0 ;
      RECT  172650.0 507600.0 173850.0 506400.0 ;
      RECT  172650.0 535200.0 173850.0 534000.0 ;
      RECT  172650.0 562800.0 173850.0 561600.0 ;
      RECT  172650.0 590400.0 173850.0 589200.0 ;
      RECT  172650.0 618000.0 173850.0 616800.0 ;
      RECT  172650.0 645600.0 173850.0 644400.0 ;
      RECT  172650.0 673200.0 173850.0 672000.0 ;
      RECT  172650.0 700800.0 173850.0 699600.0 ;
      RECT  172650.0 728400.0 173850.0 727200.0 ;
      RECT  172650.0 756000.0 173850.0 754800.0 ;
      RECT  172650.0 783600.0 173850.0 782400.0 ;
      RECT  172650.0 811200.0 173850.0 810000.0 ;
      RECT  172650.0 838800.0 173850.0 837600.0 ;
      RECT  172650.0 866400.0 173850.0 865200.0 ;
      RECT  172650.0 894000.0 173850.0 892800.0 ;
      RECT  172650.0 921600.0 173850.0 920400.0 ;
      RECT  172650.0 949200.0 173850.0 948000.0 ;
      RECT  172650.0 976800.0 173850.0 975600.0 ;
      RECT  172650.0 1004400.0 173850.0 1003200.0 ;
      RECT  172650.0 1032000.0 173850.0 1030800.0 ;
      RECT  172650.0 1059600.0 173850.0 1058400.0 ;
      RECT  172650.0 1087200.0 173850.0 1086000.0 ;
      RECT  172650.0 1114800.0 173850.0 1113600.0 ;
      RECT  172650.0 1142400.0 173850.0 1141200.0 ;
      RECT  172650.0 1170000.0 173850.0 1168800.0 ;
      RECT  172650.0 1197600.0 173850.0 1196400.0 ;
      RECT  138900.0 150450.0 137700.0 151650.0 ;
      RECT  144000.0 150300.0 142800.0 151500.0 ;
      RECT  135900.0 164250.0 134700.0 165450.0 ;
      RECT  146700.0 164100.0 145500.0 165300.0 ;
      RECT  138900.0 205650.0 137700.0 206850.0 ;
      RECT  149400.0 205500.0 148200.0 206700.0 ;
      RECT  135900.0 219450.0 134700.0 220650.0 ;
      RECT  152100.0 219300.0 150900.0 220500.0 ;
      RECT  138900.0 260850.0 137700.0 262050.0 ;
      RECT  154800.0 260700.0 153600.0 261900.0 ;
      RECT  135900.0 274650.0 134700.0 275850.0 ;
      RECT  157500.0 274500.0 156300.0 275700.0 ;
      RECT  141000.0 147600.0 139800.0 148800.0 ;
      RECT  141000.0 147600.0 139800.0 148800.0 ;
      RECT  172050.0 148800.0 173250.0 147600.0 ;
      RECT  141000.0 175200.0 139800.0 176400.0 ;
      RECT  141000.0 175200.0 139800.0 176400.0 ;
      RECT  172050.0 176400.0 173250.0 175200.0 ;
      RECT  141000.0 202800.0 139800.0 204000.0 ;
      RECT  141000.0 202800.0 139800.0 204000.0 ;
      RECT  172050.0 204000.0 173250.0 202800.0 ;
      RECT  141000.0 230400.0 139800.0 231600.0 ;
      RECT  141000.0 230400.0 139800.0 231600.0 ;
      RECT  172050.0 231600.0 173250.0 230400.0 ;
      RECT  141000.0 258000.0 139800.0 259200.0 ;
      RECT  141000.0 258000.0 139800.0 259200.0 ;
      RECT  172050.0 259200.0 173250.0 258000.0 ;
      RECT  141000.0 285600.0 139800.0 286800.0 ;
      RECT  141000.0 285600.0 139800.0 286800.0 ;
      RECT  172050.0 286800.0 173250.0 285600.0 ;
      RECT  160200.0 285750.0 159000.0 286950.0 ;
      RECT  162900.0 283650.0 161700.0 284850.0 ;
      RECT  165600.0 281550.0 164400.0 282750.0 ;
      RECT  168300.0 279450.0 167100.0 280650.0 ;
      RECT  160200.0 6600.0 159000.0 7800.0 ;
      RECT  162900.0 21000.0 161700.0 22200.0 ;
      RECT  165600.0 34200.0 164400.0 35400.0 ;
      RECT  168300.0 48600.0 167100.0 49800.0 ;
      RECT  172650.0 1200.0 173850.0 -1.15463194561e-11 ;
      RECT  172650.0 28800.0 173850.0 27600.0 ;
      RECT  172650.0 56400.0 173850.0 55200.0 ;
      RECT  118500.0 75150.0 117300.0 76350.0 ;
      RECT  78750.0 53400.0 79950.0 54600.0 ;
      RECT  118500.0 66450.0 117300.0 67650.0 ;
      RECT  81750.0 53400.0 82950.0 54600.0 ;
      RECT  118500.0 136350.0 117300.0 137550.0 ;
      RECT  144000.0 136350.0 142800.0 137550.0 ;
      RECT  118500.0 127650.0 117300.0 128850.0 ;
      RECT  146700.0 127650.0 145500.0 128850.0 ;
      RECT  118500.0 115950.0 117300.0 117150.0 ;
      RECT  149400.0 115950.0 148200.0 117150.0 ;
      RECT  118500.0 107250.0 117300.0 108450.0 ;
      RECT  152100.0 107250.0 150900.0 108450.0 ;
      RECT  118500.0 95550.0 117300.0 96750.0 ;
      RECT  154800.0 95550.0 153600.0 96750.0 ;
      RECT  118500.0 86850.0 117300.0 88050.0 ;
      RECT  157500.0 86850.0 156300.0 88050.0 ;
      RECT  120300.0 132000.0 119100.0 133200.0 ;
      RECT  173850.0 132150.0 172650.0 133350.0 ;
      RECT  120300.0 111600.0 119100.0 112800.0 ;
      RECT  173850.0 111750.0 172650.0 112950.0 ;
      RECT  120300.0 91200.0 119100.0 92400.0 ;
      RECT  173850.0 91350.0 172650.0 92550.0 ;
      RECT  120300.0 70800.0 119100.0 72000.0 ;
      RECT  173850.0 70950.0 172650.0 72150.0 ;
      RECT  189000.0 105900.0 187800.0 107100.0 ;
      RECT  183600.0 101400.0 182400.0 102600.0 ;
      RECT  186300.0 99000.0 185100.0 100200.0 ;
      RECT  189000.0 1205250.0 187800.0 1206450.0 ;
      RECT  191700.0 170700.0 190500.0 171900.0 ;
      RECT  194400.0 268800.0 193200.0 270000.0 ;
      RECT  180900.0 144300.0 179700.0 145500.0 ;
      RECT  113250.0 1198500.0 112050.0 1199700.0 ;
      RECT  180900.0 1198500.0 179700.0 1199700.0 ;
      RECT  177150.0 97050.0 175950.0 98250.0 ;
      RECT  177150.0 266850.0 175950.0 268050.0 ;
      RECT  177150.0 168750.0 175950.0 169950.0 ;
      RECT  204600.0 600.0 205500.0 2400.0 ;
      RECT  245400.0 600.0 246300.0 2400.0 ;
      RECT  286200.0 600.0 287100.0 2400.0 ;
      RECT  327000.0 600.0 327900.0 2400.0 ;
      RECT  367800.0 600.0 368700.0 2400.0 ;
      RECT  408600.0 600.0 409500.0 2400.0 ;
      RECT  449400.0 600.0 450300.0 2400.0 ;
      RECT  490200.0 600.0 491100.0 2400.0 ;
      RECT  193350.0 600.0 194250.0 1217400.0 ;
      RECT  190650.0 600.0 191550.0 1217400.0 ;
      RECT  182550.0 600.0 183450.0 1217400.0 ;
      RECT  185250.0 600.0 186150.0 1217400.0 ;
      RECT  187950.0 600.0 188850.0 1217400.0 ;
      RECT  179850.0 600.0 180750.0 1217400.0 ;
      RECT  172650.0 600.0 177150.0 1217400.0 ;
      RECT  49800.0 404400.0 1.42108547152e-11 405300.0 ;
      RECT  49800.0 407100.0 1.42108547152e-11 408000.0 ;
      RECT  49800.0 409800.0 1.42108547152e-11 410700.0 ;
      RECT  49800.0 415200.0 1.42108547152e-11 416100.0 ;
      RECT  43350.0 358050.0 36000.0 358950.0 ;
      RECT  33750.0 319650.0 32850.0 399450.0 ;
      RECT  49800.0 401700.0 47100.0 402600.0 ;
      RECT  38700.0 412500.0 36000.0 413400.0 ;
      RECT  24900.0 401700.0 22200.0 402600.0 ;
      RECT  11100.0 412500.0 8400.0 413400.0 ;
      RECT  7.1054273576e-12 316800.0 10200.0 376800.0 ;
      RECT  20400.0 316800.0 10200.0 376800.0 ;
      RECT  20400.0 316800.0 30600.0 376800.0 ;
      RECT  4500.0 374400.0 7200.0 375600.0 ;
      RECT  1800.0 372300.0 3000.0 376800.0 ;
      RECT  13200.0 374400.0 15900.0 375600.0 ;
      RECT  17400.0 372300.0 18600.0 376800.0 ;
      RECT  24900.0 374400.0 27600.0 375600.0 ;
      RECT  22200.0 372300.0 23400.0 376800.0 ;
      RECT  9600.0 316800.0 10800.0 376800.0 ;
      RECT  30000.0 316800.0 31200.0 376800.0 ;
      RECT  46650.0 432450.0 39150.0 433350.0 ;
      RECT  41700.0 427650.0 40800.0 428550.0 ;
      RECT  41700.0 432450.0 40800.0 433350.0 ;
      RECT  41250.0 427650.0 39150.0 428550.0 ;
      RECT  41700.0 428100.0 40800.0 432900.0 ;
      RECT  46650.0 432450.0 41250.0 433350.0 ;
      RECT  39150.0 427500.0 37950.0 428700.0 ;
      RECT  39150.0 432300.0 37950.0 433500.0 ;
      RECT  47850.0 432300.0 46650.0 433500.0 ;
      RECT  41850.0 432300.0 40650.0 433500.0 ;
      RECT  28800.0 430050.0 29700.0 430950.0 ;
      RECT  29250.0 430050.0 32250.0 430950.0 ;
      RECT  28800.0 430500.0 29700.0 431400.0 ;
      RECT  23700.0 430050.0 24600.0 430950.0 ;
      RECT  23700.0 428700.0 24600.0 430500.0 ;
      RECT  24150.0 430050.0 29250.0 430950.0 ;
      RECT  32250.0 429900.0 33450.0 431100.0 ;
      RECT  23550.0 428700.0 24750.0 427500.0 ;
      RECT  28650.0 432000.0 29850.0 430800.0 ;
      RECT  29550.0 444750.0 30450.0 445650.0 ;
      RECT  29550.0 447150.0 30450.0 448050.0 ;
      RECT  30000.0 444750.0 32850.0 445650.0 ;
      RECT  29550.0 445200.0 30450.0 447600.0 ;
      RECT  25350.0 447150.0 30000.0 448050.0 ;
      RECT  32850.0 444600.0 34050.0 445800.0 ;
      RECT  24150.0 447000.0 25350.0 448200.0 ;
      RECT  29400.0 448200.0 30600.0 447000.0 ;
      RECT  19050.0 442050.0 11550.0 442950.0 ;
      RECT  14100.0 437250.0 13200.0 438150.0 ;
      RECT  14100.0 442050.0 13200.0 442950.0 ;
      RECT  13650.0 437250.0 11550.0 438150.0 ;
      RECT  14100.0 437700.0 13200.0 442500.0 ;
      RECT  19050.0 442050.0 13650.0 442950.0 ;
      RECT  11550.0 437100.0 10350.0 438300.0 ;
      RECT  11550.0 441900.0 10350.0 443100.0 ;
      RECT  20250.0 441900.0 19050.0 443100.0 ;
      RECT  14250.0 441900.0 13050.0 443100.0 ;
      RECT  3000.0 377400.0 1800.0 376200.0 ;
      RECT  3000.0 416250.0 1800.0 415050.0 ;
      RECT  6450.0 376200.0 5250.0 375000.0 ;
      RECT  6450.0 405450.0 5250.0 404250.0 ;
      RECT  18600.0 377400.0 17400.0 376200.0 ;
      RECT  18600.0 408150.0 17400.0 406950.0 ;
      RECT  23400.0 377400.0 22200.0 376200.0 ;
      RECT  23400.0 410850.0 22200.0 409650.0 ;
      RECT  10800.0 377400.0 9600.0 376200.0 ;
      RECT  10800.0 402750.0 9600.0 401550.0 ;
      RECT  31200.0 377400.0 30000.0 376200.0 ;
      RECT  31200.0 402750.0 30000.0 401550.0 ;
      RECT  22650.0 486300.0 21750.0 696300.0 ;
      RECT  17250.0 486300.0 16350.0 691500.0 ;
      RECT  7050.0 486300.0 6150.0 691500.0 ;
      RECT  20400.0 490500.0 19500.0 498600.0 ;
      RECT  13650.0 490500.0 12750.0 495300.0 ;
      RECT  42750.0 530100.0 43650.0 537300.0 ;
      RECT  42750.0 537300.0 43650.0 546900.0 ;
      RECT  42750.0 546900.0 43650.0 556500.0 ;
      RECT  42750.0 558900.0 43650.0 566100.0 ;
      RECT  42750.0 566100.0 43650.0 575700.0 ;
      RECT  42750.0 575700.0 43650.0 585300.0 ;
      RECT  35550.0 587250.0 36450.0 588150.0 ;
      RECT  35550.0 578850.0 36450.0 579750.0 ;
      RECT  36000.0 587250.0 43200.0 588150.0 ;
      RECT  35550.0 579300.0 36450.0 587700.0 ;
      RECT  28800.0 578850.0 36000.0 579750.0 ;
      RECT  28350.0 569700.0 29250.0 579300.0 ;
      RECT  28350.0 560100.0 29250.0 569700.0 ;
      RECT  28350.0 550500.0 29250.0 557700.0 ;
      RECT  28350.0 540900.0 29250.0 550500.0 ;
      RECT  28350.0 531300.0 29250.0 540900.0 ;
      RECT  42600.0 536700.0 43800.0 537900.0 ;
      RECT  42600.0 546300.0 43800.0 547500.0 ;
      RECT  42600.0 555900.0 43800.0 557100.0 ;
      RECT  42600.0 565500.0 43800.0 566700.0 ;
      RECT  42600.0 575100.0 43800.0 576300.0 ;
      RECT  42600.0 584700.0 43800.0 585900.0 ;
      RECT  28200.0 578700.0 29400.0 579900.0 ;
      RECT  28200.0 569100.0 29400.0 570300.0 ;
      RECT  28200.0 559500.0 29400.0 560700.0 ;
      RECT  28200.0 549900.0 29400.0 551100.0 ;
      RECT  28200.0 540300.0 29400.0 541500.0 ;
      RECT  28200.0 530700.0 29400.0 531900.0 ;
      RECT  42600.0 529500.0 43800.0 530700.0 ;
      RECT  42600.0 558300.0 43800.0 559500.0 ;
      RECT  42600.0 587100.0 43800.0 588300.0 ;
      RECT  28200.0 557100.0 29400.0 558300.0 ;
      RECT  16800.0 509700.0 6600.0 495900.0 ;
      RECT  16800.0 509700.0 6600.0 523500.0 ;
      RECT  16800.0 537300.0 6600.0 523500.0 ;
      RECT  16800.0 537300.0 6600.0 551100.0 ;
      RECT  16800.0 564900.0 6600.0 551100.0 ;
      RECT  16800.0 564900.0 6600.0 578700.0 ;
      RECT  16800.0 592500.0 6600.0 578700.0 ;
      RECT  16800.0 592500.0 6600.0 606300.0 ;
      RECT  16800.0 620100.0 6600.0 606300.0 ;
      RECT  16800.0 620100.0 6600.0 633900.0 ;
      RECT  16800.0 647700.0 6600.0 633900.0 ;
      RECT  16800.0 647700.0 6600.0 661500.0 ;
      RECT  16800.0 675300.0 6600.0 661500.0 ;
      RECT  16800.0 675300.0 6600.0 689100.0 ;
      RECT  13800.0 510300.0 12600.0 692700.0 ;
      RECT  10800.0 509100.0 9600.0 691500.0 ;
      RECT  17400.0 509100.0 16200.0 691500.0 ;
      RECT  7200.0 509100.0 6000.0 691500.0 ;
      RECT  22350.0 511200.0 21150.0 512400.0 ;
      RECT  22350.0 534600.0 21150.0 535800.0 ;
      RECT  22350.0 538800.0 21150.0 540000.0 ;
      RECT  22350.0 562200.0 21150.0 563400.0 ;
      RECT  22350.0 566400.0 21150.0 567600.0 ;
      RECT  22350.0 589800.0 21150.0 591000.0 ;
      RECT  22350.0 594000.0 21150.0 595200.0 ;
      RECT  22350.0 617400.0 21150.0 618600.0 ;
      RECT  22350.0 621600.0 21150.0 622800.0 ;
      RECT  22350.0 645000.0 21150.0 646200.0 ;
      RECT  22350.0 649200.0 21150.0 650400.0 ;
      RECT  22350.0 672600.0 21150.0 673800.0 ;
      RECT  22350.0 676800.0 21150.0 678000.0 ;
      RECT  22200.0 524700.0 21000.0 525900.0 ;
      RECT  22800.0 485100.0 21600.0 486300.0 ;
      RECT  16200.0 485700.0 17400.0 486900.0 ;
      RECT  6000.0 485700.0 7200.0 486900.0 ;
      RECT  19350.0 498000.0 20550.0 499200.0 ;
      RECT  19350.0 489900.0 20550.0 491100.0 ;
      RECT  12600.0 489900.0 13800.0 491100.0 ;
      RECT  43950.0 400050.0 42750.0 398850.0 ;
      RECT  43950.0 359100.0 42750.0 357900.0 ;
      RECT  36600.0 359100.0 35400.0 357900.0 ;
      RECT  36600.0 418950.0 35400.0 417750.0 ;
      RECT  33900.0 320250.0 32700.0 319050.0 ;
      RECT  29850.0 400050.0 28650.0 398850.0 ;
      RECT  27150.0 405450.0 25950.0 404250.0 ;
      RECT  30600.0 442800.0 29400.0 441600.0 ;
      RECT  30600.0 442800.0 29400.0 441600.0 ;
      RECT  30600.0 418950.0 29400.0 417750.0 ;
      RECT  27900.0 445800.0 26700.0 444600.0 ;
      RECT  27900.0 445800.0 26700.0 444600.0 ;
      RECT  27900.0 416250.0 26700.0 415050.0 ;
      RECT  41850.0 418950.0 40650.0 417750.0 ;
      RECT  43800.0 416250.0 42600.0 415050.0 ;
      RECT  45750.0 408150.0 44550.0 406950.0 ;
      RECT  14250.0 418950.0 13050.0 417750.0 ;
      RECT  16200.0 408150.0 15000.0 406950.0 ;
      RECT  18150.0 410850.0 16950.0 409650.0 ;
      RECT  29850.0 437100.0 28650.0 438300.0 ;
      RECT  30600.0 454200.0 29400.0 455400.0 ;
      RECT  16200.0 476700.0 15000.0 477900.0 ;
      RECT  29400.0 456900.0 28200.0 458100.0 ;
      RECT  50400.0 402750.0 49200.0 401550.0 ;
      RECT  36600.0 413550.0 35400.0 412350.0 ;
      RECT  22800.0 402750.0 21600.0 401550.0 ;
      RECT  9000.0 413550.0 7800.0 412350.0 ;
      RECT  49800.0 457050.0 28800.0 457950.0 ;
      RECT  49800.0 476850.0 15600.0 477750.0 ;
      RECT  49800.0 437250.0 29250.0 438150.0 ;
      RECT  49800.0 454350.0 30000.0 455250.0 ;
      RECT  49800.0 417900.0 1.42108547152e-11 418800.0 ;
      RECT  49800.0 399000.0 1.42108547152e-11 399900.0 ;
      RECT  49800.0 412500.0 1.42108547152e-11 413400.0 ;
      RECT  49800.0 401700.0 1.42108547152e-11 402600.0 ;
      RECT  194400.0 456900.0 193200.0 458100.0 ;
      RECT  49500.0 457050.0 48300.0 458250.0 ;
      RECT  191700.0 476700.0 190500.0 477900.0 ;
      RECT  49500.0 476850.0 48300.0 478050.0 ;
      RECT  186300.0 437100.0 185100.0 438300.0 ;
      RECT  49500.0 437250.0 48300.0 438450.0 ;
      RECT  183600.0 454200.0 182400.0 455400.0 ;
      RECT  49500.0 454350.0 48300.0 455550.0 ;
      RECT  189000.0 417750.0 187800.0 418950.0 ;
      RECT  49500.0 417900.0 48300.0 419100.0 ;
      RECT  180900.0 398850.0 179700.0 400050.0 ;
      RECT  49500.0 399000.0 48300.0 400200.0 ;
      RECT  55650.0 412350.0 54450.0 413550.0 ;
      RECT  175500.0 401550.0 174300.0 402750.0 ;
      RECT  49500.0 401700.0 48300.0 402900.0 ;
   LAYER  metal3 ;
      RECT  49800.0 456750.0 193800.0 458250.0 ;
      RECT  49800.0 476550.0 191100.0 478050.0 ;
      RECT  49800.0 436950.0 185700.0 438450.0 ;
      RECT  49800.0 454050.0 183000.0 455550.0 ;
      RECT  49800.0 417600.0 188400.0 419100.0 ;
      RECT  49800.0 398700.0 180300.0 400200.0 ;
      RECT  49800.0 401400.0 174900.0 402900.0 ;
      RECT  200850.0 79950.0 202350.0 225150.0 ;
      RECT  241650.0 79950.0 243150.0 225150.0 ;
      RECT  282450.0 79950.0 283950.0 225150.0 ;
      RECT  323250.0 79950.0 324750.0 225150.0 ;
      RECT  364050.0 79950.0 365550.0 225150.0 ;
      RECT  404850.0 79950.0 406350.0 225150.0 ;
      RECT  445650.0 79950.0 447150.0 225150.0 ;
      RECT  486450.0 79950.0 487950.0 225150.0 ;
      RECT  204600.0 600.0 206100.0 103650.0 ;
      RECT  245400.0 600.0 246900.0 103650.0 ;
      RECT  286200.0 600.0 287700.0 103650.0 ;
      RECT  327000.0 600.0 328500.0 103650.0 ;
      RECT  367800.0 600.0 369300.0 103650.0 ;
      RECT  408600.0 600.0 410100.0 103650.0 ;
      RECT  449400.0 600.0 450900.0 103650.0 ;
      RECT  490200.0 600.0 491700.0 103650.0 ;
      RECT  140400.0 147450.0 172650.0 148950.0 ;
      RECT  140400.0 175050.0 172650.0 176550.0 ;
      RECT  140400.0 202650.0 172650.0 204150.0 ;
      RECT  140400.0 230250.0 172650.0 231750.0 ;
      RECT  140400.0 257850.0 172650.0 259350.0 ;
      RECT  140400.0 285450.0 172650.0 286950.0 ;
      RECT  78600.0 75000.0 80100.0 76500.0 ;
      RECT  79350.0 75000.0 117900.0 76500.0 ;
      RECT  78600.0 54000.0 80100.0 75750.0 ;
      RECT  81600.0 66300.0 83100.0 67800.0 ;
      RECT  82350.0 66300.0 117900.0 67800.0 ;
      RECT  81600.0 54000.0 83100.0 67050.0 ;
      RECT  200700.0 225150.0 202500.0 226950.0 ;
      RECT  241500.0 225150.0 243300.0 226950.0 ;
      RECT  282300.0 225150.0 284100.0 226950.0 ;
      RECT  323100.0 225150.0 324900.0 226950.0 ;
      RECT  363900.0 225150.0 365700.0 226950.0 ;
      RECT  404700.0 225150.0 406500.0 226950.0 ;
      RECT  445500.0 225150.0 447300.0 226950.0 ;
      RECT  486300.0 225150.0 488100.0 226950.0 ;
      RECT  204300.0 104550.0 206100.0 106350.0 ;
      RECT  245100.0 104550.0 246900.0 106350.0 ;
      RECT  285900.0 104550.0 287700.0 106350.0 ;
      RECT  326700.0 104550.0 328500.0 106350.0 ;
      RECT  367500.0 104550.0 369300.0 106350.0 ;
      RECT  408300.0 104550.0 410100.0 106350.0 ;
      RECT  449100.0 104550.0 450900.0 106350.0 ;
      RECT  489900.0 104550.0 491700.0 106350.0 ;
      RECT  60000.0 138600.0 61800.0 136800.0 ;
      RECT  60000.0 128400.0 61800.0 126600.0 ;
      RECT  60000.0 118200.0 61800.0 116400.0 ;
      RECT  60000.0 108000.0 61800.0 106200.0 ;
      RECT  60000.0 97800.0 61800.0 96000.0 ;
      RECT  60000.0 87600.0 61800.0 85800.0 ;
      RECT  60000.0 77400.0 61800.0 75600.0 ;
      RECT  60000.0 67200.0 61800.0 65400.0 ;
      RECT  200850.0 79200.0 202650.0 81000.0 ;
      RECT  241650.0 79200.0 243450.0 81000.0 ;
      RECT  282450.0 79200.0 284250.0 81000.0 ;
      RECT  323250.0 79200.0 325050.0 81000.0 ;
      RECT  364050.0 79200.0 365850.0 81000.0 ;
      RECT  404850.0 79200.0 406650.0 81000.0 ;
      RECT  445650.0 79200.0 447450.0 81000.0 ;
      RECT  486450.0 79200.0 488250.0 81000.0 ;
      RECT  204600.0 600.0 206400.0 2400.0 ;
      RECT  245400.0 600.0 247200.0 2400.0 ;
      RECT  286200.0 600.0 288000.0 2400.0 ;
      RECT  327000.0 600.0 328800.0 2400.0 ;
      RECT  367800.0 600.0 369600.0 2400.0 ;
      RECT  408600.0 600.0 410400.0 2400.0 ;
      RECT  449400.0 600.0 451200.0 2400.0 ;
      RECT  490200.0 600.0 492000.0 2400.0 ;
      RECT  141300.0 147300.0 139500.0 149100.0 ;
      RECT  171750.0 149100.0 173550.0 147300.0 ;
      RECT  141300.0 174900.0 139500.0 176700.0 ;
      RECT  171750.0 176700.0 173550.0 174900.0 ;
      RECT  141300.0 202500.0 139500.0 204300.0 ;
      RECT  171750.0 204300.0 173550.0 202500.0 ;
      RECT  141300.0 230100.0 139500.0 231900.0 ;
      RECT  171750.0 231900.0 173550.0 230100.0 ;
      RECT  141300.0 257700.0 139500.0 259500.0 ;
      RECT  171750.0 259500.0 173550.0 257700.0 ;
      RECT  141300.0 285300.0 139500.0 287100.0 ;
      RECT  171750.0 287100.0 173550.0 285300.0 ;
      RECT  118800.0 74850.0 117000.0 76650.0 ;
      RECT  78450.0 53100.0 80250.0 54900.0 ;
      RECT  118800.0 66150.0 117000.0 67950.0 ;
      RECT  81450.0 53100.0 83250.0 54900.0 ;
      RECT  52800.0 136800.0 60000.0 138300.0 ;
      RECT  52800.0 126600.0 60000.0 128100.0 ;
      RECT  52800.0 116400.0 60000.0 117900.0 ;
      RECT  52800.0 106200.0 60000.0 107700.0 ;
      RECT  52800.0 96000.0 60000.0 97500.0 ;
      RECT  52800.0 85800.0 60000.0 87300.0 ;
      RECT  52800.0 75600.0 60000.0 77100.0 ;
      RECT  52800.0 65400.0 60000.0 66900.0 ;
      RECT  3150.0 376800.0 1650.0 415650.0 ;
      RECT  6600.0 375600.0 5100.0 404850.0 ;
      RECT  18750.0 376800.0 17250.0 407550.0 ;
      RECT  23550.0 376800.0 22050.0 410250.0 ;
      RECT  10950.0 376800.0 9450.0 402150.0 ;
      RECT  31350.0 376800.0 29850.0 402150.0 ;
      RECT  36750.0 358500.0 35250.0 418350.0 ;
      RECT  30750.0 418350.0 29250.0 442200.0 ;
      RECT  28050.0 415650.0 26550.0 445200.0 ;
      RECT  4200.0 317700.0 6000.0 319500.0 ;
      RECT  14400.0 317700.0 16200.0 319500.0 ;
      RECT  24600.0 317700.0 26400.0 319500.0 ;
      RECT  3300.0 377700.0 1500.0 375900.0 ;
      RECT  3300.0 416550.0 1500.0 414750.0 ;
      RECT  6750.0 376500.0 4950.0 374700.0 ;
      RECT  6750.0 405750.0 4950.0 403950.0 ;
      RECT  18900.0 377700.0 17100.0 375900.0 ;
      RECT  18900.0 408450.0 17100.0 406650.0 ;
      RECT  23700.0 377700.0 21900.0 375900.0 ;
      RECT  23700.0 411150.0 21900.0 409350.0 ;
      RECT  11100.0 377700.0 9300.0 375900.0 ;
      RECT  11100.0 403050.0 9300.0 401250.0 ;
      RECT  31500.0 377700.0 29700.0 375900.0 ;
      RECT  31500.0 403050.0 29700.0 401250.0 ;
      RECT  36900.0 359400.0 35100.0 357600.0 ;
      RECT  36900.0 419250.0 35100.0 417450.0 ;
      RECT  30900.0 443100.0 29100.0 441300.0 ;
      RECT  30900.0 419250.0 29100.0 417450.0 ;
      RECT  28200.0 446100.0 26400.0 444300.0 ;
      RECT  28200.0 416550.0 26400.0 414750.0 ;
      RECT  16200.0 317700.0 14400.0 319500.0 ;
      RECT  26400.0 317700.0 24600.0 319500.0 ;
      RECT  6000.0 317700.0 4200.0 319500.0 ;
      RECT  194700.0 456600.0 192900.0 458400.0 ;
      RECT  49800.0 456750.0 48000.0 458550.0 ;
      RECT  192000.0 476400.0 190200.0 478200.0 ;
      RECT  49800.0 476550.0 48000.0 478350.0 ;
      RECT  186600.0 436800.0 184800.0 438600.0 ;
      RECT  49800.0 436950.0 48000.0 438750.0 ;
      RECT  183900.0 453900.0 182100.0 455700.0 ;
      RECT  49800.0 454050.0 48000.0 455850.0 ;
      RECT  189300.0 417450.0 187500.0 419250.0 ;
      RECT  49800.0 417600.0 48000.0 419400.0 ;
      RECT  181200.0 398550.0 179400.0 400350.0 ;
      RECT  49800.0 398700.0 48000.0 400500.0 ;
      RECT  175800.0 401250.0 174000.0 403050.0 ;
      RECT  49800.0 401400.0 48000.0 403200.0 ;
   END
   END    sram_1rw_8b_256w_1bank_scn3me_subm
END    LIBRARY
