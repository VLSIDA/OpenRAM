VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 215000.0 by 336100.0 ;
END  MacroSite
MACRO sram_2_16_scn4m_subm
   CLASS BLOCK ;
   SIZE 215000.0 BY 336100.0 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN DIN0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  179000.0 51800.0 179800.0 52600.0 ;
      END
   END DIN0[0]
   PIN DIN0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  200800.0 51800.0 201600.00000000003 52600.0 ;
      END
   END DIN0[1]
   PIN ADDR0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  58000.0 264700.0 58800.0 265500.0 ;
      END
   END ADDR0[0]
   PIN ADDR0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  58000.0 286700.0 58800.0 287500.0 ;
      END
   END ADDR0[1]
   PIN ADDR0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  58000.0 304700.0 58800.0 305500.0 ;
      END
   END ADDR0[2]
   PIN ADDR0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  58000.0 326700.0 58800.0 327500.0 ;
      END
   END ADDR0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  10000.0 10000.0 10799.999999999996 10799.999999999996 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  10000.0 32000.0 10799.999999999996 32800.00000000001 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  48500.0 1400.0000000000057 49099.99999999999 11200.000000000004 ;
      END
   END clk0
   PIN DOUT0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal2 ;
         RECT  172000.0 114800.00000000001 172800.0 117800.00000000001 ;
      END
   END DOUT0[0]
   PIN DOUT0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal2 ;
         RECT  178800.0 114800.00000000001 179600.00000000003 117800.00000000001 ;
      END
   END DOUT0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  174400.0 177200.0 175200.0 178000.0 ;
         LAYER metal3 ;
         RECT  181200.0 177200.0 182000.0 178000.0 ;
         LAYER metal3 ;
         RECT  174400.0 195600.00000000003 175200.0 196400.0 ;
         LAYER metal3 ;
         RECT  181200.0 195600.00000000003 182000.0 196400.0 ;
         LAYER metal3 ;
         RECT  174400.0 214000.0 175200.0 214800.0 ;
         LAYER metal3 ;
         RECT  181200.0 214000.0 182000.0 214800.0 ;
         LAYER metal3 ;
         RECT  174400.0 232400.00000000003 175200.0 233200.0 ;
         LAYER metal3 ;
         RECT  181200.0 232400.00000000003 182000.0 233200.0 ;
         LAYER metal3 ;
         RECT  174400.0 250800.0 175200.0 251600.00000000003 ;
         LAYER metal3 ;
         RECT  181200.0 250800.0 182000.0 251600.00000000003 ;
         LAYER metal3 ;
         RECT  174400.0 269200.0 175200.0 270000.0 ;
         LAYER metal3 ;
         RECT  181200.0 269200.0 182000.0 270000.0 ;
         LAYER metal3 ;
         RECT  174400.0 287600.0 175200.0 288400.00000000006 ;
         LAYER metal3 ;
         RECT  181200.0 287600.0 182000.0 288400.00000000006 ;
         LAYER metal3 ;
         RECT  174400.0 306000.0 175200.0 306800.0 ;
         LAYER metal3 ;
         RECT  181200.0 306000.0 182000.0 306800.0 ;
         LAYER metal3 ;
         RECT  174200.0 158000.0 175000.0 158800.0 ;
         LAYER metal3 ;
         RECT  181000.0 158000.0 181800.0 158800.0 ;
         LAYER metal3 ;
         RECT  176900.0 127700.0 177500.0 128300.00000000001 ;
         LAYER metal3 ;
         RECT  183700.0 127700.0 184300.0 128300.00000000001 ;
         LAYER metal3 ;
         RECT  175300.0 76500.0 175900.0 77100.00000000001 ;
         LAYER metal3 ;
         RECT  174700.0 93900.0 175300.0 94500.0 ;
         LAYER metal3 ;
         RECT  182100.00000000003 76500.0 182700.0 77100.00000000001 ;
         LAYER metal3 ;
         RECT  181500.0 93900.0 182100.00000000003 94500.0 ;
         LAYER metal3 ;
         RECT  131300.0 177600.00000000003 132100.0 178400.0 ;
         LAYER metal3 ;
         RECT  131300.0 196000.0 132100.0 196800.0 ;
         LAYER metal3 ;
         RECT  131300.0 214400.00000000003 132100.0 215200.0 ;
         LAYER metal3 ;
         RECT  131300.0 232800.0 132100.0 233600.00000000003 ;
         LAYER metal3 ;
         RECT  131300.0 251200.0 132100.0 252000.0 ;
         LAYER metal3 ;
         RECT  131300.0 269600.0 132100.0 270400.00000000006 ;
         LAYER metal3 ;
         RECT  131300.0 288000.0 132100.0 288800.0 ;
         LAYER metal3 ;
         RECT  131300.0 306400.00000000006 132100.0 307200.0 ;
         LAYER metal3 ;
         RECT  90900.0 177600.00000000003 91700.0 178400.0 ;
         LAYER metal3 ;
         RECT  108300.00000000001 177600.00000000003 109100.0 178400.0 ;
         LAYER metal3 ;
         RECT  90900.0 196000.0 91700.0 196800.0 ;
         LAYER metal3 ;
         RECT  108300.00000000001 196000.0 109100.0 196800.0 ;
         LAYER metal3 ;
         RECT  90900.0 214400.00000000003 91700.0 215200.0 ;
         LAYER metal3 ;
         RECT  108300.00000000001 214400.00000000003 109100.0 215200.0 ;
         LAYER metal3 ;
         RECT  90900.0 232800.0 91700.0 233600.00000000003 ;
         LAYER metal3 ;
         RECT  108300.00000000001 232800.0 109100.0 233600.00000000003 ;
         LAYER metal3 ;
         RECT  158800.0 177700.0 159400.0 178300.0 ;
         LAYER metal3 ;
         RECT  158800.0 196100.00000000003 159400.0 196700.0 ;
         LAYER metal3 ;
         RECT  158800.0 214500.0 159400.0 215100.00000000003 ;
         LAYER metal3 ;
         RECT  158800.0 232900.00000000003 159400.0 233500.0 ;
         LAYER metal3 ;
         RECT  158800.0 251300.0 159400.0 251900.00000000003 ;
         LAYER metal3 ;
         RECT  158800.0 269700.0 159400.0 270300.0 ;
         LAYER metal3 ;
         RECT  158800.0 288100.0 159400.0 288700.0 ;
         LAYER metal3 ;
         RECT  158800.0 306500.0 159400.0 307100.0 ;
         LAYER metal3 ;
         RECT  70400.0 21000.0 71200.0 21799.999999999996 ;
         LAYER metal3 ;
         RECT  70400.0 61000.0 71200.0 61800.00000000001 ;
         LAYER metal3 ;
         RECT  70400.0 101000.0 71200.0 101800.00000000001 ;
         LAYER metal3 ;
         RECT  70400.0 141000.0 71200.0 141800.0 ;
         LAYER metal3 ;
         RECT  33800.0 184300.0 34599.99999999999 185100.00000000003 ;
         LAYER metal3 ;
         RECT  33800.0 202700.0 34599.99999999999 203500.0 ;
         LAYER metal3 ;
         RECT  33800.0 221100.00000000003 34599.99999999999 221900.00000000003 ;
         LAYER metal3 ;
         RECT  33800.0 239500.0 34599.99999999999 240300.0 ;
         LAYER metal3 ;
         RECT  14799.999999999996 184300.0 15599.999999999995 185100.00000000003 ;
         LAYER metal3 ;
         RECT  21199.999999999996 184300.0 22000.0 185100.00000000003 ;
         LAYER metal3 ;
         RECT  14799.999999999996 202700.0 15599.999999999995 203500.0 ;
         LAYER metal3 ;
         RECT  21199.999999999996 202700.0 22000.0 203500.0 ;
         LAYER metal3 ;
         RECT  8399.99999999999 165900.0 9200.000000000004 166700.0 ;
         LAYER metal3 ;
         RECT  33800.0 165900.0 34599.99999999999 166700.0 ;
         LAYER metal3 ;
         RECT  19599.999999999993 170900.0 20400.0 171700.0 ;
         LAYER metal3 ;
         RECT  2000.0 21000.0 2799.9999999999973 21799.999999999996 ;
         LAYER metal3 ;
         RECT  60900.0 275700.0 61700.0 276500.0 ;
         LAYER metal3 ;
         RECT  60900.0 315700.0 61700.0 316500.0 ;
         LAYER metal3 ;
         RECT  181900.0 62800.00000000001 182700.0 63600.0 ;
         LAYER metal3 ;
         RECT  203700.00000000003 62800.00000000001 204500.0 63600.0 ;
         LAYER metal3 ;
         RECT  4799.999999999997 2400.0000000000055 66000.0 3599.9999999999945 ;
         LAYER metal3 ;
         RECT  74400.0 2400.0000000000055 212400.0 3599.9999999999945 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 7200.000000000003 212400.0 8399.999999999998 ;
         LAYER metal3 ;
         RECT  48000.0 12000.0 212400.0 13200.000000000004 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 16799.999999999996 212400.0 18000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 21600.0 212400.0 22799.999999999996 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 26400.0 212400.0 27600.0 ;
         LAYER metal3 ;
         RECT  69600.0 31200.000000000004 212400.0 32400.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 36000.0 39600.0 37200.0 ;
         LAYER metal3 ;
         RECT  57599.99999999999 36000.0 212400.0 37200.0 ;
         LAYER metal3 ;
         RECT  4799.999999999997 40800.0 66000.0 42000.0 ;
         LAYER metal3 ;
         RECT  74400.0 40800.0 176400.0 42000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 45600.0 212400.0 46800.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 50400.00000000001 34800.0 51600.0 ;
         LAYER metal3 ;
         RECT  62400.0 50400.00000000001 212400.0 51600.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 55200.0 212400.0 56400.00000000001 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 60000.0 212400.0 61200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 64800.0 212400.0 66000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 69600.00000000001 212400.0 70800.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 74400.0 212400.0 75600.00000000001 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 79200.0 66000.0 80400.0 ;
         LAYER metal3 ;
         RECT  74400.0 79200.0 212400.0 80400.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 84000.0 169200.0 85200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 88800.00000000001 68400.0 90000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 93600.00000000001 212400.0 94800.00000000001 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 98400.0 171600.00000000003 99600.00000000001 ;
         LAYER metal3 ;
         RECT  182400.0 98400.0 212400.0 99600.00000000001 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 103200.0 212400.0 104400.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 108000.0 212400.0 109200.0 ;
         LAYER metal3 ;
         RECT  62400.0 112800.00000000001 212400.0 114000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 117600.00000000001 212400.0 118800.00000000001 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 122400.0 66000.0 123600.00000000001 ;
         LAYER metal3 ;
         RECT  74400.0 122400.0 212400.0 123600.00000000001 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 127200.0 212400.0 128400.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 132000.0 212400.0 133200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 136800.0 212400.0 138000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 141600.00000000003 174000.0 142800.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 146400.0 212400.0 147600.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 151200.0 68400.0 152400.0 ;
         LAYER metal3 ;
         RECT  172800.0 151200.0 212400.0 152400.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 156000.0 212400.0 157200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 160800.0 66000.0 162000.0 ;
         LAYER metal3 ;
         RECT  74400.0 160800.0 212400.0 162000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 165600.00000000003 212400.0 166800.0 ;
         LAYER metal3 ;
         RECT  40800.0 170400.0 85200.0 171600.00000000003 ;
         LAYER metal3 ;
         RECT  43200.0 175200.0 212400.0 176400.0 ;
         LAYER metal3 ;
         RECT  40800.0 180000.0 70800.0 181200.0 ;
         LAYER metal3 ;
         RECT  88800.0 180000.0 166800.0 181200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 184800.0 85200.0 186000.0 ;
         LAYER metal3 ;
         RECT  163200.0 184800.0 212400.0 186000.0 ;
         LAYER metal3 ;
         RECT  40800.0 189600.00000000003 70800.0 190800.0 ;
         LAYER metal3 ;
         RECT  88800.0 189600.00000000003 166800.0 190800.0 ;
         LAYER metal3 ;
         RECT  43200.0 194400.0 109200.0 195600.00000000003 ;
         LAYER metal3 ;
         RECT  124800.00000000001 194400.0 212400.0 195600.00000000003 ;
         LAYER metal3 ;
         RECT  40800.0 199200.0 166800.0 200400.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 204000.0 85200.0 205200.0 ;
         LAYER metal3 ;
         RECT  163200.0 204000.0 212400.0 205200.0 ;
         LAYER metal3 ;
         RECT  43200.0 208800.0 166800.0 210000.0 ;
         LAYER metal3 ;
         RECT  43200.0 213600.00000000003 73200.0 214800.0 ;
         LAYER metal3 ;
         RECT  127200.0 213600.00000000003 212400.0 214800.0 ;
         LAYER metal3 ;
         RECT  40800.0 218400.00000000003 166800.0 219600.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 223200.0 75600.0 224400.00000000003 ;
         LAYER metal3 ;
         RECT  163200.0 223200.0 212400.0 224400.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 228000.0 34800.0 229200.0 ;
         LAYER metal3 ;
         RECT  43200.0 228000.0 166800.0 229200.0 ;
         LAYER metal3 ;
         RECT  43200.0 232800.0 109200.0 234000.0 ;
         LAYER metal3 ;
         RECT  129600.0 232800.0 212400.0 234000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 237600.00000000003 166800.0 238800.0 ;
         LAYER metal3 ;
         RECT  40800.0 242400.00000000003 85200.0 243600.00000000003 ;
         LAYER metal3 ;
         RECT  163200.0 242400.00000000003 212400.0 243600.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 247200.0 34800.0 248400.00000000003 ;
         LAYER metal3 ;
         RECT  43200.0 247200.0 166800.0 248400.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 252000.0 212400.0 253200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 256800.0 56400.0 258000.0 ;
         LAYER metal3 ;
         RECT  64800.0 256800.0 166800.0 258000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 261600.00000000003 46800.0 262800.0 ;
         LAYER metal3 ;
         RECT  79200.0 261600.00000000003 126000.0 262800.0 ;
         LAYER metal3 ;
         RECT  163200.0 261600.00000000003 212400.0 262800.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 266400.00000000006 63600.0 267600.0 ;
         LAYER metal3 ;
         RECT  79200.0 266400.00000000006 166800.0 267600.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 271200.0 212400.0 272400.00000000006 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 276000.0 212400.0 277200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 280800.0 126000.0 282000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 285600.0 63600.0 286800.0 ;
         LAYER metal3 ;
         RECT  81600.0 285600.0 212400.0 286800.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 290400.00000000006 166800.0 291600.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 295200.0 56400.0 296400.00000000006 ;
         LAYER metal3 ;
         RECT  64800.0 295200.0 126000.0 296400.00000000006 ;
         LAYER metal3 ;
         RECT  163200.0 295200.0 212400.0 296400.00000000006 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 300000.0 166800.0 301200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 304800.0 63600.0 306000.0 ;
         LAYER metal3 ;
         RECT  84000.0 304800.0 212400.0 306000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 309600.0 166800.0 310800.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 314400.00000000006 126000.0 315600.0 ;
         LAYER metal3 ;
         RECT  163200.0 314400.00000000006 212400.0 315600.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 319200.0 212400.0 320400.00000000006 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 324000.0 63600.0 325200.0 ;
         LAYER metal3 ;
         RECT  84000.0 324000.0 212400.0 325200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 328800.0 212400.0 330000.0 ;
         LAYER metal4 ;
         RECT  4799.999999999997 0.0 6000.0 334800.0 ;
         LAYER metal4 ;
         RECT  9599.999999999995 0.0 10799.999999999996 334800.0 ;
         LAYER metal4 ;
         RECT  14399.999999999998 0.0 15599.999999999995 334800.0 ;
         LAYER metal4 ;
         RECT  19199.999999999996 0.0 20400.0 334800.0 ;
         LAYER metal4 ;
         RECT  24000.0 0.0 25199.999999999996 334800.0 ;
         LAYER metal4 ;
         RECT  28799.999999999996 0.0 30000.0 334800.0 ;
         LAYER metal4 ;
         RECT  33599.99999999999 0.0 34800.0 334800.0 ;
         LAYER metal4 ;
         RECT  38400.0 0.0 39600.0 334800.0 ;
         LAYER metal4 ;
         RECT  43200.0 0.0 44400.0 334800.0 ;
         LAYER metal4 ;
         RECT  48000.0 0.0 49200.0 334800.0 ;
         LAYER metal4 ;
         RECT  52800.0 0.0 54000.0 334800.0 ;
         LAYER metal4 ;
         RECT  57599.99999999999 0.0 58800.0 334800.0 ;
         LAYER metal4 ;
         RECT  62400.0 0.0 63600.0 334800.0 ;
         LAYER metal4 ;
         RECT  67200.0 0.0 68400.0 334800.0 ;
         LAYER metal4 ;
         RECT  72000.0 0.0 73200.0 334800.0 ;
         LAYER metal4 ;
         RECT  76800.0 0.0 78000.0 334800.0 ;
         LAYER metal4 ;
         RECT  81600.0 0.0 82800.0 334800.0 ;
         LAYER metal4 ;
         RECT  86400.0 0.0 87600.0 334800.0 ;
         LAYER metal4 ;
         RECT  91200.0 0.0 92400.0 334800.0 ;
         LAYER metal4 ;
         RECT  96000.0 0.0 97200.0 334800.0 ;
         LAYER metal4 ;
         RECT  100800.0 0.0 102000.0 334800.0 ;
         LAYER metal4 ;
         RECT  105600.0 0.0 106800.0 334800.0 ;
         LAYER metal4 ;
         RECT  110400.0 0.0 111600.0 334800.0 ;
         LAYER metal4 ;
         RECT  115200.0 0.0 116400.0 334800.0 ;
         LAYER metal4 ;
         RECT  120000.0 0.0 121200.0 334800.0 ;
         LAYER metal4 ;
         RECT  124800.00000000001 0.0 126000.0 334800.0 ;
         LAYER metal4 ;
         RECT  129600.0 0.0 130800.00000000001 334800.0 ;
         LAYER metal4 ;
         RECT  134400.0 0.0 135600.0 334800.0 ;
         LAYER metal4 ;
         RECT  139200.0 0.0 140400.0 334800.0 ;
         LAYER metal4 ;
         RECT  144000.0 0.0 145200.0 334800.0 ;
         LAYER metal4 ;
         RECT  148800.0 0.0 150000.0 334800.0 ;
         LAYER metal4 ;
         RECT  153600.00000000003 0.0 154800.0 334800.0 ;
         LAYER metal4 ;
         RECT  158400.0 0.0 159600.00000000003 334800.0 ;
         LAYER metal4 ;
         RECT  163200.0 0.0 164400.0 334800.0 ;
         LAYER metal4 ;
         RECT  168000.0 0.0 169200.0 334800.0 ;
         LAYER metal4 ;
         RECT  172800.0 0.0 174000.0 334800.0 ;
         LAYER metal4 ;
         RECT  177600.00000000003 0.0 178800.0 334800.0 ;
         LAYER metal4 ;
         RECT  182400.0 0.0 183600.00000000003 334800.0 ;
         LAYER metal4 ;
         RECT  187200.0 0.0 188400.0 334800.0 ;
         LAYER metal4 ;
         RECT  192000.0 0.0 193200.0 334800.0 ;
         LAYER metal4 ;
         RECT  196800.0 0.0 198000.0 334800.0 ;
         LAYER metal4 ;
         RECT  201600.00000000003 0.0 202800.0 334800.0 ;
         LAYER metal4 ;
         RECT  206400.0 0.0 207600.0 334800.0 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  171000.0 172600.00000000003 171800.0 173400.0 ;
         LAYER metal3 ;
         RECT  177800.0 172600.00000000003 178600.00000000003 173400.0 ;
         LAYER metal3 ;
         RECT  184600.00000000003 172600.00000000003 185400.0 173400.0 ;
         LAYER metal3 ;
         RECT  171000.0 181800.0 171800.0 182600.00000000003 ;
         LAYER metal3 ;
         RECT  177800.0 181800.0 178600.00000000003 182600.00000000003 ;
         LAYER metal3 ;
         RECT  184600.00000000003 181800.0 185400.0 182600.00000000003 ;
         LAYER metal3 ;
         RECT  171000.0 191000.0 171800.0 191800.0 ;
         LAYER metal3 ;
         RECT  177800.0 191000.0 178600.00000000003 191800.0 ;
         LAYER metal3 ;
         RECT  184600.00000000003 191000.0 185400.0 191800.0 ;
         LAYER metal3 ;
         RECT  171000.0 200200.0 171800.0 201000.0 ;
         LAYER metal3 ;
         RECT  177800.0 200200.0 178600.00000000003 201000.0 ;
         LAYER metal3 ;
         RECT  184600.00000000003 200200.0 185400.0 201000.0 ;
         LAYER metal3 ;
         RECT  171000.0 209400.00000000003 171800.0 210200.0 ;
         LAYER metal3 ;
         RECT  177800.0 209400.00000000003 178600.00000000003 210200.0 ;
         LAYER metal3 ;
         RECT  184600.00000000003 209400.00000000003 185400.0 210200.0 ;
         LAYER metal3 ;
         RECT  171000.0 218600.00000000003 171800.0 219400.00000000003 ;
         LAYER metal3 ;
         RECT  177800.0 218600.00000000003 178600.00000000003 219400.00000000003 ;
         LAYER metal3 ;
         RECT  184600.00000000003 218600.00000000003 185400.0 219400.00000000003 ;
         LAYER metal3 ;
         RECT  171000.0 227800.0 171800.0 228600.00000000003 ;
         LAYER metal3 ;
         RECT  177800.0 227800.0 178600.00000000003 228600.00000000003 ;
         LAYER metal3 ;
         RECT  184600.00000000003 227800.0 185400.0 228600.00000000003 ;
         LAYER metal3 ;
         RECT  171000.0 237000.0 171800.0 237800.0 ;
         LAYER metal3 ;
         RECT  177800.0 237000.0 178600.00000000003 237800.0 ;
         LAYER metal3 ;
         RECT  184600.00000000003 237000.0 185400.0 237800.0 ;
         LAYER metal3 ;
         RECT  171000.0 246200.0 171800.0 247000.0 ;
         LAYER metal3 ;
         RECT  177800.0 246200.0 178600.00000000003 247000.0 ;
         LAYER metal3 ;
         RECT  184600.00000000003 246200.0 185400.0 247000.0 ;
         LAYER metal3 ;
         RECT  171000.0 255400.00000000003 171800.0 256200.0 ;
         LAYER metal3 ;
         RECT  177800.0 255400.00000000003 178600.00000000003 256200.0 ;
         LAYER metal3 ;
         RECT  184600.00000000003 255400.00000000003 185400.0 256200.0 ;
         LAYER metal3 ;
         RECT  171000.0 264600.0 171800.0 265400.00000000006 ;
         LAYER metal3 ;
         RECT  177800.0 264600.0 178600.00000000003 265400.00000000006 ;
         LAYER metal3 ;
         RECT  184600.00000000003 264600.0 185400.0 265400.00000000006 ;
         LAYER metal3 ;
         RECT  171000.0 273800.0 171800.0 274600.0 ;
         LAYER metal3 ;
         RECT  177800.0 273800.0 178600.00000000003 274600.0 ;
         LAYER metal3 ;
         RECT  184600.00000000003 273800.0 185400.0 274600.0 ;
         LAYER metal3 ;
         RECT  171000.0 283000.0 171800.0 283800.0 ;
         LAYER metal3 ;
         RECT  177800.0 283000.0 178600.00000000003 283800.0 ;
         LAYER metal3 ;
         RECT  184600.00000000003 283000.0 185400.0 283800.0 ;
         LAYER metal3 ;
         RECT  171000.0 292200.0 171800.0 293000.0 ;
         LAYER metal3 ;
         RECT  177800.0 292200.0 178600.00000000003 293000.0 ;
         LAYER metal3 ;
         RECT  184600.00000000003 292200.0 185400.0 293000.0 ;
         LAYER metal3 ;
         RECT  171000.0 301400.00000000006 171800.0 302200.0 ;
         LAYER metal3 ;
         RECT  177800.0 301400.00000000006 178600.00000000003 302200.0 ;
         LAYER metal3 ;
         RECT  184600.00000000003 301400.00000000006 185400.0 302200.0 ;
         LAYER metal3 ;
         RECT  171000.0 310600.0 171800.0 311400.00000000006 ;
         LAYER metal3 ;
         RECT  177800.0 310600.0 178600.00000000003 311400.00000000006 ;
         LAYER metal3 ;
         RECT  184600.00000000003 310600.0 185400.0 311400.00000000006 ;
         LAYER metal3 ;
         RECT  177900.0 141100.00000000003 178500.0 141700.0 ;
         LAYER metal3 ;
         RECT  184700.0 141100.00000000003 185300.0 141700.0 ;
         LAYER metal3 ;
         RECT  175300.0 83100.00000000001 175900.0 83700.0 ;
         LAYER metal3 ;
         RECT  176700.0 87500.0 177300.0 88100.00000000001 ;
         LAYER metal3 ;
         RECT  176100.00000000003 100900.0 176700.0 101500.0 ;
         LAYER metal3 ;
         RECT  182100.00000000003 83100.00000000001 182700.0 83700.0 ;
         LAYER metal3 ;
         RECT  183500.0 87500.0 184100.00000000003 88100.00000000001 ;
         LAYER metal3 ;
         RECT  182900.0 100900.0 183500.0 101500.0 ;
         LAYER metal3 ;
         RECT  131300.0 168400.0 132100.0 169200.0 ;
         LAYER metal3 ;
         RECT  131300.0 186800.0 132100.0 187600.00000000003 ;
         LAYER metal3 ;
         RECT  131300.0 205200.0 132100.0 206000.0 ;
         LAYER metal3 ;
         RECT  131300.0 223600.00000000003 132100.0 224400.00000000003 ;
         LAYER metal3 ;
         RECT  131300.0 242000.0 132100.0 242800.0 ;
         LAYER metal3 ;
         RECT  131300.0 260400.00000000003 132100.0 261200.0 ;
         LAYER metal3 ;
         RECT  131300.0 278800.0 132100.0 279600.0 ;
         LAYER metal3 ;
         RECT  131300.0 297200.0 132100.0 298000.0 ;
         LAYER metal3 ;
         RECT  131300.0 315600.0 132100.0 316400.00000000006 ;
         LAYER metal3 ;
         RECT  90900.0 168400.0 91700.0 169200.0 ;
         LAYER metal3 ;
         RECT  108300.00000000001 168400.0 109100.0 169200.0 ;
         LAYER metal3 ;
         RECT  90900.0 186800.0 91700.0 187600.00000000003 ;
         LAYER metal3 ;
         RECT  108300.00000000001 186800.0 109100.0 187600.00000000003 ;
         LAYER metal3 ;
         RECT  90900.0 205200.0 91700.0 206000.0 ;
         LAYER metal3 ;
         RECT  108300.00000000001 205200.0 109100.0 206000.0 ;
         LAYER metal3 ;
         RECT  90900.0 223600.00000000003 91700.0 224400.00000000003 ;
         LAYER metal3 ;
         RECT  108300.00000000001 223600.00000000003 109100.0 224400.00000000003 ;
         LAYER metal3 ;
         RECT  90900.0 242000.0 91700.0 242800.0 ;
         LAYER metal3 ;
         RECT  108300.00000000001 242000.0 109100.0 242800.0 ;
         LAYER metal3 ;
         RECT  158800.0 168500.0 159400.0 169100.00000000003 ;
         LAYER metal3 ;
         RECT  158800.0 186900.0 159400.0 187500.0 ;
         LAYER metal3 ;
         RECT  158800.0 205300.0 159400.0 205900.00000000003 ;
         LAYER metal3 ;
         RECT  158800.0 223700.0 159400.0 224300.0 ;
         LAYER metal3 ;
         RECT  158800.0 242100.00000000003 159400.0 242700.0 ;
         LAYER metal3 ;
         RECT  158800.0 260500.0 159400.0 261100.00000000003 ;
         LAYER metal3 ;
         RECT  158800.0 278900.00000000006 159400.0 279500.0 ;
         LAYER metal3 ;
         RECT  158800.0 297300.0 159400.0 297900.00000000006 ;
         LAYER metal3 ;
         RECT  158800.0 315700.0 159400.0 316300.0 ;
         LAYER metal3 ;
         RECT  70400.0 1000.0 71200.0 1799.9999999999973 ;
         LAYER metal3 ;
         RECT  70400.0 41000.0 71200.0 41800.0 ;
         LAYER metal3 ;
         RECT  70400.0 81000.0 71200.0 81800.00000000001 ;
         LAYER metal3 ;
         RECT  70400.0 121000.0 71200.0 121800.00000000001 ;
         LAYER metal3 ;
         RECT  70400.0 161000.0 71200.0 161800.0 ;
         LAYER metal3 ;
         RECT  30400.0 179700.0 31199.999999999996 180500.0 ;
         LAYER metal3 ;
         RECT  37199.99999999999 179700.0 38000.0 180500.0 ;
         LAYER metal3 ;
         RECT  30400.0 188900.0 31199.999999999996 189700.0 ;
         LAYER metal3 ;
         RECT  37199.99999999999 188900.0 38000.0 189700.0 ;
         LAYER metal3 ;
         RECT  30400.0 198100.00000000003 31199.999999999996 198900.00000000003 ;
         LAYER metal3 ;
         RECT  37199.99999999999 198100.00000000003 38000.0 198900.00000000003 ;
         LAYER metal3 ;
         RECT  30400.0 207300.0 31199.999999999996 208100.00000000003 ;
         LAYER metal3 ;
         RECT  37199.99999999999 207300.0 38000.0 208100.00000000003 ;
         LAYER metal3 ;
         RECT  30400.0 216500.0 31199.999999999996 217300.0 ;
         LAYER metal3 ;
         RECT  37199.99999999999 216500.0 38000.0 217300.0 ;
         LAYER metal3 ;
         RECT  30400.0 225700.0 31199.999999999996 226500.0 ;
         LAYER metal3 ;
         RECT  37199.99999999999 225700.0 38000.0 226500.0 ;
         LAYER metal3 ;
         RECT  30400.0 234900.00000000003 31199.999999999996 235700.0 ;
         LAYER metal3 ;
         RECT  37199.99999999999 234900.00000000003 38000.0 235700.0 ;
         LAYER metal3 ;
         RECT  30400.0 244100.00000000003 31199.999999999996 244900.00000000003 ;
         LAYER metal3 ;
         RECT  37199.99999999999 244100.00000000003 38000.0 244900.00000000003 ;
         LAYER metal3 ;
         RECT  14799.999999999996 175100.00000000003 15599.999999999995 175900.0 ;
         LAYER metal3 ;
         RECT  21199.999999999996 175100.00000000003 22000.0 175900.0 ;
         LAYER metal3 ;
         RECT  14799.999999999996 193500.0 15599.999999999995 194300.0 ;
         LAYER metal3 ;
         RECT  21199.999999999996 193500.0 22000.0 194300.0 ;
         LAYER metal3 ;
         RECT  14799.999999999996 211900.00000000003 15599.999999999995 212700.0 ;
         LAYER metal3 ;
         RECT  21199.999999999996 211900.00000000003 22000.0 212700.0 ;
         LAYER metal3 ;
         RECT  30400.0 170500.0 31199.999999999996 171300.0 ;
         LAYER metal3 ;
         RECT  37199.99999999999 170500.0 38000.0 171300.0 ;
         LAYER metal3 ;
         RECT  39800.0 176500.0 40600.0 177300.0 ;
         LAYER metal3 ;
         RECT  39800.0 192100.00000000003 40600.0 192900.0 ;
         LAYER metal3 ;
         RECT  39800.0 194900.0 40600.0 195700.0 ;
         LAYER metal3 ;
         RECT  39800.0 210500.0 40600.0 211300.0 ;
         LAYER metal3 ;
         RECT  39800.0 213300.0 40600.0 214100.00000000003 ;
         LAYER metal3 ;
         RECT  39800.0 228900.00000000003 40600.0 229700.0 ;
         LAYER metal3 ;
         RECT  39800.0 231700.0 40600.0 232500.0 ;
         LAYER metal3 ;
         RECT  39800.0 247300.0 40600.0 248100.00000000003 ;
         LAYER metal3 ;
         RECT  2000.0 1000.0 2799.9999999999973 1799.9999999999973 ;
         LAYER metal3 ;
         RECT  2000.0 41000.0 2799.9999999999973 41800.0 ;
         LAYER metal3 ;
         RECT  60900.0 255700.0 61700.0 256500.0 ;
         LAYER metal3 ;
         RECT  60900.0 295700.0 61700.0 296500.0 ;
         LAYER metal3 ;
         RECT  60900.0 335700.0 61700.0 336500.0 ;
         LAYER metal3 ;
         RECT  181900.0 42800.0 182700.0 43600.0 ;
         LAYER metal3 ;
         RECT  203700.00000000003 42800.0 204500.0 43600.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 4799.999999999997 212400.0 6000.0 ;
         LAYER metal3 ;
         RECT  60000.0 9600.000000000002 212400.0 10799.999999999996 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 14399.999999999998 212400.0 15600.000000000002 ;
         LAYER metal3 ;
         RECT  4799.999999999997 19200.000000000004 66000.0 20400.0 ;
         LAYER metal3 ;
         RECT  74400.0 19200.000000000004 212400.0 20400.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 24000.0 212400.0 25200.000000000004 ;
         LAYER metal3 ;
         RECT  43200.0 28799.999999999996 212400.0 30000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 33600.0 30000.0 34800.00000000001 ;
         LAYER metal3 ;
         RECT  45599.99999999999 33600.0 212400.0 34800.00000000001 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 38400.00000000001 212400.0 39600.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 43200.0 212400.0 44400.00000000001 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 48000.0 68400.0 49200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 52800.0 212400.0 54000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 57600.0 212400.0 58800.00000000001 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 62400.00000000001 66000.0 63600.0 ;
         LAYER metal3 ;
         RECT  74400.0 62400.00000000001 178800.0 63600.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 67200.0 212400.0 68400.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 72000.0 68400.0 73200.0 ;
         LAYER metal3 ;
         RECT  170400.0 72000.0 212400.0 73200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 76800.0 169200.0 78000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 81600.00000000001 212400.0 82800.00000000001 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 86400.0 212400.0 87600.00000000001 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 91200.0 68400.0 92400.0 ;
         LAYER metal3 ;
         RECT  172800.0 91200.0 212400.0 92400.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 96000.0 212400.0 97200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 100800.00000000001 66000.0 102000.0 ;
         LAYER metal3 ;
         RECT  74400.0 100800.00000000001 212400.0 102000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 105600.0 212400.0 106800.00000000001 ;
         LAYER metal3 ;
         RECT  62400.0 110400.0 212400.0 111600.00000000001 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 115200.0 212400.0 116400.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 120000.0 212400.0 121200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 124800.00000000001 212400.0 126000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 129600.00000000003 68400.0 130800.00000000001 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 134400.0 212400.0 135600.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 139200.0 66000.0 140400.0 ;
         LAYER metal3 ;
         RECT  74400.0 139200.0 212400.0 140400.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 144000.0 212400.0 145200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 148800.0 212400.0 150000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 153600.00000000003 212400.0 154800.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 158400.0 169200.0 159600.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 163200.0 212400.0 164400.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 168000.0 212400.0 169200.0 ;
         LAYER metal3 ;
         RECT  24000.0 172800.0 212400.0 174000.0 ;
         LAYER metal3 ;
         RECT  26400.0 177600.00000000003 70800.0 178800.0 ;
         LAYER metal3 ;
         RECT  36000.0 182400.0 212400.0 183600.00000000003 ;
         LAYER metal3 ;
         RECT  26400.0 187200.0 70800.0 188400.0 ;
         LAYER metal3 ;
         RECT  122400.0 187200.0 212400.0 188400.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 192000.0 212400.0 193200.0 ;
         LAYER metal3 ;
         RECT  26400.0 196800.0 85200.0 198000.0 ;
         LAYER metal3 ;
         RECT  36000.0 201600.00000000003 212400.0 202800.0 ;
         LAYER metal3 ;
         RECT  26400.0 206400.00000000003 109200.0 207600.00000000003 ;
         LAYER metal3 ;
         RECT  124800.00000000001 206400.00000000003 212400.0 207600.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 211200.0 212400.0 212400.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 216000.0 73200.0 217200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 220800.0 30000.0 222000.0 ;
         LAYER metal3 ;
         RECT  36000.0 220800.0 212400.0 222000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 225600.00000000003 75600.0 226800.0 ;
         LAYER metal3 ;
         RECT  88800.0 225600.00000000003 212400.0 226800.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 230400.00000000003 85200.0 231600.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 235200.0 212400.0 236400.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 240000.0 30000.0 241200.0 ;
         LAYER metal3 ;
         RECT  36000.0 240000.0 212400.0 241200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 244800.0 212400.0 246000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 249600.00000000003 126000.0 250800.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 254400.00000000003 212400.0 255600.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 259200.0 46800.0 260400.00000000003 ;
         LAYER metal3 ;
         RECT  79200.0 259200.0 212400.0 260400.00000000003 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 264000.0 63600.0 265200.0 ;
         LAYER metal3 ;
         RECT  79200.0 264000.0 212400.0 265200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 268800.0 126000.0 270000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 273600.0 56400.0 274800.0 ;
         LAYER metal3 ;
         RECT  64800.0 273600.0 212400.0 274800.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 278400.00000000006 212400.0 279600.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 283200.0 212400.0 284400.00000000006 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 288000.0 126000.0 289200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 292800.0 212400.0 294000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 297600.0 212400.0 298800.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 302400.00000000006 212400.0 303600.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 307200.0 126000.0 308400.00000000006 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 312000.0 212400.0 313200.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 316800.0 56400.0 318000.0 ;
         LAYER metal3 ;
         RECT  64800.0 316800.0 212400.0 318000.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 321600.0 212400.0 322800.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 326400.0 63600.0 327600.0 ;
         LAYER metal3 ;
         RECT  84000.0 326400.0 212400.0 327600.0 ;
         LAYER metal3 ;
         RECT  2399.9999999999914 331200.0 212400.0 332400.0 ;
         LAYER metal4 ;
         RECT  7200.000000000003 0.0 8399.99999999999 334800.0 ;
         LAYER metal4 ;
         RECT  12000.0 0.0 13199.999999999996 334800.0 ;
         LAYER metal4 ;
         RECT  16799.999999999996 0.0 18000.0 334800.0 ;
         LAYER metal4 ;
         RECT  21599.999999999993 0.0 22799.999999999996 334800.0 ;
         LAYER metal4 ;
         RECT  26400.0 0.0 27599.999999999993 334800.0 ;
         LAYER metal4 ;
         RECT  31199.999999999996 0.0 32400.0 334800.0 ;
         LAYER metal4 ;
         RECT  36000.0 0.0 37199.99999999999 334800.0 ;
         LAYER metal4 ;
         RECT  40800.0 0.0 42000.0 334800.0 ;
         LAYER metal4 ;
         RECT  45599.99999999999 0.0 46800.0 334800.0 ;
         LAYER metal4 ;
         RECT  50400.0 0.0 51599.99999999999 334800.0 ;
         LAYER metal4 ;
         RECT  55200.0 0.0 56400.0 334800.0 ;
         LAYER metal4 ;
         RECT  60000.0 0.0 61200.0 334800.0 ;
         LAYER metal4 ;
         RECT  64800.0 0.0 66000.0 334800.0 ;
         LAYER metal4 ;
         RECT  69600.0 0.0 70800.0 334800.0 ;
         LAYER metal4 ;
         RECT  74400.0 0.0 75600.0 334800.0 ;
         LAYER metal4 ;
         RECT  79200.0 0.0 80400.0 334800.0 ;
         LAYER metal4 ;
         RECT  84000.0 0.0 85200.0 334800.0 ;
         LAYER metal4 ;
         RECT  88800.0 0.0 90000.0 334800.0 ;
         LAYER metal4 ;
         RECT  93600.0 0.0 94800.0 334800.0 ;
         LAYER metal4 ;
         RECT  98400.0 0.0 99600.0 334800.0 ;
         LAYER metal4 ;
         RECT  103200.0 0.0 104400.0 334800.0 ;
         LAYER metal4 ;
         RECT  108000.0 0.0 109200.0 334800.0 ;
         LAYER metal4 ;
         RECT  112800.00000000001 0.0 114000.0 334800.0 ;
         LAYER metal4 ;
         RECT  117600.0 0.0 118800.00000000001 334800.0 ;
         LAYER metal4 ;
         RECT  122400.0 0.0 123600.0 334800.0 ;
         LAYER metal4 ;
         RECT  127200.0 0.0 128400.0 334800.0 ;
         LAYER metal4 ;
         RECT  132000.0 0.0 133200.0 334800.0 ;
         LAYER metal4 ;
         RECT  136800.0 0.0 138000.0 334800.0 ;
         LAYER metal4 ;
         RECT  141600.00000000003 0.0 142800.0 334800.0 ;
         LAYER metal4 ;
         RECT  146400.0 0.0 147600.00000000003 334800.0 ;
         LAYER metal4 ;
         RECT  151200.0 0.0 152400.0 334800.0 ;
         LAYER metal4 ;
         RECT  156000.0 0.0 157200.0 334800.0 ;
         LAYER metal4 ;
         RECT  160800.0 0.0 162000.0 334800.0 ;
         LAYER metal4 ;
         RECT  165600.00000000003 0.0 166800.0 334800.0 ;
         LAYER metal4 ;
         RECT  170400.0 0.0 171600.00000000003 334800.0 ;
         LAYER metal4 ;
         RECT  175200.0 0.0 176400.0 334800.0 ;
         LAYER metal4 ;
         RECT  180000.0 0.0 181200.0 334800.0 ;
         LAYER metal4 ;
         RECT  184800.0 0.0 186000.0 334800.0 ;
         LAYER metal4 ;
         RECT  189600.00000000003 0.0 190800.0 334800.0 ;
         LAYER metal4 ;
         RECT  194400.0 0.0 195600.00000000003 334800.0 ;
         LAYER metal4 ;
         RECT  199200.0 0.0 200400.0 334800.0 ;
         LAYER metal4 ;
         RECT  204000.0 0.0 205200.00000000003 334800.0 ;
         LAYER metal4 ;
         RECT  208800.0 0.0 210000.0 334800.0 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  72200.0 10299.999999999996 73600.00000000001 10899.999999999996 ;
      RECT  174800.0 65700.0 190600.00000000003 66300.0 ;
      RECT  181600.00000000003 67100.00000000001 212400.00000000003 67700.0 ;
      RECT  142500.0 172900.0 143100.0 173500.0 ;
      RECT  142500.0 171300.0 143100.0 171900.0 ;
      RECT  140400.0 172900.0 142800.0 173500.0 ;
      RECT  142500.0 171600.00000000003 143100.0 173200.0 ;
      RECT  142800.0 171300.0 145300.0 171900.0 ;
      RECT  166700.0 172900.0 167300.0 173500.0 ;
      RECT  166700.0 169500.0 167300.0 170100.0 ;
      RECT  163000.0 172900.0 167000.0 173500.0 ;
      RECT  166700.0 169800.0 167300.0 173200.00000000003 ;
      RECT  167000.0 169500.0 171000.0 170100.0 ;
      RECT  142500.0 182500.0 143100.0 183100.00000000003 ;
      RECT  142500.0 184100.00000000003 143100.0 184700.0 ;
      RECT  140400.0 182500.0 142800.0 183100.00000000003 ;
      RECT  142500.0 182800.0 143100.0 184400.0 ;
      RECT  142800.0 184100.00000000003 145300.0 184700.0 ;
      RECT  166700.0 182500.0 167300.0 183100.00000000003 ;
      RECT  166700.0 185100.00000000003 167300.0 185700.0 ;
      RECT  163000.0 182500.0 167000.0 183100.00000000003 ;
      RECT  166700.0 182800.0 167300.0 185400.0 ;
      RECT  167000.0 185100.00000000003 171000.0 185700.0 ;
      RECT  142500.0 191300.0 143100.0 191900.0 ;
      RECT  142500.0 189700.0 143100.0 190300.0 ;
      RECT  140400.0 191300.0 142800.0 191900.0 ;
      RECT  142500.0 190000.0 143100.0 191600.00000000003 ;
      RECT  142800.0 189700.0 145300.0 190300.0 ;
      RECT  166700.0 191300.0 167300.0 191900.0 ;
      RECT  166700.0 187900.0 167300.0 188500.0 ;
      RECT  163000.0 191300.0 167000.0 191900.0 ;
      RECT  166700.0 188200.0 167300.0 191600.00000000003 ;
      RECT  167000.0 187900.0 171000.0 188500.0 ;
      RECT  142500.0 200899.99999999997 143100.0 201500.0 ;
      RECT  142500.0 202500.0 143100.0 203100.00000000003 ;
      RECT  140400.0 200899.99999999997 142800.0 201500.0 ;
      RECT  142500.0 201200.0 143100.0 202800.0 ;
      RECT  142800.0 202500.0 145300.0 203100.00000000003 ;
      RECT  166700.0 200899.99999999997 167300.0 201500.0 ;
      RECT  166700.0 203500.0 167300.0 204100.00000000003 ;
      RECT  163000.0 200899.99999999997 167000.0 201500.0 ;
      RECT  166700.0 201200.0 167300.0 203800.0 ;
      RECT  167000.0 203500.0 171000.0 204100.00000000003 ;
      RECT  142500.0 209700.0 143100.0 210300.0 ;
      RECT  142500.0 208100.00000000003 143100.0 208700.0 ;
      RECT  140400.0 209700.0 142800.0 210300.0 ;
      RECT  142500.0 208399.99999999997 143100.0 210000.0 ;
      RECT  142800.0 208100.00000000003 145300.0 208700.0 ;
      RECT  166700.0 209700.0 167300.0 210300.0 ;
      RECT  166700.0 206300.0 167300.0 206899.99999999997 ;
      RECT  163000.0 209700.0 167000.0 210300.0 ;
      RECT  166700.0 206600.00000000003 167300.0 210000.0 ;
      RECT  167000.0 206300.0 171000.0 206899.99999999997 ;
      RECT  142500.0 219300.0 143100.0 219900.00000000003 ;
      RECT  142500.0 220899.99999999997 143100.0 221500.0 ;
      RECT  140400.0 219300.0 142800.0 219900.00000000003 ;
      RECT  142500.0 219600.00000000003 143100.0 221200.0 ;
      RECT  142800.0 220899.99999999997 145300.0 221500.0 ;
      RECT  166700.0 219300.0 167300.0 219900.00000000003 ;
      RECT  166700.0 221899.99999999997 167300.0 222500.0 ;
      RECT  163000.0 219300.0 167000.0 219900.00000000003 ;
      RECT  166700.0 219600.00000000003 167300.0 222200.0 ;
      RECT  167000.0 221899.99999999997 171000.0 222500.0 ;
      RECT  142500.0 228100.00000000003 143100.0 228700.0 ;
      RECT  142500.0 226500.0 143100.0 227100.00000000003 ;
      RECT  140400.0 228100.00000000003 142800.0 228700.0 ;
      RECT  142500.0 226800.0 143100.0 228400.00000000003 ;
      RECT  142800.0 226500.0 145300.0 227100.00000000003 ;
      RECT  166700.0 228100.00000000003 167300.0 228700.0 ;
      RECT  166700.0 224700.0 167300.0 225300.0 ;
      RECT  163000.0 228100.00000000003 167000.0 228700.0 ;
      RECT  166700.0 225000.0 167300.0 228400.00000000003 ;
      RECT  167000.0 224700.0 171000.0 225300.0 ;
      RECT  142500.0 237700.0 143100.0 238300.0 ;
      RECT  142500.0 239300.0 143100.0 239900.00000000003 ;
      RECT  140400.0 237700.0 142800.0 238300.0 ;
      RECT  142500.0 238000.0 143100.0 239600.00000000003 ;
      RECT  142800.0 239300.0 145300.0 239900.00000000003 ;
      RECT  166700.0 237700.0 167300.0 238300.0 ;
      RECT  166700.0 240300.0 167300.0 240900.00000000003 ;
      RECT  163000.0 237700.0 167000.0 238300.0 ;
      RECT  166700.0 238000.0 167300.0 240600.00000000003 ;
      RECT  167000.0 240300.0 171000.0 240900.00000000003 ;
      RECT  142500.0 246500.0 143100.0 247100.00000000003 ;
      RECT  142500.0 244899.99999999997 143100.0 245500.0 ;
      RECT  140400.0 246500.0 142800.0 247100.00000000003 ;
      RECT  142500.0 245200.0 143100.0 246800.0 ;
      RECT  142800.0 244899.99999999997 145300.0 245500.0 ;
      RECT  166700.0 246500.0 167300.0 247100.00000000003 ;
      RECT  166700.0 243100.00000000003 167300.0 243700.0 ;
      RECT  163000.0 246500.0 167000.0 247100.00000000003 ;
      RECT  166700.0 243399.99999999997 167300.0 246800.0 ;
      RECT  167000.0 243100.00000000003 171000.0 243700.0 ;
      RECT  142500.0 256100.00000000003 143100.0 256700.0 ;
      RECT  142500.0 257700.0 143100.0 258300.0 ;
      RECT  140400.0 256100.00000000003 142800.0 256700.0 ;
      RECT  142500.0 256399.99999999997 143100.0 258000.0 ;
      RECT  142800.0 257700.0 145300.0 258300.0 ;
      RECT  166700.0 256100.00000000003 167300.0 256700.0 ;
      RECT  166700.0 258700.0 167300.0 259300.0 ;
      RECT  163000.0 256100.00000000003 167000.0 256700.0 ;
      RECT  166700.0 256399.99999999997 167300.0 259000.0 ;
      RECT  167000.0 258700.0 171000.0 259300.0 ;
      RECT  142500.0 264900.0 143100.0 265500.0 ;
      RECT  142500.0 263300.0 143100.0 263900.00000000006 ;
      RECT  140400.0 264900.0 142800.0 265500.0 ;
      RECT  142500.0 263600.0 143100.0 265200.0 ;
      RECT  142800.0 263300.0 145300.0 263900.00000000006 ;
      RECT  166700.0 264900.0 167300.0 265500.0 ;
      RECT  166700.0 261500.0 167300.0 262100.00000000003 ;
      RECT  163000.0 264900.0 167000.0 265500.0 ;
      RECT  166700.0 261800.0 167300.0 265200.00000000006 ;
      RECT  167000.0 261500.0 171000.0 262100.00000000003 ;
      RECT  142500.0 274500.0 143100.0 275100.0 ;
      RECT  142500.0 276100.0 143100.0 276700.0 ;
      RECT  140400.0 274500.0 142800.0 275100.0 ;
      RECT  142500.0 274800.0 143100.0 276400.00000000006 ;
      RECT  142800.0 276100.0 145300.0 276700.0 ;
      RECT  166700.0 274500.0 167300.0 275100.0 ;
      RECT  166700.0 277100.0 167300.0 277700.0 ;
      RECT  163000.0 274500.0 167000.0 275100.0 ;
      RECT  166700.0 274800.0 167300.0 277400.00000000006 ;
      RECT  167000.0 277100.0 171000.0 277700.0 ;
      RECT  142500.0 283300.0 143100.0 283900.00000000006 ;
      RECT  142500.0 281700.0 143100.0 282300.0 ;
      RECT  140400.0 283300.0 142800.0 283900.00000000006 ;
      RECT  142500.0 282000.0 143100.0 283600.0 ;
      RECT  142800.0 281700.0 145300.0 282300.0 ;
      RECT  166700.0 283300.0 167300.0 283900.00000000006 ;
      RECT  166700.0 279900.0 167300.0 280500.0 ;
      RECT  163000.0 283300.0 167000.0 283900.00000000006 ;
      RECT  166700.0 280200.0 167300.0 283600.0 ;
      RECT  167000.0 279900.0 171000.0 280500.0 ;
      RECT  142500.0 292900.0 143100.0 293500.0 ;
      RECT  142500.0 294500.0 143100.0 295100.0 ;
      RECT  140400.0 292900.0 142800.0 293500.0 ;
      RECT  142500.0 293200.0 143100.0 294800.0 ;
      RECT  142800.0 294500.0 145300.0 295100.0 ;
      RECT  166700.0 292900.0 167300.0 293500.0 ;
      RECT  166700.0 295500.0 167300.0 296100.0 ;
      RECT  163000.0 292900.0 167000.0 293500.0 ;
      RECT  166700.0 293200.0 167300.0 295800.0 ;
      RECT  167000.0 295500.0 171000.0 296100.0 ;
      RECT  142500.0 301700.0 143100.0 302300.0 ;
      RECT  142500.0 300100.0 143100.0 300700.00000000006 ;
      RECT  140400.0 301700.0 142800.0 302300.0 ;
      RECT  142500.0 300400.0 143100.0 302000.0 ;
      RECT  142800.0 300100.0 145300.0 300700.00000000006 ;
      RECT  166700.0 301700.0 167300.0 302300.0 ;
      RECT  166700.0 298300.0 167300.0 298900.00000000006 ;
      RECT  163000.0 301700.0 167000.0 302300.0 ;
      RECT  166700.0 298600.0 167300.0 302000.00000000006 ;
      RECT  167000.0 298300.0 171000.0 298900.00000000006 ;
      RECT  142500.0 311300.0 143100.0 311900.00000000006 ;
      RECT  142500.0 312900.0 143100.0 313500.0 ;
      RECT  140400.0 311300.0 142800.0 311900.00000000006 ;
      RECT  142500.0 311600.0 143100.0 313200.00000000006 ;
      RECT  142800.0 312900.0 145300.0 313500.0 ;
      RECT  166700.0 311300.0 167300.0 311900.00000000006 ;
      RECT  166700.0 313900.0 167300.0 314500.0 ;
      RECT  163000.0 311300.0 167000.0 311900.00000000006 ;
      RECT  166700.0 311600.0 167300.0 314200.00000000006 ;
      RECT  167000.0 313900.0 171000.0 314500.0 ;
      RECT  169700.0 154800.0 171400.0 155399.99999999997 ;
      RECT  166900.0 75000.0 171400.0 75600.0 ;
      RECT  168300.0 144600.00000000003 171400.0 145200.0 ;
      RECT  147400.0 164300.0 165500.0 164900.0 ;
      RECT  171400.0 168400.0 178200.0 177600.00000000003 ;
      RECT  171400.0 186800.0 178200.0 177600.00000000003 ;
      RECT  171400.0 186800.0 178200.0 196000.0 ;
      RECT  171400.0 205200.0 178200.0 196000.0 ;
      RECT  171400.0 205200.0 178200.0 214400.00000000003 ;
      RECT  171400.0 223600.00000000003 178200.0 214399.99999999997 ;
      RECT  171400.0 223600.00000000003 178200.0 232800.0 ;
      RECT  171400.0 242000.0 178200.0 232800.0 ;
      RECT  171400.0 242000.0 178200.0 251200.0 ;
      RECT  171400.0 260399.99999999997 178200.0 251200.0 ;
      RECT  171400.0 260399.99999999997 178200.0 269600.0 ;
      RECT  171400.0 278800.0 178200.0 269600.0 ;
      RECT  171400.0 278800.0 178200.0 288000.0 ;
      RECT  171400.0 297200.0 178200.0 288000.0 ;
      RECT  171400.0 297200.0 178200.0 306400.0 ;
      RECT  171400.0 315600.0 178200.0 306400.00000000006 ;
      RECT  178200.0 168400.0 185000.0 177600.00000000003 ;
      RECT  178200.0 186800.0 185000.0 177600.00000000003 ;
      RECT  178200.0 186800.0 185000.0 196000.0 ;
      RECT  178200.0 205200.0 185000.0 196000.0 ;
      RECT  178200.0 205200.0 185000.0 214400.00000000003 ;
      RECT  178200.0 223600.00000000003 185000.0 214399.99999999997 ;
      RECT  178200.0 223600.00000000003 185000.0 232800.0 ;
      RECT  178200.0 242000.0 185000.0 232800.0 ;
      RECT  178200.0 242000.0 185000.0 251200.0 ;
      RECT  178200.0 260399.99999999997 185000.0 251200.0 ;
      RECT  178200.0 260399.99999999997 185000.0 269600.0 ;
      RECT  178200.0 278800.0 185000.0 269600.0 ;
      RECT  178200.0 278800.0 185000.0 288000.0 ;
      RECT  178200.0 297200.0 185000.0 288000.0 ;
      RECT  178200.0 297200.0 185000.0 306400.0 ;
      RECT  178200.0 315600.0 185000.0 306400.00000000006 ;
      RECT  171000.0 169400.0 185200.0 170200.0 ;
      RECT  171000.0 185000.0 185200.0 185800.0 ;
      RECT  171000.0 187800.0 185200.0 188600.00000000003 ;
      RECT  171000.0 203399.99999999997 185200.0 204200.0 ;
      RECT  171000.0 206200.0 185200.0 207000.0 ;
      RECT  171000.0 221800.0 185200.0 222600.00000000003 ;
      RECT  171000.0 224600.00000000003 185200.0 225399.99999999997 ;
      RECT  171000.0 240200.0 185200.0 241000.0 ;
      RECT  171000.0 243000.0 185200.0 243800.0 ;
      RECT  171000.0 258600.00000000003 185200.0 259399.99999999997 ;
      RECT  171000.0 261399.99999999997 185200.0 262200.0 ;
      RECT  171000.0 277000.0 185200.0 277800.0 ;
      RECT  171000.0 279800.0 185200.0 280600.0 ;
      RECT  171000.0 295400.0 185200.0 296200.0 ;
      RECT  171000.0 298200.0 185200.0 299000.0 ;
      RECT  171000.0 313800.0 185200.0 314600.0 ;
      RECT  171400.0 163900.0 178200.0 164500.0 ;
      RECT  174300.0 158800.0 174900.0 164200.0 ;
      RECT  174600.00000000003 153300.0 176600.00000000003 153900.0 ;
      RECT  176200.0 158100.00000000003 176600.00000000003 158700.0 ;
      RECT  172600.00000000003 153200.0 173400.0 154000.0 ;
      RECT  174200.0 153200.0 175000.0 154000.0 ;
      RECT  174200.0 153200.0 175000.0 154000.0 ;
      RECT  172600.00000000003 153200.0 173400.0 154000.0 ;
      RECT  172600.00000000003 158000.0 173400.0 158800.0 ;
      RECT  174200.0 158000.0 175000.0 158800.0 ;
      RECT  174200.0 158000.0 175000.0 158800.0 ;
      RECT  172600.00000000003 158000.0 173400.0 158800.0 ;
      RECT  174200.0 158000.0 175000.0 158800.0 ;
      RECT  175800.0 158000.0 176600.00000000003 158800.0 ;
      RECT  175800.0 158000.0 176600.00000000003 158800.0 ;
      RECT  174200.0 158000.0 175000.0 158800.0 ;
      RECT  174000.0 154700.0 173200.0 155500.0 ;
      RECT  174200.0 161600.00000000003 175000.0 162400.0 ;
      RECT  174200.0 158000.0 175000.0 158800.0 ;
      RECT  172600.00000000003 158000.0 173400.0 158800.0 ;
      RECT  172600.00000000003 153200.0 173400.0 154000.0 ;
      RECT  176200.0 158000.0 177000.0 158800.0 ;
      RECT  176200.0 153200.0 177000.0 154000.0 ;
      RECT  171400.0 154800.0 178200.0 155400.0 ;
      RECT  178200.0 163900.0 185000.0 164500.0 ;
      RECT  181100.00000000003 158800.0 181700.0 164200.0 ;
      RECT  181400.0 153300.0 183400.0 153900.0 ;
      RECT  183000.0 158100.00000000003 183400.0 158700.0 ;
      RECT  179400.0 153200.0 180200.0 154000.0 ;
      RECT  181000.0 153200.0 181800.0 154000.0 ;
      RECT  181000.0 153200.0 181800.0 154000.0 ;
      RECT  179400.0 153200.0 180200.0 154000.0 ;
      RECT  179400.0 158000.0 180200.0 158800.0 ;
      RECT  181000.0 158000.0 181800.0 158800.0 ;
      RECT  181000.0 158000.0 181800.0 158800.0 ;
      RECT  179400.0 158000.0 180200.0 158800.0 ;
      RECT  181000.0 158000.0 181800.0 158800.0 ;
      RECT  182600.00000000003 158000.0 183400.0 158800.0 ;
      RECT  182600.00000000003 158000.0 183400.0 158800.0 ;
      RECT  181000.0 158000.0 181800.0 158800.0 ;
      RECT  180800.0 154700.0 180000.0 155500.0 ;
      RECT  181000.0 161600.00000000003 181800.0 162400.0 ;
      RECT  181000.0 158000.0 181800.0 158800.0 ;
      RECT  179400.0 158000.0 180200.0 158800.0 ;
      RECT  179400.0 153200.0 180200.0 154000.0 ;
      RECT  183000.0 158000.0 183800.0 158800.0 ;
      RECT  183000.0 153200.0 183800.0 154000.0 ;
      RECT  178200.0 154800.0 185000.0 155400.0 ;
      RECT  171400.0 154800.0 185000.0 155400.0 ;
      RECT  171400.0 114800.00000000001 178200.0 147400.0 ;
      RECT  178200.0 114800.00000000001 185000.0 147400.0 ;
      RECT  171400.0 144600.00000000003 185000.0 145200.0 ;
      RECT  171400.0 70200.0 178200.0 110600.0 ;
      RECT  178200.0 70200.0 185000.0 110600.0 ;
      RECT  171400.0 75000.0 185000.0 75600.00000000001 ;
      RECT  135500.0 173300.0 136100.0 173900.0 ;
      RECT  135500.0 172900.0 136100.0 173500.0 ;
      RECT  133500.0 173300.0 135800.0 173900.0 ;
      RECT  135500.0 173200.0 136100.0 173600.00000000003 ;
      RECT  135800.0 172900.0 138100.0 173500.0 ;
      RECT  135500.0 182100.00000000003 136100.0 182700.0 ;
      RECT  135500.0 182500.0 136100.0 183100.00000000003 ;
      RECT  133500.0 182100.00000000003 135800.0 182700.0 ;
      RECT  135500.0 182400.0 136100.0 182800.0 ;
      RECT  135800.0 182500.0 138100.0 183100.00000000003 ;
      RECT  135500.0 191700.0 136100.0 192300.0 ;
      RECT  135500.0 191300.0 136100.0 191900.0 ;
      RECT  133500.0 191700.0 135800.0 192300.0 ;
      RECT  135500.0 191600.00000000003 136100.0 192000.0 ;
      RECT  135800.0 191300.0 138100.0 191900.0 ;
      RECT  135500.0 200500.0 136100.0 201100.00000000003 ;
      RECT  135500.0 200899.99999999997 136100.0 201500.0 ;
      RECT  133500.0 200500.0 135800.0 201100.00000000003 ;
      RECT  135500.0 200800.0 136100.0 201200.0 ;
      RECT  135800.0 200899.99999999997 138100.0 201500.0 ;
      RECT  135500.0 210100.00000000003 136100.0 210700.0 ;
      RECT  135500.0 209700.0 136100.0 210300.0 ;
      RECT  133500.0 210100.00000000003 135800.0 210700.0 ;
      RECT  135500.0 210000.0 136100.0 210399.99999999997 ;
      RECT  135800.0 209700.0 138100.0 210300.0 ;
      RECT  135500.0 218899.99999999997 136100.0 219500.0 ;
      RECT  135500.0 219300.0 136100.0 219899.99999999997 ;
      RECT  133500.0 218899.99999999997 135800.0 219500.0 ;
      RECT  135500.0 219200.0 136100.0 219600.00000000003 ;
      RECT  135800.0 219300.0 138100.0 219899.99999999997 ;
      RECT  135500.0 228500.0 136100.0 229100.00000000003 ;
      RECT  135500.0 228100.00000000003 136100.0 228700.0 ;
      RECT  133500.0 228500.0 135800.0 229100.00000000003 ;
      RECT  135500.0 228399.99999999997 136100.0 228800.0 ;
      RECT  135800.0 228100.00000000003 138100.0 228700.0 ;
      RECT  135500.0 237300.0 136100.0 237899.99999999997 ;
      RECT  135500.0 237700.0 136100.0 238300.0 ;
      RECT  133500.0 237300.0 135800.0 237899.99999999997 ;
      RECT  135500.0 237600.00000000003 136100.0 238000.0 ;
      RECT  135800.0 237700.0 138100.0 238300.0 ;
      RECT  135500.0 246900.00000000003 136100.0 247500.0 ;
      RECT  135500.0 246500.0 136100.0 247100.00000000003 ;
      RECT  133500.0 246900.00000000003 135800.0 247500.0 ;
      RECT  135500.0 246800.0 136100.0 247200.0 ;
      RECT  135800.0 246500.0 138100.0 247100.00000000003 ;
      RECT  135500.0 255700.0 136100.0 256300.0 ;
      RECT  135500.0 256100.00000000003 136100.0 256700.0 ;
      RECT  133500.0 255700.0 135800.0 256300.0 ;
      RECT  135500.0 256000.0 136100.0 256400.00000000003 ;
      RECT  135800.0 256100.00000000003 138100.0 256700.0 ;
      RECT  135500.0 265300.0 136100.0 265900.0 ;
      RECT  135500.0 264900.00000000006 136100.0 265500.0 ;
      RECT  133500.0 265300.0 135800.0 265900.0 ;
      RECT  135500.0 265200.0 136100.0 265600.0 ;
      RECT  135800.0 264900.00000000006 138100.0 265500.0 ;
      RECT  135500.0 274100.0 136100.0 274700.0 ;
      RECT  135500.0 274500.0 136100.0 275100.0 ;
      RECT  133500.0 274100.0 135800.0 274700.0 ;
      RECT  135500.0 274400.00000000006 136100.0 274800.0 ;
      RECT  135800.0 274500.0 138100.0 275100.0 ;
      RECT  135500.0 283700.0 136100.0 284300.0 ;
      RECT  135500.0 283300.0 136100.0 283900.0 ;
      RECT  133500.0 283700.0 135800.0 284300.0 ;
      RECT  135500.0 283600.0 136100.0 284000.0 ;
      RECT  135800.0 283300.0 138100.0 283900.0 ;
      RECT  135500.0 292500.0 136100.0 293100.0 ;
      RECT  135500.0 292900.00000000006 136100.0 293500.0 ;
      RECT  133500.0 292500.0 135800.0 293100.0 ;
      RECT  135500.0 292800.0 136100.0 293200.0 ;
      RECT  135800.0 292900.00000000006 138100.0 293500.0 ;
      RECT  135500.0 302100.0 136100.0 302700.0 ;
      RECT  135500.0 301700.0 136100.0 302300.0 ;
      RECT  133500.0 302100.0 135800.0 302700.0 ;
      RECT  135500.0 302000.0 136100.0 302400.00000000006 ;
      RECT  135800.0 301700.0 138100.0 302300.0 ;
      RECT  135500.0 310900.0 136100.0 311500.0 ;
      RECT  135500.0 311300.0 136100.0 311900.0 ;
      RECT  133500.0 310900.0 135800.0 311500.0 ;
      RECT  135500.0 311200.0 136100.0 311600.0 ;
      RECT  135800.0 311300.0 138100.0 311900.0 ;
      RECT  116300.00000000001 173300.0 128500.0 173900.0 ;
      RECT  121900.0 171900.0 130500.0 172500.0 ;
      RECT  117700.0 182100.00000000003 128500.0 182700.0 ;
      RECT  121900.0 183500.0 130500.0 184100.00000000003 ;
      RECT  119100.0 191700.0 128500.0 192300.0 ;
      RECT  121900.0 190300.0 130500.0 190900.0 ;
      RECT  120500.0 200500.0 128500.0 201100.00000000003 ;
      RECT  121900.0 201899.99999999997 130500.0 202500.0 ;
      RECT  116300.00000000001 210100.00000000003 128500.0 210700.0 ;
      RECT  123300.00000000001 208700.0 130500.0 209300.0 ;
      RECT  117700.0 218899.99999999997 128500.0 219500.0 ;
      RECT  123300.00000000001 220300.0 130500.0 220899.99999999997 ;
      RECT  119100.0 228500.0 128500.0 229100.00000000003 ;
      RECT  123300.00000000001 227100.00000000003 130500.0 227700.0 ;
      RECT  120500.0 237300.0 128500.0 237899.99999999997 ;
      RECT  123300.00000000001 238700.0 130500.0 239300.0 ;
      RECT  116300.00000000001 246900.00000000003 128500.0 247500.0 ;
      RECT  124700.0 245500.0 130500.0 246100.00000000003 ;
      RECT  117700.0 255700.0 128500.0 256300.0 ;
      RECT  124700.0 257100.00000000003 130500.0 257700.0 ;
      RECT  119100.0 265300.0 128500.0 265900.0 ;
      RECT  124700.0 263900.00000000006 130500.0 264500.0 ;
      RECT  120500.0 274100.0 128500.0 274700.0 ;
      RECT  124700.0 275500.0 130500.0 276100.0 ;
      RECT  116300.00000000001 283700.0 128500.0 284300.0 ;
      RECT  126100.0 282300.0 130500.0 282900.0 ;
      RECT  117700.0 292500.0 128500.0 293100.0 ;
      RECT  126100.0 293900.00000000006 130500.0 294500.0 ;
      RECT  119100.0 302100.0 128500.0 302700.0 ;
      RECT  126100.0 300700.0 130500.0 301300.0 ;
      RECT  120500.0 310900.0 128500.0 311500.0 ;
      RECT  126100.0 312300.0 130500.0 312900.0 ;
      RECT  126900.0 177700.0 142900.0 178300.0 ;
      RECT  126900.0 168500.0 142900.0 169100.00000000003 ;
      RECT  126900.0 196100.00000000003 142900.0 196700.0 ;
      RECT  126900.0 186900.0 142900.0 187500.0 ;
      RECT  126900.0 214500.0 142900.0 215100.00000000003 ;
      RECT  126900.0 205300.0 142900.0 205899.99999999997 ;
      RECT  126900.0 232900.00000000003 142900.0 233500.0 ;
      RECT  126900.0 223700.0 142900.0 224300.0 ;
      RECT  126900.0 251300.0 142900.0 251899.99999999997 ;
      RECT  126900.0 242100.00000000003 142900.0 242700.0 ;
      RECT  126900.0 269700.0 142900.0 270300.0 ;
      RECT  126900.0 260500.0 142900.0 261100.00000000003 ;
      RECT  126900.0 288100.0 142900.0 288700.0 ;
      RECT  126900.0 278900.00000000006 142900.0 279500.0 ;
      RECT  126900.0 306500.0 142900.0 307100.0 ;
      RECT  126900.0 297300.0 142900.0 297900.0 ;
      RECT  91600.0 172900.0 92200.0 173500.0 ;
      RECT  91600.0 175900.0 92200.0 176500.0 ;
      RECT  88800.0 172900.0 91900.0 173500.0 ;
      RECT  91600.0 173200.0 92200.0 176200.0 ;
      RECT  91900.0 175900.0 94400.0 176500.0 ;
      RECT  82700.0 172900.0 86500.0 173500.0 ;
      RECT  91600.0 182500.0 92200.0 183100.00000000003 ;
      RECT  91600.0 185100.00000000003 92200.0 185700.0 ;
      RECT  88800.0 182500.0 91900.0 183100.00000000003 ;
      RECT  91600.0 182800.0 92200.0 185400.0 ;
      RECT  91900.0 185100.00000000003 95800.00000000001 185700.0 ;
      RECT  84100.0 182500.0 86500.0 183100.00000000003 ;
      RECT  82700.0 188300.0 97200.0 188900.0 ;
      RECT  84100.0 197500.0 98600.0 198100.00000000003 ;
      RECT  94400.0 173300.0 101300.00000000001 173900.0 ;
      RECT  95800.00000000001 171900.0 103300.00000000001 172500.0 ;
      RECT  97200.0 182100.00000000003 101300.00000000001 182700.0 ;
      RECT  95800.00000000001 183500.0 103300.00000000001 184100.00000000003 ;
      RECT  94400.0 191700.0 101300.00000000001 192300.0 ;
      RECT  98600.0 190300.0 103300.0 190900.0 ;
      RECT  97200.0 200500.0 101300.00000000001 201100.00000000003 ;
      RECT  98600.0 201899.99999999997 103300.0 202500.0 ;
      RECT  108300.00000000001 173300.0 108900.0 173900.0 ;
      RECT  108300.00000000001 172900.0 108900.0 173500.0 ;
      RECT  106300.00000000001 173300.0 108600.00000000001 173900.0 ;
      RECT  108300.00000000001 173200.0 108900.0 173600.00000000003 ;
      RECT  108600.0 172900.0 110900.0 173500.0 ;
      RECT  108300.00000000001 182100.00000000003 108900.0 182700.0 ;
      RECT  108300.00000000001 182500.0 108900.0 183100.00000000003 ;
      RECT  106300.00000000001 182100.00000000003 108600.00000000001 182700.0 ;
      RECT  108300.00000000001 182400.0 108900.0 182800.0 ;
      RECT  108600.0 182500.0 110900.0 183100.00000000003 ;
      RECT  108300.00000000001 191700.0 108900.0 192300.0 ;
      RECT  108300.00000000001 191300.0 108900.0 191900.0 ;
      RECT  106300.00000000001 191700.0 108600.00000000001 192300.0 ;
      RECT  108300.00000000001 191600.00000000003 108900.0 192000.0 ;
      RECT  108600.0 191300.0 110900.0 191900.0 ;
      RECT  108300.00000000001 200500.0 108900.0 201100.00000000003 ;
      RECT  108300.00000000001 200899.99999999997 108900.0 201500.0 ;
      RECT  106300.00000000001 200500.0 108600.00000000001 201100.00000000003 ;
      RECT  108300.00000000001 200800.0 108900.0 201200.0 ;
      RECT  108600.0 200899.99999999997 110900.0 201500.0 ;
      RECT  82100.0 177700.0 115700.0 178300.0 ;
      RECT  82100.0 168500.0 115700.0 169100.00000000003 ;
      RECT  82100.0 177700.0 115700.0 178300.0 ;
      RECT  82100.0 186900.0 115700.0 187500.0 ;
      RECT  82100.0 196100.00000000003 115700.0 196700.0 ;
      RECT  82100.0 186900.0 115700.0 187500.0 ;
      RECT  82100.0 196100.00000000003 115700.0 196700.0 ;
      RECT  82100.0 205300.0 115700.0 205899.99999999997 ;
      RECT  89300.0 176700.0 90100.0 178000.0 ;
      RECT  89300.0 168800.0 90100.0 170100.00000000003 ;
      RECT  86100.0 169700.0 86900.0 168500.0 ;
      RECT  86100.0 175900.0 86900.0 178300.0 ;
      RECT  87900.0 169700.0 88500.0 175900.0 ;
      RECT  86100.0 175900.0 86900.0 176700.0 ;
      RECT  87700.0 175900.0 88500.0 176700.0 ;
      RECT  87700.0 175900.0 88500.0 176700.0 ;
      RECT  86100.0 175900.0 86900.0 176700.0 ;
      RECT  86100.0 169700.0 86900.0 170500.0 ;
      RECT  87700.0 169700.0 88500.0 170500.0 ;
      RECT  87700.0 169700.0 88500.0 170500.0 ;
      RECT  86100.0 169700.0 86900.0 170500.0 ;
      RECT  89300.0 176300.0 90100.0 177100.00000000003 ;
      RECT  89300.0 169700.0 90100.0 170500.0 ;
      RECT  86500.0 172800.0 87300.0 173600.00000000003 ;
      RECT  86500.0 172800.0 87300.0 173600.00000000003 ;
      RECT  88200.0 172900.0 88800.0 173500.0 ;
      RECT  84900.0 177700.0 91300.00000000001 178300.0 ;
      RECT  84900.0 168500.0 91300.00000000001 169100.00000000003 ;
      RECT  89300.0 179300.0 90100.0 178000.0 ;
      RECT  89300.0 187200.0 90100.0 185900.0 ;
      RECT  86100.0 186300.0 86900.0 187500.0 ;
      RECT  86100.0 180100.00000000003 86900.0 177700.0 ;
      RECT  87900.0 186300.0 88500.0 180100.00000000003 ;
      RECT  86100.0 180100.00000000003 86900.0 179300.0 ;
      RECT  87700.0 180100.00000000003 88500.0 179300.0 ;
      RECT  87700.0 180100.00000000003 88500.0 179300.0 ;
      RECT  86100.0 180100.00000000003 86900.0 179300.0 ;
      RECT  86100.0 186300.0 86900.0 185500.0 ;
      RECT  87700.0 186300.0 88500.0 185500.0 ;
      RECT  87700.0 186300.0 88500.0 185500.0 ;
      RECT  86100.0 186300.0 86900.0 185500.0 ;
      RECT  89300.0 179700.0 90100.0 178900.0 ;
      RECT  89300.0 186300.0 90100.0 185500.0 ;
      RECT  86500.0 183200.0 87300.0 182400.0 ;
      RECT  86500.0 183200.0 87300.0 182400.0 ;
      RECT  88200.0 183100.00000000003 88800.0 182500.0 ;
      RECT  84900.0 178300.0 91300.00000000001 177700.0 ;
      RECT  84900.0 187500.0 91300.00000000001 186900.0 ;
      RECT  113700.0 176700.0 114500.0 178000.0 ;
      RECT  113700.0 168800.0 114500.0 170100.00000000003 ;
      RECT  110500.0 169700.0 111300.00000000001 168500.0 ;
      RECT  110500.0 175900.0 111300.00000000001 178300.0 ;
      RECT  112300.00000000001 169700.0 112900.0 175900.0 ;
      RECT  110500.0 175900.0 111300.00000000001 176700.0 ;
      RECT  112100.00000000001 175900.0 112900.0 176700.0 ;
      RECT  112100.00000000001 175900.0 112900.0 176700.0 ;
      RECT  110500.0 175900.0 111300.00000000001 176700.0 ;
      RECT  110500.0 169700.0 111300.00000000001 170500.0 ;
      RECT  112100.00000000001 169700.0 112900.0 170500.0 ;
      RECT  112100.00000000001 169700.0 112900.0 170500.0 ;
      RECT  110500.0 169700.0 111300.00000000001 170500.0 ;
      RECT  113700.0 176300.0 114500.0 177100.00000000003 ;
      RECT  113700.0 169700.0 114500.0 170500.0 ;
      RECT  110900.0 172800.0 111700.0 173600.00000000003 ;
      RECT  110900.0 172800.0 111700.0 173600.00000000003 ;
      RECT  112600.00000000001 172900.0 113200.0 173500.0 ;
      RECT  109300.00000000001 177700.0 115700.0 178300.0 ;
      RECT  109300.00000000001 168500.0 115700.0 169100.00000000003 ;
      RECT  113700.0 179300.0 114500.0 178000.0 ;
      RECT  113700.0 187200.0 114500.0 185900.0 ;
      RECT  110500.0 186300.0 111300.00000000001 187500.0 ;
      RECT  110500.0 180100.00000000003 111300.00000000001 177700.0 ;
      RECT  112300.00000000001 186300.0 112900.0 180100.00000000003 ;
      RECT  110500.0 180100.00000000003 111300.00000000001 179300.0 ;
      RECT  112100.00000000001 180100.00000000003 112900.0 179300.0 ;
      RECT  112100.00000000001 180100.00000000003 112900.0 179300.0 ;
      RECT  110500.0 180100.00000000003 111300.00000000001 179300.0 ;
      RECT  110500.0 186300.0 111300.00000000001 185500.0 ;
      RECT  112100.00000000001 186300.0 112900.0 185500.0 ;
      RECT  112100.00000000001 186300.0 112900.0 185500.0 ;
      RECT  110500.0 186300.0 111300.00000000001 185500.0 ;
      RECT  113700.0 179700.0 114500.0 178900.0 ;
      RECT  113700.0 186300.0 114500.0 185500.0 ;
      RECT  110900.0 183200.0 111700.0 182400.0 ;
      RECT  110900.0 183200.0 111700.0 182400.0 ;
      RECT  112600.00000000001 183100.00000000003 113200.0 182500.0 ;
      RECT  109300.00000000001 178300.0 115700.0 177700.0 ;
      RECT  109300.00000000001 187500.0 115700.0 186900.0 ;
      RECT  113700.0 195100.00000000003 114500.0 196400.0 ;
      RECT  113700.0 187200.0 114500.0 188500.0 ;
      RECT  110500.0 188100.00000000003 111300.00000000001 186900.0 ;
      RECT  110500.0 194300.0 111300.00000000001 196700.0 ;
      RECT  112300.00000000001 188100.00000000003 112900.0 194300.0 ;
      RECT  110500.0 194300.0 111300.00000000001 195100.00000000003 ;
      RECT  112100.00000000001 194300.0 112900.0 195100.00000000003 ;
      RECT  112100.00000000001 194300.0 112900.0 195100.00000000003 ;
      RECT  110500.0 194300.0 111300.00000000001 195100.00000000003 ;
      RECT  110500.0 188100.00000000003 111300.00000000001 188900.0 ;
      RECT  112100.00000000001 188100.00000000003 112900.0 188900.0 ;
      RECT  112100.00000000001 188100.00000000003 112900.0 188900.0 ;
      RECT  110500.0 188100.00000000003 111300.00000000001 188900.0 ;
      RECT  113700.0 194700.0 114500.0 195500.0 ;
      RECT  113700.0 188100.00000000003 114500.0 188900.0 ;
      RECT  110900.0 191200.0 111700.0 192000.0 ;
      RECT  110900.0 191200.0 111700.0 192000.0 ;
      RECT  112600.00000000001 191300.0 113200.0 191900.0 ;
      RECT  109300.00000000001 196100.00000000003 115700.0 196700.0 ;
      RECT  109300.00000000001 186900.0 115700.0 187500.0 ;
      RECT  113700.0 197700.0 114500.0 196400.0 ;
      RECT  113700.0 205600.00000000003 114500.0 204300.0 ;
      RECT  110500.0 204700.0 111300.00000000001 205899.99999999997 ;
      RECT  110500.0 198500.0 111300.00000000001 196100.00000000003 ;
      RECT  112300.00000000001 204700.0 112900.0 198500.0 ;
      RECT  110500.0 198500.0 111300.00000000001 197700.0 ;
      RECT  112100.00000000001 198500.0 112900.0 197700.0 ;
      RECT  112100.00000000001 198500.0 112900.0 197700.0 ;
      RECT  110500.0 198500.0 111300.00000000001 197700.0 ;
      RECT  110500.0 204700.0 111300.00000000001 203899.99999999997 ;
      RECT  112100.00000000001 204700.0 112900.0 203899.99999999997 ;
      RECT  112100.00000000001 204700.0 112900.0 203899.99999999997 ;
      RECT  110500.0 204700.0 111300.00000000001 203899.99999999997 ;
      RECT  113700.0 198100.00000000003 114500.0 197300.0 ;
      RECT  113700.0 204700.0 114500.0 203899.99999999997 ;
      RECT  110900.0 201600.00000000003 111700.0 200800.0 ;
      RECT  110900.0 201600.00000000003 111700.0 200800.0 ;
      RECT  112600.00000000001 201500.0 113200.0 200899.99999999997 ;
      RECT  109300.00000000001 196700.0 115700.0 196100.00000000003 ;
      RECT  109300.00000000001 205899.99999999997 115700.0 205300.0 ;
      RECT  100900.0 170100.00000000003 101700.0 168500.0 ;
      RECT  100900.0 175900.0 101700.0 178300.0 ;
      RECT  104100.0 175900.0 104900.0 178300.0 ;
      RECT  105700.0 176700.0 106500.0 178000.0 ;
      RECT  105700.0 168800.0 106500.0 170100.00000000003 ;
      RECT  100900.0 175900.0 101700.0 176700.0 ;
      RECT  102500.0 175900.0 103300.00000000001 176700.0 ;
      RECT  102500.0 175900.0 103300.00000000001 176700.0 ;
      RECT  100900.0 175900.0 101700.0 176700.0 ;
      RECT  102500.0 175900.0 103300.00000000001 176700.0 ;
      RECT  104100.0 175900.0 104900.0 176700.0 ;
      RECT  104100.0 175900.0 104900.0 176700.0 ;
      RECT  102500.0 175900.0 103300.00000000001 176700.0 ;
      RECT  100900.0 170100.00000000003 101700.0 170900.0 ;
      RECT  102500.0 170100.00000000003 103300.00000000001 170900.0 ;
      RECT  102500.0 170100.00000000003 103300.00000000001 170900.0 ;
      RECT  100900.0 170100.00000000003 101700.0 170900.0 ;
      RECT  102500.0 170100.00000000003 103300.00000000001 170900.0 ;
      RECT  104100.0 170100.00000000003 104900.0 170900.0 ;
      RECT  104100.0 170100.00000000003 104900.0 170900.0 ;
      RECT  102500.0 170100.00000000003 103300.00000000001 170900.0 ;
      RECT  105700.0 176300.0 106500.0 177100.00000000003 ;
      RECT  105700.0 169700.0 106500.0 170500.0 ;
      RECT  104100.0 171800.0 103300.00000000001 172600.00000000003 ;
      RECT  102100.0 173200.0 101300.00000000001 174000.0 ;
      RECT  102500.0 175900.0 103300.00000000001 176700.0 ;
      RECT  104100.0 170100.00000000003 104900.0 170900.0 ;
      RECT  106300.00000000001 173200.0 105500.0 174000.0 ;
      RECT  101300.00000000001 173200.0 102100.0 174000.0 ;
      RECT  103300.00000000001 171800.0 104100.0 172600.00000000003 ;
      RECT  105500.0 173200.0 106300.00000000001 174000.0 ;
      RECT  99700.0 177700.0 109300.00000000001 178300.0 ;
      RECT  99700.0 168500.0 109300.00000000001 169100.00000000003 ;
      RECT  100900.0 185900.0 101700.0 187500.0 ;
      RECT  100900.0 180100.00000000003 101700.0 177700.0 ;
      RECT  104100.0 180100.00000000003 104900.0 177700.0 ;
      RECT  105700.0 179300.0 106500.0 178000.0 ;
      RECT  105700.0 187200.0 106500.0 185900.0 ;
      RECT  100900.0 180100.00000000003 101700.0 179300.0 ;
      RECT  102500.0 180100.00000000003 103300.00000000001 179300.0 ;
      RECT  102500.0 180100.00000000003 103300.00000000001 179300.0 ;
      RECT  100900.0 180100.00000000003 101700.0 179300.0 ;
      RECT  102500.0 180100.00000000003 103300.00000000001 179300.0 ;
      RECT  104100.0 180100.00000000003 104900.0 179300.0 ;
      RECT  104100.0 180100.00000000003 104900.0 179300.0 ;
      RECT  102500.0 180100.00000000003 103300.00000000001 179300.0 ;
      RECT  100900.0 185900.0 101700.0 185100.00000000003 ;
      RECT  102500.0 185900.0 103300.00000000001 185100.00000000003 ;
      RECT  102500.0 185900.0 103300.00000000001 185100.00000000003 ;
      RECT  100900.0 185900.0 101700.0 185100.00000000003 ;
      RECT  102500.0 185900.0 103300.00000000001 185100.00000000003 ;
      RECT  104100.0 185900.0 104900.0 185100.00000000003 ;
      RECT  104100.0 185900.0 104900.0 185100.00000000003 ;
      RECT  102500.0 185900.0 103300.00000000001 185100.00000000003 ;
      RECT  105700.0 179700.0 106500.0 178900.0 ;
      RECT  105700.0 186300.0 106500.0 185500.0 ;
      RECT  104100.0 184200.0 103300.00000000001 183400.0 ;
      RECT  102100.0 182800.0 101300.00000000001 182000.0 ;
      RECT  102500.0 180100.00000000003 103300.00000000001 179300.0 ;
      RECT  104100.0 185900.0 104900.0 185100.00000000003 ;
      RECT  106300.00000000001 182800.0 105500.0 182000.0 ;
      RECT  101300.00000000001 182800.0 102100.0 182000.0 ;
      RECT  103300.00000000001 184200.0 104100.0 183400.0 ;
      RECT  105500.0 182800.0 106300.00000000001 182000.0 ;
      RECT  99700.0 178300.0 109300.00000000001 177700.0 ;
      RECT  99700.0 187500.0 109300.00000000001 186900.0 ;
      RECT  100900.0 188500.0 101700.0 186900.0 ;
      RECT  100900.0 194300.0 101700.0 196700.0 ;
      RECT  104100.0 194300.0 104900.0 196700.0 ;
      RECT  105700.0 195100.00000000003 106500.0 196400.0 ;
      RECT  105700.0 187200.0 106500.0 188500.0 ;
      RECT  100900.0 194300.0 101700.0 195100.00000000003 ;
      RECT  102500.0 194300.0 103300.00000000001 195100.00000000003 ;
      RECT  102500.0 194300.0 103300.00000000001 195100.00000000003 ;
      RECT  100900.0 194300.0 101700.0 195100.00000000003 ;
      RECT  102500.0 194300.0 103300.00000000001 195100.00000000003 ;
      RECT  104100.0 194300.0 104900.0 195100.00000000003 ;
      RECT  104100.0 194300.0 104900.0 195100.00000000003 ;
      RECT  102500.0 194300.0 103300.00000000001 195100.00000000003 ;
      RECT  100900.0 188500.0 101700.0 189300.0 ;
      RECT  102500.0 188500.0 103300.00000000001 189300.0 ;
      RECT  102500.0 188500.0 103300.00000000001 189300.0 ;
      RECT  100900.0 188500.0 101700.0 189300.0 ;
      RECT  102500.0 188500.0 103300.00000000001 189300.0 ;
      RECT  104100.0 188500.0 104900.0 189300.0 ;
      RECT  104100.0 188500.0 104900.0 189300.0 ;
      RECT  102500.0 188500.0 103300.00000000001 189300.0 ;
      RECT  105700.0 194700.0 106500.0 195500.0 ;
      RECT  105700.0 188100.00000000003 106500.0 188900.0 ;
      RECT  104100.0 190200.0 103300.00000000001 191000.0 ;
      RECT  102100.0 191600.00000000003 101300.00000000001 192400.0 ;
      RECT  102500.0 194300.0 103300.00000000001 195100.00000000003 ;
      RECT  104100.0 188500.0 104900.0 189300.0 ;
      RECT  106300.00000000001 191600.00000000003 105500.0 192400.0 ;
      RECT  101300.00000000001 191600.00000000003 102100.0 192400.0 ;
      RECT  103300.00000000001 190200.0 104100.0 191000.0 ;
      RECT  105500.0 191600.00000000003 106300.00000000001 192400.0 ;
      RECT  99700.0 196100.00000000003 109300.00000000001 196700.0 ;
      RECT  99700.0 186900.0 109300.00000000001 187500.0 ;
      RECT  100900.0 204300.0 101700.0 205899.99999999997 ;
      RECT  100900.0 198500.0 101700.0 196100.00000000003 ;
      RECT  104100.0 198500.0 104900.0 196100.00000000003 ;
      RECT  105700.0 197700.0 106500.0 196400.0 ;
      RECT  105700.0 205600.00000000003 106500.0 204300.0 ;
      RECT  100900.0 198500.0 101700.0 197700.0 ;
      RECT  102500.0 198500.0 103300.00000000001 197700.0 ;
      RECT  102500.0 198500.0 103300.00000000001 197700.0 ;
      RECT  100900.0 198500.0 101700.0 197700.0 ;
      RECT  102500.0 198500.0 103300.00000000001 197700.0 ;
      RECT  104100.0 198500.0 104900.0 197700.0 ;
      RECT  104100.0 198500.0 104900.0 197700.0 ;
      RECT  102500.0 198500.0 103300.00000000001 197700.0 ;
      RECT  100900.0 204300.0 101700.0 203500.0 ;
      RECT  102500.0 204300.0 103300.00000000001 203500.0 ;
      RECT  102500.0 204300.0 103300.00000000001 203500.0 ;
      RECT  100900.0 204300.0 101700.0 203500.0 ;
      RECT  102500.0 204300.0 103300.00000000001 203500.0 ;
      RECT  104100.0 204300.0 104900.0 203500.0 ;
      RECT  104100.0 204300.0 104900.0 203500.0 ;
      RECT  102500.0 204300.0 103300.00000000001 203500.0 ;
      RECT  105700.0 198100.00000000003 106500.0 197300.0 ;
      RECT  105700.0 204700.0 106500.0 203899.99999999997 ;
      RECT  104100.0 202600.00000000003 103300.00000000001 201800.0 ;
      RECT  102100.0 201200.0 101300.00000000001 200400.00000000003 ;
      RECT  102500.0 198500.0 103300.00000000001 197700.0 ;
      RECT  104100.0 204300.0 104900.0 203500.0 ;
      RECT  106300.00000000001 201200.0 105500.0 200400.00000000003 ;
      RECT  101300.00000000001 201200.0 102100.0 200400.00000000003 ;
      RECT  103300.00000000001 202600.00000000003 104100.0 201800.0 ;
      RECT  105500.0 201200.0 106300.00000000001 200400.00000000003 ;
      RECT  99700.0 196700.0 109300.00000000001 196100.00000000003 ;
      RECT  99700.0 205899.99999999997 109300.00000000001 205300.0 ;
      RECT  94800.00000000001 175800.0 94000.0 176600.00000000003 ;
      RECT  83100.0 172800.0 82300.0 173600.00000000003 ;
      RECT  96200.0 185000.0 95400.0 185800.0 ;
      RECT  84500.0 182400.0 83700.0 183200.0 ;
      RECT  83100.0 188200.0 82300.0 189000.0 ;
      RECT  97600.0 188200.0 96800.0 189000.0 ;
      RECT  84500.0 197400.0 83700.0 198200.0 ;
      RECT  99000.0 197400.0 98200.0 198200.0 ;
      RECT  94800.00000000001 173200.0 94000.0 174000.0 ;
      RECT  96200.0 171800.0 95400.0 172600.00000000003 ;
      RECT  97600.0 182000.0 96800.0 182800.0 ;
      RECT  96200.0 183400.0 95400.0 184200.0 ;
      RECT  94800.00000000001 191600.00000000003 94000.0 192400.0 ;
      RECT  99000.0 190200.0 98200.0 191000.0 ;
      RECT  97600.0 200399.99999999997 96800.0 201200.0 ;
      RECT  99000.0 201800.0 98200.0 202600.00000000003 ;
      RECT  91700.0 177600.00000000003 90900.0 178400.0 ;
      RECT  109100.0 177600.00000000003 108300.0 178400.0 ;
      RECT  91700.0 168400.0 90900.0 169200.0 ;
      RECT  109100.0 168400.0 108300.0 169200.0 ;
      RECT  91700.0 177600.00000000003 90900.0 178400.0 ;
      RECT  109100.0 177600.00000000003 108300.0 178400.0 ;
      RECT  91700.0 186800.0 90900.0 187600.00000000003 ;
      RECT  109100.0 186800.0 108300.0 187600.00000000003 ;
      RECT  91700.0 196000.0 90900.0 196800.0 ;
      RECT  109100.0 196000.0 108300.0 196800.0 ;
      RECT  91700.0 186800.0 90900.0 187600.00000000003 ;
      RECT  109100.0 186800.0 108300.0 187600.00000000003 ;
      RECT  91700.0 196000.0 90900.0 196800.0 ;
      RECT  109100.0 196000.0 108300.0 196800.0 ;
      RECT  91700.0 205200.0 90900.0 206000.0 ;
      RECT  109100.0 205200.0 108300.0 206000.0 ;
      RECT  112600.0 172900.0 113200.0 173500.0 ;
      RECT  112600.0 182500.0 113200.0 183100.00000000003 ;
      RECT  112600.0 191300.0 113200.0 191900.0 ;
      RECT  112600.0 200899.99999999997 113200.0 201500.0 ;
      RECT  91600.0 209700.0 92200.0 210300.0 ;
      RECT  91600.0 212700.0 92200.0 213300.0 ;
      RECT  88800.0 209700.0 91900.0 210300.0 ;
      RECT  91600.0 210000.0 92200.0 213000.0 ;
      RECT  91900.0 212700.0 94400.0 213300.0 ;
      RECT  82700.0 209700.0 86500.0 210300.0 ;
      RECT  91600.0 219300.0 92200.0 219899.99999999997 ;
      RECT  91600.0 221899.99999999997 92200.0 222500.0 ;
      RECT  88800.0 219300.0 91900.0 219899.99999999997 ;
      RECT  91600.0 219600.00000000003 92200.0 222200.0 ;
      RECT  91900.0 221899.99999999997 95800.00000000001 222500.0 ;
      RECT  84100.0 219300.0 86500.0 219899.99999999997 ;
      RECT  82700.0 225100.00000000003 97200.0 225700.0 ;
      RECT  84100.0 234300.0 98600.0 234899.99999999997 ;
      RECT  94400.0 210100.00000000003 101300.00000000001 210700.0 ;
      RECT  95800.00000000001 208700.0 103300.00000000001 209300.0 ;
      RECT  97200.0 218899.99999999997 101300.00000000001 219500.0 ;
      RECT  95800.00000000001 220300.0 103300.00000000001 220899.99999999997 ;
      RECT  94400.0 228500.0 101300.00000000001 229100.00000000003 ;
      RECT  98600.0 227100.00000000003 103300.0 227700.0 ;
      RECT  97200.0 237300.0 101300.00000000001 237899.99999999997 ;
      RECT  98600.0 238700.0 103300.0 239300.0 ;
      RECT  108300.00000000001 210100.00000000003 108900.0 210700.0 ;
      RECT  108300.00000000001 209700.0 108900.0 210300.0 ;
      RECT  106300.00000000001 210100.00000000003 108600.00000000001 210700.0 ;
      RECT  108300.00000000001 210000.0 108900.0 210399.99999999997 ;
      RECT  108600.0 209700.0 110900.0 210300.0 ;
      RECT  108300.00000000001 218899.99999999997 108900.0 219500.0 ;
      RECT  108300.00000000001 219300.0 108900.0 219899.99999999997 ;
      RECT  106300.00000000001 218899.99999999997 108600.00000000001 219500.0 ;
      RECT  108300.00000000001 219200.0 108900.0 219600.00000000003 ;
      RECT  108600.0 219300.0 110900.0 219899.99999999997 ;
      RECT  108300.00000000001 228500.0 108900.0 229100.00000000003 ;
      RECT  108300.00000000001 228100.00000000003 108900.0 228700.0 ;
      RECT  106300.00000000001 228500.0 108600.00000000001 229100.00000000003 ;
      RECT  108300.00000000001 228399.99999999997 108900.0 228800.0 ;
      RECT  108600.0 228100.00000000003 110900.0 228700.0 ;
      RECT  108300.00000000001 237300.0 108900.0 237899.99999999997 ;
      RECT  108300.00000000001 237700.0 108900.0 238300.0 ;
      RECT  106300.00000000001 237300.0 108600.00000000001 237899.99999999997 ;
      RECT  108300.00000000001 237600.00000000003 108900.0 238000.0 ;
      RECT  108600.0 237700.0 110900.0 238300.0 ;
      RECT  82100.0 214500.0 115700.0 215100.00000000003 ;
      RECT  82100.0 205300.0 115700.0 205899.99999999997 ;
      RECT  82100.0 214500.0 115700.0 215100.00000000003 ;
      RECT  82100.0 223700.0 115700.0 224300.0 ;
      RECT  82100.0 232899.99999999997 115700.0 233500.0 ;
      RECT  82100.0 223700.0 115700.0 224300.0 ;
      RECT  82100.0 232899.99999999997 115700.0 233500.0 ;
      RECT  82100.0 242100.00000000003 115700.0 242700.0 ;
      RECT  89300.0 213500.0 90100.0 214800.0 ;
      RECT  89300.0 205600.00000000003 90100.0 206899.99999999997 ;
      RECT  86100.0 206500.0 86900.0 205300.0 ;
      RECT  86100.0 212700.0 86900.0 215100.00000000003 ;
      RECT  87900.0 206500.0 88500.0 212700.0 ;
      RECT  86100.0 212700.0 86900.0 213500.0 ;
      RECT  87700.0 212700.0 88500.0 213500.0 ;
      RECT  87700.0 212700.0 88500.0 213500.0 ;
      RECT  86100.0 212700.0 86900.0 213500.0 ;
      RECT  86100.0 206500.0 86900.0 207300.0 ;
      RECT  87700.0 206500.0 88500.0 207300.0 ;
      RECT  87700.0 206500.0 88500.0 207300.0 ;
      RECT  86100.0 206500.0 86900.0 207300.0 ;
      RECT  89300.0 213100.00000000003 90100.0 213899.99999999997 ;
      RECT  89300.0 206500.0 90100.0 207300.0 ;
      RECT  86500.0 209600.00000000003 87300.0 210399.99999999997 ;
      RECT  86500.0 209600.00000000003 87300.0 210399.99999999997 ;
      RECT  88200.0 209700.0 88800.0 210300.0 ;
      RECT  84900.0 214500.0 91300.00000000001 215100.00000000003 ;
      RECT  84900.0 205300.0 91300.00000000001 205899.99999999997 ;
      RECT  89300.0 216100.00000000003 90100.0 214800.0 ;
      RECT  89300.0 224000.0 90100.0 222700.0 ;
      RECT  86100.0 223100.00000000003 86900.0 224300.0 ;
      RECT  86100.0 216899.99999999997 86900.0 214500.0 ;
      RECT  87900.0 223100.00000000003 88500.0 216899.99999999997 ;
      RECT  86100.0 216900.00000000003 86900.0 216100.00000000003 ;
      RECT  87700.0 216900.00000000003 88500.0 216100.00000000003 ;
      RECT  87700.0 216900.00000000003 88500.0 216100.00000000003 ;
      RECT  86100.0 216900.00000000003 86900.0 216100.00000000003 ;
      RECT  86100.0 223100.00000000003 86900.0 222300.0 ;
      RECT  87700.0 223100.00000000003 88500.0 222300.0 ;
      RECT  87700.0 223100.00000000003 88500.0 222300.0 ;
      RECT  86100.0 223100.00000000003 86900.0 222300.0 ;
      RECT  89300.0 216500.0 90100.0 215700.0 ;
      RECT  89300.0 223100.00000000003 90100.0 222300.0 ;
      RECT  86500.0 220000.0 87300.0 219200.0 ;
      RECT  86500.0 220000.0 87300.0 219200.0 ;
      RECT  88200.0 219899.99999999997 88800.0 219300.0 ;
      RECT  84900.0 215100.00000000003 91300.00000000001 214500.0 ;
      RECT  84900.0 224300.0 91300.00000000001 223700.0 ;
      RECT  113700.0 213500.0 114500.0 214800.0 ;
      RECT  113700.0 205600.00000000003 114500.0 206899.99999999997 ;
      RECT  110500.0 206500.0 111300.00000000001 205300.0 ;
      RECT  110500.0 212700.0 111300.00000000001 215100.00000000003 ;
      RECT  112300.00000000001 206500.0 112900.0 212700.0 ;
      RECT  110500.0 212700.0 111300.00000000001 213500.0 ;
      RECT  112100.00000000001 212700.0 112900.0 213500.0 ;
      RECT  112100.00000000001 212700.0 112900.0 213500.0 ;
      RECT  110500.0 212700.0 111300.00000000001 213500.0 ;
      RECT  110500.0 206500.0 111300.00000000001 207300.0 ;
      RECT  112100.00000000001 206500.0 112900.0 207300.0 ;
      RECT  112100.00000000001 206500.0 112900.0 207300.0 ;
      RECT  110500.0 206500.0 111300.00000000001 207300.0 ;
      RECT  113700.0 213100.00000000003 114500.0 213899.99999999997 ;
      RECT  113700.0 206500.0 114500.0 207300.0 ;
      RECT  110900.0 209600.00000000003 111700.0 210399.99999999997 ;
      RECT  110900.0 209600.00000000003 111700.0 210399.99999999997 ;
      RECT  112600.00000000001 209700.0 113200.0 210300.0 ;
      RECT  109300.00000000001 214500.0 115700.0 215100.00000000003 ;
      RECT  109300.00000000001 205300.0 115700.0 205899.99999999997 ;
      RECT  113700.0 216100.00000000003 114500.0 214800.0 ;
      RECT  113700.0 224000.0 114500.0 222700.0 ;
      RECT  110500.0 223100.00000000003 111300.00000000001 224300.0 ;
      RECT  110500.0 216899.99999999997 111300.00000000001 214500.0 ;
      RECT  112300.00000000001 223100.00000000003 112900.0 216899.99999999997 ;
      RECT  110500.0 216900.00000000003 111300.00000000001 216100.00000000003 ;
      RECT  112100.00000000001 216900.00000000003 112900.0 216100.00000000003 ;
      RECT  112100.00000000001 216900.00000000003 112900.0 216100.00000000003 ;
      RECT  110500.0 216900.00000000003 111300.00000000001 216100.00000000003 ;
      RECT  110500.0 223100.00000000003 111300.00000000001 222300.0 ;
      RECT  112100.00000000001 223100.00000000003 112900.0 222300.0 ;
      RECT  112100.00000000001 223100.00000000003 112900.0 222300.0 ;
      RECT  110500.0 223100.00000000003 111300.00000000001 222300.0 ;
      RECT  113700.0 216500.0 114500.0 215700.0 ;
      RECT  113700.0 223100.00000000003 114500.0 222300.0 ;
      RECT  110900.0 220000.0 111700.0 219200.0 ;
      RECT  110900.0 220000.0 111700.0 219200.0 ;
      RECT  112600.00000000001 219899.99999999997 113200.0 219300.0 ;
      RECT  109300.00000000001 215100.00000000003 115700.0 214500.0 ;
      RECT  109300.00000000001 224300.0 115700.0 223700.0 ;
      RECT  113700.0 231900.00000000003 114500.0 233200.0 ;
      RECT  113700.0 224000.0 114500.0 225300.0 ;
      RECT  110500.0 224899.99999999997 111300.00000000001 223700.0 ;
      RECT  110500.0 231100.00000000003 111300.00000000001 233500.0 ;
      RECT  112300.00000000001 224899.99999999997 112900.0 231100.00000000003 ;
      RECT  110500.0 231100.00000000003 111300.00000000001 231900.00000000003 ;
      RECT  112100.00000000001 231100.00000000003 112900.0 231900.00000000003 ;
      RECT  112100.00000000001 231100.00000000003 112900.0 231900.00000000003 ;
      RECT  110500.0 231100.00000000003 111300.00000000001 231900.00000000003 ;
      RECT  110500.0 224899.99999999997 111300.00000000001 225700.0 ;
      RECT  112100.00000000001 224899.99999999997 112900.0 225700.0 ;
      RECT  112100.00000000001 224899.99999999997 112900.0 225700.0 ;
      RECT  110500.0 224899.99999999997 111300.00000000001 225700.0 ;
      RECT  113700.0 231500.0 114500.0 232300.0 ;
      RECT  113700.0 224899.99999999997 114500.0 225700.0 ;
      RECT  110900.0 228000.0 111700.0 228800.0 ;
      RECT  110900.0 228000.0 111700.0 228800.0 ;
      RECT  112600.00000000001 228100.00000000003 113200.0 228700.0 ;
      RECT  109300.00000000001 232899.99999999997 115700.0 233500.0 ;
      RECT  109300.00000000001 223700.0 115700.0 224300.0 ;
      RECT  113700.0 234500.0 114500.0 233200.0 ;
      RECT  113700.0 242399.99999999997 114500.0 241100.00000000003 ;
      RECT  110500.0 241500.0 111300.00000000001 242700.0 ;
      RECT  110500.0 235300.0 111300.00000000001 232899.99999999997 ;
      RECT  112300.00000000001 241500.0 112900.0 235300.0 ;
      RECT  110500.0 235300.0 111300.00000000001 234500.0 ;
      RECT  112100.00000000001 235300.0 112900.0 234500.0 ;
      RECT  112100.00000000001 235300.0 112900.0 234500.0 ;
      RECT  110500.0 235300.0 111300.00000000001 234500.0 ;
      RECT  110500.0 241500.0 111300.00000000001 240700.0 ;
      RECT  112100.00000000001 241500.0 112900.0 240700.0 ;
      RECT  112100.00000000001 241500.0 112900.0 240700.0 ;
      RECT  110500.0 241500.0 111300.00000000001 240700.0 ;
      RECT  113700.0 234899.99999999997 114500.0 234100.00000000003 ;
      RECT  113700.0 241500.0 114500.0 240700.0 ;
      RECT  110900.0 238399.99999999997 111700.0 237600.00000000003 ;
      RECT  110900.0 238399.99999999997 111700.0 237600.00000000003 ;
      RECT  112600.00000000001 238300.0 113200.0 237700.0 ;
      RECT  109300.00000000001 233500.0 115700.0 232899.99999999997 ;
      RECT  109300.00000000001 242700.0 115700.0 242100.00000000003 ;
      RECT  100900.0 206899.99999999997 101700.0 205300.0 ;
      RECT  100900.0 212700.0 101700.0 215100.00000000003 ;
      RECT  104100.0 212700.0 104900.0 215100.00000000003 ;
      RECT  105700.0 213500.0 106500.0 214800.0 ;
      RECT  105700.0 205600.00000000003 106500.0 206899.99999999997 ;
      RECT  100900.0 212700.0 101700.0 213500.0 ;
      RECT  102500.0 212700.0 103300.00000000001 213500.0 ;
      RECT  102500.0 212700.0 103300.00000000001 213500.0 ;
      RECT  100900.0 212700.0 101700.0 213500.0 ;
      RECT  102500.0 212700.0 103300.00000000001 213500.0 ;
      RECT  104100.0 212700.0 104900.0 213500.0 ;
      RECT  104100.0 212700.0 104900.0 213500.0 ;
      RECT  102500.0 212700.0 103300.00000000001 213500.0 ;
      RECT  100900.0 206899.99999999997 101700.0 207700.0 ;
      RECT  102500.0 206899.99999999997 103300.00000000001 207700.0 ;
      RECT  102500.0 206899.99999999997 103300.00000000001 207700.0 ;
      RECT  100900.0 206899.99999999997 101700.0 207700.0 ;
      RECT  102500.0 206899.99999999997 103300.00000000001 207700.0 ;
      RECT  104100.0 206899.99999999997 104900.0 207700.0 ;
      RECT  104100.0 206899.99999999997 104900.0 207700.0 ;
      RECT  102500.0 206899.99999999997 103300.00000000001 207700.0 ;
      RECT  105700.0 213100.00000000003 106500.0 213899.99999999997 ;
      RECT  105700.0 206500.0 106500.0 207300.0 ;
      RECT  104100.0 208600.00000000003 103300.00000000001 209399.99999999997 ;
      RECT  102100.0 210000.0 101300.00000000001 210800.0 ;
      RECT  102500.0 212700.0 103300.00000000001 213500.0 ;
      RECT  104100.0 206899.99999999997 104900.0 207700.0 ;
      RECT  106300.00000000001 210000.0 105500.0 210800.0 ;
      RECT  101300.00000000001 210000.0 102100.0 210800.0 ;
      RECT  103300.00000000001 208600.00000000003 104100.0 209399.99999999997 ;
      RECT  105500.0 210000.0 106300.00000000001 210800.0 ;
      RECT  99700.0 214500.0 109300.00000000001 215100.00000000003 ;
      RECT  99700.0 205300.0 109300.00000000001 205899.99999999997 ;
      RECT  100900.0 222700.0 101700.0 224300.0 ;
      RECT  100900.0 216899.99999999997 101700.0 214500.0 ;
      RECT  104100.0 216899.99999999997 104900.0 214500.0 ;
      RECT  105700.0 216100.00000000003 106500.0 214800.0 ;
      RECT  105700.0 224000.0 106500.0 222700.0 ;
      RECT  100900.0 216900.00000000003 101700.0 216100.00000000003 ;
      RECT  102500.0 216900.00000000003 103300.00000000001 216100.00000000003 ;
      RECT  102500.0 216900.00000000003 103300.00000000001 216100.00000000003 ;
      RECT  100900.0 216900.00000000003 101700.0 216100.00000000003 ;
      RECT  102500.0 216900.00000000003 103300.00000000001 216100.00000000003 ;
      RECT  104100.0 216900.00000000003 104900.0 216100.00000000003 ;
      RECT  104100.0 216900.00000000003 104900.0 216100.00000000003 ;
      RECT  102500.0 216900.00000000003 103300.00000000001 216100.00000000003 ;
      RECT  100900.0 222700.0 101700.0 221899.99999999997 ;
      RECT  102500.0 222700.0 103300.00000000001 221899.99999999997 ;
      RECT  102500.0 222700.0 103300.00000000001 221899.99999999997 ;
      RECT  100900.0 222700.0 101700.0 221899.99999999997 ;
      RECT  102500.0 222700.0 103300.00000000001 221899.99999999997 ;
      RECT  104100.0 222700.0 104900.0 221899.99999999997 ;
      RECT  104100.0 222700.0 104900.0 221899.99999999997 ;
      RECT  102500.0 222700.0 103300.00000000001 221899.99999999997 ;
      RECT  105700.0 216500.0 106500.0 215700.0 ;
      RECT  105700.0 223100.00000000003 106500.0 222300.0 ;
      RECT  104100.0 221000.0 103300.00000000001 220200.0 ;
      RECT  102100.0 219600.00000000003 101300.00000000001 218800.0 ;
      RECT  102500.0 216899.99999999997 103300.00000000001 216100.00000000003 ;
      RECT  104100.0 222700.0 104900.0 221899.99999999997 ;
      RECT  106300.00000000001 219600.00000000003 105500.0 218800.0 ;
      RECT  101300.00000000001 219600.00000000003 102100.0 218800.0 ;
      RECT  103300.00000000001 221000.0 104100.0 220200.0 ;
      RECT  105500.0 219600.00000000003 106300.00000000001 218800.0 ;
      RECT  99700.0 215100.00000000003 109300.00000000001 214500.0 ;
      RECT  99700.0 224300.0 109300.00000000001 223700.0 ;
      RECT  100900.0 225300.0 101700.0 223700.0 ;
      RECT  100900.0 231100.00000000003 101700.0 233500.0 ;
      RECT  104100.0 231100.00000000003 104900.0 233500.0 ;
      RECT  105700.0 231900.00000000003 106500.0 233200.0 ;
      RECT  105700.0 224000.0 106500.0 225300.0 ;
      RECT  100900.0 231100.00000000003 101700.0 231900.00000000003 ;
      RECT  102500.0 231100.00000000003 103300.00000000001 231900.00000000003 ;
      RECT  102500.0 231100.00000000003 103300.00000000001 231900.00000000003 ;
      RECT  100900.0 231100.00000000003 101700.0 231900.00000000003 ;
      RECT  102500.0 231100.00000000003 103300.00000000001 231900.00000000003 ;
      RECT  104100.0 231100.00000000003 104900.0 231900.00000000003 ;
      RECT  104100.0 231100.00000000003 104900.0 231900.00000000003 ;
      RECT  102500.0 231100.00000000003 103300.00000000001 231900.00000000003 ;
      RECT  100900.0 225300.0 101700.0 226100.00000000003 ;
      RECT  102500.0 225300.0 103300.00000000001 226100.00000000003 ;
      RECT  102500.0 225300.0 103300.00000000001 226100.00000000003 ;
      RECT  100900.0 225300.0 101700.0 226100.00000000003 ;
      RECT  102500.0 225300.0 103300.00000000001 226100.00000000003 ;
      RECT  104100.0 225300.0 104900.0 226100.00000000003 ;
      RECT  104100.0 225300.0 104900.0 226100.00000000003 ;
      RECT  102500.0 225300.0 103300.00000000001 226100.00000000003 ;
      RECT  105700.0 231500.0 106500.0 232300.0 ;
      RECT  105700.0 224899.99999999997 106500.0 225700.0 ;
      RECT  104100.0 227000.0 103300.00000000001 227800.0 ;
      RECT  102100.0 228400.00000000003 101300.00000000001 229200.0 ;
      RECT  102500.0 231100.00000000003 103300.00000000001 231900.00000000003 ;
      RECT  104100.0 225300.0 104900.0 226100.00000000003 ;
      RECT  106300.00000000001 228400.00000000003 105500.0 229200.0 ;
      RECT  101300.00000000001 228400.00000000003 102100.0 229200.0 ;
      RECT  103300.00000000001 227000.0 104100.0 227800.0 ;
      RECT  105500.0 228400.00000000003 106300.00000000001 229200.0 ;
      RECT  99700.0 232899.99999999997 109300.00000000001 233500.0 ;
      RECT  99700.0 223700.0 109300.00000000001 224300.0 ;
      RECT  100900.0 241100.00000000003 101700.0 242700.0 ;
      RECT  100900.0 235300.0 101700.0 232899.99999999997 ;
      RECT  104100.0 235300.0 104900.0 232899.99999999997 ;
      RECT  105700.0 234500.0 106500.0 233200.0 ;
      RECT  105700.0 242399.99999999997 106500.0 241100.00000000003 ;
      RECT  100900.0 235300.0 101700.0 234500.0 ;
      RECT  102500.0 235300.0 103300.00000000001 234500.0 ;
      RECT  102500.0 235300.0 103300.00000000001 234500.0 ;
      RECT  100900.0 235300.0 101700.0 234500.0 ;
      RECT  102500.0 235300.0 103300.00000000001 234500.0 ;
      RECT  104100.0 235300.0 104900.0 234500.0 ;
      RECT  104100.0 235300.0 104900.0 234500.0 ;
      RECT  102500.0 235300.0 103300.00000000001 234500.0 ;
      RECT  100900.0 241100.00000000003 101700.0 240300.0 ;
      RECT  102500.0 241100.00000000003 103300.00000000001 240300.0 ;
      RECT  102500.0 241100.00000000003 103300.00000000001 240300.0 ;
      RECT  100900.0 241100.00000000003 101700.0 240300.0 ;
      RECT  102500.0 241100.00000000003 103300.00000000001 240300.0 ;
      RECT  104100.0 241100.00000000003 104900.0 240300.0 ;
      RECT  104100.0 241100.00000000003 104900.0 240300.0 ;
      RECT  102500.0 241100.00000000003 103300.00000000001 240300.0 ;
      RECT  105700.0 234899.99999999997 106500.0 234100.00000000003 ;
      RECT  105700.0 241500.0 106500.0 240700.0 ;
      RECT  104100.0 239399.99999999997 103300.00000000001 238600.00000000003 ;
      RECT  102100.0 238000.0 101300.00000000001 237200.0 ;
      RECT  102500.0 235300.0 103300.00000000001 234500.0 ;
      RECT  104100.0 241100.00000000003 104900.0 240300.0 ;
      RECT  106300.00000000001 238000.0 105500.0 237200.0 ;
      RECT  101300.00000000001 238000.0 102100.0 237200.0 ;
      RECT  103300.00000000001 239399.99999999997 104100.0 238600.00000000003 ;
      RECT  105500.0 238000.0 106300.00000000001 237200.0 ;
      RECT  99700.0 233500.0 109300.00000000001 232899.99999999997 ;
      RECT  99700.0 242700.0 109300.00000000001 242100.00000000003 ;
      RECT  94800.00000000001 212600.00000000003 94000.0 213399.99999999997 ;
      RECT  83100.0 209600.00000000003 82300.0 210399.99999999997 ;
      RECT  96200.0 221800.0 95400.0 222600.00000000003 ;
      RECT  84500.0 219200.0 83700.0 220000.0 ;
      RECT  83100.0 225000.0 82300.0 225800.0 ;
      RECT  97600.0 225000.0 96800.0 225800.0 ;
      RECT  84500.0 234200.0 83700.0 235000.0 ;
      RECT  99000.0 234200.0 98200.0 235000.0 ;
      RECT  94800.00000000001 210000.0 94000.0 210800.0 ;
      RECT  96200.0 208600.00000000003 95400.0 209399.99999999997 ;
      RECT  97600.0 218800.0 96800.0 219600.00000000003 ;
      RECT  96200.0 220200.0 95400.0 221000.0 ;
      RECT  94800.00000000001 228399.99999999997 94000.0 229200.0 ;
      RECT  99000.0 227000.0 98200.0 227800.0 ;
      RECT  97600.0 237200.0 96800.0 238000.0 ;
      RECT  99000.0 238600.00000000003 98200.0 239399.99999999997 ;
      RECT  91700.0 214399.99999999997 90900.0 215200.0 ;
      RECT  109100.0 214399.99999999997 108300.0 215200.0 ;
      RECT  91700.0 205200.0 90900.0 206000.0 ;
      RECT  109100.0 205200.0 108300.0 206000.0 ;
      RECT  91700.0 214399.99999999997 90900.0 215200.0 ;
      RECT  109100.0 214399.99999999997 108300.0 215200.0 ;
      RECT  91700.0 223600.00000000003 90900.0 224399.99999999997 ;
      RECT  109100.0 223600.00000000003 108300.0 224399.99999999997 ;
      RECT  91700.0 232800.0 90900.0 233600.00000000003 ;
      RECT  109100.0 232800.0 108300.0 233600.00000000003 ;
      RECT  91700.0 223600.00000000003 90900.0 224399.99999999997 ;
      RECT  109100.0 223600.00000000003 108300.0 224399.99999999997 ;
      RECT  91700.0 232800.0 90900.0 233600.00000000003 ;
      RECT  109100.0 232800.0 108300.0 233600.00000000003 ;
      RECT  91700.0 242000.0 90900.0 242800.0 ;
      RECT  109100.0 242000.0 108300.0 242800.0 ;
      RECT  112600.0 209700.0 113200.0 210300.0 ;
      RECT  112600.0 219300.0 113200.0 219899.99999999997 ;
      RECT  112600.0 228100.00000000003 113200.0 228700.0 ;
      RECT  112600.0 237700.0 113200.0 238300.0 ;
      RECT  128100.00000000003 170100.00000000003 128900.0 168500.0 ;
      RECT  128100.00000000003 175900.0 128900.0 178300.0 ;
      RECT  131300.0 175900.0 132100.00000000003 178300.0 ;
      RECT  132900.0 176700.0 133700.0 178000.0 ;
      RECT  132900.0 168800.0 133700.0 170100.00000000003 ;
      RECT  128100.00000000003 175900.0 128900.0 176700.0 ;
      RECT  129699.99999999999 175900.0 130500.0 176700.0 ;
      RECT  129699.99999999999 175900.0 130500.0 176700.0 ;
      RECT  128100.00000000003 175900.0 128900.0 176700.0 ;
      RECT  129699.99999999999 175900.0 130500.0 176700.0 ;
      RECT  131300.0 175900.0 132100.00000000003 176700.0 ;
      RECT  131300.0 175900.0 132100.00000000003 176700.0 ;
      RECT  129699.99999999999 175900.0 130500.0 176700.0 ;
      RECT  128100.00000000003 170100.00000000003 128900.0 170900.0 ;
      RECT  129699.99999999999 170100.00000000003 130500.0 170900.0 ;
      RECT  129699.99999999999 170100.00000000003 130500.0 170900.0 ;
      RECT  128100.00000000003 170100.00000000003 128900.0 170900.0 ;
      RECT  129699.99999999999 170100.00000000003 130500.0 170900.0 ;
      RECT  131300.0 170100.00000000003 132100.00000000003 170900.0 ;
      RECT  131300.0 170100.00000000003 132100.00000000003 170900.0 ;
      RECT  129699.99999999999 170100.00000000003 130500.0 170900.0 ;
      RECT  132900.0 176300.0 133700.0 177100.00000000003 ;
      RECT  132900.0 169700.0 133700.0 170500.0 ;
      RECT  131300.0 171800.0 130500.0 172600.00000000003 ;
      RECT  129300.00000000001 173200.0 128500.0 174000.0 ;
      RECT  129699.99999999999 175900.0 130500.0 176700.0 ;
      RECT  131300.0 170100.00000000003 132100.00000000003 170900.0 ;
      RECT  133500.0 173200.0 132700.0 174000.0 ;
      RECT  128500.0 173200.0 129300.00000000001 174000.0 ;
      RECT  130500.0 171800.0 131300.0 172600.00000000003 ;
      RECT  132700.0 173200.0 133500.0 174000.0 ;
      RECT  126900.0 177700.0 136500.0 178300.0 ;
      RECT  126900.0 168500.0 136500.0 169100.00000000003 ;
      RECT  128100.00000000003 185900.0 128900.0 187500.0 ;
      RECT  128100.00000000003 180100.00000000003 128900.0 177700.0 ;
      RECT  131300.0 180100.00000000003 132100.00000000003 177700.0 ;
      RECT  132900.0 179300.0 133700.0 178000.0 ;
      RECT  132900.0 187200.0 133700.0 185900.0 ;
      RECT  128100.00000000003 180100.00000000003 128900.0 179300.0 ;
      RECT  129699.99999999999 180100.00000000003 130500.0 179300.0 ;
      RECT  129699.99999999999 180100.00000000003 130500.0 179300.0 ;
      RECT  128100.00000000003 180100.00000000003 128900.0 179300.0 ;
      RECT  129699.99999999999 180100.00000000003 130500.0 179300.0 ;
      RECT  131300.0 180100.00000000003 132100.00000000003 179300.0 ;
      RECT  131300.0 180100.00000000003 132100.00000000003 179300.0 ;
      RECT  129699.99999999999 180100.00000000003 130500.0 179300.0 ;
      RECT  128100.00000000003 185900.0 128900.0 185100.00000000003 ;
      RECT  129699.99999999999 185900.0 130500.0 185100.00000000003 ;
      RECT  129699.99999999999 185900.0 130500.0 185100.00000000003 ;
      RECT  128100.00000000003 185900.0 128900.0 185100.00000000003 ;
      RECT  129699.99999999999 185900.0 130500.0 185100.00000000003 ;
      RECT  131300.0 185900.0 132100.00000000003 185100.00000000003 ;
      RECT  131300.0 185900.0 132100.00000000003 185100.00000000003 ;
      RECT  129699.99999999999 185900.0 130500.0 185100.00000000003 ;
      RECT  132900.0 179700.0 133700.0 178900.0 ;
      RECT  132900.0 186300.0 133700.0 185500.0 ;
      RECT  131300.0 184200.0 130500.0 183400.0 ;
      RECT  129300.00000000001 182800.0 128500.0 182000.0 ;
      RECT  129699.99999999999 180100.00000000003 130500.0 179300.0 ;
      RECT  131300.0 185900.0 132100.00000000003 185100.00000000003 ;
      RECT  133500.0 182800.0 132700.0 182000.0 ;
      RECT  128500.0 182800.0 129300.00000000001 182000.0 ;
      RECT  130500.0 184200.0 131300.0 183400.0 ;
      RECT  132700.0 182800.0 133500.0 182000.0 ;
      RECT  126900.0 178300.0 136500.0 177700.0 ;
      RECT  126900.0 187500.0 136500.0 186900.0 ;
      RECT  128100.00000000003 188500.0 128900.0 186900.0 ;
      RECT  128100.00000000003 194300.0 128900.0 196700.0 ;
      RECT  131300.0 194300.0 132100.00000000003 196700.0 ;
      RECT  132900.0 195100.00000000003 133700.0 196400.0 ;
      RECT  132900.0 187200.0 133700.0 188500.0 ;
      RECT  128100.00000000003 194300.0 128900.0 195100.00000000003 ;
      RECT  129699.99999999999 194300.0 130500.0 195100.00000000003 ;
      RECT  129699.99999999999 194300.0 130500.0 195100.00000000003 ;
      RECT  128100.00000000003 194300.0 128900.0 195100.00000000003 ;
      RECT  129699.99999999999 194300.0 130500.0 195100.00000000003 ;
      RECT  131300.0 194300.0 132100.00000000003 195100.00000000003 ;
      RECT  131300.0 194300.0 132100.00000000003 195100.00000000003 ;
      RECT  129699.99999999999 194300.0 130500.0 195100.00000000003 ;
      RECT  128100.00000000003 188500.0 128900.0 189300.0 ;
      RECT  129699.99999999999 188500.0 130500.0 189300.0 ;
      RECT  129699.99999999999 188500.0 130500.0 189300.0 ;
      RECT  128100.00000000003 188500.0 128900.0 189300.0 ;
      RECT  129699.99999999999 188500.0 130500.0 189300.0 ;
      RECT  131300.0 188500.0 132100.00000000003 189300.0 ;
      RECT  131300.0 188500.0 132100.00000000003 189300.0 ;
      RECT  129699.99999999999 188500.0 130500.0 189300.0 ;
      RECT  132900.0 194700.0 133700.0 195500.0 ;
      RECT  132900.0 188100.00000000003 133700.0 188900.0 ;
      RECT  131300.0 190200.0 130500.0 191000.0 ;
      RECT  129300.00000000001 191600.00000000003 128500.0 192400.0 ;
      RECT  129699.99999999999 194300.0 130500.0 195100.00000000003 ;
      RECT  131300.0 188500.0 132100.00000000003 189300.0 ;
      RECT  133500.0 191600.00000000003 132700.0 192400.0 ;
      RECT  128500.0 191600.00000000003 129300.00000000001 192400.0 ;
      RECT  130500.0 190200.0 131300.0 191000.0 ;
      RECT  132700.0 191600.00000000003 133500.0 192400.0 ;
      RECT  126900.0 196100.00000000003 136500.0 196700.0 ;
      RECT  126900.0 186900.0 136500.0 187500.0 ;
      RECT  128100.00000000003 204300.0 128900.0 205899.99999999997 ;
      RECT  128100.00000000003 198500.0 128900.0 196100.00000000003 ;
      RECT  131300.0 198500.0 132100.00000000003 196100.00000000003 ;
      RECT  132900.0 197700.0 133700.0 196400.0 ;
      RECT  132900.0 205600.00000000003 133700.0 204300.0 ;
      RECT  128100.00000000003 198500.0 128900.0 197700.0 ;
      RECT  129699.99999999999 198500.0 130500.0 197700.0 ;
      RECT  129699.99999999999 198500.0 130500.0 197700.0 ;
      RECT  128100.00000000003 198500.0 128900.0 197700.0 ;
      RECT  129699.99999999999 198500.0 130500.0 197700.0 ;
      RECT  131300.0 198500.0 132100.00000000003 197700.0 ;
      RECT  131300.0 198500.0 132100.00000000003 197700.0 ;
      RECT  129699.99999999999 198500.0 130500.0 197700.0 ;
      RECT  128100.00000000003 204300.0 128900.0 203500.0 ;
      RECT  129699.99999999999 204300.0 130500.0 203500.0 ;
      RECT  129699.99999999999 204300.0 130500.0 203500.0 ;
      RECT  128100.00000000003 204300.0 128900.0 203500.0 ;
      RECT  129699.99999999999 204300.0 130500.0 203500.0 ;
      RECT  131300.0 204300.0 132100.00000000003 203500.0 ;
      RECT  131300.0 204300.0 132100.00000000003 203500.0 ;
      RECT  129699.99999999999 204300.0 130500.0 203500.0 ;
      RECT  132900.0 198100.00000000003 133700.0 197300.0 ;
      RECT  132900.0 204700.0 133700.0 203899.99999999997 ;
      RECT  131300.0 202600.00000000003 130500.0 201800.0 ;
      RECT  129300.00000000001 201200.0 128500.0 200399.99999999997 ;
      RECT  129699.99999999999 198500.0 130500.0 197700.0 ;
      RECT  131300.0 204300.0 132100.00000000003 203500.0 ;
      RECT  133500.0 201200.0 132700.0 200399.99999999997 ;
      RECT  128500.0 201200.0 129300.00000000001 200399.99999999997 ;
      RECT  130500.0 202600.00000000003 131300.0 201800.0 ;
      RECT  132700.0 201200.0 133500.0 200399.99999999997 ;
      RECT  126900.0 196700.0 136500.0 196100.00000000003 ;
      RECT  126900.0 205899.99999999997 136500.0 205300.0 ;
      RECT  128100.00000000003 206899.99999999997 128900.0 205300.0 ;
      RECT  128100.00000000003 212700.0 128900.0 215100.00000000003 ;
      RECT  131300.0 212700.0 132100.00000000003 215100.00000000003 ;
      RECT  132900.0 213500.0 133700.0 214800.0 ;
      RECT  132900.0 205600.00000000003 133700.0 206899.99999999997 ;
      RECT  128100.00000000003 212700.0 128900.0 213500.0 ;
      RECT  129699.99999999999 212700.0 130500.0 213500.0 ;
      RECT  129699.99999999999 212700.0 130500.0 213500.0 ;
      RECT  128100.00000000003 212700.0 128900.0 213500.0 ;
      RECT  129699.99999999999 212700.0 130500.0 213500.0 ;
      RECT  131300.0 212700.0 132100.00000000003 213500.0 ;
      RECT  131300.0 212700.0 132100.00000000003 213500.0 ;
      RECT  129699.99999999999 212700.0 130500.0 213500.0 ;
      RECT  128100.00000000003 206899.99999999997 128900.0 207700.0 ;
      RECT  129699.99999999999 206899.99999999997 130500.0 207700.0 ;
      RECT  129699.99999999999 206899.99999999997 130500.0 207700.0 ;
      RECT  128100.00000000003 206899.99999999997 128900.0 207700.0 ;
      RECT  129699.99999999999 206899.99999999997 130500.0 207700.0 ;
      RECT  131300.0 206899.99999999997 132100.00000000003 207700.0 ;
      RECT  131300.0 206899.99999999997 132100.00000000003 207700.0 ;
      RECT  129699.99999999999 206899.99999999997 130500.0 207700.0 ;
      RECT  132900.0 213100.00000000003 133700.0 213899.99999999997 ;
      RECT  132900.0 206500.0 133700.0 207300.0 ;
      RECT  131300.0 208600.00000000003 130500.0 209399.99999999997 ;
      RECT  129300.00000000001 210000.0 128500.0 210800.0 ;
      RECT  129699.99999999999 212700.0 130500.0 213500.0 ;
      RECT  131300.0 206899.99999999997 132100.00000000003 207700.0 ;
      RECT  133500.0 210000.0 132700.0 210800.0 ;
      RECT  128500.0 210000.0 129300.00000000001 210800.0 ;
      RECT  130500.0 208600.00000000003 131300.0 209399.99999999997 ;
      RECT  132700.0 210000.0 133500.0 210800.0 ;
      RECT  126900.0 214500.0 136500.0 215100.00000000003 ;
      RECT  126900.0 205300.0 136500.0 205899.99999999997 ;
      RECT  128100.00000000003 222700.0 128900.0 224300.0 ;
      RECT  128100.00000000003 216899.99999999997 128900.0 214500.0 ;
      RECT  131300.0 216899.99999999997 132100.00000000003 214500.0 ;
      RECT  132900.0 216100.00000000003 133700.0 214800.0 ;
      RECT  132900.0 224000.0 133700.0 222700.0 ;
      RECT  128100.00000000003 216899.99999999997 128900.0 216100.00000000003 ;
      RECT  129699.99999999999 216899.99999999997 130500.0 216100.00000000003 ;
      RECT  129699.99999999999 216899.99999999997 130500.0 216100.00000000003 ;
      RECT  128100.00000000003 216899.99999999997 128900.0 216100.00000000003 ;
      RECT  129699.99999999999 216899.99999999997 130500.0 216100.00000000003 ;
      RECT  131300.0 216899.99999999997 132100.00000000003 216100.00000000003 ;
      RECT  131300.0 216899.99999999997 132100.00000000003 216100.00000000003 ;
      RECT  129699.99999999999 216899.99999999997 130500.0 216100.00000000003 ;
      RECT  128100.00000000003 222700.0 128900.0 221899.99999999997 ;
      RECT  129699.99999999999 222700.0 130500.0 221899.99999999997 ;
      RECT  129699.99999999999 222700.0 130500.0 221899.99999999997 ;
      RECT  128100.00000000003 222700.0 128900.0 221899.99999999997 ;
      RECT  129699.99999999999 222700.0 130500.0 221899.99999999997 ;
      RECT  131300.0 222700.0 132100.00000000003 221899.99999999997 ;
      RECT  131300.0 222700.0 132100.00000000003 221899.99999999997 ;
      RECT  129699.99999999999 222700.0 130500.0 221899.99999999997 ;
      RECT  132900.0 216500.0 133700.0 215700.0 ;
      RECT  132900.0 223100.00000000003 133700.0 222300.0 ;
      RECT  131300.0 221000.0 130500.0 220200.0 ;
      RECT  129300.00000000001 219600.00000000003 128500.0 218800.0 ;
      RECT  129699.99999999999 216899.99999999997 130500.0 216100.00000000003 ;
      RECT  131300.0 222700.0 132100.00000000003 221899.99999999997 ;
      RECT  133500.0 219600.00000000003 132700.0 218800.0 ;
      RECT  128500.0 219600.00000000003 129300.00000000001 218800.0 ;
      RECT  130500.0 221000.0 131300.0 220200.0 ;
      RECT  132700.0 219600.00000000003 133500.0 218800.0 ;
      RECT  126900.0 215100.00000000003 136500.0 214500.0 ;
      RECT  126900.0 224300.0 136500.0 223700.0 ;
      RECT  128100.00000000003 225300.0 128900.0 223700.0 ;
      RECT  128100.00000000003 231100.00000000003 128900.0 233500.0 ;
      RECT  131300.0 231100.00000000003 132100.00000000003 233500.0 ;
      RECT  132900.0 231899.99999999997 133700.0 233200.0 ;
      RECT  132900.0 224000.0 133700.0 225300.0 ;
      RECT  128100.00000000003 231100.00000000003 128900.0 231899.99999999997 ;
      RECT  129699.99999999999 231100.00000000003 130500.0 231899.99999999997 ;
      RECT  129699.99999999999 231100.00000000003 130500.0 231899.99999999997 ;
      RECT  128100.00000000003 231100.00000000003 128900.0 231899.99999999997 ;
      RECT  129699.99999999999 231100.00000000003 130500.0 231899.99999999997 ;
      RECT  131300.0 231100.00000000003 132100.00000000003 231899.99999999997 ;
      RECT  131300.0 231100.00000000003 132100.00000000003 231899.99999999997 ;
      RECT  129699.99999999999 231100.00000000003 130500.0 231899.99999999997 ;
      RECT  128100.00000000003 225300.0 128900.0 226100.00000000003 ;
      RECT  129699.99999999999 225300.0 130500.0 226100.00000000003 ;
      RECT  129699.99999999999 225300.0 130500.0 226100.00000000003 ;
      RECT  128100.00000000003 225300.0 128900.0 226100.00000000003 ;
      RECT  129699.99999999999 225300.0 130500.0 226100.00000000003 ;
      RECT  131300.0 225300.0 132100.00000000003 226100.00000000003 ;
      RECT  131300.0 225300.0 132100.00000000003 226100.00000000003 ;
      RECT  129699.99999999999 225300.0 130500.0 226100.00000000003 ;
      RECT  132900.0 231500.0 133700.0 232300.0 ;
      RECT  132900.0 224899.99999999997 133700.0 225700.0 ;
      RECT  131300.0 227000.0 130500.0 227800.0 ;
      RECT  129300.00000000001 228399.99999999997 128500.0 229200.0 ;
      RECT  129699.99999999999 231100.00000000003 130500.0 231899.99999999997 ;
      RECT  131300.0 225300.0 132100.00000000003 226100.00000000003 ;
      RECT  133500.0 228399.99999999997 132700.0 229200.0 ;
      RECT  128500.0 228399.99999999997 129300.00000000001 229200.0 ;
      RECT  130500.0 227000.0 131300.0 227800.0 ;
      RECT  132700.0 228399.99999999997 133500.0 229200.0 ;
      RECT  126900.0 232899.99999999997 136500.0 233500.0 ;
      RECT  126900.0 223700.0 136500.0 224300.0 ;
      RECT  128100.00000000003 241100.00000000003 128900.0 242700.0 ;
      RECT  128100.00000000003 235300.0 128900.0 232900.00000000003 ;
      RECT  131300.0 235300.0 132100.00000000003 232900.00000000003 ;
      RECT  132900.0 234500.0 133700.0 233200.0 ;
      RECT  132900.0 242400.00000000003 133700.0 241100.00000000003 ;
      RECT  128100.00000000003 235300.0 128900.0 234500.0 ;
      RECT  129699.99999999999 235300.0 130500.0 234500.0 ;
      RECT  129699.99999999999 235300.0 130500.0 234500.0 ;
      RECT  128100.00000000003 235300.0 128900.0 234500.0 ;
      RECT  129699.99999999999 235300.0 130500.0 234500.0 ;
      RECT  131300.0 235300.0 132100.00000000003 234500.0 ;
      RECT  131300.0 235300.0 132100.00000000003 234500.0 ;
      RECT  129699.99999999999 235300.0 130500.0 234500.0 ;
      RECT  128100.00000000003 241100.00000000003 128900.0 240300.0 ;
      RECT  129699.99999999999 241100.00000000003 130500.0 240300.0 ;
      RECT  129699.99999999999 241100.00000000003 130500.0 240300.0 ;
      RECT  128100.00000000003 241100.00000000003 128900.0 240300.0 ;
      RECT  129699.99999999999 241100.00000000003 130500.0 240300.0 ;
      RECT  131300.0 241100.00000000003 132100.00000000003 240300.0 ;
      RECT  131300.0 241100.00000000003 132100.00000000003 240300.0 ;
      RECT  129699.99999999999 241100.00000000003 130500.0 240300.0 ;
      RECT  132900.0 234900.00000000003 133700.0 234100.00000000003 ;
      RECT  132900.0 241500.0 133700.0 240700.0 ;
      RECT  131300.0 239400.00000000003 130500.0 238600.00000000003 ;
      RECT  129300.00000000001 238000.0 128500.0 237200.0 ;
      RECT  129699.99999999999 235300.0 130500.0 234500.0 ;
      RECT  131300.0 241100.00000000003 132100.00000000003 240300.0 ;
      RECT  133500.0 238000.0 132700.0 237200.0 ;
      RECT  128500.0 238000.0 129300.00000000001 237200.0 ;
      RECT  130500.0 239400.00000000003 131300.0 238600.00000000003 ;
      RECT  132700.0 238000.0 133500.0 237200.0 ;
      RECT  126900.0 233500.0 136500.0 232900.00000000003 ;
      RECT  126900.0 242700.0 136500.0 242100.00000000003 ;
      RECT  128100.00000000003 243700.0 128900.0 242100.00000000003 ;
      RECT  128100.00000000003 249500.0 128900.0 251900.00000000003 ;
      RECT  131300.0 249500.0 132100.00000000003 251900.00000000003 ;
      RECT  132900.0 250300.0 133700.0 251600.00000000003 ;
      RECT  132900.0 242400.00000000003 133700.0 243700.0 ;
      RECT  128100.00000000003 249500.0 128900.0 250300.0 ;
      RECT  129699.99999999999 249500.0 130500.0 250300.0 ;
      RECT  129699.99999999999 249500.0 130500.0 250300.0 ;
      RECT  128100.00000000003 249500.0 128900.0 250300.0 ;
      RECT  129699.99999999999 249500.0 130500.0 250300.0 ;
      RECT  131300.0 249500.0 132100.00000000003 250300.0 ;
      RECT  131300.0 249500.0 132100.00000000003 250300.0 ;
      RECT  129699.99999999999 249500.0 130500.0 250300.0 ;
      RECT  128100.00000000003 243700.0 128900.0 244500.0 ;
      RECT  129699.99999999999 243700.0 130500.0 244500.0 ;
      RECT  129699.99999999999 243700.0 130500.0 244500.0 ;
      RECT  128100.00000000003 243700.0 128900.0 244500.0 ;
      RECT  129699.99999999999 243700.0 130500.0 244500.0 ;
      RECT  131300.0 243700.0 132100.00000000003 244500.0 ;
      RECT  131300.0 243700.0 132100.00000000003 244500.0 ;
      RECT  129699.99999999999 243700.0 130500.0 244500.0 ;
      RECT  132900.0 249900.00000000003 133700.0 250700.0 ;
      RECT  132900.0 243300.0 133700.0 244100.00000000003 ;
      RECT  131300.0 245400.00000000003 130500.0 246200.0 ;
      RECT  129300.00000000001 246800.0 128500.0 247600.00000000003 ;
      RECT  129699.99999999999 249500.0 130500.0 250300.0 ;
      RECT  131300.0 243700.0 132100.00000000003 244500.0 ;
      RECT  133500.0 246800.0 132700.0 247600.00000000003 ;
      RECT  128500.0 246800.0 129300.00000000001 247600.00000000003 ;
      RECT  130500.0 245400.00000000003 131300.0 246200.0 ;
      RECT  132700.0 246800.0 133500.0 247600.00000000003 ;
      RECT  126900.0 251300.0 136500.0 251900.00000000003 ;
      RECT  126900.0 242100.00000000003 136500.0 242700.0 ;
      RECT  128100.00000000003 259500.0 128900.0 261100.00000000003 ;
      RECT  128100.00000000003 253700.0 128900.0 251300.0 ;
      RECT  131300.0 253700.0 132100.00000000003 251300.0 ;
      RECT  132900.0 252899.99999999997 133700.0 251600.00000000003 ;
      RECT  132900.0 260800.0 133700.0 259500.0 ;
      RECT  128100.00000000003 253700.0 128900.0 252899.99999999997 ;
      RECT  129699.99999999999 253700.0 130500.0 252899.99999999997 ;
      RECT  129699.99999999999 253700.0 130500.0 252899.99999999997 ;
      RECT  128100.00000000003 253700.0 128900.0 252899.99999999997 ;
      RECT  129699.99999999999 253700.0 130500.0 252899.99999999997 ;
      RECT  131300.0 253700.0 132100.00000000003 252899.99999999997 ;
      RECT  131300.0 253700.0 132100.00000000003 252899.99999999997 ;
      RECT  129699.99999999999 253700.0 130500.0 252899.99999999997 ;
      RECT  128100.00000000003 259500.0 128900.0 258700.0 ;
      RECT  129699.99999999999 259500.0 130500.0 258700.0 ;
      RECT  129699.99999999999 259500.0 130500.0 258700.0 ;
      RECT  128100.00000000003 259500.0 128900.0 258700.0 ;
      RECT  129699.99999999999 259500.0 130500.0 258700.0 ;
      RECT  131300.0 259500.0 132100.00000000003 258700.0 ;
      RECT  131300.0 259500.0 132100.00000000003 258700.0 ;
      RECT  129699.99999999999 259500.0 130500.0 258700.0 ;
      RECT  132900.0 253300.0 133700.0 252500.0 ;
      RECT  132900.0 259899.99999999997 133700.0 259100.00000000003 ;
      RECT  131300.0 257800.0 130500.0 257000.0 ;
      RECT  129300.00000000001 256399.99999999997 128500.0 255600.00000000003 ;
      RECT  129699.99999999999 253700.0 130500.0 252899.99999999997 ;
      RECT  131300.0 259500.0 132100.00000000003 258700.0 ;
      RECT  133500.0 256399.99999999997 132700.0 255600.00000000003 ;
      RECT  128500.0 256399.99999999997 129300.00000000001 255600.00000000003 ;
      RECT  130500.0 257800.0 131300.0 257000.0 ;
      RECT  132700.0 256399.99999999997 133500.0 255600.00000000003 ;
      RECT  126900.0 251899.99999999997 136500.0 251300.0 ;
      RECT  126900.0 261100.00000000003 136500.0 260500.0 ;
      RECT  128100.00000000003 262100.00000000003 128900.0 260500.0 ;
      RECT  128100.00000000003 267900.0 128900.0 270300.0 ;
      RECT  131300.0 267900.0 132100.00000000003 270300.0 ;
      RECT  132900.0 268700.0 133700.0 270000.0 ;
      RECT  132900.0 260800.0 133700.0 262100.00000000003 ;
      RECT  128100.00000000003 267900.0 128900.0 268700.0 ;
      RECT  129699.99999999999 267900.0 130500.0 268700.0 ;
      RECT  129699.99999999999 267900.0 130500.0 268700.0 ;
      RECT  128100.00000000003 267900.0 128900.0 268700.0 ;
      RECT  129699.99999999999 267900.0 130500.0 268700.0 ;
      RECT  131300.0 267900.0 132100.00000000003 268700.0 ;
      RECT  131300.0 267900.0 132100.00000000003 268700.0 ;
      RECT  129699.99999999999 267900.0 130500.0 268700.0 ;
      RECT  128100.00000000003 262100.00000000003 128900.0 262900.0 ;
      RECT  129699.99999999999 262100.00000000003 130500.0 262900.0 ;
      RECT  129699.99999999999 262100.00000000003 130500.0 262900.0 ;
      RECT  128100.00000000003 262100.00000000003 128900.0 262900.0 ;
      RECT  129699.99999999999 262100.00000000003 130500.0 262900.0 ;
      RECT  131300.0 262100.00000000003 132100.00000000003 262900.0 ;
      RECT  131300.0 262100.00000000003 132100.00000000003 262900.0 ;
      RECT  129699.99999999999 262100.00000000003 130500.0 262900.0 ;
      RECT  132900.0 268300.0 133700.0 269100.0 ;
      RECT  132900.0 261700.0 133700.0 262500.0 ;
      RECT  131300.0 263800.0 130500.0 264600.0 ;
      RECT  129300.00000000001 265200.0 128500.0 266000.0 ;
      RECT  129699.99999999999 267900.0 130500.0 268700.0 ;
      RECT  131300.0 262100.00000000003 132100.00000000003 262900.0 ;
      RECT  133500.0 265200.0 132700.0 266000.0 ;
      RECT  128500.0 265200.0 129300.00000000001 266000.0 ;
      RECT  130500.0 263800.0 131300.0 264600.0 ;
      RECT  132700.0 265200.0 133500.0 266000.0 ;
      RECT  126900.0 269700.0 136500.0 270300.0 ;
      RECT  126900.0 260500.0 136500.0 261100.00000000003 ;
      RECT  128100.00000000003 277900.00000000006 128900.0 279500.0 ;
      RECT  128100.00000000003 272100.0 128900.0 269700.0 ;
      RECT  131300.0 272100.0 132100.00000000003 269700.0 ;
      RECT  132900.0 271300.0 133700.0 270000.0 ;
      RECT  132900.0 279200.0 133700.0 277900.00000000006 ;
      RECT  128100.00000000003 272100.0 128900.0 271300.0 ;
      RECT  129699.99999999999 272100.0 130500.0 271300.0 ;
      RECT  129699.99999999999 272100.0 130500.0 271300.0 ;
      RECT  128100.00000000003 272100.0 128900.0 271300.0 ;
      RECT  129699.99999999999 272100.0 130500.0 271300.0 ;
      RECT  131300.0 272100.0 132100.00000000003 271300.0 ;
      RECT  131300.0 272100.0 132100.00000000003 271300.0 ;
      RECT  129699.99999999999 272100.0 130500.0 271300.0 ;
      RECT  128100.00000000003 277900.00000000006 128900.0 277100.0 ;
      RECT  129699.99999999999 277900.00000000006 130500.0 277100.0 ;
      RECT  129699.99999999999 277900.00000000006 130500.0 277100.0 ;
      RECT  128100.00000000003 277900.00000000006 128900.0 277100.0 ;
      RECT  129699.99999999999 277900.00000000006 130500.0 277100.0 ;
      RECT  131300.0 277900.00000000006 132100.00000000003 277100.0 ;
      RECT  131300.0 277900.00000000006 132100.00000000003 277100.0 ;
      RECT  129699.99999999999 277900.00000000006 130500.0 277100.0 ;
      RECT  132900.0 271700.0 133700.0 270900.00000000006 ;
      RECT  132900.0 278300.0 133700.0 277500.0 ;
      RECT  131300.0 276200.0 130500.0 275400.00000000006 ;
      RECT  129300.00000000001 274800.0 128500.0 274000.0 ;
      RECT  129699.99999999999 272100.0 130500.0 271300.0 ;
      RECT  131300.0 277900.00000000006 132100.00000000003 277100.0 ;
      RECT  133500.0 274800.0 132700.0 274000.0 ;
      RECT  128500.0 274800.0 129300.00000000001 274000.0 ;
      RECT  130500.0 276200.0 131300.0 275400.00000000006 ;
      RECT  132700.0 274800.0 133500.0 274000.0 ;
      RECT  126900.0 270300.0 136500.0 269700.0 ;
      RECT  126900.0 279500.0 136500.0 278900.00000000006 ;
      RECT  128100.00000000003 280500.0 128900.0 278900.00000000006 ;
      RECT  128100.00000000003 286300.0 128900.0 288700.0 ;
      RECT  131300.0 286300.0 132100.00000000003 288700.0 ;
      RECT  132900.0 287100.0 133700.0 288400.00000000006 ;
      RECT  132900.0 279200.0 133700.0 280500.0 ;
      RECT  128100.00000000003 286300.0 128900.0 287100.0 ;
      RECT  129699.99999999999 286300.0 130500.0 287100.0 ;
      RECT  129699.99999999999 286300.0 130500.0 287100.0 ;
      RECT  128100.00000000003 286300.0 128900.0 287100.0 ;
      RECT  129699.99999999999 286300.0 130500.0 287100.0 ;
      RECT  131300.0 286300.0 132100.00000000003 287100.0 ;
      RECT  131300.0 286300.0 132100.00000000003 287100.0 ;
      RECT  129699.99999999999 286300.0 130500.0 287100.0 ;
      RECT  128100.00000000003 280500.0 128900.0 281300.0 ;
      RECT  129699.99999999999 280500.0 130500.0 281300.0 ;
      RECT  129699.99999999999 280500.0 130500.0 281300.0 ;
      RECT  128100.00000000003 280500.0 128900.0 281300.0 ;
      RECT  129699.99999999999 280500.0 130500.0 281300.0 ;
      RECT  131300.0 280500.0 132100.00000000003 281300.0 ;
      RECT  131300.0 280500.0 132100.00000000003 281300.0 ;
      RECT  129699.99999999999 280500.0 130500.0 281300.0 ;
      RECT  132900.0 286700.0 133700.0 287500.0 ;
      RECT  132900.0 280100.0 133700.0 280900.00000000006 ;
      RECT  131300.0 282200.0 130500.0 283000.0 ;
      RECT  129300.00000000001 283600.0 128500.0 284400.00000000006 ;
      RECT  129699.99999999999 286300.0 130500.0 287100.0 ;
      RECT  131300.0 280500.0 132100.00000000003 281300.0 ;
      RECT  133500.0 283600.0 132700.0 284400.00000000006 ;
      RECT  128500.0 283600.0 129300.00000000001 284400.00000000006 ;
      RECT  130500.0 282200.0 131300.0 283000.0 ;
      RECT  132700.0 283600.0 133500.0 284400.00000000006 ;
      RECT  126900.0 288100.0 136500.0 288700.0 ;
      RECT  126900.0 278900.00000000006 136500.0 279500.0 ;
      RECT  128100.00000000003 296300.0 128900.0 297900.00000000006 ;
      RECT  128100.00000000003 290500.0 128900.0 288100.0 ;
      RECT  131300.0 290500.0 132100.00000000003 288100.0 ;
      RECT  132900.0 289700.0 133700.0 288400.00000000006 ;
      RECT  132900.0 297600.0 133700.0 296300.0 ;
      RECT  128100.00000000003 290500.0 128900.0 289700.0 ;
      RECT  129699.99999999999 290500.0 130500.0 289700.0 ;
      RECT  129699.99999999999 290500.0 130500.0 289700.0 ;
      RECT  128100.00000000003 290500.0 128900.0 289700.0 ;
      RECT  129699.99999999999 290500.0 130500.0 289700.0 ;
      RECT  131300.0 290500.0 132100.00000000003 289700.0 ;
      RECT  131300.0 290500.0 132100.00000000003 289700.0 ;
      RECT  129699.99999999999 290500.0 130500.0 289700.0 ;
      RECT  128100.00000000003 296300.0 128900.0 295500.0 ;
      RECT  129699.99999999999 296300.0 130500.0 295500.0 ;
      RECT  129699.99999999999 296300.0 130500.0 295500.0 ;
      RECT  128100.00000000003 296300.0 128900.0 295500.0 ;
      RECT  129699.99999999999 296300.0 130500.0 295500.0 ;
      RECT  131300.0 296300.0 132100.00000000003 295500.0 ;
      RECT  131300.0 296300.0 132100.00000000003 295500.0 ;
      RECT  129699.99999999999 296300.0 130500.0 295500.0 ;
      RECT  132900.0 290100.0 133700.0 289300.0 ;
      RECT  132900.0 296700.0 133700.0 295900.00000000006 ;
      RECT  131300.0 294600.0 130500.0 293800.0 ;
      RECT  129300.00000000001 293200.0 128500.0 292400.00000000006 ;
      RECT  129699.99999999999 290500.0 130500.0 289700.0 ;
      RECT  131300.0 296300.0 132100.00000000003 295500.0 ;
      RECT  133500.0 293200.0 132700.0 292400.00000000006 ;
      RECT  128500.0 293200.0 129300.00000000001 292400.00000000006 ;
      RECT  130500.0 294600.0 131300.0 293800.0 ;
      RECT  132700.0 293200.0 133500.0 292400.00000000006 ;
      RECT  126900.0 288700.0 136500.0 288100.0 ;
      RECT  126900.0 297900.00000000006 136500.0 297300.0 ;
      RECT  128100.00000000003 298900.00000000006 128900.0 297300.0 ;
      RECT  128100.00000000003 304700.0 128900.0 307100.0 ;
      RECT  131300.0 304700.0 132100.00000000003 307100.0 ;
      RECT  132900.0 305500.0 133700.0 306800.0 ;
      RECT  132900.0 297600.0 133700.0 298900.00000000006 ;
      RECT  128100.00000000003 304700.0 128900.0 305500.0 ;
      RECT  129699.99999999999 304700.0 130500.0 305500.0 ;
      RECT  129699.99999999999 304700.0 130500.0 305500.0 ;
      RECT  128100.00000000003 304700.0 128900.0 305500.0 ;
      RECT  129699.99999999999 304700.0 130500.0 305500.0 ;
      RECT  131300.0 304700.0 132100.00000000003 305500.0 ;
      RECT  131300.0 304700.0 132100.00000000003 305500.0 ;
      RECT  129699.99999999999 304700.0 130500.0 305500.0 ;
      RECT  128100.00000000003 298900.00000000006 128900.0 299700.0 ;
      RECT  129699.99999999999 298900.00000000006 130500.0 299700.0 ;
      RECT  129699.99999999999 298900.00000000006 130500.0 299700.0 ;
      RECT  128100.00000000003 298900.00000000006 128900.0 299700.0 ;
      RECT  129699.99999999999 298900.00000000006 130500.0 299700.0 ;
      RECT  131300.0 298900.00000000006 132100.00000000003 299700.0 ;
      RECT  131300.0 298900.00000000006 132100.00000000003 299700.0 ;
      RECT  129699.99999999999 298900.00000000006 130500.0 299700.0 ;
      RECT  132900.0 305100.0 133700.0 305900.00000000006 ;
      RECT  132900.0 298500.0 133700.0 299300.0 ;
      RECT  131300.0 300600.0 130500.0 301400.00000000006 ;
      RECT  129300.00000000001 302000.0 128500.0 302800.0 ;
      RECT  129699.99999999999 304700.0 130500.0 305500.0 ;
      RECT  131300.0 298900.00000000006 132100.00000000003 299700.0 ;
      RECT  133500.0 302000.0 132700.0 302800.0 ;
      RECT  128500.0 302000.0 129300.00000000001 302800.0 ;
      RECT  130500.0 300600.0 131300.0 301400.00000000006 ;
      RECT  132700.0 302000.0 133500.0 302800.0 ;
      RECT  126900.0 306500.0 136500.0 307100.0 ;
      RECT  126900.0 297300.0 136500.0 297900.00000000006 ;
      RECT  128100.00000000003 314700.0 128900.0 316300.0 ;
      RECT  128100.00000000003 308900.00000000006 128900.0 306500.0 ;
      RECT  131300.0 308900.00000000006 132100.00000000003 306500.0 ;
      RECT  132900.0 308100.0 133700.0 306800.0 ;
      RECT  132900.0 316000.0 133700.0 314700.0 ;
      RECT  128100.00000000003 308900.00000000006 128900.0 308100.0 ;
      RECT  129699.99999999999 308900.00000000006 130500.0 308100.0 ;
      RECT  129699.99999999999 308900.00000000006 130500.0 308100.0 ;
      RECT  128100.00000000003 308900.00000000006 128900.0 308100.0 ;
      RECT  129699.99999999999 308900.00000000006 130500.0 308100.0 ;
      RECT  131300.0 308900.00000000006 132100.00000000003 308100.0 ;
      RECT  131300.0 308900.00000000006 132100.00000000003 308100.0 ;
      RECT  129699.99999999999 308900.00000000006 130500.0 308100.0 ;
      RECT  128100.00000000003 314700.0 128900.0 313900.00000000006 ;
      RECT  129699.99999999999 314700.0 130500.0 313900.00000000006 ;
      RECT  129699.99999999999 314700.0 130500.0 313900.00000000006 ;
      RECT  128100.00000000003 314700.0 128900.0 313900.00000000006 ;
      RECT  129699.99999999999 314700.0 130500.0 313900.00000000006 ;
      RECT  131300.0 314700.0 132100.00000000003 313900.00000000006 ;
      RECT  131300.0 314700.0 132100.00000000003 313900.00000000006 ;
      RECT  129699.99999999999 314700.0 130500.0 313900.00000000006 ;
      RECT  132900.0 308500.0 133700.0 307700.0 ;
      RECT  132900.0 315100.0 133700.0 314300.0 ;
      RECT  131300.0 313000.0 130500.0 312200.0 ;
      RECT  129300.00000000001 311600.0 128500.0 310800.0 ;
      RECT  129699.99999999999 308900.00000000006 130500.0 308100.0 ;
      RECT  131300.0 314700.0 132100.00000000003 313900.00000000006 ;
      RECT  133500.0 311600.0 132700.0 310800.0 ;
      RECT  128500.0 311600.0 129300.00000000001 310800.0 ;
      RECT  130500.0 313000.0 131300.0 312200.0 ;
      RECT  132700.0 311600.0 133500.0 310800.0 ;
      RECT  126900.0 307100.0 136500.0 306500.0 ;
      RECT  126900.0 316300.0 136500.0 315700.0 ;
      RECT  140900.0 176700.0 141700.0 178000.0 ;
      RECT  140900.0 168800.0 141700.0 170100.00000000003 ;
      RECT  137700.0 169700.0 138500.0 168500.0 ;
      RECT  137700.0 175900.0 138500.0 178300.0 ;
      RECT  139500.0 169700.0 140100.0 175900.0 ;
      RECT  137700.0 175900.0 138500.0 176700.0 ;
      RECT  139300.0 175900.0 140100.0 176700.0 ;
      RECT  139300.0 175900.0 140100.0 176700.0 ;
      RECT  137700.0 175900.0 138500.0 176700.0 ;
      RECT  137700.0 169700.0 138500.0 170500.0 ;
      RECT  139300.0 169700.0 140100.0 170500.0 ;
      RECT  139300.0 169700.0 140100.0 170500.0 ;
      RECT  137700.0 169700.0 138500.0 170500.0 ;
      RECT  140900.0 176300.0 141700.0 177100.00000000003 ;
      RECT  140900.0 169700.0 141700.0 170500.0 ;
      RECT  138100.0 172800.0 138900.0 173600.00000000003 ;
      RECT  138100.0 172800.0 138900.0 173600.00000000003 ;
      RECT  139800.0 172900.0 140400.0 173500.0 ;
      RECT  136500.0 177700.0 142900.0 178300.0 ;
      RECT  136500.0 168500.0 142900.0 169100.00000000003 ;
      RECT  140900.0 179300.0 141700.0 178000.0 ;
      RECT  140900.0 187200.0 141700.0 185900.0 ;
      RECT  137700.0 186300.0 138500.0 187500.0 ;
      RECT  137700.0 180100.00000000003 138500.0 177700.0 ;
      RECT  139500.0 186300.0 140100.0 180100.00000000003 ;
      RECT  137700.0 180100.00000000003 138500.0 179300.0 ;
      RECT  139300.0 180100.00000000003 140100.0 179300.0 ;
      RECT  139300.0 180100.00000000003 140100.0 179300.0 ;
      RECT  137700.0 180100.00000000003 138500.0 179300.0 ;
      RECT  137700.0 186300.0 138500.0 185500.0 ;
      RECT  139300.0 186300.0 140100.0 185500.0 ;
      RECT  139300.0 186300.0 140100.0 185500.0 ;
      RECT  137700.0 186300.0 138500.0 185500.0 ;
      RECT  140900.0 179700.0 141700.0 178900.0 ;
      RECT  140900.0 186300.0 141700.0 185500.0 ;
      RECT  138100.0 183200.0 138900.0 182400.0 ;
      RECT  138100.0 183200.0 138900.0 182400.0 ;
      RECT  139800.0 183100.00000000003 140400.0 182500.0 ;
      RECT  136500.0 178300.0 142900.0 177700.0 ;
      RECT  136500.0 187500.0 142900.0 186900.0 ;
      RECT  140900.0 195100.00000000003 141700.0 196400.0 ;
      RECT  140900.0 187200.0 141700.0 188500.0 ;
      RECT  137700.0 188100.00000000003 138500.0 186900.0 ;
      RECT  137700.0 194300.0 138500.0 196700.0 ;
      RECT  139500.0 188100.00000000003 140100.0 194300.0 ;
      RECT  137700.0 194300.0 138500.0 195100.00000000003 ;
      RECT  139300.0 194300.0 140100.0 195100.00000000003 ;
      RECT  139300.0 194300.0 140100.0 195100.00000000003 ;
      RECT  137700.0 194300.0 138500.0 195100.00000000003 ;
      RECT  137700.0 188100.00000000003 138500.0 188900.0 ;
      RECT  139300.0 188100.00000000003 140100.0 188900.0 ;
      RECT  139300.0 188100.00000000003 140100.0 188900.0 ;
      RECT  137700.0 188100.00000000003 138500.0 188900.0 ;
      RECT  140900.0 194700.0 141700.0 195500.0 ;
      RECT  140900.0 188100.00000000003 141700.0 188900.0 ;
      RECT  138100.0 191200.0 138900.0 192000.0 ;
      RECT  138100.0 191200.0 138900.0 192000.0 ;
      RECT  139800.0 191300.0 140400.0 191900.0 ;
      RECT  136500.0 196100.00000000003 142900.0 196700.0 ;
      RECT  136500.0 186900.0 142900.0 187500.0 ;
      RECT  140900.0 197700.0 141700.0 196400.0 ;
      RECT  140900.0 205600.00000000003 141700.0 204300.0 ;
      RECT  137700.0 204700.0 138500.0 205899.99999999997 ;
      RECT  137700.0 198500.0 138500.0 196100.00000000003 ;
      RECT  139500.0 204700.0 140100.0 198500.0 ;
      RECT  137700.0 198500.0 138500.0 197700.0 ;
      RECT  139300.0 198500.0 140100.0 197700.0 ;
      RECT  139300.0 198500.0 140100.0 197700.0 ;
      RECT  137700.0 198500.0 138500.0 197700.0 ;
      RECT  137700.0 204700.0 138500.0 203899.99999999997 ;
      RECT  139300.0 204700.0 140100.0 203899.99999999997 ;
      RECT  139300.0 204700.0 140100.0 203899.99999999997 ;
      RECT  137700.0 204700.0 138500.0 203899.99999999997 ;
      RECT  140900.0 198100.00000000003 141700.0 197300.0 ;
      RECT  140900.0 204700.0 141700.0 203899.99999999997 ;
      RECT  138100.0 201600.00000000003 138900.0 200800.0 ;
      RECT  138100.0 201600.00000000003 138900.0 200800.0 ;
      RECT  139800.0 201500.0 140400.0 200899.99999999997 ;
      RECT  136500.0 196700.0 142900.0 196100.00000000003 ;
      RECT  136500.0 205899.99999999997 142900.0 205300.0 ;
      RECT  140900.0 213500.0 141700.0 214800.0 ;
      RECT  140900.0 205600.00000000003 141700.0 206899.99999999997 ;
      RECT  137700.0 206500.0 138500.0 205300.0 ;
      RECT  137700.0 212700.0 138500.0 215100.00000000003 ;
      RECT  139500.0 206500.0 140100.0 212700.0 ;
      RECT  137700.0 212700.0 138500.0 213500.0 ;
      RECT  139300.0 212700.0 140100.0 213500.0 ;
      RECT  139300.0 212700.0 140100.0 213500.0 ;
      RECT  137700.0 212700.0 138500.0 213500.0 ;
      RECT  137700.0 206500.0 138500.0 207300.0 ;
      RECT  139300.0 206500.0 140100.0 207300.0 ;
      RECT  139300.0 206500.0 140100.0 207300.0 ;
      RECT  137700.0 206500.0 138500.0 207300.0 ;
      RECT  140900.0 213100.00000000003 141700.0 213899.99999999997 ;
      RECT  140900.0 206500.0 141700.0 207300.0 ;
      RECT  138100.0 209600.00000000003 138900.0 210399.99999999997 ;
      RECT  138100.0 209600.00000000003 138900.0 210399.99999999997 ;
      RECT  139800.0 209700.0 140400.0 210300.0 ;
      RECT  136500.0 214500.0 142900.0 215100.00000000003 ;
      RECT  136500.0 205300.0 142900.0 205899.99999999997 ;
      RECT  140900.0 216100.00000000003 141700.0 214800.0 ;
      RECT  140900.0 224000.0 141700.0 222700.0 ;
      RECT  137700.0 223100.00000000003 138500.0 224300.0 ;
      RECT  137700.0 216899.99999999997 138500.0 214500.0 ;
      RECT  139500.0 223100.00000000003 140100.0 216899.99999999997 ;
      RECT  137700.0 216899.99999999997 138500.0 216100.00000000003 ;
      RECT  139300.0 216899.99999999997 140100.0 216100.00000000003 ;
      RECT  139300.0 216899.99999999997 140100.0 216100.00000000003 ;
      RECT  137700.0 216899.99999999997 138500.0 216100.00000000003 ;
      RECT  137700.0 223100.00000000003 138500.0 222300.0 ;
      RECT  139300.0 223100.00000000003 140100.0 222300.0 ;
      RECT  139300.0 223100.00000000003 140100.0 222300.0 ;
      RECT  137700.0 223100.00000000003 138500.0 222300.0 ;
      RECT  140900.0 216500.0 141700.0 215700.0 ;
      RECT  140900.0 223100.00000000003 141700.0 222300.0 ;
      RECT  138100.0 220000.0 138900.0 219200.0 ;
      RECT  138100.0 220000.0 138900.0 219200.0 ;
      RECT  139800.0 219899.99999999997 140400.0 219300.0 ;
      RECT  136500.0 215100.00000000003 142900.0 214500.0 ;
      RECT  136500.0 224300.0 142900.0 223700.0 ;
      RECT  140900.0 231899.99999999997 141700.0 233200.0 ;
      RECT  140900.0 224000.0 141700.0 225300.0 ;
      RECT  137700.0 224899.99999999997 138500.0 223700.0 ;
      RECT  137700.0 231100.00000000003 138500.0 233500.0 ;
      RECT  139500.0 224899.99999999997 140100.0 231100.00000000003 ;
      RECT  137700.0 231100.00000000003 138500.0 231899.99999999997 ;
      RECT  139300.0 231100.00000000003 140100.0 231899.99999999997 ;
      RECT  139300.0 231100.00000000003 140100.0 231899.99999999997 ;
      RECT  137700.0 231100.00000000003 138500.0 231899.99999999997 ;
      RECT  137700.0 224899.99999999997 138500.0 225700.0 ;
      RECT  139300.0 224899.99999999997 140100.0 225700.0 ;
      RECT  139300.0 224899.99999999997 140100.0 225700.0 ;
      RECT  137700.0 224899.99999999997 138500.0 225700.0 ;
      RECT  140900.0 231500.0 141700.0 232300.0 ;
      RECT  140900.0 224899.99999999997 141700.0 225700.0 ;
      RECT  138100.0 228000.0 138900.0 228800.0 ;
      RECT  138100.0 228000.0 138900.0 228800.0 ;
      RECT  139800.0 228100.00000000003 140400.0 228700.0 ;
      RECT  136500.0 232899.99999999997 142900.0 233500.0 ;
      RECT  136500.0 223700.0 142900.0 224300.0 ;
      RECT  140900.0 234500.0 141700.0 233200.0 ;
      RECT  140900.0 242400.00000000003 141700.0 241100.00000000003 ;
      RECT  137700.0 241500.0 138500.0 242700.0 ;
      RECT  137700.0 235300.0 138500.0 232900.00000000003 ;
      RECT  139500.0 241500.0 140100.0 235300.0 ;
      RECT  137700.0 235300.0 138500.0 234500.0 ;
      RECT  139300.0 235300.0 140100.0 234500.0 ;
      RECT  139300.0 235300.0 140100.0 234500.0 ;
      RECT  137700.0 235300.0 138500.0 234500.0 ;
      RECT  137700.0 241500.0 138500.0 240700.0 ;
      RECT  139300.0 241500.0 140100.0 240700.0 ;
      RECT  139300.0 241500.0 140100.0 240700.0 ;
      RECT  137700.0 241500.0 138500.0 240700.0 ;
      RECT  140900.0 234900.00000000003 141700.0 234100.00000000003 ;
      RECT  140900.0 241500.0 141700.0 240700.0 ;
      RECT  138100.0 238400.00000000003 138900.0 237600.00000000003 ;
      RECT  138100.0 238400.00000000003 138900.0 237600.00000000003 ;
      RECT  139800.0 238300.0 140400.0 237700.0 ;
      RECT  136500.0 233500.0 142900.0 232900.00000000003 ;
      RECT  136500.0 242700.0 142900.0 242100.00000000003 ;
      RECT  140900.0 250300.0 141700.0 251600.00000000003 ;
      RECT  140900.0 242400.00000000003 141700.0 243700.0 ;
      RECT  137700.0 243300.0 138500.0 242100.00000000003 ;
      RECT  137700.0 249500.0 138500.0 251900.00000000003 ;
      RECT  139500.0 243300.0 140100.0 249500.0 ;
      RECT  137700.0 249500.0 138500.0 250300.0 ;
      RECT  139300.0 249500.0 140100.0 250300.0 ;
      RECT  139300.0 249500.0 140100.0 250300.0 ;
      RECT  137700.0 249500.0 138500.0 250300.0 ;
      RECT  137700.0 243300.0 138500.0 244100.00000000003 ;
      RECT  139300.0 243300.0 140100.0 244100.00000000003 ;
      RECT  139300.0 243300.0 140100.0 244100.00000000003 ;
      RECT  137700.0 243300.0 138500.0 244100.00000000003 ;
      RECT  140900.0 249900.00000000003 141700.0 250700.0 ;
      RECT  140900.0 243300.0 141700.0 244100.00000000003 ;
      RECT  138100.0 246400.00000000003 138900.0 247200.0 ;
      RECT  138100.0 246400.00000000003 138900.0 247200.0 ;
      RECT  139800.0 246500.0 140400.0 247100.00000000003 ;
      RECT  136500.0 251300.0 142900.0 251900.00000000003 ;
      RECT  136500.0 242100.00000000003 142900.0 242700.0 ;
      RECT  140900.0 252899.99999999997 141700.0 251600.00000000003 ;
      RECT  140900.0 260800.0 141700.0 259500.0 ;
      RECT  137700.0 259899.99999999997 138500.0 261100.00000000003 ;
      RECT  137700.0 253700.0 138500.0 251300.0 ;
      RECT  139500.0 259899.99999999997 140100.0 253700.0 ;
      RECT  137700.0 253700.0 138500.0 252899.99999999997 ;
      RECT  139300.0 253700.0 140100.0 252899.99999999997 ;
      RECT  139300.0 253700.0 140100.0 252899.99999999997 ;
      RECT  137700.0 253700.0 138500.0 252899.99999999997 ;
      RECT  137700.0 259899.99999999997 138500.0 259100.00000000003 ;
      RECT  139300.0 259899.99999999997 140100.0 259100.00000000003 ;
      RECT  139300.0 259899.99999999997 140100.0 259100.00000000003 ;
      RECT  137700.0 259899.99999999997 138500.0 259100.00000000003 ;
      RECT  140900.0 253300.0 141700.0 252500.0 ;
      RECT  140900.0 259899.99999999997 141700.0 259100.00000000003 ;
      RECT  138100.0 256800.0 138900.0 256000.0 ;
      RECT  138100.0 256800.0 138900.0 256000.0 ;
      RECT  139800.0 256700.0 140400.0 256100.00000000003 ;
      RECT  136500.0 251899.99999999997 142900.0 251300.0 ;
      RECT  136500.0 261100.00000000003 142900.0 260500.0 ;
      RECT  140900.0 268700.0 141700.0 270000.0 ;
      RECT  140900.0 260800.0 141700.0 262100.00000000003 ;
      RECT  137700.0 261700.0 138500.0 260500.0 ;
      RECT  137700.0 267900.0 138500.0 270300.0 ;
      RECT  139500.0 261700.0 140100.0 267900.0 ;
      RECT  137700.0 267900.0 138500.0 268700.0 ;
      RECT  139300.0 267900.0 140100.0 268700.0 ;
      RECT  139300.0 267900.0 140100.0 268700.0 ;
      RECT  137700.0 267900.0 138500.0 268700.0 ;
      RECT  137700.0 261700.0 138500.0 262500.0 ;
      RECT  139300.0 261700.0 140100.0 262500.0 ;
      RECT  139300.0 261700.0 140100.0 262500.0 ;
      RECT  137700.0 261700.0 138500.0 262500.0 ;
      RECT  140900.0 268300.0 141700.0 269100.0 ;
      RECT  140900.0 261700.0 141700.0 262500.0 ;
      RECT  138100.0 264800.0 138900.0 265600.0 ;
      RECT  138100.0 264800.0 138900.0 265600.0 ;
      RECT  139800.0 264900.0 140400.0 265500.0 ;
      RECT  136500.0 269700.0 142900.0 270300.0 ;
      RECT  136500.0 260500.0 142900.0 261100.00000000003 ;
      RECT  140900.0 271300.0 141700.0 270000.0 ;
      RECT  140900.0 279200.0 141700.0 277900.00000000006 ;
      RECT  137700.0 278300.0 138500.0 279500.0 ;
      RECT  137700.0 272100.0 138500.0 269700.0 ;
      RECT  139500.0 278300.0 140100.0 272100.0 ;
      RECT  137700.0 272100.0 138500.0 271300.0 ;
      RECT  139300.0 272100.0 140100.0 271300.0 ;
      RECT  139300.0 272100.0 140100.0 271300.0 ;
      RECT  137700.0 272100.0 138500.0 271300.0 ;
      RECT  137700.0 278300.0 138500.0 277500.0 ;
      RECT  139300.0 278300.0 140100.0 277500.0 ;
      RECT  139300.0 278300.0 140100.0 277500.0 ;
      RECT  137700.0 278300.0 138500.0 277500.0 ;
      RECT  140900.0 271700.0 141700.0 270900.00000000006 ;
      RECT  140900.0 278300.0 141700.0 277500.0 ;
      RECT  138100.0 275200.0 138900.0 274400.00000000006 ;
      RECT  138100.0 275200.0 138900.0 274400.00000000006 ;
      RECT  139800.0 275100.0 140400.0 274500.0 ;
      RECT  136500.0 270300.0 142900.0 269700.0 ;
      RECT  136500.0 279500.0 142900.0 278900.00000000006 ;
      RECT  140900.0 287100.0 141700.0 288400.00000000006 ;
      RECT  140900.0 279200.0 141700.0 280500.0 ;
      RECT  137700.0 280100.0 138500.0 278900.00000000006 ;
      RECT  137700.0 286300.0 138500.0 288700.0 ;
      RECT  139500.0 280100.0 140100.0 286300.0 ;
      RECT  137700.0 286300.0 138500.0 287100.0 ;
      RECT  139300.0 286300.0 140100.0 287100.0 ;
      RECT  139300.0 286300.0 140100.0 287100.0 ;
      RECT  137700.0 286300.0 138500.0 287100.0 ;
      RECT  137700.0 280100.0 138500.0 280900.00000000006 ;
      RECT  139300.0 280100.0 140100.0 280900.00000000006 ;
      RECT  139300.0 280100.0 140100.0 280900.00000000006 ;
      RECT  137700.0 280100.0 138500.0 280900.00000000006 ;
      RECT  140900.0 286700.0 141700.0 287500.0 ;
      RECT  140900.0 280100.0 141700.0 280900.00000000006 ;
      RECT  138100.0 283200.0 138900.0 284000.0 ;
      RECT  138100.0 283200.0 138900.0 284000.0 ;
      RECT  139800.0 283300.0 140400.0 283900.00000000006 ;
      RECT  136500.0 288100.0 142900.0 288700.0 ;
      RECT  136500.0 278900.00000000006 142900.0 279500.0 ;
      RECT  140900.0 289700.0 141700.0 288400.00000000006 ;
      RECT  140900.0 297600.0 141700.0 296300.0 ;
      RECT  137700.0 296700.0 138500.0 297900.00000000006 ;
      RECT  137700.0 290500.0 138500.0 288100.0 ;
      RECT  139500.0 296700.0 140100.0 290500.0 ;
      RECT  137700.0 290500.0 138500.0 289700.0 ;
      RECT  139300.0 290500.0 140100.0 289700.0 ;
      RECT  139300.0 290500.0 140100.0 289700.0 ;
      RECT  137700.0 290500.0 138500.0 289700.0 ;
      RECT  137700.0 296700.0 138500.0 295900.00000000006 ;
      RECT  139300.0 296700.0 140100.0 295900.00000000006 ;
      RECT  139300.0 296700.0 140100.0 295900.00000000006 ;
      RECT  137700.0 296700.0 138500.0 295900.00000000006 ;
      RECT  140900.0 290100.0 141700.0 289300.0 ;
      RECT  140900.0 296700.0 141700.0 295900.00000000006 ;
      RECT  138100.0 293600.0 138900.0 292800.0 ;
      RECT  138100.0 293600.0 138900.0 292800.0 ;
      RECT  139800.0 293500.0 140400.0 292900.00000000006 ;
      RECT  136500.0 288700.0 142900.0 288100.0 ;
      RECT  136500.0 297900.00000000006 142900.0 297300.0 ;
      RECT  140900.0 305500.0 141700.0 306800.0 ;
      RECT  140900.0 297600.0 141700.0 298900.00000000006 ;
      RECT  137700.0 298500.0 138500.0 297300.0 ;
      RECT  137700.0 304700.0 138500.0 307100.0 ;
      RECT  139500.0 298500.0 140100.0 304700.0 ;
      RECT  137700.0 304700.0 138500.0 305500.0 ;
      RECT  139300.0 304700.0 140100.0 305500.0 ;
      RECT  139300.0 304700.0 140100.0 305500.0 ;
      RECT  137700.0 304700.0 138500.0 305500.0 ;
      RECT  137700.0 298500.0 138500.0 299300.0 ;
      RECT  139300.0 298500.0 140100.0 299300.0 ;
      RECT  139300.0 298500.0 140100.0 299300.0 ;
      RECT  137700.0 298500.0 138500.0 299300.0 ;
      RECT  140900.0 305100.0 141700.0 305900.00000000006 ;
      RECT  140900.0 298500.0 141700.0 299300.0 ;
      RECT  138100.0 301600.0 138900.0 302400.00000000006 ;
      RECT  138100.0 301600.0 138900.0 302400.00000000006 ;
      RECT  139800.0 301700.0 140400.0 302300.0 ;
      RECT  136500.0 306500.0 142900.0 307100.0 ;
      RECT  136500.0 297300.0 142900.0 297900.00000000006 ;
      RECT  140900.0 308100.0 141700.0 306800.0 ;
      RECT  140900.0 316000.0 141700.0 314700.0 ;
      RECT  137700.0 315100.0 138500.0 316300.0 ;
      RECT  137700.0 308900.00000000006 138500.0 306500.0 ;
      RECT  139500.0 315100.0 140100.0 308900.00000000006 ;
      RECT  137700.0 308900.00000000006 138500.0 308100.0 ;
      RECT  139300.0 308900.00000000006 140100.0 308100.0 ;
      RECT  139300.0 308900.00000000006 140100.0 308100.0 ;
      RECT  137700.0 308900.00000000006 138500.0 308100.0 ;
      RECT  137700.0 315100.0 138500.0 314300.0 ;
      RECT  139300.0 315100.0 140100.0 314300.0 ;
      RECT  139300.0 315100.0 140100.0 314300.0 ;
      RECT  137700.0 315100.0 138500.0 314300.0 ;
      RECT  140900.0 308500.0 141700.0 307700.0 ;
      RECT  140900.0 315100.0 141700.0 314300.0 ;
      RECT  138100.0 312000.0 138900.0 311200.0 ;
      RECT  138100.0 312000.0 138900.0 311200.0 ;
      RECT  139800.0 311900.00000000006 140400.0 311300.0 ;
      RECT  136500.0 307100.0 142900.0 306500.0 ;
      RECT  136500.0 316300.0 142900.0 315700.0 ;
      RECT  113300.00000000001 172800.0 112500.0 173600.00000000003 ;
      RECT  113300.00000000001 182400.0 112500.0 183200.0 ;
      RECT  113300.00000000001 191200.0 112500.0 192000.0 ;
      RECT  113300.00000000001 200800.0 112500.0 201600.00000000003 ;
      RECT  113300.00000000001 209600.00000000003 112500.0 210399.99999999997 ;
      RECT  113300.00000000001 219200.0 112500.0 220000.0 ;
      RECT  113300.00000000001 228000.0 112500.0 228800.0 ;
      RECT  113300.00000000001 237600.00000000003 112500.0 238399.99999999997 ;
      RECT  116700.0 173200.0 115900.0 174000.0 ;
      RECT  122300.00000000001 171800.0 121500.0 172600.00000000003 ;
      RECT  118100.0 182000.0 117300.00000000001 182800.0 ;
      RECT  122300.00000000001 183400.0 121500.0 184200.0 ;
      RECT  119500.0 191600.00000000003 118700.0 192400.0 ;
      RECT  122300.00000000001 190200.0 121500.0 191000.0 ;
      RECT  120900.0 200399.99999999997 120100.00000000001 201200.0 ;
      RECT  122300.00000000001 201800.0 121500.0 202600.00000000003 ;
      RECT  116700.0 210000.0 115900.0 210800.0 ;
      RECT  123700.0 208600.00000000003 122900.0 209399.99999999997 ;
      RECT  118100.0 218800.0 117300.00000000001 219600.00000000003 ;
      RECT  123700.0 220200.0 122900.0 221000.0 ;
      RECT  119500.0 228399.99999999997 118700.0 229200.0 ;
      RECT  123700.0 227000.0 122900.0 227800.0 ;
      RECT  120900.0 237200.0 120100.00000000001 238000.0 ;
      RECT  123700.0 238600.00000000003 122900.0 239399.99999999997 ;
      RECT  116700.0 246800.0 115900.0 247600.00000000003 ;
      RECT  125100.0 245400.00000000003 124300.00000000001 246200.0 ;
      RECT  118100.0 255600.00000000003 117300.00000000001 256400.00000000003 ;
      RECT  125100.0 257000.0 124300.00000000001 257800.0 ;
      RECT  119500.0 265200.0 118700.0 266000.0 ;
      RECT  125100.0 263800.0 124300.00000000001 264600.0 ;
      RECT  120900.0 274000.0 120100.00000000001 274800.0 ;
      RECT  125100.0 275400.00000000006 124300.00000000001 276200.0 ;
      RECT  116700.0 283600.0 115900.0 284400.00000000006 ;
      RECT  126500.0 282200.0 125700.0 283000.0 ;
      RECT  118100.0 292400.00000000006 117300.00000000001 293200.0 ;
      RECT  126500.0 293800.0 125700.0 294600.0 ;
      RECT  119500.0 302000.0 118700.0 302800.0 ;
      RECT  126500.0 300600.0 125700.0 301400.00000000006 ;
      RECT  120900.0 310800.0 120100.00000000001 311600.0 ;
      RECT  126500.0 312200.0 125700.0 313000.0 ;
      RECT  132100.00000000003 177600.00000000003 131300.0 178400.0 ;
      RECT  132100.00000000003 168400.0 131300.0 169200.0 ;
      RECT  132100.00000000003 177600.00000000003 131300.0 178400.0 ;
      RECT  132100.00000000003 186800.0 131300.0 187600.00000000003 ;
      RECT  132100.00000000003 196000.0 131300.0 196800.0 ;
      RECT  132100.00000000003 186800.0 131300.0 187600.00000000003 ;
      RECT  132100.00000000003 196000.0 131300.0 196800.0 ;
      RECT  132100.00000000003 205200.0 131300.0 206000.0 ;
      RECT  132100.00000000003 214399.99999999997 131300.0 215200.0 ;
      RECT  132100.00000000003 205200.0 131300.0 206000.0 ;
      RECT  132100.00000000003 214399.99999999997 131300.0 215200.0 ;
      RECT  132100.00000000003 223600.00000000003 131300.0 224399.99999999997 ;
      RECT  132100.00000000003 232800.0 131300.0 233600.00000000003 ;
      RECT  132100.00000000003 223600.00000000003 131300.0 224399.99999999997 ;
      RECT  132100.00000000003 232800.0 131300.0 233600.00000000003 ;
      RECT  132100.00000000003 242000.0 131300.0 242800.0 ;
      RECT  132100.00000000003 251200.0 131300.0 252000.0 ;
      RECT  132100.00000000003 242000.0 131300.0 242800.0 ;
      RECT  132100.00000000003 251200.0 131300.0 252000.0 ;
      RECT  132100.00000000003 260400.00000000003 131300.0 261200.0 ;
      RECT  132100.00000000003 269600.0 131300.0 270400.00000000006 ;
      RECT  132100.00000000003 260400.00000000003 131300.0 261200.0 ;
      RECT  132100.00000000003 269600.0 131300.0 270400.00000000006 ;
      RECT  132100.00000000003 278800.0 131300.0 279600.0 ;
      RECT  132100.00000000003 288000.0 131300.0 288800.0 ;
      RECT  132100.00000000003 278800.0 131300.0 279600.0 ;
      RECT  132100.00000000003 288000.0 131300.0 288800.0 ;
      RECT  132100.00000000003 297200.0 131300.0 298000.0 ;
      RECT  132100.00000000003 306400.0 131300.0 307200.0 ;
      RECT  132100.00000000003 297200.0 131300.0 298000.0 ;
      RECT  132100.00000000003 306400.0 131300.0 307200.0 ;
      RECT  132100.00000000003 315600.0 131300.0 316400.00000000006 ;
      RECT  139800.0 172900.0 140400.0 173500.0 ;
      RECT  139800.0 182500.0 140400.0 183100.00000000003 ;
      RECT  139800.0 191300.0 140400.0 191900.0 ;
      RECT  139800.0 200899.99999999997 140400.0 201500.0 ;
      RECT  139800.0 209700.0 140400.0 210300.0 ;
      RECT  139800.0 219300.0 140400.0 219899.99999999997 ;
      RECT  139800.0 228100.00000000003 140400.0 228700.0 ;
      RECT  139800.0 237700.0 140400.0 238300.0 ;
      RECT  139800.0 246500.0 140400.0 247100.00000000003 ;
      RECT  139800.0 256100.00000000003 140400.0 256700.0 ;
      RECT  139800.0 264900.00000000006 140400.0 265500.0 ;
      RECT  139800.0 274500.0 140400.0 275100.0 ;
      RECT  139800.0 283300.0 140400.0 283900.00000000006 ;
      RECT  139800.0 292900.00000000006 140400.0 293500.0 ;
      RECT  139800.0 301700.0 140400.0 302300.0 ;
      RECT  139800.0 311300.0 140400.0 311900.0 ;
      RECT  147400.0 173300.0 151100.0 173900.0 ;
      RECT  158100.0 173300.0 158700.0 173900.0 ;
      RECT  158100.0 172900.0 158700.0 173500.0 ;
      RECT  156100.0 173300.0 158400.0 173900.0 ;
      RECT  158100.0 173200.0 158700.0 173600.00000000003 ;
      RECT  158400.0 172900.0 160700.0 173500.0 ;
      RECT  147400.0 182100.00000000003 151100.0 182700.0 ;
      RECT  158100.0 182100.00000000003 158700.0 182700.0 ;
      RECT  158100.0 182500.0 158700.0 183100.00000000003 ;
      RECT  156100.0 182100.00000000003 158400.0 182700.0 ;
      RECT  158100.0 182400.0 158700.0 182800.0 ;
      RECT  158400.0 182500.0 160700.0 183100.00000000003 ;
      RECT  147400.0 191700.0 151100.0 192300.0 ;
      RECT  158100.0 191700.0 158700.0 192300.0 ;
      RECT  158100.0 191300.0 158700.0 191900.0 ;
      RECT  156100.0 191700.0 158400.0 192300.0 ;
      RECT  158100.0 191600.00000000003 158700.0 192000.0 ;
      RECT  158400.0 191300.0 160700.0 191900.0 ;
      RECT  147400.0 200500.0 151100.0 201100.00000000003 ;
      RECT  158100.0 200500.0 158700.0 201100.00000000003 ;
      RECT  158100.0 200899.99999999997 158700.0 201500.0 ;
      RECT  156100.0 200500.0 158400.0 201100.00000000003 ;
      RECT  158100.0 200800.0 158700.0 201200.0 ;
      RECT  158400.0 200899.99999999997 160700.0 201500.0 ;
      RECT  147400.0 210100.00000000003 151100.0 210700.0 ;
      RECT  158100.0 210100.00000000003 158700.0 210700.0 ;
      RECT  158100.0 209700.0 158700.0 210300.0 ;
      RECT  156100.0 210100.00000000003 158400.0 210700.0 ;
      RECT  158100.0 210000.0 158700.0 210399.99999999997 ;
      RECT  158400.0 209700.0 160700.0 210300.0 ;
      RECT  147400.0 218899.99999999997 151100.0 219500.0 ;
      RECT  158100.0 218899.99999999997 158700.0 219500.0 ;
      RECT  158100.0 219300.0 158700.0 219899.99999999997 ;
      RECT  156100.0 218899.99999999997 158400.0 219500.0 ;
      RECT  158100.0 219200.0 158700.0 219600.00000000003 ;
      RECT  158400.0 219300.0 160700.0 219899.99999999997 ;
      RECT  147400.0 228500.0 151100.0 229100.00000000003 ;
      RECT  158100.0 228500.0 158700.0 229100.00000000003 ;
      RECT  158100.0 228100.00000000003 158700.0 228700.0 ;
      RECT  156100.0 228500.0 158400.0 229100.00000000003 ;
      RECT  158100.0 228399.99999999997 158700.0 228800.0 ;
      RECT  158400.0 228100.00000000003 160700.0 228700.0 ;
      RECT  147400.0 237300.0 151100.0 237899.99999999997 ;
      RECT  158100.0 237300.0 158700.0 237899.99999999997 ;
      RECT  158100.0 237700.0 158700.0 238300.0 ;
      RECT  156100.0 237300.0 158400.0 237899.99999999997 ;
      RECT  158100.0 237600.00000000003 158700.0 238000.0 ;
      RECT  158400.0 237700.0 160700.0 238300.0 ;
      RECT  147400.0 246900.00000000003 151100.0 247500.0 ;
      RECT  158100.0 246900.00000000003 158700.0 247500.0 ;
      RECT  158100.0 246500.0 158700.0 247100.00000000003 ;
      RECT  156100.0 246900.00000000003 158400.0 247500.0 ;
      RECT  158100.0 246800.0 158700.0 247200.0 ;
      RECT  158400.0 246500.0 160700.0 247100.00000000003 ;
      RECT  147400.0 255700.0 151100.0 256300.0 ;
      RECT  158100.0 255700.0 158700.0 256300.0 ;
      RECT  158100.0 256100.00000000003 158700.0 256700.0 ;
      RECT  156100.0 255700.0 158400.0 256300.0 ;
      RECT  158100.0 256000.0 158700.0 256400.00000000003 ;
      RECT  158400.0 256100.00000000003 160700.0 256700.0 ;
      RECT  147400.0 265300.0 151100.0 265900.0 ;
      RECT  158100.0 265300.0 158700.0 265900.0 ;
      RECT  158100.0 264900.00000000006 158700.0 265500.0 ;
      RECT  156100.0 265300.0 158400.0 265900.0 ;
      RECT  158100.0 265200.0 158700.0 265600.0 ;
      RECT  158400.0 264900.00000000006 160700.0 265500.0 ;
      RECT  147400.0 274100.0 151100.0 274700.0 ;
      RECT  158100.0 274100.0 158700.0 274700.0 ;
      RECT  158100.0 274500.0 158700.0 275100.0 ;
      RECT  156100.0 274100.0 158400.0 274700.0 ;
      RECT  158100.0 274400.00000000006 158700.0 274800.0 ;
      RECT  158400.0 274500.0 160700.0 275100.0 ;
      RECT  147400.0 283700.0 151100.0 284300.0 ;
      RECT  158100.0 283700.0 158700.0 284300.0 ;
      RECT  158100.0 283300.0 158700.0 283900.0 ;
      RECT  156100.0 283700.0 158400.0 284300.0 ;
      RECT  158100.0 283600.0 158700.0 284000.0 ;
      RECT  158400.0 283300.0 160700.0 283900.0 ;
      RECT  147400.0 292500.0 151100.0 293100.0 ;
      RECT  158100.0 292500.0 158700.0 293100.0 ;
      RECT  158100.0 292900.00000000006 158700.0 293500.0 ;
      RECT  156100.0 292500.0 158400.0 293100.0 ;
      RECT  158100.0 292800.0 158700.0 293200.0 ;
      RECT  158400.0 292900.00000000006 160700.0 293500.0 ;
      RECT  147400.0 302100.0 151100.0 302700.0 ;
      RECT  158100.0 302100.0 158700.0 302700.0 ;
      RECT  158100.0 301700.0 158700.0 302300.0 ;
      RECT  156100.0 302100.0 158400.0 302700.0 ;
      RECT  158100.0 302000.0 158700.0 302400.00000000006 ;
      RECT  158400.0 301700.0 160700.0 302300.0 ;
      RECT  147400.0 310900.0 151100.0 311500.0 ;
      RECT  158100.0 310900.0 158700.0 311500.0 ;
      RECT  158100.0 311300.0 158700.0 311900.0 ;
      RECT  156100.0 310900.0 158400.0 311500.0 ;
      RECT  158100.0 311200.0 158700.0 311600.0 ;
      RECT  158400.0 311300.0 160700.0 311900.0 ;
      RECT  150700.0 170100.00000000003 151500.0 168500.0 ;
      RECT  150700.0 175900.0 151500.0 178300.0 ;
      RECT  153900.0 175900.0 154700.0 178300.0 ;
      RECT  155500.0 176700.0 156300.0 178000.0 ;
      RECT  155500.0 168800.0 156300.0 170100.00000000003 ;
      RECT  150700.0 175900.0 151500.0 176700.0 ;
      RECT  152300.0 175900.0 153100.0 176700.0 ;
      RECT  152300.0 175900.0 153100.0 176700.0 ;
      RECT  150700.0 175900.0 151500.0 176700.0 ;
      RECT  152300.0 175900.0 153100.0 176700.0 ;
      RECT  153900.0 175900.0 154700.0 176700.0 ;
      RECT  153900.0 175900.0 154700.0 176700.0 ;
      RECT  152300.0 175900.0 153100.0 176700.0 ;
      RECT  150700.0 170100.00000000003 151500.0 170900.0 ;
      RECT  152300.0 170100.00000000003 153100.0 170900.0 ;
      RECT  152300.0 170100.00000000003 153100.0 170900.0 ;
      RECT  150700.0 170100.00000000003 151500.0 170900.0 ;
      RECT  152300.0 170100.00000000003 153100.0 170900.0 ;
      RECT  153900.0 170100.00000000003 154700.0 170900.0 ;
      RECT  153900.0 170100.00000000003 154700.0 170900.0 ;
      RECT  152300.0 170100.00000000003 153100.0 170900.0 ;
      RECT  155500.0 176300.0 156300.0 177100.00000000003 ;
      RECT  155500.0 169700.0 156300.0 170500.0 ;
      RECT  153900.0 171800.0 153100.0 172600.00000000003 ;
      RECT  151900.0 173200.0 151100.0 174000.0 ;
      RECT  152300.0 175900.0 153100.0 176700.0 ;
      RECT  153900.0 170100.00000000003 154700.0 170900.0 ;
      RECT  156100.0 173200.0 155300.0 174000.0 ;
      RECT  151100.0 173200.0 151900.0 174000.0 ;
      RECT  153100.0 171800.0 153900.0 172600.00000000003 ;
      RECT  155300.0 173200.0 156100.0 174000.0 ;
      RECT  149500.0 177700.0 159100.0 178300.0 ;
      RECT  149500.0 168500.0 159100.0 169100.00000000003 ;
      RECT  163500.0 176700.0 164300.0 178000.0 ;
      RECT  163500.0 168800.0 164300.0 170100.00000000003 ;
      RECT  160300.0 169700.0 161100.0 168500.0 ;
      RECT  160300.0 175900.0 161100.0 178300.0 ;
      RECT  162100.0 169700.0 162700.0 175900.0 ;
      RECT  160300.0 175900.0 161100.0 176700.0 ;
      RECT  161900.0 175900.0 162700.0 176700.0 ;
      RECT  161900.0 175900.0 162700.0 176700.0 ;
      RECT  160300.0 175900.0 161100.0 176700.0 ;
      RECT  160300.0 169700.0 161100.0 170500.0 ;
      RECT  161900.0 169700.0 162700.0 170500.0 ;
      RECT  161900.0 169700.0 162700.0 170500.0 ;
      RECT  160300.0 169700.0 161100.0 170500.0 ;
      RECT  163500.0 176300.0 164300.0 177100.00000000003 ;
      RECT  163500.0 169700.0 164300.0 170500.0 ;
      RECT  160700.0 172800.0 161500.0 173600.00000000003 ;
      RECT  160700.0 172800.0 161500.0 173600.00000000003 ;
      RECT  162400.0 172900.0 163000.0 173500.0 ;
      RECT  159100.0 177700.0 165500.0 178300.0 ;
      RECT  159100.0 168500.0 165500.0 169100.00000000003 ;
      RECT  150700.0 185900.0 151500.0 187500.0 ;
      RECT  150700.0 180100.00000000003 151500.0 177700.0 ;
      RECT  153900.0 180100.00000000003 154700.0 177700.0 ;
      RECT  155500.0 179300.0 156300.0 178000.0 ;
      RECT  155500.0 187200.0 156300.0 185900.0 ;
      RECT  150700.0 180100.00000000003 151500.0 179300.0 ;
      RECT  152300.0 180100.00000000003 153100.0 179300.0 ;
      RECT  152300.0 180100.00000000003 153100.0 179300.0 ;
      RECT  150700.0 180100.00000000003 151500.0 179300.0 ;
      RECT  152300.0 180100.00000000003 153100.0 179300.0 ;
      RECT  153900.0 180100.00000000003 154700.0 179300.0 ;
      RECT  153900.0 180100.00000000003 154700.0 179300.0 ;
      RECT  152300.0 180100.00000000003 153100.0 179300.0 ;
      RECT  150700.0 185900.0 151500.0 185100.00000000003 ;
      RECT  152300.0 185900.0 153100.0 185100.00000000003 ;
      RECT  152300.0 185900.0 153100.0 185100.00000000003 ;
      RECT  150700.0 185900.0 151500.0 185100.00000000003 ;
      RECT  152300.0 185900.0 153100.0 185100.00000000003 ;
      RECT  153900.0 185900.0 154700.0 185100.00000000003 ;
      RECT  153900.0 185900.0 154700.0 185100.00000000003 ;
      RECT  152300.0 185900.0 153100.0 185100.00000000003 ;
      RECT  155500.0 179700.0 156300.0 178900.0 ;
      RECT  155500.0 186300.0 156300.0 185500.0 ;
      RECT  153900.0 184200.0 153100.0 183400.0 ;
      RECT  151900.0 182800.0 151100.0 182000.0 ;
      RECT  152300.0 180100.00000000003 153100.0 179300.0 ;
      RECT  153900.0 185900.0 154700.0 185100.00000000003 ;
      RECT  156100.0 182800.0 155300.0 182000.0 ;
      RECT  151100.0 182800.0 151900.0 182000.0 ;
      RECT  153100.0 184200.0 153900.0 183400.0 ;
      RECT  155300.0 182800.0 156100.0 182000.0 ;
      RECT  149500.0 178300.0 159100.0 177700.0 ;
      RECT  149500.0 187500.0 159100.0 186900.0 ;
      RECT  163500.0 179300.0 164300.0 178000.0 ;
      RECT  163500.0 187200.0 164300.0 185900.0 ;
      RECT  160300.0 186300.0 161100.0 187500.0 ;
      RECT  160300.0 180100.00000000003 161100.0 177700.0 ;
      RECT  162100.0 186300.0 162700.0 180100.00000000003 ;
      RECT  160300.0 180100.00000000003 161100.0 179300.0 ;
      RECT  161900.0 180100.00000000003 162700.0 179300.0 ;
      RECT  161900.0 180100.00000000003 162700.0 179300.0 ;
      RECT  160300.0 180100.00000000003 161100.0 179300.0 ;
      RECT  160300.0 186300.0 161100.0 185500.0 ;
      RECT  161900.0 186300.0 162700.0 185500.0 ;
      RECT  161900.0 186300.0 162700.0 185500.0 ;
      RECT  160300.0 186300.0 161100.0 185500.0 ;
      RECT  163500.0 179700.0 164300.0 178900.0 ;
      RECT  163500.0 186300.0 164300.0 185500.0 ;
      RECT  160700.0 183200.0 161500.0 182400.0 ;
      RECT  160700.0 183200.0 161500.0 182400.0 ;
      RECT  162400.0 183100.00000000003 163000.0 182500.0 ;
      RECT  159100.0 178300.0 165500.0 177700.0 ;
      RECT  159100.0 187500.0 165500.0 186900.0 ;
      RECT  150700.0 188500.0 151500.0 186900.0 ;
      RECT  150700.0 194300.0 151500.0 196700.0 ;
      RECT  153900.0 194300.0 154700.0 196700.0 ;
      RECT  155500.0 195100.00000000003 156300.0 196400.0 ;
      RECT  155500.0 187200.0 156300.0 188500.0 ;
      RECT  150700.0 194300.0 151500.0 195100.00000000003 ;
      RECT  152300.0 194300.0 153100.0 195100.00000000003 ;
      RECT  152300.0 194300.0 153100.0 195100.00000000003 ;
      RECT  150700.0 194300.0 151500.0 195100.00000000003 ;
      RECT  152300.0 194300.0 153100.0 195100.00000000003 ;
      RECT  153900.0 194300.0 154700.0 195100.00000000003 ;
      RECT  153900.0 194300.0 154700.0 195100.00000000003 ;
      RECT  152300.0 194300.0 153100.0 195100.00000000003 ;
      RECT  150700.0 188500.0 151500.0 189300.0 ;
      RECT  152300.0 188500.0 153100.0 189300.0 ;
      RECT  152300.0 188500.0 153100.0 189300.0 ;
      RECT  150700.0 188500.0 151500.0 189300.0 ;
      RECT  152300.0 188500.0 153100.0 189300.0 ;
      RECT  153900.0 188500.0 154700.0 189300.0 ;
      RECT  153900.0 188500.0 154700.0 189300.0 ;
      RECT  152300.0 188500.0 153100.0 189300.0 ;
      RECT  155500.0 194700.0 156300.0 195500.0 ;
      RECT  155500.0 188100.00000000003 156300.0 188900.0 ;
      RECT  153900.0 190200.0 153100.0 191000.0 ;
      RECT  151900.0 191600.00000000003 151100.0 192400.0 ;
      RECT  152300.0 194300.0 153100.0 195100.00000000003 ;
      RECT  153900.0 188500.0 154700.0 189300.0 ;
      RECT  156100.0 191600.00000000003 155300.0 192400.0 ;
      RECT  151100.0 191600.00000000003 151900.0 192400.0 ;
      RECT  153100.0 190200.0 153900.0 191000.0 ;
      RECT  155300.0 191600.00000000003 156100.0 192400.0 ;
      RECT  149500.0 196100.00000000003 159100.0 196700.0 ;
      RECT  149500.0 186900.0 159100.0 187500.0 ;
      RECT  163500.0 195100.00000000003 164300.0 196400.0 ;
      RECT  163500.0 187200.0 164300.0 188500.0 ;
      RECT  160300.0 188100.00000000003 161100.0 186900.0 ;
      RECT  160300.0 194300.0 161100.0 196700.0 ;
      RECT  162100.0 188100.00000000003 162700.0 194300.0 ;
      RECT  160300.0 194300.0 161100.0 195100.00000000003 ;
      RECT  161900.0 194300.0 162700.0 195100.00000000003 ;
      RECT  161900.0 194300.0 162700.0 195100.00000000003 ;
      RECT  160300.0 194300.0 161100.0 195100.00000000003 ;
      RECT  160300.0 188100.00000000003 161100.0 188900.0 ;
      RECT  161900.0 188100.00000000003 162700.0 188900.0 ;
      RECT  161900.0 188100.00000000003 162700.0 188900.0 ;
      RECT  160300.0 188100.00000000003 161100.0 188900.0 ;
      RECT  163500.0 194700.0 164300.0 195500.0 ;
      RECT  163500.0 188100.00000000003 164300.0 188900.0 ;
      RECT  160700.0 191200.0 161500.0 192000.0 ;
      RECT  160700.0 191200.0 161500.0 192000.0 ;
      RECT  162400.0 191300.0 163000.0 191900.0 ;
      RECT  159100.0 196100.00000000003 165500.0 196700.0 ;
      RECT  159100.0 186900.0 165500.0 187500.0 ;
      RECT  150700.0 204300.0 151500.0 205899.99999999997 ;
      RECT  150700.0 198500.0 151500.0 196100.00000000003 ;
      RECT  153900.0 198500.0 154700.0 196100.00000000003 ;
      RECT  155500.0 197700.0 156300.0 196400.0 ;
      RECT  155500.0 205600.00000000003 156300.0 204300.0 ;
      RECT  150700.0 198500.0 151500.0 197700.0 ;
      RECT  152300.0 198500.0 153100.0 197700.0 ;
      RECT  152300.0 198500.0 153100.0 197700.0 ;
      RECT  150700.0 198500.0 151500.0 197700.0 ;
      RECT  152300.0 198500.0 153100.0 197700.0 ;
      RECT  153900.0 198500.0 154700.0 197700.0 ;
      RECT  153900.0 198500.0 154700.0 197700.0 ;
      RECT  152300.0 198500.0 153100.0 197700.0 ;
      RECT  150700.0 204300.0 151500.0 203500.0 ;
      RECT  152300.0 204300.0 153100.0 203500.0 ;
      RECT  152300.0 204300.0 153100.0 203500.0 ;
      RECT  150700.0 204300.0 151500.0 203500.0 ;
      RECT  152300.0 204300.0 153100.0 203500.0 ;
      RECT  153900.0 204300.0 154700.0 203500.0 ;
      RECT  153900.0 204300.0 154700.0 203500.0 ;
      RECT  152300.0 204300.0 153100.0 203500.0 ;
      RECT  155500.0 198100.00000000003 156300.0 197300.0 ;
      RECT  155500.0 204700.0 156300.0 203899.99999999997 ;
      RECT  153900.0 202600.00000000003 153100.0 201800.0 ;
      RECT  151900.0 201200.0 151100.0 200399.99999999997 ;
      RECT  152300.0 198500.0 153100.0 197700.0 ;
      RECT  153900.0 204300.0 154700.0 203500.0 ;
      RECT  156100.0 201200.0 155300.0 200399.99999999997 ;
      RECT  151100.0 201200.0 151900.0 200399.99999999997 ;
      RECT  153100.0 202600.00000000003 153900.0 201800.0 ;
      RECT  155300.0 201200.0 156100.0 200399.99999999997 ;
      RECT  149500.0 196700.0 159100.0 196100.00000000003 ;
      RECT  149500.0 205899.99999999997 159100.0 205300.0 ;
      RECT  163500.0 197700.0 164300.0 196400.0 ;
      RECT  163500.0 205600.00000000003 164300.0 204300.0 ;
      RECT  160300.0 204700.0 161100.0 205899.99999999997 ;
      RECT  160300.0 198500.0 161100.0 196100.00000000003 ;
      RECT  162100.0 204700.0 162700.0 198500.0 ;
      RECT  160300.0 198500.0 161100.0 197700.0 ;
      RECT  161900.0 198500.0 162700.0 197700.0 ;
      RECT  161900.0 198500.0 162700.0 197700.0 ;
      RECT  160300.0 198500.0 161100.0 197700.0 ;
      RECT  160300.0 204700.0 161100.0 203899.99999999997 ;
      RECT  161900.0 204700.0 162700.0 203899.99999999997 ;
      RECT  161900.0 204700.0 162700.0 203899.99999999997 ;
      RECT  160300.0 204700.0 161100.0 203899.99999999997 ;
      RECT  163500.0 198100.00000000003 164300.0 197300.0 ;
      RECT  163500.0 204700.0 164300.0 203899.99999999997 ;
      RECT  160700.0 201600.00000000003 161500.0 200800.0 ;
      RECT  160700.0 201600.00000000003 161500.0 200800.0 ;
      RECT  162400.0 201500.0 163000.0 200899.99999999997 ;
      RECT  159100.0 196700.0 165500.0 196100.00000000003 ;
      RECT  159100.0 205899.99999999997 165500.0 205300.0 ;
      RECT  150700.0 206899.99999999997 151500.0 205300.0 ;
      RECT  150700.0 212700.0 151500.0 215100.00000000003 ;
      RECT  153900.0 212700.0 154700.0 215100.00000000003 ;
      RECT  155500.0 213500.0 156300.0 214800.0 ;
      RECT  155500.0 205600.00000000003 156300.0 206899.99999999997 ;
      RECT  150700.0 212700.0 151500.0 213500.0 ;
      RECT  152300.0 212700.0 153100.0 213500.0 ;
      RECT  152300.0 212700.0 153100.0 213500.0 ;
      RECT  150700.0 212700.0 151500.0 213500.0 ;
      RECT  152300.0 212700.0 153100.0 213500.0 ;
      RECT  153900.0 212700.0 154700.0 213500.0 ;
      RECT  153900.0 212700.0 154700.0 213500.0 ;
      RECT  152300.0 212700.0 153100.0 213500.0 ;
      RECT  150700.0 206899.99999999997 151500.0 207700.0 ;
      RECT  152300.0 206899.99999999997 153100.0 207700.0 ;
      RECT  152300.0 206899.99999999997 153100.0 207700.0 ;
      RECT  150700.0 206899.99999999997 151500.0 207700.0 ;
      RECT  152300.0 206899.99999999997 153100.0 207700.0 ;
      RECT  153900.0 206899.99999999997 154700.0 207700.0 ;
      RECT  153900.0 206899.99999999997 154700.0 207700.0 ;
      RECT  152300.0 206899.99999999997 153100.0 207700.0 ;
      RECT  155500.0 213100.00000000003 156300.0 213899.99999999997 ;
      RECT  155500.0 206500.0 156300.0 207300.0 ;
      RECT  153900.0 208600.00000000003 153100.0 209399.99999999997 ;
      RECT  151900.0 210000.0 151100.0 210800.0 ;
      RECT  152300.0 212700.0 153100.0 213500.0 ;
      RECT  153900.0 206899.99999999997 154700.0 207700.0 ;
      RECT  156100.0 210000.0 155300.0 210800.0 ;
      RECT  151100.0 210000.0 151900.0 210800.0 ;
      RECT  153100.0 208600.00000000003 153900.0 209399.99999999997 ;
      RECT  155300.0 210000.0 156100.0 210800.0 ;
      RECT  149500.0 214500.0 159100.0 215100.00000000003 ;
      RECT  149500.0 205300.0 159100.0 205899.99999999997 ;
      RECT  163500.0 213500.0 164300.0 214800.0 ;
      RECT  163500.0 205600.00000000003 164300.0 206899.99999999997 ;
      RECT  160300.0 206500.0 161100.0 205300.0 ;
      RECT  160300.0 212700.0 161100.0 215100.00000000003 ;
      RECT  162100.0 206500.0 162700.0 212700.0 ;
      RECT  160300.0 212700.0 161100.0 213500.0 ;
      RECT  161900.0 212700.0 162700.0 213500.0 ;
      RECT  161900.0 212700.0 162700.0 213500.0 ;
      RECT  160300.0 212700.0 161100.0 213500.0 ;
      RECT  160300.0 206500.0 161100.0 207300.0 ;
      RECT  161900.0 206500.0 162700.0 207300.0 ;
      RECT  161900.0 206500.0 162700.0 207300.0 ;
      RECT  160300.0 206500.0 161100.0 207300.0 ;
      RECT  163500.0 213100.00000000003 164300.0 213899.99999999997 ;
      RECT  163500.0 206500.0 164300.0 207300.0 ;
      RECT  160700.0 209600.00000000003 161500.0 210399.99999999997 ;
      RECT  160700.0 209600.00000000003 161500.0 210399.99999999997 ;
      RECT  162400.0 209700.0 163000.0 210300.0 ;
      RECT  159100.0 214500.0 165500.0 215100.00000000003 ;
      RECT  159100.0 205300.0 165500.0 205899.99999999997 ;
      RECT  150700.0 222700.0 151500.0 224300.0 ;
      RECT  150700.0 216899.99999999997 151500.0 214500.0 ;
      RECT  153900.0 216899.99999999997 154700.0 214500.0 ;
      RECT  155500.0 216100.00000000003 156300.0 214800.0 ;
      RECT  155500.0 224000.0 156300.0 222700.0 ;
      RECT  150700.0 216899.99999999997 151500.0 216100.00000000003 ;
      RECT  152300.0 216899.99999999997 153100.0 216100.00000000003 ;
      RECT  152300.0 216899.99999999997 153100.0 216100.00000000003 ;
      RECT  150700.0 216899.99999999997 151500.0 216100.00000000003 ;
      RECT  152300.0 216899.99999999997 153100.0 216100.00000000003 ;
      RECT  153900.0 216899.99999999997 154700.0 216100.00000000003 ;
      RECT  153900.0 216899.99999999997 154700.0 216100.00000000003 ;
      RECT  152300.0 216899.99999999997 153100.0 216100.00000000003 ;
      RECT  150700.0 222700.0 151500.0 221899.99999999997 ;
      RECT  152300.0 222700.0 153100.0 221899.99999999997 ;
      RECT  152300.0 222700.0 153100.0 221899.99999999997 ;
      RECT  150700.0 222700.0 151500.0 221899.99999999997 ;
      RECT  152300.0 222700.0 153100.0 221899.99999999997 ;
      RECT  153900.0 222700.0 154700.0 221899.99999999997 ;
      RECT  153900.0 222700.0 154700.0 221899.99999999997 ;
      RECT  152300.0 222700.0 153100.0 221899.99999999997 ;
      RECT  155500.0 216500.0 156300.0 215700.0 ;
      RECT  155500.0 223100.00000000003 156300.0 222300.0 ;
      RECT  153900.0 221000.0 153100.0 220200.0 ;
      RECT  151900.0 219600.00000000003 151100.0 218800.0 ;
      RECT  152300.0 216899.99999999997 153100.0 216100.00000000003 ;
      RECT  153900.0 222700.0 154700.0 221899.99999999997 ;
      RECT  156100.0 219600.00000000003 155300.0 218800.0 ;
      RECT  151100.0 219600.00000000003 151900.0 218800.0 ;
      RECT  153100.0 221000.0 153900.0 220200.0 ;
      RECT  155300.0 219600.00000000003 156100.0 218800.0 ;
      RECT  149500.0 215100.00000000003 159100.0 214500.0 ;
      RECT  149500.0 224300.0 159100.0 223700.0 ;
      RECT  163500.0 216100.00000000003 164300.0 214800.0 ;
      RECT  163500.0 224000.0 164300.0 222700.0 ;
      RECT  160300.0 223100.00000000003 161100.0 224300.0 ;
      RECT  160300.0 216899.99999999997 161100.0 214500.0 ;
      RECT  162100.0 223100.00000000003 162700.0 216899.99999999997 ;
      RECT  160300.0 216899.99999999997 161100.0 216100.00000000003 ;
      RECT  161900.0 216899.99999999997 162700.0 216100.00000000003 ;
      RECT  161900.0 216899.99999999997 162700.0 216100.00000000003 ;
      RECT  160300.0 216899.99999999997 161100.0 216100.00000000003 ;
      RECT  160300.0 223100.00000000003 161100.0 222300.0 ;
      RECT  161900.0 223100.00000000003 162700.0 222300.0 ;
      RECT  161900.0 223100.00000000003 162700.0 222300.0 ;
      RECT  160300.0 223100.00000000003 161100.0 222300.0 ;
      RECT  163500.0 216500.0 164300.0 215700.0 ;
      RECT  163500.0 223100.00000000003 164300.0 222300.0 ;
      RECT  160700.0 220000.0 161500.0 219200.0 ;
      RECT  160700.0 220000.0 161500.0 219200.0 ;
      RECT  162400.0 219899.99999999997 163000.0 219300.0 ;
      RECT  159100.0 215100.00000000003 165500.0 214500.0 ;
      RECT  159100.0 224300.0 165500.0 223700.0 ;
      RECT  150700.0 225300.0 151500.0 223700.0 ;
      RECT  150700.0 231100.00000000003 151500.0 233500.0 ;
      RECT  153900.0 231100.00000000003 154700.0 233500.0 ;
      RECT  155500.0 231899.99999999997 156300.0 233200.0 ;
      RECT  155500.0 224000.0 156300.0 225300.0 ;
      RECT  150700.0 231100.00000000003 151500.0 231899.99999999997 ;
      RECT  152300.0 231100.00000000003 153100.0 231899.99999999997 ;
      RECT  152300.0 231100.00000000003 153100.0 231899.99999999997 ;
      RECT  150700.0 231100.00000000003 151500.0 231899.99999999997 ;
      RECT  152300.0 231100.00000000003 153100.0 231899.99999999997 ;
      RECT  153900.0 231100.00000000003 154700.0 231899.99999999997 ;
      RECT  153900.0 231100.00000000003 154700.0 231899.99999999997 ;
      RECT  152300.0 231100.00000000003 153100.0 231899.99999999997 ;
      RECT  150700.0 225300.0 151500.0 226100.00000000003 ;
      RECT  152300.0 225300.0 153100.0 226100.00000000003 ;
      RECT  152300.0 225300.0 153100.0 226100.00000000003 ;
      RECT  150700.0 225300.0 151500.0 226100.00000000003 ;
      RECT  152300.0 225300.0 153100.0 226100.00000000003 ;
      RECT  153900.0 225300.0 154700.0 226100.00000000003 ;
      RECT  153900.0 225300.0 154700.0 226100.00000000003 ;
      RECT  152300.0 225300.0 153100.0 226100.00000000003 ;
      RECT  155500.0 231500.0 156300.0 232300.0 ;
      RECT  155500.0 224899.99999999997 156300.0 225700.0 ;
      RECT  153900.0 227000.0 153100.0 227800.0 ;
      RECT  151900.0 228399.99999999997 151100.0 229200.0 ;
      RECT  152300.0 231100.00000000003 153100.0 231899.99999999997 ;
      RECT  153900.0 225300.0 154700.0 226100.00000000003 ;
      RECT  156100.0 228399.99999999997 155300.0 229200.0 ;
      RECT  151100.0 228399.99999999997 151900.0 229200.0 ;
      RECT  153100.0 227000.0 153900.0 227800.0 ;
      RECT  155300.0 228399.99999999997 156100.0 229200.0 ;
      RECT  149500.0 232899.99999999997 159100.0 233500.0 ;
      RECT  149500.0 223700.0 159100.0 224300.0 ;
      RECT  163500.0 231899.99999999997 164300.0 233200.0 ;
      RECT  163500.0 224000.0 164300.0 225300.0 ;
      RECT  160300.0 224899.99999999997 161100.0 223700.0 ;
      RECT  160300.0 231100.00000000003 161100.0 233500.0 ;
      RECT  162100.0 224899.99999999997 162700.0 231100.00000000003 ;
      RECT  160300.0 231100.00000000003 161100.0 231899.99999999997 ;
      RECT  161900.0 231100.00000000003 162700.0 231899.99999999997 ;
      RECT  161900.0 231100.00000000003 162700.0 231899.99999999997 ;
      RECT  160300.0 231100.00000000003 161100.0 231899.99999999997 ;
      RECT  160300.0 224899.99999999997 161100.0 225700.0 ;
      RECT  161900.0 224899.99999999997 162700.0 225700.0 ;
      RECT  161900.0 224899.99999999997 162700.0 225700.0 ;
      RECT  160300.0 224899.99999999997 161100.0 225700.0 ;
      RECT  163500.0 231500.0 164300.0 232300.0 ;
      RECT  163500.0 224899.99999999997 164300.0 225700.0 ;
      RECT  160700.0 228000.0 161500.0 228800.0 ;
      RECT  160700.0 228000.0 161500.0 228800.0 ;
      RECT  162400.0 228100.00000000003 163000.0 228700.0 ;
      RECT  159100.0 232899.99999999997 165500.0 233500.0 ;
      RECT  159100.0 223700.0 165500.0 224300.0 ;
      RECT  150700.0 241100.00000000003 151500.0 242700.0 ;
      RECT  150700.0 235300.0 151500.0 232900.00000000003 ;
      RECT  153900.0 235300.0 154700.0 232900.00000000003 ;
      RECT  155500.0 234500.0 156300.0 233200.0 ;
      RECT  155500.0 242400.00000000003 156300.0 241100.00000000003 ;
      RECT  150700.0 235300.0 151500.0 234500.0 ;
      RECT  152300.0 235300.0 153100.0 234500.0 ;
      RECT  152300.0 235300.0 153100.0 234500.0 ;
      RECT  150700.0 235300.0 151500.0 234500.0 ;
      RECT  152300.0 235300.0 153100.0 234500.0 ;
      RECT  153900.0 235300.0 154700.0 234500.0 ;
      RECT  153900.0 235300.0 154700.0 234500.0 ;
      RECT  152300.0 235300.0 153100.0 234500.0 ;
      RECT  150700.0 241100.00000000003 151500.0 240300.0 ;
      RECT  152300.0 241100.00000000003 153100.0 240300.0 ;
      RECT  152300.0 241100.00000000003 153100.0 240300.0 ;
      RECT  150700.0 241100.00000000003 151500.0 240300.0 ;
      RECT  152300.0 241100.00000000003 153100.0 240300.0 ;
      RECT  153900.0 241100.00000000003 154700.0 240300.0 ;
      RECT  153900.0 241100.00000000003 154700.0 240300.0 ;
      RECT  152300.0 241100.00000000003 153100.0 240300.0 ;
      RECT  155500.0 234900.00000000003 156300.0 234100.00000000003 ;
      RECT  155500.0 241500.0 156300.0 240700.0 ;
      RECT  153900.0 239400.00000000003 153100.0 238600.00000000003 ;
      RECT  151900.0 238000.0 151100.0 237200.0 ;
      RECT  152300.0 235300.0 153100.0 234500.0 ;
      RECT  153900.0 241100.00000000003 154700.0 240300.0 ;
      RECT  156100.0 238000.0 155300.0 237200.0 ;
      RECT  151100.0 238000.0 151900.0 237200.0 ;
      RECT  153100.0 239400.00000000003 153900.0 238600.00000000003 ;
      RECT  155300.0 238000.0 156100.0 237200.0 ;
      RECT  149500.0 233500.0 159100.0 232900.00000000003 ;
      RECT  149500.0 242700.0 159100.0 242100.00000000003 ;
      RECT  163500.0 234500.0 164300.0 233200.0 ;
      RECT  163500.0 242400.00000000003 164300.0 241100.00000000003 ;
      RECT  160300.0 241500.0 161100.0 242700.0 ;
      RECT  160300.0 235300.0 161100.0 232900.00000000003 ;
      RECT  162100.0 241500.0 162700.0 235300.0 ;
      RECT  160300.0 235300.0 161100.0 234500.0 ;
      RECT  161900.0 235300.0 162700.0 234500.0 ;
      RECT  161900.0 235300.0 162700.0 234500.0 ;
      RECT  160300.0 235300.0 161100.0 234500.0 ;
      RECT  160300.0 241500.0 161100.0 240700.0 ;
      RECT  161900.0 241500.0 162700.0 240700.0 ;
      RECT  161900.0 241500.0 162700.0 240700.0 ;
      RECT  160300.0 241500.0 161100.0 240700.0 ;
      RECT  163500.0 234900.00000000003 164300.0 234100.00000000003 ;
      RECT  163500.0 241500.0 164300.0 240700.0 ;
      RECT  160700.0 238400.00000000003 161500.0 237600.00000000003 ;
      RECT  160700.0 238400.00000000003 161500.0 237600.00000000003 ;
      RECT  162400.0 238300.0 163000.0 237700.0 ;
      RECT  159100.0 233500.0 165500.0 232900.00000000003 ;
      RECT  159100.0 242700.0 165500.0 242100.00000000003 ;
      RECT  150700.0 243700.0 151500.0 242100.00000000003 ;
      RECT  150700.0 249500.0 151500.0 251900.00000000003 ;
      RECT  153900.0 249500.0 154700.0 251900.00000000003 ;
      RECT  155500.0 250300.0 156300.0 251600.00000000003 ;
      RECT  155500.0 242400.00000000003 156300.0 243700.0 ;
      RECT  150700.0 249500.0 151500.0 250300.0 ;
      RECT  152300.0 249500.0 153100.0 250300.0 ;
      RECT  152300.0 249500.0 153100.0 250300.0 ;
      RECT  150700.0 249500.0 151500.0 250300.0 ;
      RECT  152300.0 249500.0 153100.0 250300.0 ;
      RECT  153900.0 249500.0 154700.0 250300.0 ;
      RECT  153900.0 249500.0 154700.0 250300.0 ;
      RECT  152300.0 249500.0 153100.0 250300.0 ;
      RECT  150700.0 243700.0 151500.0 244500.0 ;
      RECT  152300.0 243700.0 153100.0 244500.0 ;
      RECT  152300.0 243700.0 153100.0 244500.0 ;
      RECT  150700.0 243700.0 151500.0 244500.0 ;
      RECT  152300.0 243700.0 153100.0 244500.0 ;
      RECT  153900.0 243700.0 154700.0 244500.0 ;
      RECT  153900.0 243700.0 154700.0 244500.0 ;
      RECT  152300.0 243700.0 153100.0 244500.0 ;
      RECT  155500.0 249900.00000000003 156300.0 250700.0 ;
      RECT  155500.0 243300.0 156300.0 244100.00000000003 ;
      RECT  153900.0 245400.00000000003 153100.0 246200.0 ;
      RECT  151900.0 246800.0 151100.0 247600.00000000003 ;
      RECT  152300.0 249500.0 153100.0 250300.0 ;
      RECT  153900.0 243700.0 154700.0 244500.0 ;
      RECT  156100.0 246800.0 155300.0 247600.00000000003 ;
      RECT  151100.0 246800.0 151900.0 247600.00000000003 ;
      RECT  153100.0 245400.00000000003 153900.0 246200.0 ;
      RECT  155300.0 246800.0 156100.0 247600.00000000003 ;
      RECT  149500.0 251300.0 159100.0 251900.00000000003 ;
      RECT  149500.0 242100.00000000003 159100.0 242700.0 ;
      RECT  163500.0 250300.0 164300.0 251600.00000000003 ;
      RECT  163500.0 242400.00000000003 164300.0 243700.0 ;
      RECT  160300.0 243300.0 161100.0 242100.00000000003 ;
      RECT  160300.0 249500.0 161100.0 251900.00000000003 ;
      RECT  162100.0 243300.0 162700.0 249500.0 ;
      RECT  160300.0 249500.0 161100.0 250300.0 ;
      RECT  161900.0 249500.0 162700.0 250300.0 ;
      RECT  161900.0 249500.0 162700.0 250300.0 ;
      RECT  160300.0 249500.0 161100.0 250300.0 ;
      RECT  160300.0 243300.0 161100.0 244100.00000000003 ;
      RECT  161900.0 243300.0 162700.0 244100.00000000003 ;
      RECT  161900.0 243300.0 162700.0 244100.00000000003 ;
      RECT  160300.0 243300.0 161100.0 244100.00000000003 ;
      RECT  163500.0 249900.00000000003 164300.0 250700.0 ;
      RECT  163500.0 243300.0 164300.0 244100.00000000003 ;
      RECT  160700.0 246400.00000000003 161500.0 247200.0 ;
      RECT  160700.0 246400.00000000003 161500.0 247200.0 ;
      RECT  162400.0 246500.0 163000.0 247100.00000000003 ;
      RECT  159100.0 251300.0 165500.0 251900.00000000003 ;
      RECT  159100.0 242100.00000000003 165500.0 242700.0 ;
      RECT  150700.0 259500.0 151500.0 261100.00000000003 ;
      RECT  150700.0 253700.0 151500.0 251300.0 ;
      RECT  153900.0 253700.0 154700.0 251300.0 ;
      RECT  155500.0 252899.99999999997 156300.0 251600.00000000003 ;
      RECT  155500.0 260800.0 156300.0 259500.0 ;
      RECT  150700.0 253700.0 151500.0 252899.99999999997 ;
      RECT  152300.0 253700.0 153100.0 252899.99999999997 ;
      RECT  152300.0 253700.0 153100.0 252899.99999999997 ;
      RECT  150700.0 253700.0 151500.0 252899.99999999997 ;
      RECT  152300.0 253700.0 153100.0 252899.99999999997 ;
      RECT  153900.0 253700.0 154700.0 252899.99999999997 ;
      RECT  153900.0 253700.0 154700.0 252899.99999999997 ;
      RECT  152300.0 253700.0 153100.0 252899.99999999997 ;
      RECT  150700.0 259500.0 151500.0 258700.0 ;
      RECT  152300.0 259500.0 153100.0 258700.0 ;
      RECT  152300.0 259500.0 153100.0 258700.0 ;
      RECT  150700.0 259500.0 151500.0 258700.0 ;
      RECT  152300.0 259500.0 153100.0 258700.0 ;
      RECT  153900.0 259500.0 154700.0 258700.0 ;
      RECT  153900.0 259500.0 154700.0 258700.0 ;
      RECT  152300.0 259500.0 153100.0 258700.0 ;
      RECT  155500.0 253300.0 156300.0 252500.0 ;
      RECT  155500.0 259899.99999999997 156300.0 259100.00000000003 ;
      RECT  153900.0 257800.0 153100.0 257000.0 ;
      RECT  151900.0 256399.99999999997 151100.0 255600.00000000003 ;
      RECT  152300.0 253700.0 153100.0 252899.99999999997 ;
      RECT  153900.0 259500.0 154700.0 258700.0 ;
      RECT  156100.0 256399.99999999997 155300.0 255600.00000000003 ;
      RECT  151100.0 256399.99999999997 151900.0 255600.00000000003 ;
      RECT  153100.0 257800.0 153900.0 257000.0 ;
      RECT  155300.0 256399.99999999997 156100.0 255600.00000000003 ;
      RECT  149500.0 251899.99999999997 159100.0 251300.0 ;
      RECT  149500.0 261100.00000000003 159100.0 260500.0 ;
      RECT  163500.0 252899.99999999997 164300.0 251600.00000000003 ;
      RECT  163500.0 260800.0 164300.0 259500.0 ;
      RECT  160300.0 259899.99999999997 161100.0 261100.00000000003 ;
      RECT  160300.0 253700.0 161100.0 251300.0 ;
      RECT  162100.0 259899.99999999997 162700.0 253700.0 ;
      RECT  160300.0 253700.0 161100.0 252899.99999999997 ;
      RECT  161900.0 253700.0 162700.0 252899.99999999997 ;
      RECT  161900.0 253700.0 162700.0 252899.99999999997 ;
      RECT  160300.0 253700.0 161100.0 252899.99999999997 ;
      RECT  160300.0 259899.99999999997 161100.0 259100.00000000003 ;
      RECT  161900.0 259899.99999999997 162700.0 259100.00000000003 ;
      RECT  161900.0 259899.99999999997 162700.0 259100.00000000003 ;
      RECT  160300.0 259899.99999999997 161100.0 259100.00000000003 ;
      RECT  163500.0 253300.0 164300.0 252500.0 ;
      RECT  163500.0 259899.99999999997 164300.0 259100.00000000003 ;
      RECT  160700.0 256800.0 161500.0 256000.0 ;
      RECT  160700.0 256800.0 161500.0 256000.0 ;
      RECT  162400.0 256700.0 163000.0 256100.00000000003 ;
      RECT  159100.0 251899.99999999997 165500.0 251300.0 ;
      RECT  159100.0 261100.00000000003 165500.0 260500.0 ;
      RECT  150700.0 262100.00000000003 151500.0 260500.0 ;
      RECT  150700.0 267900.0 151500.0 270300.0 ;
      RECT  153900.0 267900.0 154700.0 270300.0 ;
      RECT  155500.0 268700.0 156300.0 270000.0 ;
      RECT  155500.0 260800.0 156300.0 262100.00000000003 ;
      RECT  150700.0 267900.0 151500.0 268700.0 ;
      RECT  152300.0 267900.0 153100.0 268700.0 ;
      RECT  152300.0 267900.0 153100.0 268700.0 ;
      RECT  150700.0 267900.0 151500.0 268700.0 ;
      RECT  152300.0 267900.0 153100.0 268700.0 ;
      RECT  153900.0 267900.0 154700.0 268700.0 ;
      RECT  153900.0 267900.0 154700.0 268700.0 ;
      RECT  152300.0 267900.0 153100.0 268700.0 ;
      RECT  150700.0 262100.00000000003 151500.0 262900.0 ;
      RECT  152300.0 262100.00000000003 153100.0 262900.0 ;
      RECT  152300.0 262100.00000000003 153100.0 262900.0 ;
      RECT  150700.0 262100.00000000003 151500.0 262900.0 ;
      RECT  152300.0 262100.00000000003 153100.0 262900.0 ;
      RECT  153900.0 262100.00000000003 154700.0 262900.0 ;
      RECT  153900.0 262100.00000000003 154700.0 262900.0 ;
      RECT  152300.0 262100.00000000003 153100.0 262900.0 ;
      RECT  155500.0 268300.0 156300.0 269100.0 ;
      RECT  155500.0 261700.0 156300.0 262500.0 ;
      RECT  153900.0 263800.0 153100.0 264600.0 ;
      RECT  151900.0 265200.0 151100.0 266000.0 ;
      RECT  152300.0 267900.0 153100.0 268700.0 ;
      RECT  153900.0 262100.00000000003 154700.0 262900.0 ;
      RECT  156100.0 265200.0 155300.0 266000.0 ;
      RECT  151100.0 265200.0 151900.0 266000.0 ;
      RECT  153100.0 263800.0 153900.0 264600.0 ;
      RECT  155300.0 265200.0 156100.0 266000.0 ;
      RECT  149500.0 269700.0 159100.0 270300.0 ;
      RECT  149500.0 260500.0 159100.0 261100.00000000003 ;
      RECT  163500.0 268700.0 164300.0 270000.0 ;
      RECT  163500.0 260800.0 164300.0 262100.00000000003 ;
      RECT  160300.0 261700.0 161100.0 260500.0 ;
      RECT  160300.0 267900.0 161100.0 270300.0 ;
      RECT  162100.0 261700.0 162700.0 267900.0 ;
      RECT  160300.0 267900.0 161100.0 268700.0 ;
      RECT  161900.0 267900.0 162700.0 268700.0 ;
      RECT  161900.0 267900.0 162700.0 268700.0 ;
      RECT  160300.0 267900.0 161100.0 268700.0 ;
      RECT  160300.0 261700.0 161100.0 262500.0 ;
      RECT  161900.0 261700.0 162700.0 262500.0 ;
      RECT  161900.0 261700.0 162700.0 262500.0 ;
      RECT  160300.0 261700.0 161100.0 262500.0 ;
      RECT  163500.0 268300.0 164300.0 269100.0 ;
      RECT  163500.0 261700.0 164300.0 262500.0 ;
      RECT  160700.0 264800.0 161500.0 265600.0 ;
      RECT  160700.0 264800.0 161500.0 265600.0 ;
      RECT  162400.0 264900.0 163000.0 265500.0 ;
      RECT  159100.0 269700.0 165500.0 270300.0 ;
      RECT  159100.0 260500.0 165500.0 261100.00000000003 ;
      RECT  150700.0 277900.00000000006 151500.0 279500.0 ;
      RECT  150700.0 272100.0 151500.0 269700.0 ;
      RECT  153900.0 272100.0 154700.0 269700.0 ;
      RECT  155500.0 271300.0 156300.0 270000.0 ;
      RECT  155500.0 279200.0 156300.0 277900.00000000006 ;
      RECT  150700.0 272100.0 151500.0 271300.0 ;
      RECT  152300.0 272100.0 153100.0 271300.0 ;
      RECT  152300.0 272100.0 153100.0 271300.0 ;
      RECT  150700.0 272100.0 151500.0 271300.0 ;
      RECT  152300.0 272100.0 153100.0 271300.0 ;
      RECT  153900.0 272100.0 154700.0 271300.0 ;
      RECT  153900.0 272100.0 154700.0 271300.0 ;
      RECT  152300.0 272100.0 153100.0 271300.0 ;
      RECT  150700.0 277900.00000000006 151500.0 277100.0 ;
      RECT  152300.0 277900.00000000006 153100.0 277100.0 ;
      RECT  152300.0 277900.00000000006 153100.0 277100.0 ;
      RECT  150700.0 277900.00000000006 151500.0 277100.0 ;
      RECT  152300.0 277900.00000000006 153100.0 277100.0 ;
      RECT  153900.0 277900.00000000006 154700.0 277100.0 ;
      RECT  153900.0 277900.00000000006 154700.0 277100.0 ;
      RECT  152300.0 277900.00000000006 153100.0 277100.0 ;
      RECT  155500.0 271700.0 156300.0 270900.00000000006 ;
      RECT  155500.0 278300.0 156300.0 277500.0 ;
      RECT  153900.0 276200.0 153100.0 275400.00000000006 ;
      RECT  151900.0 274800.0 151100.0 274000.0 ;
      RECT  152300.0 272100.0 153100.0 271300.0 ;
      RECT  153900.0 277900.00000000006 154700.0 277100.0 ;
      RECT  156100.0 274800.0 155300.0 274000.0 ;
      RECT  151100.0 274800.0 151900.0 274000.0 ;
      RECT  153100.0 276200.0 153900.0 275400.00000000006 ;
      RECT  155300.0 274800.0 156100.0 274000.0 ;
      RECT  149500.0 270300.0 159100.0 269700.0 ;
      RECT  149500.0 279500.0 159100.0 278900.00000000006 ;
      RECT  163500.0 271300.0 164300.0 270000.0 ;
      RECT  163500.0 279200.0 164300.0 277900.00000000006 ;
      RECT  160300.0 278300.0 161100.0 279500.0 ;
      RECT  160300.0 272100.0 161100.0 269700.0 ;
      RECT  162100.0 278300.0 162700.0 272100.0 ;
      RECT  160300.0 272100.0 161100.0 271300.0 ;
      RECT  161900.0 272100.0 162700.0 271300.0 ;
      RECT  161900.0 272100.0 162700.0 271300.0 ;
      RECT  160300.0 272100.0 161100.0 271300.0 ;
      RECT  160300.0 278300.0 161100.0 277500.0 ;
      RECT  161900.0 278300.0 162700.0 277500.0 ;
      RECT  161900.0 278300.0 162700.0 277500.0 ;
      RECT  160300.0 278300.0 161100.0 277500.0 ;
      RECT  163500.0 271700.0 164300.0 270900.00000000006 ;
      RECT  163500.0 278300.0 164300.0 277500.0 ;
      RECT  160700.0 275200.0 161500.0 274400.00000000006 ;
      RECT  160700.0 275200.0 161500.0 274400.00000000006 ;
      RECT  162400.0 275100.0 163000.0 274500.0 ;
      RECT  159100.0 270300.0 165500.0 269700.0 ;
      RECT  159100.0 279500.0 165500.0 278900.00000000006 ;
      RECT  150700.0 280500.0 151500.0 278900.00000000006 ;
      RECT  150700.0 286300.0 151500.0 288700.0 ;
      RECT  153900.0 286300.0 154700.0 288700.0 ;
      RECT  155500.0 287100.0 156300.0 288400.00000000006 ;
      RECT  155500.0 279200.0 156300.0 280500.0 ;
      RECT  150700.0 286300.0 151500.0 287100.0 ;
      RECT  152300.0 286300.0 153100.0 287100.0 ;
      RECT  152300.0 286300.0 153100.0 287100.0 ;
      RECT  150700.0 286300.0 151500.0 287100.0 ;
      RECT  152300.0 286300.0 153100.0 287100.0 ;
      RECT  153900.0 286300.0 154700.0 287100.0 ;
      RECT  153900.0 286300.0 154700.0 287100.0 ;
      RECT  152300.0 286300.0 153100.0 287100.0 ;
      RECT  150700.0 280500.0 151500.0 281300.0 ;
      RECT  152300.0 280500.0 153100.0 281300.0 ;
      RECT  152300.0 280500.0 153100.0 281300.0 ;
      RECT  150700.0 280500.0 151500.0 281300.0 ;
      RECT  152300.0 280500.0 153100.0 281300.0 ;
      RECT  153900.0 280500.0 154700.0 281300.0 ;
      RECT  153900.0 280500.0 154700.0 281300.0 ;
      RECT  152300.0 280500.0 153100.0 281300.0 ;
      RECT  155500.0 286700.0 156300.0 287500.0 ;
      RECT  155500.0 280100.0 156300.0 280900.00000000006 ;
      RECT  153900.0 282200.0 153100.0 283000.0 ;
      RECT  151900.0 283600.0 151100.0 284400.00000000006 ;
      RECT  152300.0 286300.0 153100.0 287100.0 ;
      RECT  153900.0 280500.0 154700.0 281300.0 ;
      RECT  156100.0 283600.0 155300.0 284400.00000000006 ;
      RECT  151100.0 283600.0 151900.0 284400.00000000006 ;
      RECT  153100.0 282200.0 153900.0 283000.0 ;
      RECT  155300.0 283600.0 156100.0 284400.00000000006 ;
      RECT  149500.0 288100.0 159100.0 288700.0 ;
      RECT  149500.0 278900.00000000006 159100.0 279500.0 ;
      RECT  163500.0 287100.0 164300.0 288400.00000000006 ;
      RECT  163500.0 279200.0 164300.0 280500.0 ;
      RECT  160300.0 280100.0 161100.0 278900.00000000006 ;
      RECT  160300.0 286300.0 161100.0 288700.0 ;
      RECT  162100.0 280100.0 162700.0 286300.0 ;
      RECT  160300.0 286300.0 161100.0 287100.0 ;
      RECT  161900.0 286300.0 162700.0 287100.0 ;
      RECT  161900.0 286300.0 162700.0 287100.0 ;
      RECT  160300.0 286300.0 161100.0 287100.0 ;
      RECT  160300.0 280100.0 161100.0 280900.00000000006 ;
      RECT  161900.0 280100.0 162700.0 280900.00000000006 ;
      RECT  161900.0 280100.0 162700.0 280900.00000000006 ;
      RECT  160300.0 280100.0 161100.0 280900.00000000006 ;
      RECT  163500.0 286700.0 164300.0 287500.0 ;
      RECT  163500.0 280100.0 164300.0 280900.00000000006 ;
      RECT  160700.0 283200.0 161500.0 284000.0 ;
      RECT  160700.0 283200.0 161500.0 284000.0 ;
      RECT  162400.0 283300.0 163000.0 283900.00000000006 ;
      RECT  159100.0 288100.0 165500.0 288700.0 ;
      RECT  159100.0 278900.00000000006 165500.0 279500.0 ;
      RECT  150700.0 296300.0 151500.0 297900.00000000006 ;
      RECT  150700.0 290500.0 151500.0 288100.0 ;
      RECT  153900.0 290500.0 154700.0 288100.0 ;
      RECT  155500.0 289700.0 156300.0 288400.00000000006 ;
      RECT  155500.0 297600.0 156300.0 296300.0 ;
      RECT  150700.0 290500.0 151500.0 289700.0 ;
      RECT  152300.0 290500.0 153100.0 289700.0 ;
      RECT  152300.0 290500.0 153100.0 289700.0 ;
      RECT  150700.0 290500.0 151500.0 289700.0 ;
      RECT  152300.0 290500.0 153100.0 289700.0 ;
      RECT  153900.0 290500.0 154700.0 289700.0 ;
      RECT  153900.0 290500.0 154700.0 289700.0 ;
      RECT  152300.0 290500.0 153100.0 289700.0 ;
      RECT  150700.0 296300.0 151500.0 295500.0 ;
      RECT  152300.0 296300.0 153100.0 295500.0 ;
      RECT  152300.0 296300.0 153100.0 295500.0 ;
      RECT  150700.0 296300.0 151500.0 295500.0 ;
      RECT  152300.0 296300.0 153100.0 295500.0 ;
      RECT  153900.0 296300.0 154700.0 295500.0 ;
      RECT  153900.0 296300.0 154700.0 295500.0 ;
      RECT  152300.0 296300.0 153100.0 295500.0 ;
      RECT  155500.0 290100.0 156300.0 289300.0 ;
      RECT  155500.0 296700.0 156300.0 295900.00000000006 ;
      RECT  153900.0 294600.0 153100.0 293800.0 ;
      RECT  151900.0 293200.0 151100.0 292400.00000000006 ;
      RECT  152300.0 290500.0 153100.0 289700.0 ;
      RECT  153900.0 296300.0 154700.0 295500.0 ;
      RECT  156100.0 293200.0 155300.0 292400.00000000006 ;
      RECT  151100.0 293200.0 151900.0 292400.00000000006 ;
      RECT  153100.0 294600.0 153900.0 293800.0 ;
      RECT  155300.0 293200.0 156100.0 292400.00000000006 ;
      RECT  149500.0 288700.0 159100.0 288100.0 ;
      RECT  149500.0 297900.00000000006 159100.0 297300.0 ;
      RECT  163500.0 289700.0 164300.0 288400.00000000006 ;
      RECT  163500.0 297600.0 164300.0 296300.0 ;
      RECT  160300.0 296700.0 161100.0 297900.00000000006 ;
      RECT  160300.0 290500.0 161100.0 288100.0 ;
      RECT  162100.0 296700.0 162700.0 290500.0 ;
      RECT  160300.0 290500.0 161100.0 289700.0 ;
      RECT  161900.0 290500.0 162700.0 289700.0 ;
      RECT  161900.0 290500.0 162700.0 289700.0 ;
      RECT  160300.0 290500.0 161100.0 289700.0 ;
      RECT  160300.0 296700.0 161100.0 295900.00000000006 ;
      RECT  161900.0 296700.0 162700.0 295900.00000000006 ;
      RECT  161900.0 296700.0 162700.0 295900.00000000006 ;
      RECT  160300.0 296700.0 161100.0 295900.00000000006 ;
      RECT  163500.0 290100.0 164300.0 289300.0 ;
      RECT  163500.0 296700.0 164300.0 295900.00000000006 ;
      RECT  160700.0 293600.0 161500.0 292800.0 ;
      RECT  160700.0 293600.0 161500.0 292800.0 ;
      RECT  162400.0 293500.0 163000.0 292900.00000000006 ;
      RECT  159100.0 288700.0 165500.0 288100.0 ;
      RECT  159100.0 297900.00000000006 165500.0 297300.0 ;
      RECT  150700.0 298900.00000000006 151500.0 297300.0 ;
      RECT  150700.0 304700.0 151500.0 307100.0 ;
      RECT  153900.0 304700.0 154700.0 307100.0 ;
      RECT  155500.0 305500.0 156300.0 306800.0 ;
      RECT  155500.0 297600.0 156300.0 298900.00000000006 ;
      RECT  150700.0 304700.0 151500.0 305500.0 ;
      RECT  152300.0 304700.0 153100.0 305500.0 ;
      RECT  152300.0 304700.0 153100.0 305500.0 ;
      RECT  150700.0 304700.0 151500.0 305500.0 ;
      RECT  152300.0 304700.0 153100.0 305500.0 ;
      RECT  153900.0 304700.0 154700.0 305500.0 ;
      RECT  153900.0 304700.0 154700.0 305500.0 ;
      RECT  152300.0 304700.0 153100.0 305500.0 ;
      RECT  150700.0 298900.00000000006 151500.0 299700.0 ;
      RECT  152300.0 298900.00000000006 153100.0 299700.0 ;
      RECT  152300.0 298900.00000000006 153100.0 299700.0 ;
      RECT  150700.0 298900.00000000006 151500.0 299700.0 ;
      RECT  152300.0 298900.00000000006 153100.0 299700.0 ;
      RECT  153900.0 298900.00000000006 154700.0 299700.0 ;
      RECT  153900.0 298900.00000000006 154700.0 299700.0 ;
      RECT  152300.0 298900.00000000006 153100.0 299700.0 ;
      RECT  155500.0 305100.0 156300.0 305900.00000000006 ;
      RECT  155500.0 298500.0 156300.0 299300.0 ;
      RECT  153900.0 300600.0 153100.0 301400.00000000006 ;
      RECT  151900.0 302000.0 151100.0 302800.0 ;
      RECT  152300.0 304700.0 153100.0 305500.0 ;
      RECT  153900.0 298900.00000000006 154700.0 299700.0 ;
      RECT  156100.0 302000.0 155300.0 302800.0 ;
      RECT  151100.0 302000.0 151900.0 302800.0 ;
      RECT  153100.0 300600.0 153900.0 301400.00000000006 ;
      RECT  155300.0 302000.0 156100.0 302800.0 ;
      RECT  149500.0 306500.0 159100.0 307100.0 ;
      RECT  149500.0 297300.0 159100.0 297900.00000000006 ;
      RECT  163500.0 305500.0 164300.0 306800.0 ;
      RECT  163500.0 297600.0 164300.0 298900.00000000006 ;
      RECT  160300.0 298500.0 161100.0 297300.0 ;
      RECT  160300.0 304700.0 161100.0 307100.0 ;
      RECT  162100.0 298500.0 162700.0 304700.0 ;
      RECT  160300.0 304700.0 161100.0 305500.0 ;
      RECT  161900.0 304700.0 162700.0 305500.0 ;
      RECT  161900.0 304700.0 162700.0 305500.0 ;
      RECT  160300.0 304700.0 161100.0 305500.0 ;
      RECT  160300.0 298500.0 161100.0 299300.0 ;
      RECT  161900.0 298500.0 162700.0 299300.0 ;
      RECT  161900.0 298500.0 162700.0 299300.0 ;
      RECT  160300.0 298500.0 161100.0 299300.0 ;
      RECT  163500.0 305100.0 164300.0 305900.00000000006 ;
      RECT  163500.0 298500.0 164300.0 299300.0 ;
      RECT  160700.0 301600.0 161500.0 302400.00000000006 ;
      RECT  160700.0 301600.0 161500.0 302400.00000000006 ;
      RECT  162400.0 301700.0 163000.0 302300.0 ;
      RECT  159100.0 306500.0 165500.0 307100.0 ;
      RECT  159100.0 297300.0 165500.0 297900.00000000006 ;
      RECT  150700.0 314700.0 151500.0 316300.0 ;
      RECT  150700.0 308900.00000000006 151500.0 306500.0 ;
      RECT  153900.0 308900.00000000006 154700.0 306500.0 ;
      RECT  155500.0 308100.0 156300.0 306800.0 ;
      RECT  155500.0 316000.0 156300.0 314700.0 ;
      RECT  150700.0 308900.00000000006 151500.0 308100.0 ;
      RECT  152300.0 308900.00000000006 153100.0 308100.0 ;
      RECT  152300.0 308900.00000000006 153100.0 308100.0 ;
      RECT  150700.0 308900.00000000006 151500.0 308100.0 ;
      RECT  152300.0 308900.00000000006 153100.0 308100.0 ;
      RECT  153900.0 308900.00000000006 154700.0 308100.0 ;
      RECT  153900.0 308900.00000000006 154700.0 308100.0 ;
      RECT  152300.0 308900.00000000006 153100.0 308100.0 ;
      RECT  150700.0 314700.0 151500.0 313900.00000000006 ;
      RECT  152300.0 314700.0 153100.0 313900.00000000006 ;
      RECT  152300.0 314700.0 153100.0 313900.00000000006 ;
      RECT  150700.0 314700.0 151500.0 313900.00000000006 ;
      RECT  152300.0 314700.0 153100.0 313900.00000000006 ;
      RECT  153900.0 314700.0 154700.0 313900.00000000006 ;
      RECT  153900.0 314700.0 154700.0 313900.00000000006 ;
      RECT  152300.0 314700.0 153100.0 313900.00000000006 ;
      RECT  155500.0 308500.0 156300.0 307700.0 ;
      RECT  155500.0 315100.0 156300.0 314300.0 ;
      RECT  153900.0 313000.0 153100.0 312200.0 ;
      RECT  151900.0 311600.0 151100.0 310800.0 ;
      RECT  152300.0 308900.00000000006 153100.0 308100.0 ;
      RECT  153900.0 314700.0 154700.0 313900.00000000006 ;
      RECT  156100.0 311600.0 155300.0 310800.0 ;
      RECT  151100.0 311600.0 151900.0 310800.0 ;
      RECT  153100.0 313000.0 153900.0 312200.0 ;
      RECT  155300.0 311600.0 156100.0 310800.0 ;
      RECT  149500.0 307100.0 159100.0 306500.0 ;
      RECT  149500.0 316300.0 159100.0 315700.0 ;
      RECT  163500.0 308100.0 164300.0 306800.0 ;
      RECT  163500.0 316000.0 164300.0 314700.0 ;
      RECT  160300.0 315100.0 161100.0 316300.0 ;
      RECT  160300.0 308900.00000000006 161100.0 306500.0 ;
      RECT  162100.0 315100.0 162700.0 308900.00000000006 ;
      RECT  160300.0 308900.00000000006 161100.0 308100.0 ;
      RECT  161900.0 308900.00000000006 162700.0 308100.0 ;
      RECT  161900.0 308900.00000000006 162700.0 308100.0 ;
      RECT  160300.0 308900.00000000006 161100.0 308100.0 ;
      RECT  160300.0 315100.0 161100.0 314300.0 ;
      RECT  161900.0 315100.0 162700.0 314300.0 ;
      RECT  161900.0 315100.0 162700.0 314300.0 ;
      RECT  160300.0 315100.0 161100.0 314300.0 ;
      RECT  163500.0 308500.0 164300.0 307700.0 ;
      RECT  163500.0 315100.0 164300.0 314300.0 ;
      RECT  160700.0 312000.0 161500.0 311200.0 ;
      RECT  160700.0 312000.0 161500.0 311200.0 ;
      RECT  162400.0 311900.00000000006 163000.0 311300.0 ;
      RECT  159100.0 307100.0 165500.0 306500.0 ;
      RECT  159100.0 316300.0 165500.0 315700.0 ;
      RECT  147000.0 173200.0 147800.0 174000.0 ;
      RECT  148300.0 171200.0 149100.0 172000.0 ;
      RECT  153100.0 171800.0 152300.0 172600.00000000003 ;
      RECT  147000.0 182000.0 147800.0 182800.0 ;
      RECT  148300.0 184000.0 149100.0 184800.0 ;
      RECT  153100.0 183400.0 152300.0 184200.0 ;
      RECT  147000.0 191600.00000000003 147800.0 192400.0 ;
      RECT  148300.0 189600.00000000003 149100.0 190400.0 ;
      RECT  153100.0 190200.0 152300.0 191000.0 ;
      RECT  147000.0 200399.99999999997 147800.0 201200.0 ;
      RECT  148300.0 202399.99999999997 149100.0 203200.0 ;
      RECT  153100.0 201800.0 152300.0 202600.00000000003 ;
      RECT  147000.0 210000.0 147800.0 210800.0 ;
      RECT  148300.0 208000.0 149100.0 208800.0 ;
      RECT  153100.0 208600.00000000003 152300.0 209399.99999999997 ;
      RECT  147000.0 218800.0 147800.0 219600.00000000003 ;
      RECT  148300.0 220800.0 149100.0 221600.00000000003 ;
      RECT  153100.0 220200.0 152300.0 221000.0 ;
      RECT  147000.0 228399.99999999997 147800.0 229200.0 ;
      RECT  148300.0 226399.99999999997 149100.0 227200.0 ;
      RECT  153100.0 227000.0 152300.0 227800.0 ;
      RECT  147000.0 237200.0 147800.0 238000.0 ;
      RECT  148300.0 239200.0 149100.0 240000.0 ;
      RECT  153100.0 238600.00000000003 152300.0 239399.99999999997 ;
      RECT  147000.0 246800.0 147800.0 247600.00000000003 ;
      RECT  148300.0 244800.0 149100.0 245600.00000000003 ;
      RECT  153100.0 245400.00000000003 152300.0 246200.0 ;
      RECT  147000.0 255600.00000000003 147800.0 256400.00000000003 ;
      RECT  148300.0 257600.00000000003 149100.0 258400.00000000003 ;
      RECT  153100.0 257000.0 152300.0 257800.0 ;
      RECT  147000.0 265200.0 147800.0 266000.0 ;
      RECT  148300.0 263200.0 149100.0 264000.0 ;
      RECT  153100.0 263800.0 152300.0 264600.0 ;
      RECT  147000.0 274000.0 147800.0 274800.0 ;
      RECT  148300.0 276000.0 149100.0 276800.0 ;
      RECT  153100.0 275400.00000000006 152300.0 276200.0 ;
      RECT  147000.0 283600.0 147800.0 284400.00000000006 ;
      RECT  148300.0 281600.0 149100.0 282400.00000000006 ;
      RECT  153100.0 282200.0 152300.0 283000.0 ;
      RECT  147000.0 292400.00000000006 147800.0 293200.0 ;
      RECT  148300.0 294400.00000000006 149100.0 295200.0 ;
      RECT  153100.0 293800.0 152300.0 294600.0 ;
      RECT  147000.0 302000.0 147800.0 302800.0 ;
      RECT  148300.0 300000.0 149100.0 300800.0 ;
      RECT  153100.0 300600.0 152300.0 301400.00000000006 ;
      RECT  147000.0 310800.0 147800.0 311600.0 ;
      RECT  148300.0 312800.0 149100.0 313600.0 ;
      RECT  153100.0 312200.0 152300.0 313000.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 168400.0 158700.0 169200.0 ;
      RECT  159500.0 168400.0 158700.0 169200.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 315600.0 158700.0 316400.00000000006 ;
      RECT  159500.0 315600.0 158700.0 316400.00000000006 ;
      RECT  145300.0 171300.0 148700.0 171900.0 ;
      RECT  145300.0 184100.00000000003 148700.0 184700.0 ;
      RECT  145300.0 189700.0 148700.0 190300.0 ;
      RECT  145300.0 202500.0 148700.0 203100.00000000003 ;
      RECT  145300.0 208100.00000000003 148700.0 208700.0 ;
      RECT  145300.0 220899.99999999997 148700.0 221500.0 ;
      RECT  145300.0 226500.0 148700.0 227100.00000000003 ;
      RECT  145300.0 239300.0 148700.0 239900.00000000003 ;
      RECT  145300.0 244900.00000000003 148700.0 245500.0 ;
      RECT  145300.0 257700.0 148700.0 258300.0 ;
      RECT  145300.0 263300.0 148700.0 263900.00000000006 ;
      RECT  145300.0 276100.0 148700.0 276700.0 ;
      RECT  145300.0 281700.0 148700.0 282300.0 ;
      RECT  145300.0 294500.0 148700.0 295100.0 ;
      RECT  145300.0 300100.0 148700.0 300700.0 ;
      RECT  145300.0 312900.0 148700.0 313500.0 ;
      RECT  162400.0 172900.0 163000.0 173500.0 ;
      RECT  162400.0 182500.0 163000.0 183100.00000000003 ;
      RECT  162400.0 191300.0 163000.0 191900.0 ;
      RECT  162400.0 200899.99999999997 163000.0 201500.0 ;
      RECT  162400.0 209700.0 163000.0 210300.0 ;
      RECT  162400.0 219300.0 163000.0 219899.99999999997 ;
      RECT  162400.0 228100.00000000003 163000.0 228700.0 ;
      RECT  162400.0 237700.0 163000.0 238300.0 ;
      RECT  162400.0 246500.0 163000.0 247100.00000000003 ;
      RECT  162400.0 256100.00000000003 163000.0 256700.0 ;
      RECT  162400.0 264900.00000000006 163000.0 265500.0 ;
      RECT  162400.0 274500.0 163000.0 275100.0 ;
      RECT  162400.0 283300.0 163000.0 283900.00000000006 ;
      RECT  162400.0 292900.00000000006 163000.0 293500.0 ;
      RECT  162400.0 301700.0 163000.0 302300.0 ;
      RECT  162400.0 311300.0 163000.0 311900.0 ;
      RECT  170100.00000000003 154700.0 169300.0 155500.0 ;
      RECT  167300.0 74900.0 166500.0 75700.0 ;
      RECT  168700.0 144500.0 167900.0 145300.0 ;
      RECT  147800.0 164200.0 147000.0 165000.0 ;
      RECT  165900.0 164200.0 165100.00000000003 165000.0 ;
      RECT  5499.999999999991 43900.00000000001 41499.99999999999 44500.00000000001 ;
      RECT  37299.99999999999 71900.0 48799.99999999999 72500.0 ;
      RECT  40099.99999999999 90700.00000000001 48800.0 91300.00000000001 ;
      RECT  37299.99999999999 116300.00000000001 48799.99999999999 116900.0 ;
      RECT  42899.99999999999 117700.00000000001 50799.99999999999 118300.00000000001 ;
      RECT  38699.99999999999 125900.0 48800.0 126500.0 ;
      RECT  42899.99999999999 124500.00000000001 50799.99999999999 125100.00000000001 ;
      RECT  59999.99999999999 130300.00000000001 64399.99999999999 130900.0 ;
      RECT  11599.999999999993 151500.0 48400.0 152100.0 ;
      RECT  41499.99999999999 31300.000000000007 48800.0 31900.00000000001 ;
      RECT  56899.99999999999 31300.000000000007 57499.99999999999 31900.00000000001 ;
      RECT  50399.99999999999 31300.000000000007 57199.999999999985 31900.00000000001 ;
      RECT  56899.99999999999 31600.000000000007 57499.99999999999 38000.00000000001 ;
      RECT  41499.99999999999 45900.00000000001 48800.0 46500.00000000001 ;
      RECT  44300.0 44500.00000000001 50800.0 45100.00000000001 ;
      RECT  59599.99999999999 21100.000000000007 70800.0 21700.00000000001 ;
      RECT  59599.99999999999 1100.0000000000057 70800.0 1700.0000000000057 ;
      RECT  69199.99999999999 21100.000000000007 70799.99999999999 21700.00000000001 ;
      RECT  69199.99999999999 41100.00000000001 70799.99999999999 41700.00000000001 ;
      RECT  62800.0 61100.00000000001 70800.0 61700.00000000001 ;
      RECT  62800.0 41100.00000000001 70800.0 41700.00000000001 ;
      RECT  64399.99999999999 61100.00000000001 70800.0 61700.00000000001 ;
      RECT  64399.99999999999 81100.00000000001 70800.0 81700.0 ;
      RECT  61199.99999999999 101100.00000000001 70800.0 101700.0 ;
      RECT  61199.99999999999 81100.00000000001 70800.0 81700.0 ;
      RECT  62800.0 101100.00000000001 70800.0 101700.0 ;
      RECT  62800.0 121100.00000000001 70800.0 121700.0 ;
      RECT  61199.99999999999 141100.00000000003 70800.0 141700.00000000003 ;
      RECT  61199.99999999999 161100.00000000003 70800.0 161700.00000000003 ;
      RECT  29899.999999999993 10700.000000000007 30499.999999999993 11300.000000000005 ;
      RECT  29899.999999999993 10300.000000000005 30499.999999999993 10900.000000000005 ;
      RECT  27799.999999999993 10700.000000000007 30199.999999999996 11300.000000000005 ;
      RECT  29899.999999999993 10600.000000000007 30499.999999999993 11000.000000000007 ;
      RECT  30199.999999999993 10300.000000000005 32599.999999999993 10900.000000000005 ;
      RECT  35299.99999999999 10300.000000000005 35899.99999999999 10900.000000000005 ;
      RECT  34199.999999999985 10300.000000000005 35599.99999999999 10900.000000000005 ;
      RECT  35299.99999999999 9200.000000000007 35899.99999999999 10600.000000000007 ;
      RECT  29899.999999999993 11000.000000000007 30499.999999999993 12400.000000000007 ;
      RECT  2399.9999999999914 1400.0000000000057 24199.999999999993 21400.000000000007 ;
      RECT  28599.999999999993 20100.000000000004 29399.999999999993 21400.000000000007 ;
      RECT  28599.999999999993 1400.0000000000057 29399.999999999993 2700.0000000000055 ;
      RECT  25399.999999999993 2700.0000000000055 26199.999999999993 1100.0000000000057 ;
      RECT  25399.999999999993 18500.000000000007 26199.999999999993 21700.000000000007 ;
      RECT  27199.999999999993 2700.0000000000055 27799.999999999993 18500.000000000007 ;
      RECT  25399.999999999993 18500.000000000007 26199.999999999993 19300.000000000004 ;
      RECT  26999.999999999993 18500.000000000007 27799.999999999993 19300.000000000004 ;
      RECT  26999.999999999993 18500.000000000007 27799.999999999993 19300.000000000004 ;
      RECT  25399.999999999993 18500.000000000007 26199.999999999993 19300.000000000004 ;
      RECT  25399.999999999993 2700.0000000000055 26199.999999999993 3500.000000000006 ;
      RECT  26999.999999999993 2700.0000000000055 27799.999999999993 3500.000000000006 ;
      RECT  26999.999999999993 2700.0000000000055 27799.999999999993 3500.000000000006 ;
      RECT  25399.999999999993 2700.0000000000055 26199.999999999993 3500.000000000006 ;
      RECT  28599.999999999993 19700.000000000007 29399.999999999993 20500.000000000007 ;
      RECT  28599.999999999993 2300.0000000000055 29399.999999999993 3100.000000000006 ;
      RECT  25799.999999999993 10600.000000000007 26599.999999999993 11400.000000000007 ;
      RECT  25799.999999999993 10600.000000000007 26599.999999999993 11400.000000000005 ;
      RECT  27499.999999999993 10700.000000000007 28099.999999999993 11300.000000000005 ;
      RECT  24199.999999999993 21100.000000000007 30599.999999999993 21700.000000000007 ;
      RECT  24199.999999999993 1100.0000000000057 30599.999999999993 1700.0000000000057 ;
      RECT  34999.99999999999 20100.000000000004 35800.0 21400.000000000007 ;
      RECT  34999.99999999999 1400.0000000000057 35800.0 2700.0000000000055 ;
      RECT  31799.999999999993 3500.000000000006 32599.999999999993 1100.0000000000055 ;
      RECT  31799.999999999993 16900.000000000007 32599.999999999993 21700.000000000007 ;
      RECT  33599.99999999999 3500.000000000006 34199.99999999999 16900.000000000007 ;
      RECT  31799.999999999993 16900.000000000007 32599.999999999993 17700.000000000007 ;
      RECT  33399.99999999999 16900.000000000007 34199.99999999999 17700.000000000007 ;
      RECT  33399.99999999999 16900.000000000007 34199.99999999999 17700.000000000007 ;
      RECT  31799.999999999993 16900.000000000007 32599.999999999993 17700.000000000007 ;
      RECT  31799.999999999993 3500.000000000006 32599.999999999993 4300.000000000006 ;
      RECT  33399.99999999999 3500.000000000006 34199.99999999999 4300.000000000006 ;
      RECT  33399.99999999999 3500.000000000006 34199.99999999999 4300.000000000006 ;
      RECT  31799.999999999993 3500.000000000006 32599.999999999993 4300.000000000006 ;
      RECT  34999.99999999999 19700.000000000007 35800.0 20500.000000000007 ;
      RECT  34999.99999999999 2300.0000000000055 35800.0 3100.000000000006 ;
      RECT  32199.999999999996 10200.000000000007 32999.99999999999 11000.000000000007 ;
      RECT  32199.999999999996 10200.000000000007 32999.99999999999 11000.000000000007 ;
      RECT  33899.99999999999 10300.000000000005 34499.99999999999 10900.000000000005 ;
      RECT  30599.999999999993 21100.000000000007 36999.99999999999 21700.000000000007 ;
      RECT  30599.999999999993 1100.0000000000057 36999.99999999999 1700.0000000000057 ;
      RECT  25799.999999999993 10600.000000000007 26599.999999999993 11400.000000000007 ;
      RECT  35199.99999999999 8800.000000000005 35999.99999999999 9600.000000000007 ;
      RECT  29799.999999999993 12000.000000000007 30599.999999999993 12800.000000000007 ;
      RECT  2399.9999999999914 20800.000000000007 36999.99999999999 22000.000000000007 ;
      RECT  2399.9999999999914 800.0000000000056 36999.99999999999 2000.0000000000057 ;
      RECT  29899.999999999993 32100.000000000007 30499.999999999993 31500.000000000007 ;
      RECT  29899.999999999993 32500.000000000007 30499.999999999993 31900.000000000007 ;
      RECT  27799.999999999993 32100.000000000007 30199.999999999996 31500.000000000007 ;
      RECT  29899.999999999993 32200.000000000004 30499.999999999993 31800.000000000004 ;
      RECT  30199.999999999993 32500.000000000007 32599.999999999993 31900.000000000007 ;
      RECT  35299.99999999999 32500.000000000007 35899.99999999999 31900.000000000007 ;
      RECT  34199.999999999985 32500.000000000007 35599.99999999999 31900.000000000007 ;
      RECT  35299.99999999999 33600.00000000001 35899.99999999999 32200.000000000004 ;
      RECT  29899.999999999993 31800.000000000004 30499.999999999993 30400.000000000007 ;
      RECT  2399.9999999999914 41400.00000000001 24199.999999999993 21400.000000000007 ;
      RECT  28599.999999999993 22700.000000000007 29399.999999999993 21400.000000000007 ;
      RECT  28599.999999999993 41400.00000000001 29399.999999999993 40100.00000000001 ;
      RECT  25399.999999999993 40100.00000000001 26199.999999999993 41700.0 ;
      RECT  25399.999999999993 24300.000000000004 26199.999999999993 21100.000000000004 ;
      RECT  27199.999999999993 40100.00000000001 27799.999999999993 24300.000000000004 ;
      RECT  25399.999999999993 24300.000000000004 26199.999999999993 23500.000000000007 ;
      RECT  26999.999999999993 24300.000000000004 27799.999999999993 23500.000000000007 ;
      RECT  26999.999999999993 24300.000000000004 27799.999999999993 23500.000000000007 ;
      RECT  25399.999999999993 24300.000000000004 26199.999999999993 23500.000000000007 ;
      RECT  25399.999999999993 40100.00000000001 26199.999999999993 39300.00000000001 ;
      RECT  26999.999999999993 40100.00000000001 27799.999999999993 39300.00000000001 ;
      RECT  26999.999999999993 40100.00000000001 27799.999999999993 39300.00000000001 ;
      RECT  25399.999999999993 40100.00000000001 26199.999999999993 39300.00000000001 ;
      RECT  28599.999999999993 23100.000000000004 29399.999999999993 22300.000000000004 ;
      RECT  28599.999999999993 40500.00000000001 29399.999999999993 39700.0 ;
      RECT  25799.999999999993 32200.000000000004 26599.999999999993 31400.000000000007 ;
      RECT  25799.999999999993 32200.000000000004 26599.999999999993 31400.000000000007 ;
      RECT  27499.999999999993 32100.000000000007 28099.999999999993 31500.000000000007 ;
      RECT  24199.999999999993 21700.000000000004 30599.999999999993 21100.000000000004 ;
      RECT  24199.999999999993 41700.0 30599.999999999993 41100.00000000001 ;
      RECT  34999.99999999999 22700.000000000007 35800.0 21400.000000000007 ;
      RECT  34999.99999999999 41400.00000000001 35800.0 40100.00000000001 ;
      RECT  31799.999999999993 39300.00000000001 32599.999999999993 41700.0 ;
      RECT  31799.999999999993 25900.000000000007 32599.999999999993 21100.000000000004 ;
      RECT  33599.99999999999 39300.00000000001 34199.99999999999 25900.000000000007 ;
      RECT  31799.999999999993 25900.000000000007 32599.999999999993 25100.000000000004 ;
      RECT  33399.99999999999 25900.000000000007 34199.99999999999 25100.000000000004 ;
      RECT  33399.99999999999 25900.000000000007 34199.99999999999 25100.000000000004 ;
      RECT  31799.999999999993 25900.000000000007 32599.999999999993 25100.000000000004 ;
      RECT  31799.999999999993 39300.00000000001 32599.999999999993 38500.00000000001 ;
      RECT  33399.99999999999 39300.00000000001 34199.99999999999 38500.00000000001 ;
      RECT  33399.99999999999 39300.00000000001 34199.99999999999 38500.00000000001 ;
      RECT  31799.999999999993 39300.00000000001 32599.999999999993 38500.00000000001 ;
      RECT  34999.99999999999 23100.000000000004 35800.0 22300.000000000004 ;
      RECT  34999.99999999999 40500.00000000001 35800.0 39700.0 ;
      RECT  32199.999999999996 32600.000000000007 32999.99999999999 31800.000000000004 ;
      RECT  32199.999999999996 32600.000000000007 32999.99999999999 31800.000000000004 ;
      RECT  33899.99999999999 32500.000000000007 34499.99999999999 31900.000000000007 ;
      RECT  30599.999999999993 21700.000000000004 36999.99999999999 21100.000000000004 ;
      RECT  30599.999999999993 41700.0 36999.99999999999 41100.00000000001 ;
      RECT  25799.999999999993 32200.000000000004 26599.999999999993 31400.000000000007 ;
      RECT  35199.99999999999 34000.00000000001 35999.99999999999 33200.0 ;
      RECT  29799.999999999993 30800.000000000004 30599.999999999993 30000.000000000004 ;
      RECT  2399.9999999999914 22000.000000000004 36999.99999999999 20800.000000000004 ;
      RECT  2399.9999999999914 42000.00000000001 36999.99999999999 40800.00000000001 ;
      RECT  2799.9999999999914 21000.000000000007 1999.9999999999916 21800.000000000007 ;
      RECT  2799.9999999999914 1000.0000000000058 1999.9999999999916 1800.0000000000057 ;
      RECT  2799.9999999999914 21000.000000000007 1999.9999999999916 21800.000000000007 ;
      RECT  2799.9999999999914 41000.00000000001 1999.9999999999916 41800.00000000001 ;
      RECT  50099.99999999999 10300.000000000005 50699.99999999999 10900.000000000005 ;
      RECT  50099.99999999999 10600.000000000007 50699.99999999999 11200.000000000007 ;
      RECT  50400.0 10300.000000000005 55199.99999999999 10900.000000000005 ;
      RECT  51199.99999999999 20100.000000000004 52000.0 21400.000000000007 ;
      RECT  51199.99999999999 1400.0000000000057 52000.0 2700.0000000000055 ;
      RECT  48000.0 2300.0000000000055 48800.0 1100.0000000000055 ;
      RECT  48000.0 19300.000000000007 48800.0 21700.00000000001 ;
      RECT  49800.0 2300.0000000000055 50400.0 19300.000000000004 ;
      RECT  48000.0 19300.000000000004 48800.0 20100.000000000004 ;
      RECT  49599.99999999999 19300.000000000004 50400.0 20100.000000000004 ;
      RECT  49599.99999999999 19300.000000000004 50400.0 20100.000000000004 ;
      RECT  48000.0 19300.000000000004 48800.0 20100.000000000004 ;
      RECT  48000.0 2300.0000000000055 48800.0 3100.000000000006 ;
      RECT  49599.99999999999 2300.0000000000055 50400.0 3100.000000000006 ;
      RECT  49599.99999999999 2300.0000000000055 50400.0 3100.0000000000055 ;
      RECT  48000.0 2300.0000000000055 48800.0 3100.0000000000055 ;
      RECT  51199.99999999999 19700.000000000007 52000.0 20500.000000000007 ;
      RECT  51199.99999999999 2300.0000000000055 52000.0 3100.000000000006 ;
      RECT  48400.0 10800.000000000005 49199.99999999999 11600.000000000007 ;
      RECT  48400.0 10800.000000000005 49199.99999999999 11600.000000000007 ;
      RECT  50099.99999999999 10900.000000000005 50699.99999999999 11500.000000000007 ;
      RECT  46800.0 21100.000000000007 53199.99999999999 21700.000000000007 ;
      RECT  46800.0 1100.0000000000057 53199.99999999999 1700.0000000000057 ;
      RECT  57599.99999999999 20100.000000000004 58400.0 21400.000000000007 ;
      RECT  57599.99999999999 1400.0000000000057 58400.0 2700.0000000000055 ;
      RECT  54400.0 3500.000000000006 55199.99999999999 1100.0000000000055 ;
      RECT  54400.0 16900.000000000007 55199.99999999999 21700.000000000007 ;
      RECT  56199.99999999999 3500.000000000006 56800.0 16900.000000000007 ;
      RECT  54400.0 16900.000000000007 55199.99999999999 17700.000000000007 ;
      RECT  56000.0 16900.000000000007 56800.0 17700.000000000007 ;
      RECT  56000.0 16900.000000000007 56800.0 17700.000000000007 ;
      RECT  54400.0 16900.000000000007 55199.99999999999 17700.000000000007 ;
      RECT  54400.0 3500.000000000006 55199.99999999999 4300.000000000006 ;
      RECT  56000.0 3500.000000000006 56800.0 4300.000000000006 ;
      RECT  56000.0 3500.000000000006 56800.0 4300.000000000006 ;
      RECT  54400.0 3500.000000000006 55199.99999999999 4300.000000000006 ;
      RECT  57599.99999999999 19700.000000000007 58400.0 20500.000000000007 ;
      RECT  57599.99999999999 2300.0000000000055 58400.0 3100.000000000006 ;
      RECT  54800.0 10200.000000000007 55599.99999999999 11000.000000000007 ;
      RECT  54800.0 10200.000000000007 55599.99999999999 11000.000000000007 ;
      RECT  56500.0 10300.000000000005 57099.99999999999 10900.000000000005 ;
      RECT  53199.99999999999 21100.000000000007 59599.99999999999 21700.000000000007 ;
      RECT  53199.99999999999 1100.0000000000057 59599.99999999999 1700.0000000000057 ;
      RECT  48400.0 10800.000000000005 49199.99999999999 11600.000000000007 ;
      RECT  56500.0 10300.000000000005 57099.99999999999 10900.000000000005 ;
      RECT  46800.0 21100.000000000007 59599.99999999999 21700.000000000007 ;
      RECT  46800.0 1100.0000000000057 59599.99999999999 1700.0000000000057 ;
      RECT  51199.99999999999 22700.000000000007 52000.0 21400.000000000007 ;
      RECT  51199.99999999999 41400.00000000001 52000.0 40100.00000000001 ;
      RECT  48000.0 40500.00000000001 48800.0 41700.0 ;
      RECT  48000.0 23500.000000000004 48800.0 21100.0 ;
      RECT  49800.0 40500.00000000001 50400.0 23500.000000000007 ;
      RECT  48000.0 23500.000000000007 48800.0 22700.000000000007 ;
      RECT  49599.99999999999 23500.000000000007 50400.0 22700.000000000007 ;
      RECT  49599.99999999999 23500.000000000007 50400.0 22700.000000000007 ;
      RECT  48000.0 23500.000000000007 48800.0 22700.000000000007 ;
      RECT  48000.0 40500.00000000001 48800.0 39700.0 ;
      RECT  49599.99999999999 40500.00000000001 50400.0 39700.0 ;
      RECT  49599.99999999999 40500.00000000001 50400.0 39700.0 ;
      RECT  48000.0 40500.00000000001 48800.0 39700.0 ;
      RECT  51199.99999999999 23100.000000000004 52000.0 22300.000000000004 ;
      RECT  51199.99999999999 40500.00000000001 52000.0 39700.0 ;
      RECT  48400.0 32000.000000000007 49199.99999999999 31200.000000000004 ;
      RECT  48400.0 32000.000000000007 49199.99999999999 31200.000000000004 ;
      RECT  50099.99999999999 31900.000000000007 50699.99999999999 31300.000000000004 ;
      RECT  46800.0 21700.000000000004 53199.99999999999 21100.000000000004 ;
      RECT  46800.0 41700.0 53199.99999999999 41100.00000000001 ;
      RECT  61800.0 36900.00000000001 62399.99999999999 36300.00000000001 ;
      RECT  61800.0 32500.000000000007 62399.99999999999 31900.000000000007 ;
      RECT  59400.0 36900.00000000001 62099.99999999999 36300.00000000001 ;
      RECT  61800.0 36600.00000000001 62399.99999999999 32200.000000000004 ;
      RECT  62099.99999999999 32500.000000000007 64800.0 31900.000000000007 ;
      RECT  54400.0 40100.00000000001 55199.99999999999 41700.0 ;
      RECT  54400.0 23500.000000000004 55199.99999999999 21100.0 ;
      RECT  57599.99999999999 23500.000000000004 58400.0 21100.0 ;
      RECT  59199.99999999999 22700.000000000007 59999.99999999999 21400.000000000007 ;
      RECT  59199.99999999999 41400.00000000001 59999.99999999999 40100.00000000001 ;
      RECT  54400.0 23500.000000000007 55199.99999999999 22700.000000000007 ;
      RECT  55999.99999999999 23500.000000000007 56800.0 22700.000000000007 ;
      RECT  55999.99999999999 23500.000000000007 56800.0 22700.000000000007 ;
      RECT  54400.0 23500.000000000007 55199.99999999999 22700.000000000007 ;
      RECT  55999.99999999999 23500.000000000007 56800.0 22700.000000000007 ;
      RECT  57599.99999999999 23500.000000000007 58400.0 22700.000000000007 ;
      RECT  57599.99999999999 23500.000000000007 58400.0 22700.000000000007 ;
      RECT  55999.99999999999 23500.000000000007 56800.0 22700.000000000007 ;
      RECT  54400.0 40100.00000000001 55199.99999999999 39300.00000000001 ;
      RECT  55999.99999999999 40100.00000000001 56800.0 39300.00000000001 ;
      RECT  55999.99999999999 40100.00000000001 56800.0 39300.00000000001 ;
      RECT  54400.0 40100.00000000001 55199.99999999999 39300.00000000001 ;
      RECT  55999.99999999999 40100.00000000001 56800.0 39300.00000000001 ;
      RECT  57599.99999999999 40100.00000000001 58400.0 39300.00000000001 ;
      RECT  57599.99999999999 40100.00000000001 58400.0 39300.00000000001 ;
      RECT  55999.99999999999 40100.00000000001 56800.0 39300.00000000001 ;
      RECT  59199.99999999999 23100.000000000004 59999.99999999999 22300.000000000004 ;
      RECT  59199.99999999999 40500.00000000001 59999.99999999999 39700.0 ;
      RECT  57599.99999999999 38400.00000000001 56800.0 37600.00000000001 ;
      RECT  55599.99999999999 37000.00000000001 54800.0 36200.0 ;
      RECT  55999.99999999999 23500.000000000004 56800.0 22700.000000000004 ;
      RECT  57599.99999999999 40100.00000000001 58400.0 39300.00000000001 ;
      RECT  59800.0 37000.00000000001 59000.0 36200.0 ;
      RECT  54800.0 37000.00000000001 55599.99999999999 36200.0 ;
      RECT  56800.0 38400.00000000001 57599.99999999999 37600.00000000001 ;
      RECT  59000.0 37000.00000000001 59800.0 36200.0 ;
      RECT  53199.99999999999 21700.000000000004 62800.0 21100.000000000004 ;
      RECT  53199.99999999999 41700.0 62800.0 41100.00000000001 ;
      RECT  67200.0 22700.000000000007 68000.0 21400.000000000007 ;
      RECT  67200.0 41400.00000000001 68000.0 40100.00000000001 ;
      RECT  64000.0 39300.00000000001 64800.0 41700.0 ;
      RECT  64000.0 25900.000000000007 64800.0 21100.000000000004 ;
      RECT  65800.0 39300.00000000001 66399.99999999999 25900.000000000007 ;
      RECT  64000.0 25900.000000000007 64800.0 25100.000000000004 ;
      RECT  65600.0 25900.000000000007 66399.99999999999 25100.000000000004 ;
      RECT  65600.0 25900.000000000007 66399.99999999999 25100.000000000004 ;
      RECT  64000.0 25900.000000000007 64800.0 25100.000000000004 ;
      RECT  64000.0 39300.00000000001 64800.0 38500.00000000001 ;
      RECT  65600.0 39300.00000000001 66399.99999999999 38500.00000000001 ;
      RECT  65600.0 39300.00000000001 66399.99999999999 38500.00000000001 ;
      RECT  64000.0 39300.00000000001 64800.0 38500.00000000001 ;
      RECT  67200.0 23100.000000000004 68000.0 22300.000000000004 ;
      RECT  67200.0 40500.00000000001 68000.0 39700.0 ;
      RECT  64400.00000000001 32600.000000000007 65199.999999999985 31800.000000000004 ;
      RECT  64400.00000000001 32600.000000000007 65199.999999999985 31800.000000000004 ;
      RECT  66100.0 32500.000000000007 66700.0 31900.000000000007 ;
      RECT  62800.0 21700.000000000004 69200.0 21100.000000000004 ;
      RECT  62800.0 41700.0 69200.0 41100.00000000001 ;
      RECT  54800.0 37000.00000000001 55599.99999999999 36200.0 ;
      RECT  56800.0 38400.00000000001 57599.99999999999 37600.00000000001 ;
      RECT  66100.0 32500.000000000007 66700.0 31900.000000000007 ;
      RECT  53199.99999999999 21700.000000000004 69200.0 21100.000000000004 ;
      RECT  53199.99999999999 41700.0 69200.0 41100.00000000001 ;
      RECT  55400.0 45900.00000000001 56000.0 46500.00000000001 ;
      RECT  55400.0 50300.00000000001 56000.0 50900.00000000001 ;
      RECT  53000.0 45900.00000000001 55699.99999999999 46500.00000000001 ;
      RECT  55400.0 46200.0 56000.0 50600.00000000001 ;
      RECT  55699.99999999999 50300.00000000001 58400.0 50900.00000000001 ;
      RECT  48000.0 42700.0 48800.0 41100.00000000001 ;
      RECT  48000.0 59300.000000000015 48800.0 61700.00000000001 ;
      RECT  51199.99999999999 59300.000000000015 52000.0 61700.00000000001 ;
      RECT  52800.0 60100.00000000001 53599.99999999999 61400.00000000001 ;
      RECT  52800.0 41400.00000000001 53599.99999999999 42700.0 ;
      RECT  48000.0 59300.00000000001 48800.0 60100.00000000001 ;
      RECT  49599.99999999999 59300.00000000001 50400.0 60100.00000000001 ;
      RECT  49599.99999999999 59300.00000000001 50400.0 60100.00000000001 ;
      RECT  48000.0 59300.00000000001 48800.0 60100.00000000001 ;
      RECT  49599.99999999999 59300.00000000001 50400.0 60100.00000000001 ;
      RECT  51199.99999999999 59300.00000000001 52000.0 60100.00000000001 ;
      RECT  51199.99999999999 59300.00000000001 52000.0 60100.00000000001 ;
      RECT  49599.99999999999 59300.00000000001 50400.0 60100.00000000001 ;
      RECT  48000.0 42700.0 48800.0 43500.00000000001 ;
      RECT  49599.99999999999 42700.0 50400.0 43500.00000000001 ;
      RECT  49599.99999999999 42700.0 50400.0 43500.00000000001 ;
      RECT  48000.0 42700.0 48800.0 43500.00000000001 ;
      RECT  49599.99999999999 42700.0 50400.0 43500.00000000001 ;
      RECT  51199.99999999999 42700.0 52000.0 43500.00000000001 ;
      RECT  51199.99999999999 42700.0 52000.0 43500.00000000001 ;
      RECT  49599.99999999999 42700.0 50400.0 43500.00000000001 ;
      RECT  52800.0 59700.0 53599.99999999999 60500.00000000001 ;
      RECT  52800.0 42300.00000000001 53599.99999999999 43100.00000000001 ;
      RECT  51199.99999999999 44400.00000000001 50400.0 45200.0 ;
      RECT  49199.99999999999 45800.00000000001 48400.0 46600.00000000001 ;
      RECT  49599.99999999999 59300.000000000015 50400.0 60100.00000000001 ;
      RECT  51199.99999999999 42700.0 52000.0 43500.00000000001 ;
      RECT  53400.0 45800.00000000001 52599.99999999999 46600.00000000001 ;
      RECT  48400.0 45800.00000000001 49199.99999999999 46600.00000000001 ;
      RECT  50400.0 44400.00000000001 51199.99999999999 45200.0 ;
      RECT  52599.99999999999 45800.00000000001 53400.0 46600.00000000001 ;
      RECT  46800.0 61100.00000000001 56400.0 61700.0 ;
      RECT  46800.0 41100.00000000001 56400.0 41700.0 ;
      RECT  60800.0 60100.00000000001 61599.99999999999 61400.00000000001 ;
      RECT  60800.0 41400.00000000001 61599.99999999999 42700.0 ;
      RECT  57599.99999999999 43500.00000000001 58400.0 41100.00000000001 ;
      RECT  57599.99999999999 56900.00000000001 58400.0 61700.0 ;
      RECT  59400.0 43500.00000000001 60000.0 56900.00000000001 ;
      RECT  57599.99999999999 56900.00000000001 58400.0 57700.0 ;
      RECT  59200.0 56900.00000000001 60000.0 57700.0 ;
      RECT  59200.0 56900.00000000001 60000.0 57700.0 ;
      RECT  57599.99999999999 56900.00000000001 58400.0 57700.0 ;
      RECT  57599.99999999999 43500.00000000001 58400.0 44300.00000000001 ;
      RECT  59200.0 43500.00000000001 60000.0 44300.00000000001 ;
      RECT  59200.0 43500.00000000001 60000.0 44300.00000000001 ;
      RECT  57599.99999999999 43500.00000000001 58400.0 44300.00000000001 ;
      RECT  60800.0 59700.0 61599.99999999999 60500.00000000001 ;
      RECT  60800.0 42300.00000000001 61599.99999999999 43100.00000000001 ;
      RECT  58000.0 50200.0 58800.0 51000.00000000001 ;
      RECT  58000.0 50200.0 58800.0 51000.00000000001 ;
      RECT  59700.0 50300.00000000001 60300.0 50900.00000000001 ;
      RECT  56400.0 61100.00000000001 62800.0 61700.0 ;
      RECT  56400.0 41100.00000000001 62800.0 41700.0 ;
      RECT  48400.0 45800.00000000001 49199.99999999999 46600.00000000001 ;
      RECT  50400.0 44400.00000000001 51199.99999999999 45200.0 ;
      RECT  59699.99999999999 50300.00000000001 60300.0 50900.00000000001 ;
      RECT  46800.0 61100.00000000001 62800.0 61700.0 ;
      RECT  46800.0 41100.00000000001 62800.0 41700.0 ;
      RECT  50400.0 72500.0 55199.99999999999 71900.0 ;
      RECT  51199.99999999999 62700.0 52000.0 61400.00000000001 ;
      RECT  51199.99999999999 81400.0 52000.0 80100.00000000001 ;
      RECT  48000.0 79300.00000000001 48800.0 81700.0 ;
      RECT  48000.0 65900.0 48800.0 61100.00000000001 ;
      RECT  49800.0 79300.00000000001 50400.0 65900.0 ;
      RECT  48000.0 65900.0 48800.0 65100.00000000001 ;
      RECT  49599.99999999999 65900.0 50400.0 65100.00000000001 ;
      RECT  49599.99999999999 65900.0 50400.0 65100.00000000001 ;
      RECT  48000.0 65900.0 48800.0 65100.00000000001 ;
      RECT  48000.0 79300.00000000001 48800.0 78500.0 ;
      RECT  49599.99999999999 79300.00000000001 50400.0 78500.0 ;
      RECT  49599.99999999999 79300.00000000001 50400.0 78500.0 ;
      RECT  48000.0 79300.00000000001 48800.0 78500.0 ;
      RECT  51199.99999999999 63100.00000000001 52000.0 62300.00000000001 ;
      RECT  51199.99999999999 80500.0 52000.0 79700.0 ;
      RECT  48400.0 72600.00000000001 49199.99999999999 71800.00000000001 ;
      RECT  48400.0 72600.00000000001 49199.99999999999 71800.00000000001 ;
      RECT  50099.99999999999 72500.0 50699.99999999999 71900.0 ;
      RECT  46800.0 61700.0 53199.99999999999 61100.00000000001 ;
      RECT  46800.0 81700.0 53199.99999999999 81100.00000000001 ;
      RECT  62400.0 62700.0 63200.0 61400.00000000001 ;
      RECT  62400.0 81400.0 63200.0 80100.00000000001 ;
      RECT  54500.0 80500.0 61500.0 81700.0 ;
      RECT  54500.0 64500.0 61500.0 61100.0 ;
      RECT  59300.0 77900.0 59900.0 67100.00000000001 ;
      RECT  54500.0 65500.0 55099.99999999999 64200.0 ;
      RECT  57699.99999999999 65500.0 58300.0 64200.0 ;
      RECT  60900.0 65500.0 61500.0 64200.0 ;
      RECT  56099.99999999999 66800.00000000001 56699.99999999999 65500.0 ;
      RECT  59300.0 66800.00000000001 59900.0 65500.0 ;
      RECT  54400.0 65900.0 55199.99999999999 65100.00000000001 ;
      RECT  57599.99999999999 65900.0 58400.0 65100.00000000001 ;
      RECT  60800.0 65900.0 61599.99999999999 65100.00000000001 ;
      RECT  56000.0 65900.0 56800.0 65100.00000000001 ;
      RECT  59199.99999999999 65900.0 60000.0 65100.00000000001 ;
      RECT  56099.99999999999 67100.00000000001 59900.0 66500.0 ;
      RECT  54500.0 64500.0 61500.0 63900.00000000001 ;
      RECT  54500.0 80200.0 55099.99999999999 78900.0 ;
      RECT  57699.99999999999 80200.0 58300.0 78900.0 ;
      RECT  60900.0 80200.0 61500.0 78900.0 ;
      RECT  56099.99999999999 78900.0 56699.99999999999 77600.00000000001 ;
      RECT  59300.0 78900.0 59900.0 77600.00000000001 ;
      RECT  54400.0 79300.00000000001 55199.99999999999 78500.0 ;
      RECT  57599.99999999999 79300.00000000001 58400.0 78500.0 ;
      RECT  60800.0 79300.00000000001 61599.99999999999 78500.0 ;
      RECT  56000.0 79300.00000000001 56800.0 78500.0 ;
      RECT  59199.99999999999 79300.00000000001 60000.0 78500.0 ;
      RECT  56099.99999999999 77900.0 59900.0 77300.00000000001 ;
      RECT  54500.0 80500.0 61500.0 79900.0 ;
      RECT  62400.0 63100.00000000001 63200.0 62300.00000000001 ;
      RECT  62400.0 80500.0 63200.0 79700.0 ;
      RECT  54800.0 72600.00000000001 55599.99999999999 71800.00000000001 ;
      RECT  54800.0 72600.00000000001 55599.99999999999 71800.00000000001 ;
      RECT  59599.99999999999 72500.0 60199.99999999999 71900.0 ;
      RECT  53199.99999999999 61700.0 64400.00000000001 61100.00000000001 ;
      RECT  53199.99999999999 81700.0 64400.00000000001 81100.00000000001 ;
      RECT  48400.0 72600.00000000001 49199.99999999999 71800.00000000001 ;
      RECT  59599.99999999999 72500.0 60199.99999999999 71900.0 ;
      RECT  46800.0 61700.0 64400.00000000001 61100.00000000001 ;
      RECT  46800.0 81700.0 64400.00000000001 81100.00000000001 ;
      RECT  50099.99999999999 90300.00000000001 50699.99999999999 90900.0 ;
      RECT  50099.99999999999 90600.00000000001 50699.99999999999 91000.0 ;
      RECT  50400.0 90300.00000000001 55199.99999999999 90900.0 ;
      RECT  51199.99999999999 100100.00000000001 52000.0 101400.0 ;
      RECT  51199.99999999999 81400.0 52000.0 82700.0 ;
      RECT  48000.0 82700.0 48800.0 81100.00000000001 ;
      RECT  48000.0 98500.0 48800.0 101700.0 ;
      RECT  49800.0 82700.0 50400.0 98500.0 ;
      RECT  48000.0 98500.0 48800.0 99300.00000000001 ;
      RECT  49599.99999999999 98500.0 50400.0 99300.00000000001 ;
      RECT  49599.99999999999 98500.0 50400.0 99300.00000000001 ;
      RECT  48000.0 98500.0 48800.0 99300.00000000001 ;
      RECT  48000.0 82700.0 48800.0 83500.0 ;
      RECT  49599.99999999999 82700.0 50400.0 83500.0 ;
      RECT  49599.99999999999 82700.0 50400.0 83500.0 ;
      RECT  48000.0 82700.0 48800.0 83500.0 ;
      RECT  51199.99999999999 99700.0 52000.0 100500.0 ;
      RECT  51199.99999999999 82300.00000000001 52000.0 83100.00000000001 ;
      RECT  48400.0 90600.00000000001 49199.99999999999 91400.0 ;
      RECT  48400.0 90600.00000000001 49199.99999999999 91400.0 ;
      RECT  50099.99999999999 90700.0 50699.99999999999 91300.00000000001 ;
      RECT  46800.0 101100.00000000001 53199.99999999999 101700.0 ;
      RECT  46800.0 81100.00000000001 53199.99999999999 81700.0 ;
      RECT  59199.99999999999 100100.00000000001 60000.0 101400.0 ;
      RECT  59199.99999999999 81400.0 60000.0 82700.0 ;
      RECT  54500.0 82300.00000000001 58300.0 81100.00000000001 ;
      RECT  54500.0 98300.00000000001 58300.0 101700.00000000001 ;
      RECT  56199.99999999999 83500.0 56800.0 96900.0 ;
      RECT  54500.0 97300.00000000001 55099.99999999999 98600.00000000001 ;
      RECT  57699.99999999999 97300.00000000001 58300.0 98600.00000000001 ;
      RECT  54400.0 96900.0 55199.99999999999 97700.0 ;
      RECT  57599.99999999999 96900.0 58400.0 97700.0 ;
      RECT  56000.0 96900.0 56800.0 97700.0 ;
      RECT  56000.0 96900.0 56800.0 97700.0 ;
      RECT  54500.0 98300.00000000001 58300.0 98900.0 ;
      RECT  54500.0 82600.00000000001 55099.99999999999 83900.0 ;
      RECT  57699.99999999999 82600.00000000001 58300.0 83900.0 ;
      RECT  54400.0 83500.0 55199.99999999999 84300.00000000001 ;
      RECT  57599.99999999999 83500.0 58400.0 84300.00000000001 ;
      RECT  56000.0 83500.0 56800.0 84300.00000000001 ;
      RECT  56000.0 83500.0 56800.0 84300.00000000001 ;
      RECT  54500.0 82300.00000000001 58300.0 82900.0 ;
      RECT  59199.99999999999 99700.0 60000.0 100500.0 ;
      RECT  59199.99999999999 82300.00000000001 60000.0 83100.00000000001 ;
      RECT  54800.0 90200.0 55599.99999999999 91000.0 ;
      RECT  54800.0 90200.0 55599.99999999999 91000.0 ;
      RECT  56500.0 90300.00000000001 57099.99999999999 90900.0 ;
      RECT  53199.99999999999 101100.00000000001 61199.99999999999 101700.0 ;
      RECT  53199.99999999999 81100.00000000001 61199.99999999999 81700.0 ;
      RECT  48400.0 90600.00000000001 49199.99999999999 91400.0 ;
      RECT  56500.0 90300.00000000001 57099.99999999999 90900.0 ;
      RECT  46800.0 101100.00000000001 61199.99999999999 101700.0 ;
      RECT  46800.0 81100.00000000001 61199.99999999999 81700.0 ;
      RECT  55400.0 116900.0 56000.0 116300.00000000001 ;
      RECT  55400.0 112500.0 56000.0 111900.0 ;
      RECT  53000.0 116900.0 55699.99999999999 116300.00000000001 ;
      RECT  55400.0 116600.00000000001 56000.0 112200.0 ;
      RECT  55699.99999999999 112500.0 58400.0 111900.0 ;
      RECT  48000.0 120100.00000000001 48800.0 121700.0 ;
      RECT  48000.0 103500.0 48800.0 101100.0 ;
      RECT  51199.99999999999 103500.0 52000.0 101100.0 ;
      RECT  52800.0 102700.0 53599.99999999999 101400.0 ;
      RECT  52800.0 121400.0 53599.99999999999 120100.00000000001 ;
      RECT  48000.0 103500.0 48800.0 102700.0 ;
      RECT  49599.99999999999 103500.0 50400.0 102700.0 ;
      RECT  49599.99999999999 103500.0 50400.0 102700.0 ;
      RECT  48000.0 103500.0 48800.0 102700.0 ;
      RECT  49599.99999999999 103500.0 50400.0 102700.0 ;
      RECT  51199.99999999999 103500.0 52000.0 102700.0 ;
      RECT  51199.99999999999 103500.0 52000.0 102700.0 ;
      RECT  49599.99999999999 103500.0 50400.0 102700.0 ;
      RECT  48000.0 120100.00000000001 48800.0 119300.00000000001 ;
      RECT  49599.99999999999 120100.00000000001 50400.0 119300.00000000001 ;
      RECT  49599.99999999999 120100.00000000001 50400.0 119300.00000000001 ;
      RECT  48000.0 120100.00000000001 48800.0 119300.00000000001 ;
      RECT  49599.99999999999 120100.00000000001 50400.0 119300.00000000001 ;
      RECT  51199.99999999999 120100.00000000001 52000.0 119300.00000000001 ;
      RECT  51199.99999999999 120100.00000000001 52000.0 119300.00000000001 ;
      RECT  49599.99999999999 120100.00000000001 50400.0 119300.00000000001 ;
      RECT  52800.0 103100.00000000001 53599.99999999999 102300.00000000001 ;
      RECT  52800.0 120500.0 53599.99999999999 119700.0 ;
      RECT  51199.99999999999 118400.0 50400.0 117600.00000000001 ;
      RECT  49199.99999999999 117000.0 48400.0 116200.0 ;
      RECT  49599.99999999999 103500.0 50400.0 102700.0 ;
      RECT  51199.99999999999 120100.00000000001 52000.0 119300.00000000001 ;
      RECT  53400.0 117000.0 52599.99999999999 116200.0 ;
      RECT  48400.0 117000.0 49199.99999999999 116200.0 ;
      RECT  50400.0 118400.0 51199.99999999999 117600.00000000001 ;
      RECT  52599.99999999999 117000.0 53400.0 116200.0 ;
      RECT  46800.0 101700.0 56400.0 101100.00000000001 ;
      RECT  46800.0 121700.0 56400.0 121100.00000000001 ;
      RECT  60800.0 102700.0 61599.99999999999 101400.0 ;
      RECT  60800.0 121400.0 61599.99999999999 120100.00000000001 ;
      RECT  57599.99999999999 119300.00000000001 58400.0 121700.0 ;
      RECT  57599.99999999999 105900.0 58400.0 101100.00000000001 ;
      RECT  59400.0 119300.00000000001 60000.0 105900.0 ;
      RECT  57599.99999999999 105900.0 58400.0 105100.00000000001 ;
      RECT  59200.0 105900.0 60000.0 105100.00000000001 ;
      RECT  59200.0 105900.0 60000.0 105100.00000000001 ;
      RECT  57599.99999999999 105900.0 58400.0 105100.00000000001 ;
      RECT  57599.99999999999 119300.00000000001 58400.0 118500.0 ;
      RECT  59200.0 119300.00000000001 60000.0 118500.0 ;
      RECT  59200.0 119300.00000000001 60000.0 118500.0 ;
      RECT  57599.99999999999 119300.00000000001 58400.0 118500.0 ;
      RECT  60800.0 103100.00000000001 61599.99999999999 102300.00000000001 ;
      RECT  60800.0 120500.0 61599.99999999999 119700.0 ;
      RECT  58000.0 112600.00000000001 58800.0 111800.00000000001 ;
      RECT  58000.0 112600.00000000001 58800.0 111800.00000000001 ;
      RECT  59700.0 112500.0 60300.0 111900.0 ;
      RECT  56400.0 101700.0 62800.0 101100.00000000001 ;
      RECT  56400.0 121700.0 62800.0 121100.00000000001 ;
      RECT  48400.0 117000.0 49199.99999999999 116200.0 ;
      RECT  50400.0 118400.0 51199.99999999999 117600.00000000001 ;
      RECT  59699.99999999999 112500.0 60300.0 111900.0 ;
      RECT  46800.0 101700.0 62800.0 101100.00000000001 ;
      RECT  46800.0 121700.0 62800.0 121100.00000000001 ;
      RECT  55400.0 125900.0 56000.0 126500.0 ;
      RECT  55400.0 130300.00000000001 56000.0 130900.0 ;
      RECT  53000.0 125900.0 55699.99999999999 126500.0 ;
      RECT  55400.0 126200.0 56000.0 130600.0 ;
      RECT  55699.99999999999 130300.00000000001 58400.0 130900.0 ;
      RECT  48000.0 122700.0 48800.0 121100.00000000001 ;
      RECT  48000.0 139300.0 48800.0 141700.00000000003 ;
      RECT  51199.99999999999 139300.0 52000.0 141700.00000000003 ;
      RECT  52800.0 140100.0 53599.99999999999 141400.0 ;
      RECT  52800.0 121400.0 53599.99999999999 122700.0 ;
      RECT  48000.0 139300.0 48800.0 140100.0 ;
      RECT  49599.99999999999 139300.0 50400.0 140100.0 ;
      RECT  49599.99999999999 139300.0 50400.0 140100.0 ;
      RECT  48000.0 139300.0 48800.0 140100.0 ;
      RECT  49599.99999999999 139300.0 50400.0 140100.0 ;
      RECT  51199.99999999999 139300.0 52000.0 140100.0 ;
      RECT  51199.99999999999 139300.0 52000.0 140100.0 ;
      RECT  49599.99999999999 139300.0 50400.0 140100.0 ;
      RECT  48000.0 122700.0 48800.0 123500.0 ;
      RECT  49599.99999999999 122700.0 50400.0 123500.0 ;
      RECT  49599.99999999999 122700.0 50400.0 123500.0 ;
      RECT  48000.0 122700.0 48800.0 123500.0 ;
      RECT  49599.99999999999 122700.0 50400.0 123500.0 ;
      RECT  51199.99999999999 122700.0 52000.0 123500.0 ;
      RECT  51199.99999999999 122700.0 52000.0 123500.0 ;
      RECT  49599.99999999999 122700.0 50400.0 123500.0 ;
      RECT  52800.0 139700.00000000003 53599.99999999999 140500.0 ;
      RECT  52800.0 122300.00000000001 53599.99999999999 123100.00000000001 ;
      RECT  51199.99999999999 124400.0 50400.0 125200.0 ;
      RECT  49199.99999999999 125800.00000000001 48400.0 126600.00000000001 ;
      RECT  49599.99999999999 139300.0 50400.0 140100.0 ;
      RECT  51199.99999999999 122700.0 52000.0 123500.0 ;
      RECT  53400.0 125800.00000000001 52599.99999999999 126600.00000000001 ;
      RECT  48400.0 125800.00000000001 49199.99999999999 126600.00000000001 ;
      RECT  50400.0 124400.0 51199.99999999999 125200.0 ;
      RECT  52599.99999999999 125800.00000000001 53400.0 126600.00000000001 ;
      RECT  46800.0 141100.0 56400.0 141700.00000000003 ;
      RECT  46800.0 121100.00000000001 56400.0 121700.0 ;
      RECT  60800.0 140100.0 61599.99999999999 141400.0 ;
      RECT  60800.0 121400.0 61599.99999999999 122700.0 ;
      RECT  57599.99999999999 123500.0 58400.0 121100.00000000001 ;
      RECT  57599.99999999999 136900.0 58400.0 141700.00000000003 ;
      RECT  59400.0 123500.0 60000.0 136900.0 ;
      RECT  57599.99999999999 136900.0 58400.0 137700.00000000003 ;
      RECT  59200.0 136900.0 60000.0 137700.00000000003 ;
      RECT  59200.0 136900.0 60000.0 137700.00000000003 ;
      RECT  57599.99999999999 136900.0 58400.0 137700.00000000003 ;
      RECT  57599.99999999999 123500.0 58400.0 124300.00000000001 ;
      RECT  59200.0 123500.0 60000.0 124300.00000000001 ;
      RECT  59200.0 123500.0 60000.0 124300.00000000001 ;
      RECT  57599.99999999999 123500.0 58400.0 124300.00000000001 ;
      RECT  60800.0 139700.00000000003 61599.99999999999 140500.0 ;
      RECT  60800.0 122300.00000000001 61599.99999999999 123100.00000000001 ;
      RECT  58000.0 130200.00000000001 58800.0 131000.0 ;
      RECT  58000.0 130200.00000000001 58800.0 131000.0 ;
      RECT  59700.0 130300.00000000001 60300.0 130900.0 ;
      RECT  56400.0 141100.0 62800.0 141700.00000000003 ;
      RECT  56400.0 121100.00000000001 62800.0 121700.0 ;
      RECT  48400.0 125800.00000000001 49199.99999999999 126600.00000000001 ;
      RECT  50400.0 124400.0 51199.99999999999 125200.0 ;
      RECT  59699.99999999999 130300.00000000001 60300.0 130900.0 ;
      RECT  46800.0 141100.0 62800.0 141700.00000000003 ;
      RECT  46800.0 121100.00000000001 62800.0 121700.0 ;
      RECT  68800.0 140100.0 69600.0 141400.0 ;
      RECT  68800.0 121400.0 69600.0 122700.0 ;
      RECT  64099.99999999999 122300.00000000001 67899.99999999999 121100.00000000001 ;
      RECT  64099.99999999999 138300.0 67899.99999999999 141700.00000000003 ;
      RECT  65800.0 123500.0 66399.99999999999 136900.0 ;
      RECT  64099.99999999999 137300.0 64699.999999999985 138600.0 ;
      RECT  67300.0 137300.0 67899.99999999999 138600.0 ;
      RECT  64000.0 136900.0 64800.0 137700.00000000003 ;
      RECT  67200.0 136900.0 68000.0 137700.00000000003 ;
      RECT  65600.0 136900.0 66399.99999999999 137700.00000000003 ;
      RECT  65600.0 136900.0 66399.99999999999 137700.00000000003 ;
      RECT  64099.99999999999 138300.0 67899.99999999999 138900.0 ;
      RECT  64099.99999999999 122600.00000000001 64699.999999999985 123900.0 ;
      RECT  67300.0 122600.00000000001 67899.99999999999 123900.0 ;
      RECT  64000.0 123500.0 64800.0 124300.00000000001 ;
      RECT  67200.0 123500.0 68000.0 124300.00000000001 ;
      RECT  65600.0 123500.0 66399.99999999999 124300.00000000001 ;
      RECT  65600.0 123500.0 66399.99999999999 124300.00000000001 ;
      RECT  64099.99999999999 122300.00000000001 67899.99999999999 122900.0 ;
      RECT  68800.0 139700.00000000003 69600.0 140500.0 ;
      RECT  68800.0 122300.00000000001 69600.0 123100.00000000001 ;
      RECT  64400.00000000001 130200.00000000001 65199.999999999985 131000.0 ;
      RECT  64400.00000000001 130200.00000000001 65199.999999999985 131000.0 ;
      RECT  66100.0 130300.00000000001 66700.0 130900.0 ;
      RECT  62800.0 141100.0 70800.0 141700.00000000003 ;
      RECT  62800.0 121100.00000000001 70800.0 121700.0 ;
      RECT  50099.99999999999 152500.0 50699.99999999999 151900.0 ;
      RECT  50099.99999999999 152200.00000000003 50699.99999999999 151800.0 ;
      RECT  50400.0 152500.0 55199.99999999999 151900.0 ;
      RECT  51199.99999999999 142700.00000000003 52000.0 141400.0 ;
      RECT  51199.99999999999 161400.0 52000.0 160100.0 ;
      RECT  48000.0 160100.0 48800.0 161700.00000000003 ;
      RECT  48000.0 144300.0 48800.0 141100.0 ;
      RECT  49800.0 160100.0 50400.0 144300.0 ;
      RECT  48000.0 144300.0 48800.0 143500.0 ;
      RECT  49599.99999999999 144300.0 50400.0 143500.0 ;
      RECT  49599.99999999999 144300.0 50400.0 143500.0 ;
      RECT  48000.0 144300.0 48800.0 143500.0 ;
      RECT  48000.0 160100.0 48800.0 159300.0 ;
      RECT  49599.99999999999 160100.0 50400.0 159300.0 ;
      RECT  49599.99999999999 160100.0 50400.0 159300.0 ;
      RECT  48000.0 160100.0 48800.0 159300.0 ;
      RECT  51199.99999999999 143100.0 52000.0 142300.0 ;
      RECT  51199.99999999999 160500.0 52000.0 159700.00000000003 ;
      RECT  48400.0 152200.00000000003 49199.99999999999 151400.0 ;
      RECT  48400.0 152200.00000000003 49199.99999999999 151400.0 ;
      RECT  50099.99999999999 152100.0 50699.99999999999 151500.0 ;
      RECT  46800.0 141700.00000000003 53199.99999999999 141100.0 ;
      RECT  46800.0 161700.00000000003 53199.99999999999 161100.0 ;
      RECT  59199.99999999999 142700.00000000003 60000.0 141400.0 ;
      RECT  59199.99999999999 161400.0 60000.0 160100.0 ;
      RECT  54500.0 160500.0 58300.0 161700.00000000003 ;
      RECT  54500.0 144500.0 58300.0 141100.0 ;
      RECT  56199.99999999999 159300.0 56800.0 145900.0 ;
      RECT  54500.0 145500.0 55099.99999999999 144200.00000000003 ;
      RECT  57699.99999999999 145500.0 58300.0 144200.00000000003 ;
      RECT  54400.0 145900.0 55199.99999999999 145100.0 ;
      RECT  57599.99999999999 145900.0 58400.0 145100.0 ;
      RECT  56000.0 145900.0 56800.0 145100.0 ;
      RECT  56000.0 145900.0 56800.0 145100.0 ;
      RECT  54500.0 144500.0 58300.0 143900.0 ;
      RECT  54500.0 160200.00000000003 55099.99999999999 158900.0 ;
      RECT  57699.99999999999 160200.00000000003 58300.0 158900.0 ;
      RECT  54400.0 159300.0 55199.99999999999 158500.0 ;
      RECT  57599.99999999999 159300.0 58400.0 158500.0 ;
      RECT  56000.0 159300.0 56800.0 158500.0 ;
      RECT  56000.0 159300.0 56800.0 158500.0 ;
      RECT  54500.0 160500.0 58300.0 159900.0 ;
      RECT  59199.99999999999 143100.0 60000.0 142300.0 ;
      RECT  59199.99999999999 160500.0 60000.0 159700.00000000003 ;
      RECT  54800.0 152600.0 55599.99999999999 151800.0 ;
      RECT  54800.0 152600.0 55599.99999999999 151800.0 ;
      RECT  56500.0 152500.0 57099.99999999999 151900.0 ;
      RECT  53199.99999999999 141700.00000000003 61199.99999999999 141100.0 ;
      RECT  53199.99999999999 161700.00000000003 61199.99999999999 161100.0 ;
      RECT  48400.0 152200.00000000003 49199.99999999999 151400.0 ;
      RECT  56500.0 152500.0 57099.99999999999 151900.0 ;
      RECT  46800.0 141700.00000000003 61199.99999999999 141100.0 ;
      RECT  46800.0 161700.00000000003 61199.99999999999 161100.0 ;
      RECT  37800.0 176500.00000000003 40199.99999999999 177300.0 ;
      RECT  37800.0 192100.00000000003 40199.99999999999 192900.0 ;
      RECT  37800.0 194900.0 40199.99999999999 195700.00000000003 ;
      RECT  37800.0 210500.00000000003 40199.99999999999 211300.0 ;
      RECT  37800.0 213300.0 40199.99999999999 214100.00000000003 ;
      RECT  37800.0 228900.0 40199.99999999999 229700.00000000003 ;
      RECT  37800.0 231700.00000000003 40199.99999999999 232500.00000000003 ;
      RECT  37800.0 247300.0 40199.99999999999 248100.0 ;
      RECT  29199.999999999993 173800.0 29799.999999999993 174400.0 ;
      RECT  29199.999999999993 173200.00000000003 29799.999999999993 173800.0 ;
      RECT  29499.999999999993 173800.0 30399.999999999993 174400.0 ;
      RECT  29199.999999999993 173500.00000000003 29799.999999999993 174100.00000000003 ;
      RECT  19199.999999999993 173200.00000000003 29499.999999999993 173800.0 ;
      RECT  18099.999999999993 170800.0 18699.999999999993 171400.0 ;
      RECT  18099.999999999993 171100.00000000003 18699.999999999993 171300.0 ;
      RECT  13199.999999999993 170800.0 18399.999999999993 171400.0 ;
      RECT  10799.99999999999 167600.00000000003 9999.99999999999 166300.0 ;
      RECT  10799.999999999993 175500.00000000003 9999.999999999993 174200.00000000003 ;
      RECT  13999.999999999993 174600.00000000003 13199.999999999993 175800.0 ;
      RECT  13999.99999999999 168400.0 13199.99999999999 166000.00000000003 ;
      RECT  12199.999999999993 174600.00000000003 11599.99999999999 168400.0 ;
      RECT  13999.99999999999 168400.0 13199.999999999993 167600.00000000003 ;
      RECT  12399.99999999999 168400.0 11599.99999999999 167600.00000000003 ;
      RECT  12399.99999999999 168400.0 11599.99999999999 167600.00000000003 ;
      RECT  13999.99999999999 168400.0 13199.999999999993 167600.00000000003 ;
      RECT  13999.999999999993 174600.00000000003 13199.999999999993 173800.0 ;
      RECT  12399.99999999999 174600.00000000003 11599.99999999999 173800.0 ;
      RECT  12399.99999999999 174600.00000000003 11599.999999999993 173800.0 ;
      RECT  13999.999999999993 174600.00000000003 13199.999999999993 173800.0 ;
      RECT  10799.99999999999 168000.00000000003 9999.99999999999 167200.00000000003 ;
      RECT  10799.999999999993 174600.00000000003 9999.999999999993 173800.0 ;
      RECT  13599.99999999999 171500.00000000003 12799.999999999993 170700.00000000003 ;
      RECT  13599.99999999999 171500.00000000003 12799.999999999993 170700.00000000003 ;
      RECT  11899.99999999999 171400.0 11299.999999999993 170800.0 ;
      RECT  15199.99999999999 166600.00000000003 8799.99999999999 166000.00000000003 ;
      RECT  15199.999999999993 175800.0 8799.999999999993 175200.00000000003 ;
      RECT  17999.999999999993 170900.0 18799.999999999993 171700.00000000003 ;
      RECT  19599.999999999993 170900.0 20399.999999999993 171700.00000000003 ;
      RECT  19599.999999999993 170900.0 20399.999999999993 171700.00000000003 ;
      RECT  17999.999999999993 170900.0 18799.999999999993 171700.00000000003 ;
      RECT  6799.999999999992 183400.0 7599.999999999992 184700.00000000003 ;
      RECT  6799.999999999992 175500.00000000003 7599.999999999992 176800.0 ;
      RECT  3599.999999999992 176400.0 4399.999999999992 175200.00000000003 ;
      RECT  3599.999999999992 182600.00000000003 4399.999999999992 185000.00000000003 ;
      RECT  5399.999999999992 176400.0 5999.999999999991 182600.00000000003 ;
      RECT  3599.999999999992 182600.00000000003 4399.999999999992 183400.0 ;
      RECT  5199.999999999992 182600.00000000003 5999.999999999992 183400.0 ;
      RECT  5199.999999999992 182600.00000000003 5999.999999999991 183400.0 ;
      RECT  3599.999999999992 182600.00000000003 4399.999999999992 183400.0 ;
      RECT  3599.999999999992 176400.0 4399.999999999992 177200.00000000003 ;
      RECT  5199.999999999992 176400.0 5999.999999999992 177200.00000000003 ;
      RECT  5199.999999999992 176400.0 5999.999999999991 177200.00000000003 ;
      RECT  3599.999999999992 176400.0 4399.999999999992 177200.00000000003 ;
      RECT  6799.999999999992 183000.00000000003 7599.999999999992 183800.0 ;
      RECT  6799.999999999992 176400.0 7599.999999999992 177200.00000000003 ;
      RECT  3999.9999999999914 179500.00000000003 4799.999999999992 180300.0 ;
      RECT  3999.9999999999914 179500.00000000003 4799.999999999992 180300.0 ;
      RECT  5699.999999999992 179600.00000000003 6299.999999999992 180200.00000000003 ;
      RECT  2399.9999999999914 184400.0 8799.999999999993 185000.00000000003 ;
      RECT  2399.9999999999914 175200.00000000003 8799.999999999993 175800.0 ;
      RECT  13199.999999999993 183400.0 13999.999999999993 184700.00000000003 ;
      RECT  13199.999999999993 175500.00000000003 13999.999999999993 176800.0 ;
      RECT  9999.999999999993 176400.0 10799.999999999993 175200.00000000003 ;
      RECT  9999.999999999993 182600.00000000003 10799.999999999993 185000.00000000003 ;
      RECT  11799.999999999993 176400.0 12399.99999999999 182600.00000000003 ;
      RECT  9999.999999999993 182600.00000000003 10799.999999999993 183400.0 ;
      RECT  11599.999999999993 182600.00000000003 12399.99999999999 183400.0 ;
      RECT  11599.999999999993 182600.00000000003 12399.99999999999 183400.0 ;
      RECT  9999.999999999993 182600.00000000003 10799.999999999993 183400.0 ;
      RECT  9999.999999999993 176400.0 10799.999999999993 177200.00000000003 ;
      RECT  11599.999999999993 176400.0 12399.99999999999 177200.00000000003 ;
      RECT  11599.999999999993 176400.0 12399.99999999999 177200.00000000003 ;
      RECT  9999.999999999993 176400.0 10799.999999999993 177200.00000000003 ;
      RECT  13199.999999999993 183000.00000000003 13999.999999999993 183800.0 ;
      RECT  13199.999999999993 176400.0 13999.999999999993 177200.00000000003 ;
      RECT  10399.99999999999 179500.00000000003 11199.999999999993 180300.0 ;
      RECT  10399.99999999999 179500.00000000003 11199.999999999993 180300.0 ;
      RECT  12099.999999999993 179600.00000000003 12699.999999999993 180200.00000000003 ;
      RECT  8799.999999999993 184400.0 15199.999999999993 185000.00000000003 ;
      RECT  8799.999999999993 175200.00000000003 15199.999999999993 175800.0 ;
      RECT  19599.999999999993 183400.0 20399.999999999993 184700.00000000003 ;
      RECT  19599.999999999993 175500.00000000003 20399.999999999993 176800.0 ;
      RECT  16399.999999999993 176400.0 17199.999999999993 175200.00000000003 ;
      RECT  16399.999999999993 182600.00000000003 17199.999999999993 185000.00000000003 ;
      RECT  18199.999999999993 176400.0 18799.999999999993 182600.00000000003 ;
      RECT  16399.999999999993 182600.00000000003 17199.999999999993 183400.0 ;
      RECT  17999.999999999993 182600.00000000003 18799.999999999993 183400.0 ;
      RECT  17999.999999999993 182600.00000000003 18799.999999999993 183400.0 ;
      RECT  16399.999999999993 182600.00000000003 17199.999999999993 183400.0 ;
      RECT  16399.999999999993 176400.0 17199.999999999993 177200.00000000003 ;
      RECT  17999.999999999993 176400.0 18799.999999999993 177200.00000000003 ;
      RECT  17999.999999999993 176400.0 18799.999999999993 177200.00000000003 ;
      RECT  16399.999999999993 176400.0 17199.999999999993 177200.00000000003 ;
      RECT  19599.999999999993 183000.00000000003 20399.999999999993 183800.0 ;
      RECT  19599.999999999993 176400.0 20399.999999999993 177200.00000000003 ;
      RECT  16799.99999999999 179500.00000000003 17599.999999999993 180300.0 ;
      RECT  16799.99999999999 179500.00000000003 17599.999999999993 180300.0 ;
      RECT  18499.999999999993 179600.00000000003 19099.999999999993 180200.00000000003 ;
      RECT  15199.999999999993 184400.0 21599.999999999993 185000.00000000003 ;
      RECT  15199.999999999993 175200.00000000003 21599.999999999993 175800.0 ;
      RECT  25999.999999999993 183400.0 26799.999999999993 184700.00000000003 ;
      RECT  25999.999999999993 175500.00000000003 26799.999999999993 176800.0 ;
      RECT  22799.999999999993 176400.0 23599.999999999993 175200.00000000003 ;
      RECT  22799.999999999993 182600.00000000003 23599.999999999993 185000.00000000003 ;
      RECT  24599.999999999993 176400.0 25199.999999999996 182600.00000000003 ;
      RECT  22799.999999999993 182600.00000000003 23599.999999999993 183400.0 ;
      RECT  24399.999999999996 182600.00000000003 25199.999999999996 183400.0 ;
      RECT  24399.999999999996 182600.00000000003 25199.999999999996 183400.0 ;
      RECT  22799.999999999993 182600.00000000003 23599.999999999993 183400.0 ;
      RECT  22799.999999999993 176400.0 23599.999999999993 177200.00000000003 ;
      RECT  24399.999999999996 176400.0 25199.999999999996 177200.00000000003 ;
      RECT  24399.999999999996 176400.0 25199.999999999996 177200.00000000003 ;
      RECT  22799.999999999993 176400.0 23599.999999999993 177200.00000000003 ;
      RECT  25999.999999999993 183000.00000000003 26799.999999999993 183800.0 ;
      RECT  25999.999999999993 176400.0 26799.999999999993 177200.00000000003 ;
      RECT  23199.999999999996 179500.00000000003 23999.999999999993 180300.0 ;
      RECT  23199.999999999996 179500.00000000003 23999.999999999993 180300.0 ;
      RECT  24899.999999999996 179600.00000000003 25499.999999999993 180200.00000000003 ;
      RECT  21599.999999999993 184400.0 27999.999999999993 185000.00000000003 ;
      RECT  21599.999999999993 175200.00000000003 27999.999999999993 175800.0 ;
      RECT  6799.999999999992 186000.00000000003 7599.999999999992 184700.00000000003 ;
      RECT  6799.999999999992 193900.0 7599.999999999992 192600.00000000003 ;
      RECT  3599.999999999992 193000.00000000003 4399.999999999992 194200.00000000003 ;
      RECT  3599.999999999992 186800.0 4399.999999999992 184400.0 ;
      RECT  5399.999999999992 193000.00000000003 5999.999999999991 186800.0 ;
      RECT  3599.999999999992 186800.0 4399.999999999992 186000.00000000003 ;
      RECT  5199.999999999992 186800.0 5999.999999999992 186000.00000000003 ;
      RECT  5199.999999999992 186800.0 5999.999999999991 186000.00000000003 ;
      RECT  3599.999999999992 186800.0 4399.999999999992 186000.00000000003 ;
      RECT  3599.999999999992 193000.00000000003 4399.999999999992 192200.00000000003 ;
      RECT  5199.999999999992 193000.00000000003 5999.999999999992 192200.00000000003 ;
      RECT  5199.999999999992 193000.00000000003 5999.999999999991 192200.00000000003 ;
      RECT  3599.999999999992 193000.00000000003 4399.999999999992 192200.00000000003 ;
      RECT  6799.999999999992 186400.0 7599.999999999992 185600.00000000003 ;
      RECT  6799.999999999992 193000.00000000003 7599.999999999992 192200.00000000003 ;
      RECT  3999.9999999999914 189900.0 4799.999999999992 189100.00000000003 ;
      RECT  3999.9999999999914 189900.0 4799.999999999992 189100.00000000003 ;
      RECT  5699.999999999992 189800.0 6299.999999999992 189200.00000000003 ;
      RECT  2399.9999999999914 185000.00000000003 8799.999999999993 184400.0 ;
      RECT  2399.9999999999914 194200.00000000003 8799.999999999993 193600.00000000003 ;
      RECT  13199.999999999993 186000.00000000003 13999.999999999993 184700.00000000003 ;
      RECT  13199.999999999993 193900.0 13999.999999999993 192600.00000000003 ;
      RECT  9999.999999999993 193000.00000000003 10799.999999999993 194200.00000000003 ;
      RECT  9999.999999999993 186800.0 10799.999999999993 184400.0 ;
      RECT  11799.999999999993 193000.00000000003 12399.99999999999 186800.0 ;
      RECT  9999.999999999993 186800.0 10799.999999999993 186000.00000000003 ;
      RECT  11599.999999999993 186800.0 12399.99999999999 186000.00000000003 ;
      RECT  11599.999999999993 186800.0 12399.99999999999 186000.00000000003 ;
      RECT  9999.999999999993 186800.0 10799.999999999993 186000.00000000003 ;
      RECT  9999.999999999993 193000.00000000003 10799.999999999993 192200.00000000003 ;
      RECT  11599.999999999993 193000.00000000003 12399.99999999999 192200.00000000003 ;
      RECT  11599.999999999993 193000.00000000003 12399.99999999999 192200.00000000003 ;
      RECT  9999.999999999993 193000.00000000003 10799.999999999993 192200.00000000003 ;
      RECT  13199.999999999993 186400.0 13999.999999999993 185600.00000000003 ;
      RECT  13199.999999999993 193000.00000000003 13999.999999999993 192200.00000000003 ;
      RECT  10399.99999999999 189900.0 11199.999999999993 189100.00000000003 ;
      RECT  10399.99999999999 189900.0 11199.999999999993 189100.00000000003 ;
      RECT  12099.999999999993 189800.0 12699.999999999993 189200.00000000003 ;
      RECT  8799.999999999993 185000.00000000003 15199.999999999993 184400.0 ;
      RECT  8799.999999999993 194200.00000000003 15199.999999999993 193600.00000000003 ;
      RECT  19599.999999999993 186000.00000000003 20399.999999999993 184700.00000000003 ;
      RECT  19599.999999999993 193900.0 20399.999999999993 192600.00000000003 ;
      RECT  16399.999999999993 193000.00000000003 17199.999999999993 194200.00000000003 ;
      RECT  16399.999999999993 186800.0 17199.999999999993 184400.0 ;
      RECT  18199.999999999993 193000.00000000003 18799.999999999993 186800.0 ;
      RECT  16399.999999999993 186800.0 17199.999999999993 186000.00000000003 ;
      RECT  17999.999999999993 186800.0 18799.999999999993 186000.00000000003 ;
      RECT  17999.999999999993 186800.0 18799.999999999993 186000.00000000003 ;
      RECT  16399.999999999993 186800.0 17199.999999999993 186000.00000000003 ;
      RECT  16399.999999999993 193000.00000000003 17199.999999999993 192200.00000000003 ;
      RECT  17999.999999999993 193000.00000000003 18799.999999999993 192200.00000000003 ;
      RECT  17999.999999999993 193000.00000000003 18799.999999999993 192200.00000000003 ;
      RECT  16399.999999999993 193000.00000000003 17199.999999999993 192200.00000000003 ;
      RECT  19599.999999999993 186400.0 20399.999999999993 185600.00000000003 ;
      RECT  19599.999999999993 193000.00000000003 20399.999999999993 192200.00000000003 ;
      RECT  16799.99999999999 189900.0 17599.999999999993 189100.00000000003 ;
      RECT  16799.99999999999 189900.0 17599.999999999993 189100.00000000003 ;
      RECT  18499.999999999993 189800.0 19099.999999999993 189200.00000000003 ;
      RECT  15199.999999999993 185000.00000000003 21599.999999999993 184400.0 ;
      RECT  15199.999999999993 194200.00000000003 21599.999999999993 193600.00000000003 ;
      RECT  25999.999999999993 186000.00000000003 26799.999999999993 184700.00000000003 ;
      RECT  25999.999999999993 193900.0 26799.999999999993 192600.00000000003 ;
      RECT  22799.999999999993 193000.00000000003 23599.999999999993 194200.00000000003 ;
      RECT  22799.999999999993 186800.0 23599.999999999993 184400.0 ;
      RECT  24599.999999999993 193000.00000000003 25199.999999999996 186800.0 ;
      RECT  22799.999999999993 186800.0 23599.999999999993 186000.00000000003 ;
      RECT  24399.999999999996 186800.0 25199.999999999996 186000.00000000003 ;
      RECT  24399.999999999996 186800.0 25199.999999999996 186000.00000000003 ;
      RECT  22799.999999999993 186800.0 23599.999999999993 186000.00000000003 ;
      RECT  22799.999999999993 193000.00000000003 23599.999999999993 192200.00000000003 ;
      RECT  24399.999999999996 193000.00000000003 25199.999999999996 192200.00000000003 ;
      RECT  24399.999999999996 193000.00000000003 25199.999999999996 192200.00000000003 ;
      RECT  22799.999999999993 193000.00000000003 23599.999999999993 192200.00000000003 ;
      RECT  25999.999999999993 186400.0 26799.999999999993 185600.00000000003 ;
      RECT  25999.999999999993 193000.00000000003 26799.999999999993 192200.00000000003 ;
      RECT  23199.999999999996 189900.0 23999.999999999993 189100.00000000003 ;
      RECT  23199.999999999996 189900.0 23999.999999999993 189100.00000000003 ;
      RECT  24899.999999999996 189800.0 25499.999999999993 189200.00000000003 ;
      RECT  21599.999999999993 185000.00000000003 27999.999999999993 184400.0 ;
      RECT  21599.999999999993 194200.00000000003 27999.999999999993 193600.00000000003 ;
      RECT  6799.999999999992 201800.00000000003 7599.999999999992 203100.00000000003 ;
      RECT  6799.999999999992 193900.0 7599.999999999992 195200.00000000003 ;
      RECT  3599.999999999992 194800.0 4399.999999999992 193600.00000000003 ;
      RECT  3599.999999999992 201000.00000000003 4399.999999999992 203400.0 ;
      RECT  5399.999999999992 194800.0 5999.999999999991 201000.00000000003 ;
      RECT  3599.999999999992 201000.00000000003 4399.999999999992 201800.00000000003 ;
      RECT  5199.999999999992 201000.00000000003 5999.999999999992 201800.00000000003 ;
      RECT  5199.999999999992 201000.00000000003 5999.999999999991 201800.00000000003 ;
      RECT  3599.999999999992 201000.00000000003 4399.999999999992 201800.00000000003 ;
      RECT  3599.999999999992 194800.0 4399.999999999992 195600.00000000003 ;
      RECT  5199.999999999992 194800.0 5999.999999999992 195600.00000000003 ;
      RECT  5199.999999999992 194800.0 5999.999999999991 195600.00000000003 ;
      RECT  3599.999999999992 194800.0 4399.999999999992 195600.00000000003 ;
      RECT  6799.999999999992 201400.0 7599.999999999992 202200.00000000003 ;
      RECT  6799.999999999992 194800.0 7599.999999999992 195600.00000000003 ;
      RECT  3999.9999999999914 197900.0 4799.999999999992 198700.00000000003 ;
      RECT  3999.9999999999914 197900.0 4799.999999999992 198700.00000000003 ;
      RECT  5699.999999999992 198000.00000000003 6299.999999999992 198600.00000000003 ;
      RECT  2399.9999999999914 202800.00000000003 8799.999999999993 203400.0 ;
      RECT  2399.9999999999914 193600.00000000003 8799.999999999993 194200.00000000003 ;
      RECT  13199.999999999993 201800.00000000003 13999.999999999993 203100.00000000003 ;
      RECT  13199.999999999993 193900.0 13999.999999999993 195200.00000000003 ;
      RECT  9999.999999999993 194800.0 10799.999999999993 193600.00000000003 ;
      RECT  9999.999999999993 201000.00000000003 10799.999999999993 203400.0 ;
      RECT  11799.999999999993 194800.0 12399.99999999999 201000.00000000003 ;
      RECT  9999.999999999993 201000.00000000003 10799.999999999993 201800.00000000003 ;
      RECT  11599.999999999993 201000.00000000003 12399.99999999999 201800.00000000003 ;
      RECT  11599.999999999993 201000.00000000003 12399.99999999999 201800.00000000003 ;
      RECT  9999.999999999993 201000.00000000003 10799.999999999993 201800.00000000003 ;
      RECT  9999.999999999993 194800.0 10799.999999999993 195600.00000000003 ;
      RECT  11599.999999999993 194800.0 12399.99999999999 195600.00000000003 ;
      RECT  11599.999999999993 194800.0 12399.99999999999 195600.00000000003 ;
      RECT  9999.999999999993 194800.0 10799.999999999993 195600.00000000003 ;
      RECT  13199.999999999993 201400.0 13999.999999999993 202200.00000000003 ;
      RECT  13199.999999999993 194800.0 13999.999999999993 195600.00000000003 ;
      RECT  10399.99999999999 197900.0 11199.999999999993 198700.00000000003 ;
      RECT  10399.99999999999 197900.0 11199.999999999993 198700.00000000003 ;
      RECT  12099.999999999993 198000.00000000003 12699.999999999993 198600.00000000003 ;
      RECT  8799.999999999993 202800.00000000003 15199.999999999993 203400.0 ;
      RECT  8799.999999999993 193600.00000000003 15199.999999999993 194200.00000000003 ;
      RECT  19599.999999999993 201800.00000000003 20399.999999999993 203100.00000000003 ;
      RECT  19599.999999999993 193900.0 20399.999999999993 195200.00000000003 ;
      RECT  16399.999999999993 194800.0 17199.999999999993 193600.00000000003 ;
      RECT  16399.999999999993 201000.00000000003 17199.999999999993 203400.0 ;
      RECT  18199.999999999993 194800.0 18799.999999999993 201000.00000000003 ;
      RECT  16399.999999999993 201000.00000000003 17199.999999999993 201800.00000000003 ;
      RECT  17999.999999999993 201000.00000000003 18799.999999999993 201800.00000000003 ;
      RECT  17999.999999999993 201000.00000000003 18799.999999999993 201800.00000000003 ;
      RECT  16399.999999999993 201000.00000000003 17199.999999999993 201800.00000000003 ;
      RECT  16399.999999999993 194800.0 17199.999999999993 195600.00000000003 ;
      RECT  17999.999999999993 194800.0 18799.999999999993 195600.00000000003 ;
      RECT  17999.999999999993 194800.0 18799.999999999993 195600.00000000003 ;
      RECT  16399.999999999993 194800.0 17199.999999999993 195600.00000000003 ;
      RECT  19599.999999999993 201400.0 20399.999999999993 202200.00000000003 ;
      RECT  19599.999999999993 194800.0 20399.999999999993 195600.00000000003 ;
      RECT  16799.99999999999 197900.0 17599.999999999993 198700.00000000003 ;
      RECT  16799.99999999999 197900.0 17599.999999999993 198700.00000000003 ;
      RECT  18499.999999999993 198000.00000000003 19099.999999999993 198600.00000000003 ;
      RECT  15199.999999999993 202800.00000000003 21599.999999999993 203400.0 ;
      RECT  15199.999999999993 193600.00000000003 21599.999999999993 194200.00000000003 ;
      RECT  25999.999999999993 201800.00000000003 26799.999999999993 203100.00000000003 ;
      RECT  25999.999999999993 193900.0 26799.999999999993 195200.00000000003 ;
      RECT  22799.999999999993 194800.0 23599.999999999993 193600.00000000003 ;
      RECT  22799.999999999993 201000.00000000003 23599.999999999993 203400.0 ;
      RECT  24599.999999999993 194800.0 25199.999999999996 201000.00000000003 ;
      RECT  22799.999999999993 201000.00000000003 23599.999999999993 201800.00000000003 ;
      RECT  24399.999999999996 201000.00000000003 25199.999999999996 201800.00000000003 ;
      RECT  24399.999999999996 201000.00000000003 25199.999999999996 201800.00000000003 ;
      RECT  22799.999999999993 201000.00000000003 23599.999999999993 201800.00000000003 ;
      RECT  22799.999999999993 194800.0 23599.999999999993 195600.00000000003 ;
      RECT  24399.999999999996 194800.0 25199.999999999996 195600.00000000003 ;
      RECT  24399.999999999996 194800.0 25199.999999999996 195600.00000000003 ;
      RECT  22799.999999999993 194800.0 23599.999999999993 195600.00000000003 ;
      RECT  25999.999999999993 201400.0 26799.999999999993 202200.00000000003 ;
      RECT  25999.999999999993 194800.0 26799.999999999993 195600.00000000003 ;
      RECT  23199.999999999996 197900.0 23999.999999999993 198700.00000000003 ;
      RECT  23199.999999999996 197900.0 23999.999999999993 198700.00000000003 ;
      RECT  24899.999999999996 198000.00000000003 25499.999999999993 198600.00000000003 ;
      RECT  21599.999999999993 202800.00000000003 27999.999999999993 203400.0 ;
      RECT  21599.999999999993 193600.00000000003 27999.999999999993 194200.00000000003 ;
      RECT  6799.999999999992 204400.0 7599.999999999992 203100.00000000003 ;
      RECT  6799.999999999992 212300.00000000003 7599.999999999992 211000.00000000003 ;
      RECT  3599.999999999992 211400.0 4399.999999999992 212600.00000000003 ;
      RECT  3599.999999999992 205200.00000000003 4399.999999999992 202800.00000000003 ;
      RECT  5399.999999999992 211400.0 5999.999999999991 205200.00000000003 ;
      RECT  3599.999999999992 205200.00000000003 4399.999999999992 204400.0 ;
      RECT  5199.999999999992 205200.00000000003 5999.999999999992 204400.0 ;
      RECT  5199.999999999992 205200.00000000003 5999.999999999991 204400.0 ;
      RECT  3599.999999999992 205200.00000000003 4399.999999999992 204400.0 ;
      RECT  3599.999999999992 211400.0 4399.999999999992 210600.00000000003 ;
      RECT  5199.999999999992 211400.0 5999.999999999992 210600.00000000003 ;
      RECT  5199.999999999992 211400.0 5999.999999999991 210600.00000000003 ;
      RECT  3599.999999999992 211400.0 4399.999999999992 210600.00000000003 ;
      RECT  6799.999999999992 204800.00000000003 7599.999999999992 204000.00000000003 ;
      RECT  6799.999999999992 211400.0 7599.999999999992 210600.00000000003 ;
      RECT  3999.9999999999914 208300.00000000003 4799.999999999992 207500.00000000003 ;
      RECT  3999.9999999999914 208300.00000000003 4799.999999999992 207500.00000000003 ;
      RECT  5699.999999999992 208200.00000000003 6299.999999999992 207600.00000000003 ;
      RECT  2399.9999999999914 203400.0 8799.999999999993 202800.00000000003 ;
      RECT  2399.9999999999914 212600.00000000003 8799.999999999993 212000.00000000003 ;
      RECT  13199.999999999993 204400.0 13999.999999999993 203100.00000000003 ;
      RECT  13199.999999999993 212300.00000000003 13999.999999999993 211000.00000000003 ;
      RECT  9999.999999999993 211400.0 10799.999999999993 212600.00000000003 ;
      RECT  9999.999999999993 205200.00000000003 10799.999999999993 202800.00000000003 ;
      RECT  11799.999999999993 211400.0 12399.99999999999 205200.00000000003 ;
      RECT  9999.999999999993 205200.00000000003 10799.999999999993 204400.0 ;
      RECT  11599.999999999993 205200.00000000003 12399.99999999999 204400.0 ;
      RECT  11599.999999999993 205200.00000000003 12399.99999999999 204400.0 ;
      RECT  9999.999999999993 205200.00000000003 10799.999999999993 204400.0 ;
      RECT  9999.999999999993 211400.0 10799.999999999993 210600.00000000003 ;
      RECT  11599.999999999993 211400.0 12399.99999999999 210600.00000000003 ;
      RECT  11599.999999999993 211400.0 12399.99999999999 210600.00000000003 ;
      RECT  9999.999999999993 211400.0 10799.999999999993 210600.00000000003 ;
      RECT  13199.999999999993 204800.00000000003 13999.999999999993 204000.00000000003 ;
      RECT  13199.999999999993 211400.0 13999.999999999993 210600.00000000003 ;
      RECT  10399.99999999999 208300.00000000003 11199.999999999993 207500.00000000003 ;
      RECT  10399.99999999999 208300.00000000003 11199.999999999993 207500.00000000003 ;
      RECT  12099.999999999993 208200.00000000003 12699.999999999993 207600.00000000003 ;
      RECT  8799.999999999993 203400.0 15199.999999999993 202800.00000000003 ;
      RECT  8799.999999999993 212600.00000000003 15199.999999999993 212000.00000000003 ;
      RECT  19599.999999999993 204400.0 20399.999999999993 203100.00000000003 ;
      RECT  19599.999999999993 212300.00000000003 20399.999999999993 211000.00000000003 ;
      RECT  16399.999999999993 211400.0 17199.999999999993 212600.00000000003 ;
      RECT  16399.999999999993 205200.00000000003 17199.999999999993 202800.00000000003 ;
      RECT  18199.999999999993 211400.0 18799.999999999993 205200.00000000003 ;
      RECT  16399.999999999993 205200.00000000003 17199.999999999993 204400.0 ;
      RECT  17999.999999999993 205200.00000000003 18799.999999999993 204400.0 ;
      RECT  17999.999999999993 205200.00000000003 18799.999999999993 204400.0 ;
      RECT  16399.999999999993 205200.00000000003 17199.999999999993 204400.0 ;
      RECT  16399.999999999993 211400.0 17199.999999999993 210600.00000000003 ;
      RECT  17999.999999999993 211400.0 18799.999999999993 210600.00000000003 ;
      RECT  17999.999999999993 211400.0 18799.999999999993 210600.00000000003 ;
      RECT  16399.999999999993 211400.0 17199.999999999993 210600.00000000003 ;
      RECT  19599.999999999993 204800.00000000003 20399.999999999993 204000.00000000003 ;
      RECT  19599.999999999993 211400.0 20399.999999999993 210600.00000000003 ;
      RECT  16799.99999999999 208300.00000000003 17599.999999999993 207500.00000000003 ;
      RECT  16799.99999999999 208300.00000000003 17599.999999999993 207500.00000000003 ;
      RECT  18499.999999999993 208200.00000000003 19099.999999999993 207600.00000000003 ;
      RECT  15199.999999999993 203400.0 21599.999999999993 202800.00000000003 ;
      RECT  15199.999999999993 212600.00000000003 21599.999999999993 212000.00000000003 ;
      RECT  25999.999999999993 204400.0 26799.999999999993 203100.00000000003 ;
      RECT  25999.999999999993 212300.00000000003 26799.999999999993 211000.00000000003 ;
      RECT  22799.999999999993 211400.0 23599.999999999993 212600.00000000003 ;
      RECT  22799.999999999993 205200.00000000003 23599.999999999993 202800.00000000003 ;
      RECT  24599.999999999993 211400.0 25199.999999999996 205200.00000000003 ;
      RECT  22799.999999999993 205200.00000000003 23599.999999999993 204400.0 ;
      RECT  24399.999999999996 205200.00000000003 25199.999999999996 204400.0 ;
      RECT  24399.999999999996 205200.00000000003 25199.999999999996 204400.0 ;
      RECT  22799.999999999993 205200.00000000003 23599.999999999993 204400.0 ;
      RECT  22799.999999999993 211400.0 23599.999999999993 210600.00000000003 ;
      RECT  24399.999999999996 211400.0 25199.999999999996 210600.00000000003 ;
      RECT  24399.999999999996 211400.0 25199.999999999996 210600.00000000003 ;
      RECT  22799.999999999993 211400.0 23599.999999999993 210600.00000000003 ;
      RECT  25999.999999999993 204800.00000000003 26799.999999999993 204000.00000000003 ;
      RECT  25999.999999999993 211400.0 26799.999999999993 210600.00000000003 ;
      RECT  23199.999999999996 208300.00000000003 23999.999999999993 207500.00000000003 ;
      RECT  23199.999999999996 208300.00000000003 23999.999999999993 207500.00000000003 ;
      RECT  24899.999999999996 208200.00000000003 25499.999999999993 207600.00000000003 ;
      RECT  21599.999999999993 203400.0 27999.999999999993 202800.00000000003 ;
      RECT  21599.999999999993 212600.00000000003 27999.999999999993 212000.00000000003 ;
      RECT  10399.99999999999 179500.00000000003 11199.999999999993 180300.0 ;
      RECT  16799.99999999999 179500.00000000003 17599.999999999993 180300.0 ;
      RECT  23199.999999999993 179500.00000000003 23999.999999999993 180300.0 ;
      RECT  3999.9999999999914 179500.00000000003 4799.999999999992 180300.0 ;
      RECT  5599.999999999992 179500.00000000003 6399.999999999992 180300.0 ;
      RECT  10399.99999999999 189100.00000000003 11199.999999999993 189900.0 ;
      RECT  16799.99999999999 189100.00000000003 17599.999999999993 189900.0 ;
      RECT  23199.999999999993 189100.00000000003 23999.999999999993 189900.0 ;
      RECT  3999.9999999999914 189100.00000000003 4799.999999999992 189900.0 ;
      RECT  5599.999999999992 189100.00000000003 6399.999999999992 189900.0 ;
      RECT  10399.99999999999 197900.0 11199.999999999993 198700.00000000003 ;
      RECT  16799.99999999999 197900.0 17599.999999999993 198700.00000000003 ;
      RECT  23199.999999999993 197900.0 23999.999999999993 198700.00000000003 ;
      RECT  3999.9999999999914 197900.0 4799.999999999992 198700.00000000003 ;
      RECT  5599.999999999992 197900.0 6399.999999999992 198700.00000000003 ;
      RECT  10399.99999999999 207500.00000000003 11199.999999999993 208300.0 ;
      RECT  16799.99999999999 207500.00000000003 17599.999999999993 208300.0 ;
      RECT  23199.999999999993 207500.00000000003 23999.999999999993 208300.0 ;
      RECT  3999.9999999999914 207500.00000000003 4799.999999999992 208300.0 ;
      RECT  5599.999999999992 207500.00000000003 6399.999999999992 208300.0 ;
      RECT  15599.999999999993 184300.0 14799.999999999993 185100.00000000003 ;
      RECT  15599.999999999993 175100.00000000003 14799.999999999993 175900.0 ;
      RECT  21999.999999999993 184300.0 21199.999999999993 185100.00000000003 ;
      RECT  21999.999999999993 175100.00000000003 21199.999999999993 175900.0 ;
      RECT  15599.999999999993 202700.00000000003 14799.999999999993 203500.00000000003 ;
      RECT  15599.999999999993 193500.00000000003 14799.999999999993 194300.0 ;
      RECT  21999.999999999993 202700.00000000003 21199.999999999993 203500.00000000003 ;
      RECT  21999.999999999993 193500.00000000003 21199.999999999993 194300.0 ;
      RECT  15599.999999999993 211900.0 14799.999999999993 212700.00000000003 ;
      RECT  21999.999999999993 211900.0 21199.999999999993 212700.00000000003 ;
      RECT  3999.9999999999914 179500.00000000003 4799.999999999992 180300.0 ;
      RECT  23199.999999999993 207500.00000000003 23999.999999999993 208300.0 ;
      RECT  30799.999999999993 175500.00000000003 37599.99999999999 166300.0 ;
      RECT  30799.999999999993 175500.00000000003 37599.99999999999 184700.00000000003 ;
      RECT  30799.999999999993 193900.0 37599.99999999999 184700.00000000003 ;
      RECT  30799.999999999993 193900.0 37599.99999999999 203100.00000000003 ;
      RECT  30799.999999999993 212300.00000000003 37599.99999999999 203100.00000000003 ;
      RECT  30799.999999999993 212300.00000000003 37599.99999999999 221500.00000000003 ;
      RECT  30799.999999999993 230700.00000000003 37599.99999999999 221500.00000000003 ;
      RECT  30799.999999999993 230700.00000000003 37599.99999999999 239900.0 ;
      RECT  30799.999999999993 249100.00000000003 37599.99999999999 239900.0 ;
      RECT  30399.999999999996 176500.00000000003 37800.0 177300.0 ;
      RECT  30399.999999999996 192100.00000000003 37800.0 192900.0 ;
      RECT  30399.999999999996 194900.0 37800.0 195700.00000000003 ;
      RECT  30399.999999999996 210500.00000000003 37800.0 211300.00000000003 ;
      RECT  30399.999999999996 213300.00000000003 37800.0 214100.00000000003 ;
      RECT  30399.999999999996 228900.0 37800.0 229700.00000000003 ;
      RECT  30399.999999999996 231700.00000000003 37800.0 232500.00000000003 ;
      RECT  30399.999999999996 247300.0 37800.0 248100.00000000003 ;
      RECT  9199.999999999993 165900.0 8399.99999999999 166700.00000000003 ;
      RECT  31199.999999999993 170500.00000000003 30399.999999999993 171300.0 ;
      RECT  37999.99999999999 170500.00000000003 37199.99999999999 171300.0 ;
      RECT  40599.99999999999 176500.00000000003 39800.0 177300.0 ;
      RECT  40599.99999999999 192100.00000000003 39800.0 192900.0 ;
      RECT  40599.99999999999 194900.0 39800.0 195700.00000000003 ;
      RECT  40599.99999999999 210500.00000000003 39800.0 211300.0 ;
      RECT  40599.99999999999 213300.0 39800.0 214100.00000000003 ;
      RECT  40599.99999999999 228900.0 39800.0 229700.00000000003 ;
      RECT  40599.99999999999 231700.00000000003 39800.0 232500.00000000003 ;
      RECT  40599.99999999999 247300.0 39800.0 248100.0 ;
      RECT  18799.999999999993 173100.00000000003 19599.999999999993 173900.0 ;
      RECT  18799.999999999993 173100.00000000003 19599.999999999993 173900.0 ;
      RECT  19599.999999999993 170900.0 20399.999999999996 171700.00000000003 ;
      RECT  17999.999999999993 170900.0 18799.999999999993 171700.00000000003 ;
      RECT  11199.999999999993 170700.00000000003 11999.999999999993 171500.00000000003 ;
      RECT  5899.999999999992 43800.000000000015 5099.999999999992 44600.00000000001 ;
      RECT  41899.99999999999 43800.000000000015 41099.99999999999 44600.00000000001 ;
      RECT  37699.99999999999 71800.00000000001 36900.0 72600.00000000001 ;
      RECT  40499.99999999999 90600.00000000001 39699.99999999999 91400.0 ;
      RECT  37699.99999999999 116200.00000000001 36900.0 117000.00000000001 ;
      RECT  43300.0 117600.00000000001 42500.0 118400.0 ;
      RECT  60399.99999999999 111800.00000000001 59599.99999999999 112600.00000000001 ;
      RECT  39099.99999999999 125800.00000000001 38300.0 126600.00000000001 ;
      RECT  43300.0 124400.0 42500.0 125200.0 ;
      RECT  11999.999999999993 151400.0 11199.999999999993 152200.00000000003 ;
      RECT  48399.99999999999 10800.000000000005 49199.999999999985 11600.000000000007 ;
      RECT  56399.99999999999 10200.000000000007 57199.999999999985 11000.000000000007 ;
      RECT  41899.99999999999 31200.000000000007 41099.99999999999 32000.000000000007 ;
      RECT  54800.0 36200.00000000001 55599.99999999999 37000.00000000001 ;
      RECT  66000.0 31800.000000000007 66800.0 32600.000000000007 ;
      RECT  41899.99999999999 45800.000000000015 41099.99999999999 46600.00000000001 ;
      RECT  44699.99999999999 44400.00000000001 43900.0 45200.0 ;
      RECT  59599.99999999999 50200.00000000001 60399.99999999999 51000.00000000001 ;
      RECT  71199.99999999999 21000.000000000007 70399.99999999999 21800.000000000007 ;
      RECT  71199.99999999999 1000.0000000000058 70399.99999999999 1800.0000000000057 ;
      RECT  71199.99999999999 21000.000000000007 70399.99999999999 21800.000000000007 ;
      RECT  71199.99999999999 41000.00000000001 70399.99999999999 41800.00000000001 ;
      RECT  71199.99999999999 61000.00000000001 70399.99999999999 61800.00000000001 ;
      RECT  71199.99999999999 41000.00000000001 70399.99999999999 41800.00000000001 ;
      RECT  71199.99999999999 61000.00000000001 70399.99999999999 61800.00000000001 ;
      RECT  71199.99999999999 81000.00000000001 70399.99999999999 81800.00000000001 ;
      RECT  71199.99999999999 101000.00000000001 70399.99999999999 101800.00000000001 ;
      RECT  71199.99999999999 81000.00000000001 70399.99999999999 81800.00000000001 ;
      RECT  71199.99999999999 101000.00000000001 70399.99999999999 101800.00000000001 ;
      RECT  71199.99999999999 121000.00000000001 70399.99999999999 121800.00000000001 ;
      RECT  71199.99999999999 141000.0 70399.99999999999 141800.0 ;
      RECT  71199.99999999999 121000.00000000001 70399.99999999999 121800.00000000001 ;
      RECT  71199.99999999999 141000.0 70399.99999999999 141800.0 ;
      RECT  71199.99999999999 161000.00000000003 70399.99999999999 161800.00000000003 ;
      RECT  56800.0 151900.0 72199.99999999999 152500.0 ;
      RECT  56800.0 90300.00000000001 72199.99999999999 90900.0 ;
      RECT  66399.99999999999 130300.00000000001 72199.99999999999 130900.0 ;
      RECT  59899.99999999999 71900.0 72199.99999999999 72500.00000000001 ;
      RECT  56800.0 10300.000000000005 72199.99999999999 10900.000000000005 ;
      RECT  50400.0 256100.00000000003 72200.0 276100.0 ;
      RECT  50400.0 296100.0 72200.0 276100.0 ;
      RECT  50400.0 296100.0 72200.0 316100.0 ;
      RECT  50400.0 336100.0 72200.0 316100.0 ;
      RECT  61700.0 275700.00000000006 60900.0 276500.0 ;
      RECT  61700.0 255700.00000000003 60900.0 256500.0 ;
      RECT  61700.0 275700.00000000006 60900.0 276500.0 ;
      RECT  61700.0 295700.00000000006 60900.0 296500.0 ;
      RECT  61700.0 315700.00000000006 60900.0 316500.0 ;
      RECT  61700.0 295700.00000000006 60900.0 296500.0 ;
      RECT  61700.0 315700.00000000006 60900.0 316500.0 ;
      RECT  61700.0 335700.00000000006 60900.0 336500.0 ;
      RECT  171400.0 43200.0 193200.00000000003 63200.0 ;
      RECT  193200.00000000003 43200.0 215000.0 63200.0 ;
      RECT  182700.00000000003 62800.00000000001 181900.0 63600.00000000001 ;
      RECT  182700.00000000003 42800.00000000001 181900.0 43600.0 ;
      RECT  204500.0 62800.00000000001 203700.00000000003 63600.00000000001 ;
      RECT  204500.0 42800.00000000001 203700.00000000003 43600.0 ;
      RECT  74000.0 10200.000000000004 73200.0 11000.000000000004 ;
      RECT  72600.0 151800.0 71800.0 152600.00000000003 ;
      RECT  72600.0 90200.0 71800.0 91000.0 ;
      RECT  72600.0 130199.99999999999 71800.0 131000.0 ;
      RECT  72600.0 71800.0 71800.0 72600.0 ;
      RECT  174400.0 65600.00000000001 175200.00000000003 66400.0 ;
      RECT  190200.0 65600.00000000001 191000.0 66400.0 ;
      RECT  181200.0 67000.0 182000.0 67800.0 ;
      RECT  212000.0 67000.0 212800.0 67800.0 ;
   LAYER  metal2 ;
      RECT  73300.0 10600.000000000002 73899.99999999999 261500.0 ;
      RECT  73200.0 10600.000000000002 74000.0 48600.0 ;
      RECT  73300.0 10600.000000000002 73899.99999999999 48600.0 ;
      RECT  168000.0 117900.0 168600.0 152200.00000000003 ;
      RECT  166600.00000000003 90600.00000000001 167200.00000000003 117900.0 ;
      RECT  169400.0 117900.0 170000.0 130600.0 ;
      RECT  165200.0 72200.0 165799.99999999997 117900.0 ;
      RECT  75100.0 205600.00000000003 75699.99999999999 265900.00000000006 ;
      RECT  76500.0 205600.00000000003 77100.0 286300.0 ;
      RECT  77900.0 205600.00000000003 78500.0 305900.00000000006 ;
      RECT  79300.0 205600.00000000003 79899.99999999999 326300.0 ;
      RECT  174500.0 66000.0 175100.0 71200.0 ;
      RECT  190300.0 53000.0 190900.0 66000.0 ;
      RECT  181300.0 67400.0 181900.0 71200.0 ;
      RECT  212100.0 53000.0 212700.0 67400.0 ;
      RECT  173500.0 111700.0 174100.0 112300.00000000001 ;
      RECT  173500.0 109600.0 174100.0 112000.0 ;
      RECT  173500.0 112000.0 174100.0 135900.0 ;
      RECT  175500.0 113100.0 176100.0 113700.0 ;
      RECT  175500.0 108100.0 176100.0 113400.0 ;
      RECT  175500.0 113400.0 176100.0 135900.0 ;
      RECT  180300.0 111700.0 180900.0 112300.00000000001 ;
      RECT  180300.0 109600.0 180900.0 112000.0 ;
      RECT  180300.0 112000.0 180900.0 135900.0 ;
      RECT  182300.0 113100.0 182900.0 113700.0 ;
      RECT  182300.0 108100.0 182900.0 113400.0 ;
      RECT  182300.0 113400.0 182900.0 135900.0 ;
      RECT  172700.0 148500.0 174100.00000000003 149100.0 ;
      RECT  173500.0 135900.0 174100.0 148800.0 ;
      RECT  172700.0 148800.0 173300.0 157899.99999999997 ;
      RECT  175500.0 149900.0 176900.0 150500.0 ;
      RECT  175500.0 135900.0 176100.0 150200.0 ;
      RECT  176300.0 150200.0 176900.0 157900.0 ;
      RECT  179500.0 148500.0 180900.0 149100.0 ;
      RECT  180300.0 135900.0 180900.0 148800.0 ;
      RECT  179500.0 148800.0 180100.0 157899.99999999997 ;
      RECT  182300.0 149900.0 183700.00000000003 150500.0 ;
      RECT  182300.0 135900.0 182900.0 150200.0 ;
      RECT  183100.00000000003 150200.0 183700.0 157900.0 ;
      RECT  172700.0 164200.0 173300.0 166100.00000000003 ;
      RECT  172700.0 166100.00000000003 173300.0 168000.0 ;
      RECT  176300.0 164200.0 176900.0 166100.00000000003 ;
      RECT  176300.0 166100.00000000003 176900.0 168800.0 ;
      RECT  179500.0 164200.0 180100.0 166100.00000000003 ;
      RECT  179500.0 166100.00000000003 180100.0 168000.0 ;
      RECT  183100.00000000003 164200.0 183700.0 166100.00000000003 ;
      RECT  183100.00000000003 166100.00000000003 183700.0 168800.0 ;
      RECT  147100.00000000003 164600.00000000003 147700.0 168800.0 ;
      RECT  171400.0 168400.0 178200.0 177600.00000000003 ;
      RECT  171400.0 186800.0 178200.0 177600.00000000003 ;
      RECT  171400.0 186800.0 178200.0 196000.0 ;
      RECT  171400.0 205200.0 178200.0 196000.0 ;
      RECT  171400.0 205200.0 178200.0 214400.00000000003 ;
      RECT  171400.0 223600.00000000003 178200.0 214399.99999999997 ;
      RECT  171400.0 223600.00000000003 178200.0 232800.0 ;
      RECT  171400.0 242000.0 178200.0 232800.0 ;
      RECT  171400.0 242000.0 178200.0 251200.0 ;
      RECT  171400.0 260399.99999999997 178200.0 251200.0 ;
      RECT  171400.0 260399.99999999997 178200.0 269600.0 ;
      RECT  171400.0 278800.0 178200.0 269600.0 ;
      RECT  171400.0 278800.0 178200.0 288000.0 ;
      RECT  171400.0 297200.0 178200.0 288000.0 ;
      RECT  171400.0 297200.0 178200.0 306400.0 ;
      RECT  171400.0 315600.0 178200.0 306400.00000000006 ;
      RECT  178200.0 168400.0 185000.0 177600.00000000003 ;
      RECT  178200.0 186800.0 185000.0 177600.00000000003 ;
      RECT  178200.0 186800.0 185000.0 196000.0 ;
      RECT  178200.0 205200.0 185000.0 196000.0 ;
      RECT  178200.0 205200.0 185000.0 214400.00000000003 ;
      RECT  178200.0 223600.00000000003 185000.0 214399.99999999997 ;
      RECT  178200.0 223600.00000000003 185000.0 232800.0 ;
      RECT  178200.0 242000.0 185000.0 232800.0 ;
      RECT  178200.0 242000.0 185000.0 251200.0 ;
      RECT  178200.0 260399.99999999997 185000.0 251200.0 ;
      RECT  178200.0 260399.99999999997 185000.0 269600.0 ;
      RECT  178200.0 278800.0 185000.0 269600.0 ;
      RECT  178200.0 278800.0 185000.0 288000.0 ;
      RECT  178200.0 297200.0 185000.0 288000.0 ;
      RECT  178200.0 297200.0 185000.0 306400.0 ;
      RECT  178200.0 315600.0 185000.0 306400.00000000006 ;
      RECT  174400.0 177200.0 175200.0 178000.0 ;
      RECT  171000.0 172600.00000000003 171800.0 173400.0 ;
      RECT  177800.0 172600.00000000003 178600.00000000003 173400.0 ;
      RECT  181200.0 177200.0 182000.0 178000.0 ;
      RECT  177800.0 172600.00000000003 178600.00000000003 173400.0 ;
      RECT  184600.00000000003 172600.00000000003 185400.0 173400.0 ;
      RECT  174400.0 177200.0 175200.0 178000.0 ;
      RECT  171000.0 181800.0 171800.0 182600.00000000003 ;
      RECT  177800.0 181800.0 178600.00000000003 182600.00000000003 ;
      RECT  181200.0 177200.0 182000.0 178000.0 ;
      RECT  177800.0 181800.0 178600.00000000003 182600.00000000003 ;
      RECT  184600.00000000003 181800.0 185400.0 182600.00000000003 ;
      RECT  174400.0 195600.00000000003 175200.0 196400.0 ;
      RECT  171000.0 191000.0 171800.0 191800.0 ;
      RECT  177800.0 191000.0 178600.00000000003 191800.0 ;
      RECT  181200.0 195600.00000000003 182000.0 196400.0 ;
      RECT  177800.0 191000.0 178600.00000000003 191800.0 ;
      RECT  184600.00000000003 191000.0 185400.0 191800.0 ;
      RECT  174400.0 195600.00000000003 175200.0 196400.0 ;
      RECT  171000.0 200200.0 171800.0 201000.0 ;
      RECT  177800.0 200200.0 178600.00000000003 201000.0 ;
      RECT  181200.0 195600.00000000003 182000.0 196400.0 ;
      RECT  177800.0 200200.0 178600.00000000003 201000.0 ;
      RECT  184600.00000000003 200200.0 185400.0 201000.0 ;
      RECT  174400.0 214000.0 175200.0 214800.0 ;
      RECT  171000.0 209399.99999999997 171800.0 210200.0 ;
      RECT  177800.0 209399.99999999997 178600.00000000003 210200.0 ;
      RECT  181200.0 214000.0 182000.0 214800.0 ;
      RECT  177800.0 209399.99999999997 178600.00000000003 210200.0 ;
      RECT  184600.00000000003 209399.99999999997 185400.0 210200.0 ;
      RECT  174400.0 214000.0 175200.0 214800.0 ;
      RECT  171000.0 218600.00000000003 171800.0 219399.99999999997 ;
      RECT  177800.0 218600.00000000003 178600.00000000003 219399.99999999997 ;
      RECT  181200.0 214000.0 182000.0 214800.0 ;
      RECT  177800.0 218600.00000000003 178600.00000000003 219399.99999999997 ;
      RECT  184600.00000000003 218600.00000000003 185400.0 219399.99999999997 ;
      RECT  174400.0 232399.99999999997 175200.0 233200.0 ;
      RECT  171000.0 227800.0 171800.0 228600.00000000003 ;
      RECT  177800.0 227800.0 178600.00000000003 228600.00000000003 ;
      RECT  181200.0 232399.99999999997 182000.0 233200.0 ;
      RECT  177800.0 227800.0 178600.00000000003 228600.00000000003 ;
      RECT  184600.00000000003 227800.0 185400.0 228600.00000000003 ;
      RECT  174400.0 232399.99999999997 175200.0 233200.0 ;
      RECT  171000.0 237000.0 171800.0 237800.0 ;
      RECT  177800.0 237000.0 178600.00000000003 237800.0 ;
      RECT  181200.0 232399.99999999997 182000.0 233200.0 ;
      RECT  177800.0 237000.0 178600.00000000003 237800.0 ;
      RECT  184600.00000000003 237000.0 185400.0 237800.0 ;
      RECT  174400.0 250800.0 175200.0 251600.00000000003 ;
      RECT  171000.0 246200.0 171800.0 247000.0 ;
      RECT  177800.0 246200.0 178600.00000000003 247000.0 ;
      RECT  181200.0 250800.0 182000.0 251600.00000000003 ;
      RECT  177800.0 246200.0 178600.00000000003 247000.0 ;
      RECT  184600.00000000003 246200.0 185400.0 247000.0 ;
      RECT  174400.0 250800.0 175200.0 251600.00000000003 ;
      RECT  171000.0 255399.99999999997 171800.0 256200.0 ;
      RECT  177800.0 255399.99999999997 178600.00000000003 256200.0 ;
      RECT  181200.0 250800.0 182000.0 251600.00000000003 ;
      RECT  177800.0 255399.99999999997 178600.00000000003 256200.0 ;
      RECT  184600.00000000003 255399.99999999997 185400.0 256200.0 ;
      RECT  174400.0 269200.0 175200.0 270000.0 ;
      RECT  171000.0 264600.0 171800.0 265400.0 ;
      RECT  177800.0 264600.0 178600.00000000003 265400.0 ;
      RECT  181200.0 269200.0 182000.0 270000.0 ;
      RECT  177800.0 264600.0 178600.00000000003 265400.0 ;
      RECT  184600.00000000003 264600.0 185400.0 265400.0 ;
      RECT  174400.0 269200.0 175200.0 270000.0 ;
      RECT  171000.0 273800.0 171800.0 274600.0 ;
      RECT  177800.0 273800.0 178600.00000000003 274600.0 ;
      RECT  181200.0 269200.0 182000.0 270000.0 ;
      RECT  177800.0 273800.0 178600.00000000003 274600.0 ;
      RECT  184600.00000000003 273800.0 185400.0 274600.0 ;
      RECT  174400.0 287600.0 175200.0 288400.0 ;
      RECT  171000.0 283000.0 171800.0 283800.0 ;
      RECT  177800.0 283000.0 178600.00000000003 283800.0 ;
      RECT  181200.0 287600.0 182000.0 288400.0 ;
      RECT  177800.0 283000.0 178600.00000000003 283800.0 ;
      RECT  184600.00000000003 283000.0 185400.0 283800.0 ;
      RECT  174400.0 287600.0 175200.0 288400.0 ;
      RECT  171000.0 292200.0 171800.0 293000.0 ;
      RECT  177800.0 292200.0 178600.00000000003 293000.0 ;
      RECT  181200.0 287600.0 182000.0 288400.0 ;
      RECT  177800.0 292200.0 178600.00000000003 293000.0 ;
      RECT  184600.00000000003 292200.0 185400.0 293000.0 ;
      RECT  174400.0 306000.0 175200.0 306800.0 ;
      RECT  171000.0 301400.0 171800.0 302200.0 ;
      RECT  177800.0 301400.0 178600.00000000003 302200.0 ;
      RECT  181200.0 306000.0 182000.0 306800.0 ;
      RECT  177800.0 301400.0 178600.00000000003 302200.0 ;
      RECT  184600.00000000003 301400.0 185400.0 302200.0 ;
      RECT  174400.0 306000.0 175200.0 306800.0 ;
      RECT  171000.0 310600.0 171800.0 311400.00000000006 ;
      RECT  177800.0 310600.0 178600.00000000003 311400.00000000006 ;
      RECT  181200.0 306000.0 182000.0 306800.0 ;
      RECT  177800.0 310600.0 178600.00000000003 311400.00000000006 ;
      RECT  184600.00000000003 310600.0 185400.0 311400.00000000006 ;
      RECT  172600.00000000003 168000.0 173400.0 317000.0 ;
      RECT  176200.0 168800.0 177000.0 317800.0 ;
      RECT  179400.0 168000.0 180200.0 317000.0 ;
      RECT  183000.0 168800.0 183800.0 317800.0 ;
      RECT  174200.0 158000.0 175000.0 158800.0 ;
      RECT  174200.0 158000.0 175000.0 158800.0 ;
      RECT  172600.00000000003 158000.0 173400.0 158800.0 ;
      RECT  172600.00000000003 153200.0 173400.0 154000.0 ;
      RECT  176200.0 158000.0 177000.0 158800.0 ;
      RECT  176200.0 153200.0 177000.0 154000.0 ;
      RECT  172700.0 151600.00000000003 173300.0 164200.0 ;
      RECT  176300.0 151600.00000000003 176900.0 164200.0 ;
      RECT  181000.0 158000.0 181800.0 158800.0 ;
      RECT  181000.0 158000.0 181800.0 158800.0 ;
      RECT  179400.0 158000.0 180200.0 158800.0 ;
      RECT  179400.0 153200.0 180200.0 154000.0 ;
      RECT  183000.0 158000.0 183800.0 158800.0 ;
      RECT  183000.0 153200.0 183800.0 154000.0 ;
      RECT  179500.0 151600.00000000003 180100.00000000003 164200.0 ;
      RECT  183100.00000000003 151600.00000000003 183700.0 164200.0 ;
      RECT  172700.0 151600.00000000003 173300.0 164200.0 ;
      RECT  176300.0 151600.00000000003 176900.0 164200.0 ;
      RECT  179500.0 151600.00000000003 180100.00000000003 164200.0 ;
      RECT  183100.00000000003 151600.00000000003 183700.0 164200.0 ;
      RECT  171400.0 114800.00000000001 178200.0 147400.0 ;
      RECT  178200.0 114800.00000000001 185000.0 147400.0 ;
      RECT  177800.0 141000.0 178600.00000000003 141800.0 ;
      RECT  176800.0 127600.00000000001 177600.00000000003 128400.0 ;
      RECT  184600.00000000003 141000.0 185400.0 141800.0 ;
      RECT  183600.00000000003 127600.00000000001 184400.0 128400.0 ;
      RECT  172000.0 114800.00000000001 172800.0 117800.00000000001 ;
      RECT  173400.0 124400.0 174200.0 147400.0 ;
      RECT  175400.0 124400.0 176200.0 147400.0 ;
      RECT  178800.0 114800.00000000001 179600.00000000003 117800.00000000001 ;
      RECT  180200.0 124400.0 181000.0 147400.0 ;
      RECT  182200.0 124400.0 183000.0 147400.0 ;
      RECT  171400.0 70200.0 178200.0 110600.0 ;
      RECT  178200.0 70200.0 185000.0 110600.0 ;
      RECT  175200.0 76400.0 176000.0 77200.0 ;
      RECT  174600.00000000003 93800.00000000001 175400.0 94600.00000000001 ;
      RECT  175200.0 83000.0 176000.0 83800.00000000001 ;
      RECT  176600.00000000003 87400.0 177400.0 88200.0 ;
      RECT  176000.0 100800.00000000001 176800.0 101600.00000000001 ;
      RECT  182000.0 76400.0 182800.0 77200.0 ;
      RECT  181400.0 93800.00000000001 182200.0 94600.00000000001 ;
      RECT  182000.0 83000.0 182800.0 83800.00000000001 ;
      RECT  183400.0 87400.0 184200.0 88200.0 ;
      RECT  182800.0 100800.00000000001 183600.00000000003 101600.00000000001 ;
      RECT  174400.0 70200.0 175200.0 72200.0 ;
      RECT  181200.0 70200.0 182000.0 72200.0 ;
      RECT  173400.0 108600.00000000001 174200.0 110600.00000000001 ;
      RECT  175400.0 105600.0 176200.0 110600.00000000001 ;
      RECT  180200.0 108600.00000000001 181000.0 110600.00000000001 ;
      RECT  182200.0 105600.0 183000.0 110600.00000000001 ;
      RECT  112600.0 173500.0 113200.0 177800.0 ;
      RECT  112600.0 183100.00000000003 113200.0 187400.0 ;
      RECT  112600.0 191900.0 113200.0 196200.0 ;
      RECT  112600.0 201500.0 113200.0 205800.0 ;
      RECT  112600.0 210300.0 113200.0 214600.00000000003 ;
      RECT  112600.0 219899.99999999997 113200.0 224200.0 ;
      RECT  112600.0 228700.0 113200.0 233000.0 ;
      RECT  112600.0 238300.0 113200.0 242600.00000000003 ;
      RECT  94100.0 170000.0 94700.0 205600.00000000003 ;
      RECT  95500.0 170000.0 96100.0 205600.00000000003 ;
      RECT  96900.0 170000.0 97500.0 205600.00000000003 ;
      RECT  98300.0 170000.0 98900.0 205600.00000000003 ;
      RECT  105600.0 176000.0 106200.0 176600.00000000003 ;
      RECT  105600.0 170200.0 106200.0 170800.0 ;
      RECT  102900.0 176000.0 105900.0 176600.00000000003 ;
      RECT  105600.0 173600.00000000003 106200.0 176300.0 ;
      RECT  105600.0 170500.0 106200.0 173600.00000000003 ;
      RECT  104500.0 170200.0 105900.0 170800.0 ;
      RECT  102500.0 175900.0 103300.00000000001 176700.0 ;
      RECT  104100.0 170100.00000000003 104900.0 170900.0 ;
      RECT  106300.00000000001 173200.0 105500.0 174000.0 ;
      RECT  105600.0 180000.0 106200.0 179400.0 ;
      RECT  105600.0 185800.0 106200.0 185200.0 ;
      RECT  102900.0 180000.0 105900.0 179400.0 ;
      RECT  105600.0 182400.0 106200.0 179700.0 ;
      RECT  105600.0 185500.0 106200.0 182400.0 ;
      RECT  104500.0 185800.0 105900.0 185200.0 ;
      RECT  102500.0 180100.00000000003 103300.00000000001 179300.0 ;
      RECT  104100.0 185900.0 104900.0 185100.00000000003 ;
      RECT  106300.00000000001 182800.0 105500.0 182000.0 ;
      RECT  105600.0 194400.0 106200.0 195000.0 ;
      RECT  105600.0 188600.00000000003 106200.0 189200.0 ;
      RECT  102900.0 194400.0 105900.0 195000.0 ;
      RECT  105600.0 192000.0 106200.0 194700.0 ;
      RECT  105600.0 188900.0 106200.0 192000.0 ;
      RECT  104500.0 188600.00000000003 105900.0 189200.0 ;
      RECT  102500.0 194300.0 103300.00000000001 195100.00000000003 ;
      RECT  104100.0 188500.0 104900.0 189300.0 ;
      RECT  106300.00000000001 191600.00000000003 105500.0 192400.0 ;
      RECT  105600.0 198400.00000000003 106200.0 197800.0 ;
      RECT  105600.0 204200.0 106200.0 203600.00000000003 ;
      RECT  102900.0 198400.00000000003 105900.0 197800.0 ;
      RECT  105600.0 200800.0 106200.0 198100.00000000003 ;
      RECT  105600.0 203899.99999999997 106200.0 200800.0 ;
      RECT  104500.0 204200.0 105900.0 203600.00000000003 ;
      RECT  102500.0 198500.0 103300.00000000001 197700.0 ;
      RECT  104100.0 204300.0 104900.0 203500.0 ;
      RECT  106300.00000000001 201200.0 105500.0 200400.00000000003 ;
      RECT  94800.00000000001 175800.0 94000.0 176600.00000000003 ;
      RECT  83100.0 172800.0 82300.0 173600.00000000003 ;
      RECT  96200.0 185000.0 95400.0 185800.0 ;
      RECT  84500.0 182400.0 83700.0 183200.0 ;
      RECT  83100.0 188200.0 82300.0 189000.0 ;
      RECT  97600.0 188200.0 96800.0 189000.0 ;
      RECT  84500.0 197400.0 83700.0 198200.0 ;
      RECT  99000.0 197400.0 98200.0 198200.0 ;
      RECT  94800.00000000001 173200.0 94000.0 174000.0 ;
      RECT  96200.0 171800.0 95400.0 172600.00000000003 ;
      RECT  97600.0 182000.0 96800.0 182800.0 ;
      RECT  96200.0 183400.0 95400.0 184200.0 ;
      RECT  94800.00000000001 191600.00000000003 94000.0 192400.0 ;
      RECT  99000.0 190200.0 98200.0 191000.0 ;
      RECT  97600.0 200399.99999999997 96800.0 201200.0 ;
      RECT  99000.0 201800.0 98200.0 202600.00000000003 ;
      RECT  91700.0 177600.00000000003 90900.0 178400.0 ;
      RECT  91700.0 177600.00000000003 90900.0 178400.0 ;
      RECT  109100.0 177600.00000000003 108300.0 178400.0 ;
      RECT  109100.0 177600.00000000003 108300.0 178400.0 ;
      RECT  91700.0 168400.0 90900.0 169200.0 ;
      RECT  91700.0 168400.0 90900.0 169200.0 ;
      RECT  109100.0 168400.0 108300.0 169200.0 ;
      RECT  109100.0 168400.0 108300.0 169200.0 ;
      RECT  91700.0 177600.00000000003 90900.0 178400.0 ;
      RECT  91700.0 177600.00000000003 90900.0 178400.0 ;
      RECT  109100.0 177600.00000000003 108300.0 178400.0 ;
      RECT  109100.0 177600.00000000003 108300.0 178400.0 ;
      RECT  91700.0 186800.0 90900.0 187600.00000000003 ;
      RECT  91700.0 186800.0 90900.0 187600.00000000003 ;
      RECT  109100.0 186800.0 108300.0 187600.00000000003 ;
      RECT  109100.0 186800.0 108300.0 187600.00000000003 ;
      RECT  91700.0 196000.0 90900.0 196800.0 ;
      RECT  91700.0 196000.0 90900.0 196800.0 ;
      RECT  109100.0 196000.0 108300.0 196800.0 ;
      RECT  109100.0 196000.0 108300.0 196800.0 ;
      RECT  91700.0 186800.0 90900.0 187600.00000000003 ;
      RECT  91700.0 186800.0 90900.0 187600.00000000003 ;
      RECT  109100.0 186800.0 108300.0 187600.00000000003 ;
      RECT  109100.0 186800.0 108300.0 187600.00000000003 ;
      RECT  91700.0 196000.0 90900.0 196800.0 ;
      RECT  91700.0 196000.0 90900.0 196800.0 ;
      RECT  109100.0 196000.0 108300.0 196800.0 ;
      RECT  109100.0 196000.0 108300.0 196800.0 ;
      RECT  91700.0 205200.0 90900.0 206000.0 ;
      RECT  91700.0 205200.0 90900.0 206000.0 ;
      RECT  109100.0 205200.0 108300.0 206000.0 ;
      RECT  109100.0 205200.0 108300.0 206000.0 ;
      RECT  82400.0 170000.0 83000.0 205600.00000000003 ;
      RECT  83800.0 170000.0 84400.0 205600.00000000003 ;
      RECT  94100.0 206800.0 94700.0 242399.99999999997 ;
      RECT  95500.0 206800.0 96100.0 242399.99999999997 ;
      RECT  96900.0 206800.0 97500.0 242399.99999999997 ;
      RECT  98300.0 206800.0 98900.0 242399.99999999997 ;
      RECT  105600.0 212800.0 106200.0 213399.99999999997 ;
      RECT  105600.0 207000.0 106200.0 207600.00000000003 ;
      RECT  102900.0 212800.0 105900.0 213399.99999999997 ;
      RECT  105600.0 210399.99999999997 106200.0 213100.00000000003 ;
      RECT  105600.0 207300.0 106200.0 210399.99999999997 ;
      RECT  104500.0 207000.0 105900.0 207600.00000000003 ;
      RECT  102500.0 212700.0 103300.00000000001 213500.0 ;
      RECT  104100.0 206899.99999999997 104900.0 207700.0 ;
      RECT  106300.00000000001 210000.0 105500.0 210800.0 ;
      RECT  105600.0 216800.0 106200.0 216200.0 ;
      RECT  105600.0 222600.00000000003 106200.0 222000.0 ;
      RECT  102900.0 216800.0 105900.0 216200.0 ;
      RECT  105600.0 219200.0 106200.0 216500.0 ;
      RECT  105600.0 222300.0 106200.0 219200.0 ;
      RECT  104500.0 222600.00000000003 105900.0 222000.0 ;
      RECT  102500.0 216899.99999999997 103300.00000000001 216100.00000000003 ;
      RECT  104100.0 222700.0 104900.0 221899.99999999997 ;
      RECT  106300.00000000001 219600.00000000003 105500.0 218800.0 ;
      RECT  105600.0 231200.0 106200.0 231800.0 ;
      RECT  105600.0 225399.99999999997 106200.0 226000.0 ;
      RECT  102900.0 231200.0 105900.0 231800.0 ;
      RECT  105600.0 228800.0 106200.0 231500.0 ;
      RECT  105600.0 225700.0 106200.0 228800.0 ;
      RECT  104500.0 225399.99999999997 105900.0 226000.0 ;
      RECT  102500.0 231100.00000000003 103300.00000000001 231900.00000000003 ;
      RECT  104100.0 225300.0 104900.0 226100.00000000003 ;
      RECT  106300.00000000001 228400.00000000003 105500.0 229200.0 ;
      RECT  105600.0 235200.0 106200.0 234600.00000000003 ;
      RECT  105600.0 241000.0 106200.0 240399.99999999997 ;
      RECT  102900.0 235200.0 105900.0 234600.00000000003 ;
      RECT  105600.0 237600.00000000003 106200.0 234899.99999999997 ;
      RECT  105600.0 240700.0 106200.0 237600.00000000003 ;
      RECT  104500.0 241000.0 105900.0 240399.99999999997 ;
      RECT  102500.0 235300.0 103300.00000000001 234500.0 ;
      RECT  104100.0 241100.00000000003 104900.0 240300.0 ;
      RECT  106300.00000000001 238000.0 105500.0 237200.0 ;
      RECT  94800.00000000001 212600.00000000003 94000.0 213399.99999999997 ;
      RECT  83100.0 209600.00000000003 82300.0 210399.99999999997 ;
      RECT  96200.0 221800.0 95400.0 222600.00000000003 ;
      RECT  84500.0 219200.0 83700.0 220000.0 ;
      RECT  83100.0 225000.0 82300.0 225800.0 ;
      RECT  97600.0 225000.0 96800.0 225800.0 ;
      RECT  84500.0 234200.0 83700.0 235000.0 ;
      RECT  99000.0 234200.0 98200.0 235000.0 ;
      RECT  94800.00000000001 210000.0 94000.0 210800.0 ;
      RECT  96200.0 208600.00000000003 95400.0 209399.99999999997 ;
      RECT  97600.0 218800.0 96800.0 219600.00000000003 ;
      RECT  96200.0 220200.0 95400.0 221000.0 ;
      RECT  94800.00000000001 228399.99999999997 94000.0 229200.0 ;
      RECT  99000.0 227000.0 98200.0 227800.0 ;
      RECT  97600.0 237200.0 96800.0 238000.0 ;
      RECT  99000.0 238600.00000000003 98200.0 239399.99999999997 ;
      RECT  91700.0 214399.99999999997 90900.0 215200.0 ;
      RECT  91700.0 214399.99999999997 90900.0 215200.0 ;
      RECT  109100.0 214399.99999999997 108300.0 215200.0 ;
      RECT  109100.0 214399.99999999997 108300.0 215200.0 ;
      RECT  91700.0 205200.0 90900.0 206000.0 ;
      RECT  91700.0 205200.0 90900.0 206000.0 ;
      RECT  109100.0 205200.0 108300.0 206000.0 ;
      RECT  109100.0 205200.0 108300.0 206000.0 ;
      RECT  91700.0 214399.99999999997 90900.0 215200.0 ;
      RECT  91700.0 214399.99999999997 90900.0 215200.0 ;
      RECT  109100.0 214399.99999999997 108300.0 215200.0 ;
      RECT  109100.0 214399.99999999997 108300.0 215200.0 ;
      RECT  91700.0 223600.00000000003 90900.0 224399.99999999997 ;
      RECT  91700.0 223600.00000000003 90900.0 224399.99999999997 ;
      RECT  109100.0 223600.00000000003 108300.0 224399.99999999997 ;
      RECT  109100.0 223600.00000000003 108300.0 224399.99999999997 ;
      RECT  91700.0 232800.0 90900.0 233600.00000000003 ;
      RECT  91700.0 232800.0 90900.0 233600.00000000003 ;
      RECT  109100.0 232800.0 108300.0 233600.00000000003 ;
      RECT  109100.0 232800.0 108300.0 233600.00000000003 ;
      RECT  91700.0 223600.00000000003 90900.0 224399.99999999997 ;
      RECT  91700.0 223600.00000000003 90900.0 224399.99999999997 ;
      RECT  109100.0 223600.00000000003 108300.0 224399.99999999997 ;
      RECT  109100.0 223600.00000000003 108300.0 224399.99999999997 ;
      RECT  91700.0 232800.0 90900.0 233600.00000000003 ;
      RECT  91700.0 232800.0 90900.0 233600.00000000003 ;
      RECT  109100.0 232800.0 108300.0 233600.00000000003 ;
      RECT  109100.0 232800.0 108300.0 233600.00000000003 ;
      RECT  91700.0 242000.0 90900.0 242800.0 ;
      RECT  91700.0 242000.0 90900.0 242800.0 ;
      RECT  109100.0 242000.0 108300.0 242800.0 ;
      RECT  109100.0 242000.0 108300.0 242800.0 ;
      RECT  82400.0 206800.0 83000.0 242399.99999999997 ;
      RECT  83800.0 206800.0 84400.0 242399.99999999997 ;
      RECT  132800.0 176000.0 133400.0 176600.00000000003 ;
      RECT  132800.0 170200.0 133400.0 170800.0 ;
      RECT  130100.00000000003 176000.0 133100.00000000003 176600.00000000003 ;
      RECT  132800.0 173600.00000000003 133400.0 176300.0 ;
      RECT  132800.0 170500.0 133400.0 173600.00000000003 ;
      RECT  131700.0 170200.0 133100.00000000003 170800.0 ;
      RECT  129699.99999999999 175900.0 130500.0 176700.0 ;
      RECT  131300.0 170100.00000000003 132100.00000000003 170900.0 ;
      RECT  133500.0 173200.0 132700.0 174000.0 ;
      RECT  132800.0 180000.0 133400.0 179400.0 ;
      RECT  132800.0 185800.0 133400.0 185200.0 ;
      RECT  130100.00000000003 180000.0 133100.00000000003 179400.0 ;
      RECT  132800.0 182400.0 133400.0 179700.0 ;
      RECT  132800.0 185500.0 133400.0 182400.0 ;
      RECT  131700.0 185800.0 133100.00000000003 185200.0 ;
      RECT  129699.99999999999 180100.00000000003 130500.0 179300.0 ;
      RECT  131300.0 185900.0 132100.00000000003 185100.00000000003 ;
      RECT  133500.0 182800.0 132700.0 182000.0 ;
      RECT  132800.0 194400.0 133400.0 195000.0 ;
      RECT  132800.0 188600.00000000003 133400.0 189200.0 ;
      RECT  130100.00000000003 194400.0 133100.00000000003 195000.0 ;
      RECT  132800.0 192000.0 133400.0 194700.0 ;
      RECT  132800.0 188900.0 133400.0 192000.0 ;
      RECT  131700.0 188600.00000000003 133100.00000000003 189200.0 ;
      RECT  129699.99999999999 194300.0 130500.0 195100.00000000003 ;
      RECT  131300.0 188500.0 132100.00000000003 189300.0 ;
      RECT  133500.0 191600.00000000003 132700.0 192400.0 ;
      RECT  132800.0 198400.00000000003 133400.0 197800.0 ;
      RECT  132800.0 204200.0 133400.0 203600.00000000003 ;
      RECT  130100.00000000003 198400.00000000003 133100.00000000003 197800.0 ;
      RECT  132800.0 200800.0 133400.0 198100.00000000003 ;
      RECT  132800.0 203899.99999999997 133400.0 200800.0 ;
      RECT  131700.0 204200.0 133100.00000000003 203600.00000000003 ;
      RECT  129699.99999999999 198500.0 130500.0 197700.0 ;
      RECT  131300.0 204300.0 132100.00000000003 203500.0 ;
      RECT  133500.0 201200.0 132700.0 200399.99999999997 ;
      RECT  132800.0 212800.0 133400.0 213399.99999999997 ;
      RECT  132800.0 207000.0 133400.0 207600.00000000003 ;
      RECT  130100.00000000003 212800.0 133100.00000000003 213399.99999999997 ;
      RECT  132800.0 210399.99999999997 133400.0 213100.00000000003 ;
      RECT  132800.0 207300.0 133400.0 210399.99999999997 ;
      RECT  131700.0 207000.0 133100.00000000003 207600.00000000003 ;
      RECT  129699.99999999999 212700.0 130500.0 213500.0 ;
      RECT  131300.0 206899.99999999997 132100.00000000003 207700.0 ;
      RECT  133500.0 210000.0 132700.0 210800.0 ;
      RECT  132800.0 216800.0 133400.0 216200.0 ;
      RECT  132800.0 222600.00000000003 133400.0 222000.0 ;
      RECT  130100.00000000003 216800.0 133100.00000000003 216200.0 ;
      RECT  132800.0 219200.0 133400.0 216500.0 ;
      RECT  132800.0 222300.0 133400.0 219200.0 ;
      RECT  131700.0 222600.00000000003 133100.00000000003 222000.0 ;
      RECT  129699.99999999999 216899.99999999997 130500.0 216100.00000000003 ;
      RECT  131300.0 222700.0 132100.00000000003 221899.99999999997 ;
      RECT  133500.0 219600.00000000003 132700.0 218800.0 ;
      RECT  132800.0 231200.0 133400.0 231800.0 ;
      RECT  132800.0 225399.99999999997 133400.0 226000.0 ;
      RECT  130100.00000000003 231200.0 133100.00000000003 231800.0 ;
      RECT  132800.0 228800.0 133400.0 231500.0 ;
      RECT  132800.0 225700.0 133400.0 228800.0 ;
      RECT  131700.0 225399.99999999997 133100.00000000003 226000.0 ;
      RECT  129699.99999999999 231100.00000000003 130500.0 231899.99999999997 ;
      RECT  131300.0 225300.0 132100.00000000003 226100.00000000003 ;
      RECT  133500.0 228399.99999999997 132700.0 229200.0 ;
      RECT  132800.0 235200.0 133400.0 234600.00000000003 ;
      RECT  132800.0 241000.0 133400.0 240400.00000000003 ;
      RECT  130100.00000000003 235200.0 133100.00000000003 234600.00000000003 ;
      RECT  132800.0 237600.00000000003 133400.0 234900.00000000003 ;
      RECT  132800.0 240700.0 133400.0 237600.00000000003 ;
      RECT  131700.0 241000.0 133100.00000000003 240400.00000000003 ;
      RECT  129699.99999999999 235300.0 130500.0 234500.0 ;
      RECT  131300.0 241100.00000000003 132100.00000000003 240300.0 ;
      RECT  133500.0 238000.0 132700.0 237200.0 ;
      RECT  132800.0 249600.00000000003 133400.0 250200.0 ;
      RECT  132800.0 243800.0 133400.0 244400.00000000003 ;
      RECT  130100.00000000003 249600.00000000003 133100.00000000003 250200.0 ;
      RECT  132800.0 247200.0 133400.0 249900.00000000003 ;
      RECT  132800.0 244100.00000000003 133400.0 247200.0 ;
      RECT  131700.0 243800.0 133100.00000000003 244400.00000000003 ;
      RECT  129699.99999999999 249500.0 130500.0 250300.0 ;
      RECT  131300.0 243700.0 132100.00000000003 244500.0 ;
      RECT  133500.0 246800.0 132700.0 247600.00000000003 ;
      RECT  132800.0 253600.00000000003 133400.0 253000.0 ;
      RECT  132800.0 259399.99999999997 133400.0 258800.0 ;
      RECT  130100.00000000003 253600.00000000003 133100.00000000003 253000.0 ;
      RECT  132800.0 256000.0 133400.0 253300.0 ;
      RECT  132800.0 259100.00000000003 133400.0 256000.0 ;
      RECT  131700.0 259399.99999999997 133100.00000000003 258800.0 ;
      RECT  129699.99999999999 253700.0 130500.0 252899.99999999997 ;
      RECT  131300.0 259500.0 132100.00000000003 258700.0 ;
      RECT  133500.0 256399.99999999997 132700.0 255600.00000000003 ;
      RECT  132800.0 268000.0 133400.0 268600.0 ;
      RECT  132800.0 262200.0 133400.0 262800.0 ;
      RECT  130100.00000000003 268000.0 133100.00000000003 268600.0 ;
      RECT  132800.0 265600.0 133400.0 268300.0 ;
      RECT  132800.0 262500.0 133400.0 265600.0 ;
      RECT  131700.0 262200.0 133100.00000000003 262800.0 ;
      RECT  129699.99999999999 267900.0 130500.0 268700.0 ;
      RECT  131300.0 262100.00000000003 132100.00000000003 262900.0 ;
      RECT  133500.0 265200.0 132700.0 266000.0 ;
      RECT  132800.0 272000.0 133400.0 271400.00000000006 ;
      RECT  132800.0 277800.0 133400.0 277200.0 ;
      RECT  130100.00000000003 272000.0 133100.00000000003 271400.00000000006 ;
      RECT  132800.0 274400.00000000006 133400.0 271700.0 ;
      RECT  132800.0 277500.0 133400.0 274400.00000000006 ;
      RECT  131700.0 277800.0 133100.00000000003 277200.0 ;
      RECT  129699.99999999999 272100.0 130500.0 271300.0 ;
      RECT  131300.0 277900.00000000006 132100.00000000003 277100.0 ;
      RECT  133500.0 274800.0 132700.0 274000.0 ;
      RECT  132800.0 286400.00000000006 133400.0 287000.0 ;
      RECT  132800.0 280600.0 133400.0 281200.0 ;
      RECT  130100.00000000003 286400.00000000006 133100.00000000003 287000.0 ;
      RECT  132800.0 284000.0 133400.0 286700.0 ;
      RECT  132800.0 280900.00000000006 133400.0 284000.0 ;
      RECT  131700.0 280600.0 133100.00000000003 281200.0 ;
      RECT  129699.99999999999 286300.0 130500.0 287100.0 ;
      RECT  131300.0 280500.0 132100.00000000003 281300.0 ;
      RECT  133500.0 283600.0 132700.0 284400.00000000006 ;
      RECT  132800.0 290400.00000000006 133400.0 289800.0 ;
      RECT  132800.0 296200.0 133400.0 295600.0 ;
      RECT  130100.00000000003 290400.00000000006 133100.00000000003 289800.0 ;
      RECT  132800.0 292800.0 133400.0 290100.0 ;
      RECT  132800.0 295900.00000000006 133400.0 292800.0 ;
      RECT  131700.0 296200.0 133100.00000000003 295600.0 ;
      RECT  129699.99999999999 290500.0 130500.0 289700.0 ;
      RECT  131300.0 296300.0 132100.00000000003 295500.0 ;
      RECT  133500.0 293200.0 132700.0 292400.00000000006 ;
      RECT  132800.0 304800.0 133400.0 305400.00000000006 ;
      RECT  132800.0 299000.0 133400.0 299600.0 ;
      RECT  130100.00000000003 304800.0 133100.00000000003 305400.00000000006 ;
      RECT  132800.0 302400.00000000006 133400.0 305100.0 ;
      RECT  132800.0 299300.0 133400.0 302400.00000000006 ;
      RECT  131700.0 299000.0 133100.00000000003 299600.0 ;
      RECT  129699.99999999999 304700.0 130500.0 305500.0 ;
      RECT  131300.0 298900.00000000006 132100.00000000003 299700.0 ;
      RECT  133500.0 302000.0 132700.0 302800.0 ;
      RECT  132800.0 308800.0 133400.0 308200.0 ;
      RECT  132800.0 314600.0 133400.0 314000.0 ;
      RECT  130100.00000000003 308800.0 133100.00000000003 308200.0 ;
      RECT  132800.0 311200.0 133400.0 308500.0 ;
      RECT  132800.0 314300.0 133400.0 311200.0 ;
      RECT  131700.0 314600.0 133100.00000000003 314000.0 ;
      RECT  129699.99999999999 308900.00000000006 130500.0 308100.0 ;
      RECT  131300.0 314700.0 132100.00000000003 313900.00000000006 ;
      RECT  133500.0 311600.0 132700.0 310800.0 ;
      RECT  83100.0 178800.0 82300.0 179600.00000000003 ;
      RECT  75800.0 178800.0 75000.0 179600.00000000003 ;
      RECT  84500.0 188000.0 83700.0 188800.0 ;
      RECT  77200.0 188000.0 76400.0 188800.0 ;
      RECT  83100.0 215600.00000000003 82300.0 216399.99999999997 ;
      RECT  78600.0 215600.00000000003 77800.0 216399.99999999997 ;
      RECT  84500.0 224800.0 83700.0 225600.00000000003 ;
      RECT  80000.0 224800.0 79200.0 225600.00000000003 ;
      RECT  113300.00000000001 172800.0 112500.0 173600.00000000003 ;
      RECT  113300.00000000001 177400.0 112500.0 178200.0 ;
      RECT  116700.0 177400.0 115900.0 178200.0 ;
      RECT  113300.00000000001 182400.0 112500.0 183200.0 ;
      RECT  113300.00000000001 187000.0 112500.0 187800.0 ;
      RECT  118100.0 187000.0 117300.00000000001 187800.0 ;
      RECT  113300.00000000001 191200.0 112500.0 192000.0 ;
      RECT  113300.00000000001 195800.0 112500.0 196600.00000000003 ;
      RECT  119500.0 195800.0 118700.0 196600.00000000003 ;
      RECT  113300.00000000001 200800.0 112500.0 201600.00000000003 ;
      RECT  113300.00000000001 205399.99999999997 112500.0 206200.0 ;
      RECT  120900.0 205399.99999999997 120100.00000000001 206200.0 ;
      RECT  113300.00000000001 209600.00000000003 112500.0 210399.99999999997 ;
      RECT  113300.00000000001 214200.0 112500.0 215000.0 ;
      RECT  122300.00000000001 214200.0 121500.0 215000.0 ;
      RECT  113300.00000000001 219200.0 112500.0 220000.0 ;
      RECT  113300.00000000001 223800.0 112500.0 224600.00000000003 ;
      RECT  123700.0 223800.0 122900.0 224600.00000000003 ;
      RECT  113300.00000000001 228000.0 112500.0 228800.0 ;
      RECT  113300.00000000001 232600.00000000003 112500.0 233399.99999999997 ;
      RECT  125100.0 232600.00000000003 124300.00000000001 233399.99999999997 ;
      RECT  113300.00000000001 237600.00000000003 112500.0 238399.99999999997 ;
      RECT  113300.00000000001 242200.0 112500.0 243000.0 ;
      RECT  126500.0 242200.0 125700.0 243000.0 ;
      RECT  116700.0 173200.0 115900.0 174000.0 ;
      RECT  122300.00000000001 171800.0 121500.0 172600.00000000003 ;
      RECT  118100.0 182000.0 117300.00000000001 182800.0 ;
      RECT  122300.00000000001 183400.0 121500.0 184200.0 ;
      RECT  119500.0 191600.00000000003 118700.0 192400.0 ;
      RECT  122300.00000000001 190200.0 121500.0 191000.0 ;
      RECT  120900.0 200399.99999999997 120100.00000000001 201200.0 ;
      RECT  122300.00000000001 201800.0 121500.0 202600.00000000003 ;
      RECT  116700.0 210000.0 115900.0 210800.0 ;
      RECT  123700.0 208600.00000000003 122900.0 209399.99999999997 ;
      RECT  118100.0 218800.0 117300.00000000001 219600.00000000003 ;
      RECT  123700.0 220200.0 122900.0 221000.0 ;
      RECT  119500.0 228399.99999999997 118700.0 229200.0 ;
      RECT  123700.0 227000.0 122900.0 227800.0 ;
      RECT  120900.0 237200.0 120100.00000000001 238000.0 ;
      RECT  123700.0 238600.00000000003 122900.0 239399.99999999997 ;
      RECT  116700.0 246800.0 115900.0 247600.00000000003 ;
      RECT  125100.0 245400.00000000003 124300.00000000001 246200.0 ;
      RECT  118100.0 255600.00000000003 117300.00000000001 256400.00000000003 ;
      RECT  125100.0 257000.0 124300.00000000001 257800.0 ;
      RECT  119500.0 265200.0 118700.0 266000.0 ;
      RECT  125100.0 263800.0 124300.00000000001 264600.0 ;
      RECT  120900.0 274000.0 120100.00000000001 274800.0 ;
      RECT  125100.0 275400.00000000006 124300.00000000001 276200.0 ;
      RECT  116700.0 283600.0 115900.0 284400.00000000006 ;
      RECT  126500.0 282200.0 125700.0 283000.0 ;
      RECT  118100.0 292400.00000000006 117300.00000000001 293200.0 ;
      RECT  126500.0 293800.0 125700.0 294600.0 ;
      RECT  119500.0 302000.0 118700.0 302800.0 ;
      RECT  126500.0 300600.0 125700.0 301400.00000000006 ;
      RECT  120900.0 310800.0 120100.00000000001 311600.0 ;
      RECT  126500.0 312200.0 125700.0 313000.0 ;
      RECT  132100.00000000003 177600.00000000003 131300.0 178400.0 ;
      RECT  132100.00000000003 177600.00000000003 131300.0 178400.0 ;
      RECT  132100.00000000003 168400.0 131300.0 169200.0 ;
      RECT  132100.00000000003 168400.0 131300.0 169200.0 ;
      RECT  132100.00000000003 177600.00000000003 131300.0 178400.0 ;
      RECT  132100.00000000003 177600.00000000003 131300.0 178400.0 ;
      RECT  132100.00000000003 186800.0 131300.0 187600.00000000003 ;
      RECT  132100.00000000003 186800.0 131300.0 187600.00000000003 ;
      RECT  132100.00000000003 196000.0 131300.0 196800.0 ;
      RECT  132100.00000000003 196000.0 131300.0 196800.0 ;
      RECT  132100.00000000003 186800.0 131300.0 187600.00000000003 ;
      RECT  132100.00000000003 186800.0 131300.0 187600.00000000003 ;
      RECT  132100.00000000003 196000.0 131300.0 196800.0 ;
      RECT  132100.00000000003 196000.0 131300.0 196800.0 ;
      RECT  132100.00000000003 205200.0 131300.0 206000.0 ;
      RECT  132100.00000000003 205200.0 131300.0 206000.0 ;
      RECT  132100.00000000003 214399.99999999997 131300.0 215200.0 ;
      RECT  132100.00000000003 214399.99999999997 131300.0 215200.0 ;
      RECT  132100.00000000003 205200.0 131300.0 206000.0 ;
      RECT  132100.00000000003 205200.0 131300.0 206000.0 ;
      RECT  132100.00000000003 214399.99999999997 131300.0 215200.0 ;
      RECT  132100.00000000003 214399.99999999997 131300.0 215200.0 ;
      RECT  132100.00000000003 223600.00000000003 131300.0 224399.99999999997 ;
      RECT  132100.00000000003 223600.00000000003 131300.0 224399.99999999997 ;
      RECT  132100.00000000003 232800.0 131300.0 233600.00000000003 ;
      RECT  132100.00000000003 232800.0 131300.0 233600.00000000003 ;
      RECT  132100.00000000003 223600.00000000003 131300.0 224399.99999999997 ;
      RECT  132100.00000000003 223600.00000000003 131300.0 224399.99999999997 ;
      RECT  132100.00000000003 232800.0 131300.0 233600.00000000003 ;
      RECT  132100.00000000003 232800.0 131300.0 233600.00000000003 ;
      RECT  132100.00000000003 242000.0 131300.0 242800.0 ;
      RECT  132100.00000000003 242000.0 131300.0 242800.0 ;
      RECT  132100.00000000003 251200.0 131300.0 252000.0 ;
      RECT  132100.00000000003 251200.0 131300.0 252000.0 ;
      RECT  132100.00000000003 242000.0 131300.0 242800.0 ;
      RECT  132100.00000000003 242000.0 131300.0 242800.0 ;
      RECT  132100.00000000003 251200.0 131300.0 252000.0 ;
      RECT  132100.00000000003 251200.0 131300.0 252000.0 ;
      RECT  132100.00000000003 260400.00000000003 131300.0 261200.0 ;
      RECT  132100.00000000003 260400.00000000003 131300.0 261200.0 ;
      RECT  132100.00000000003 269600.0 131300.0 270400.00000000006 ;
      RECT  132100.00000000003 269600.0 131300.0 270400.00000000006 ;
      RECT  132100.00000000003 260400.00000000003 131300.0 261200.0 ;
      RECT  132100.00000000003 260400.00000000003 131300.0 261200.0 ;
      RECT  132100.00000000003 269600.0 131300.0 270400.00000000006 ;
      RECT  132100.00000000003 269600.0 131300.0 270400.00000000006 ;
      RECT  132100.00000000003 278800.0 131300.0 279600.0 ;
      RECT  132100.00000000003 278800.0 131300.0 279600.0 ;
      RECT  132100.00000000003 288000.0 131300.0 288800.0 ;
      RECT  132100.00000000003 288000.0 131300.0 288800.0 ;
      RECT  132100.00000000003 278800.0 131300.0 279600.0 ;
      RECT  132100.00000000003 278800.0 131300.0 279600.0 ;
      RECT  132100.00000000003 288000.0 131300.0 288800.0 ;
      RECT  132100.00000000003 288000.0 131300.0 288800.0 ;
      RECT  132100.00000000003 297200.0 131300.0 298000.0 ;
      RECT  132100.00000000003 297200.0 131300.0 298000.0 ;
      RECT  132100.00000000003 306400.0 131300.0 307200.0 ;
      RECT  132100.00000000003 306400.0 131300.0 307200.0 ;
      RECT  132100.00000000003 297200.0 131300.0 298000.0 ;
      RECT  132100.00000000003 297200.0 131300.0 298000.0 ;
      RECT  132100.00000000003 306400.0 131300.0 307200.0 ;
      RECT  132100.00000000003 306400.0 131300.0 307200.0 ;
      RECT  132100.00000000003 315600.0 131300.0 316400.00000000006 ;
      RECT  132100.00000000003 315600.0 131300.0 316400.00000000006 ;
      RECT  75100.0 168800.0 75700.0 242400.00000000003 ;
      RECT  76500.0 168800.0 77100.0 242400.00000000003 ;
      RECT  77900.0 168800.0 78500.0 242400.00000000003 ;
      RECT  79300.00000000001 168800.0 79900.0 242400.00000000003 ;
      RECT  148400.0 171900.0 149000.0 172500.0 ;
      RECT  148400.0 171600.00000000003 149000.0 172200.0 ;
      RECT  148700.0 171900.0 153100.0 172500.0 ;
      RECT  148400.0 183500.0 149000.0 184100.00000000003 ;
      RECT  148400.0 183800.0 149000.0 184400.0 ;
      RECT  148700.0 183500.0 153100.0 184100.00000000003 ;
      RECT  148400.0 190300.0 149000.0 190900.0 ;
      RECT  148400.0 190000.0 149000.0 190600.00000000003 ;
      RECT  148700.0 190300.0 153100.0 190900.0 ;
      RECT  148400.0 201899.99999999997 149000.0 202500.0 ;
      RECT  148400.0 202200.0 149000.0 202800.0 ;
      RECT  148700.0 201899.99999999997 153100.0 202500.0 ;
      RECT  148400.0 208700.0 149000.0 209300.0 ;
      RECT  148400.0 208399.99999999997 149000.0 209000.0 ;
      RECT  148700.0 208700.0 153100.0 209300.0 ;
      RECT  148400.0 220300.0 149000.0 220899.99999999997 ;
      RECT  148400.0 220600.00000000003 149000.0 221200.0 ;
      RECT  148700.0 220300.0 153100.0 220899.99999999997 ;
      RECT  148400.0 227100.00000000003 149000.0 227700.0 ;
      RECT  148400.0 226800.0 149000.0 227399.99999999997 ;
      RECT  148700.0 227100.00000000003 153100.0 227700.0 ;
      RECT  148400.0 238700.0 149000.0 239300.0 ;
      RECT  148400.0 239000.0 149000.0 239600.00000000003 ;
      RECT  148700.0 238700.0 153100.0 239300.0 ;
      RECT  148400.0 245500.0 149000.0 246100.00000000003 ;
      RECT  148400.0 245200.0 149000.0 245800.0 ;
      RECT  148700.0 245500.0 153100.0 246100.00000000003 ;
      RECT  148400.0 257100.00000000003 149000.0 257700.0 ;
      RECT  148400.0 257400.00000000003 149000.0 258000.0 ;
      RECT  148700.0 257100.00000000003 153100.0 257700.0 ;
      RECT  148400.0 263900.00000000006 149000.0 264500.0 ;
      RECT  148400.0 263600.0 149000.0 264200.0 ;
      RECT  148700.0 263900.00000000006 153100.0 264500.0 ;
      RECT  148400.0 275500.0 149000.0 276100.0 ;
      RECT  148400.0 275800.0 149000.0 276400.0 ;
      RECT  148700.0 275500.0 153100.0 276100.0 ;
      RECT  148400.0 282300.0 149000.0 282900.0 ;
      RECT  148400.0 282000.0 149000.0 282600.0 ;
      RECT  148700.0 282300.0 153100.0 282900.0 ;
      RECT  148400.0 293900.00000000006 149000.0 294500.0 ;
      RECT  148400.0 294200.0 149000.0 294800.0 ;
      RECT  148700.0 293900.00000000006 153100.0 294500.0 ;
      RECT  148400.0 300700.0 149000.0 301300.0 ;
      RECT  148400.0 300400.0 149000.0 301000.0 ;
      RECT  148700.0 300700.0 153100.0 301300.0 ;
      RECT  148400.0 312300.0 149000.0 312900.0 ;
      RECT  148400.0 312600.0 149000.0 313200.0 ;
      RECT  148700.0 312300.0 153100.0 312900.0 ;
      RECT  155400.0 176000.0 156000.0 176600.00000000003 ;
      RECT  155400.0 170200.0 156000.0 170800.0 ;
      RECT  152700.0 176000.0 155700.0 176600.00000000003 ;
      RECT  155400.0 173600.00000000003 156000.0 176300.0 ;
      RECT  155400.0 170500.0 156000.0 173600.00000000003 ;
      RECT  154300.0 170200.0 155700.0 170800.0 ;
      RECT  152300.0 175900.0 153100.0 176700.0 ;
      RECT  153900.0 170100.00000000003 154700.0 170900.0 ;
      RECT  156100.0 173200.0 155300.0 174000.0 ;
      RECT  155400.0 180000.0 156000.0 179400.0 ;
      RECT  155400.0 185800.0 156000.0 185200.0 ;
      RECT  152700.0 180000.0 155700.0 179400.0 ;
      RECT  155400.0 182400.0 156000.0 179700.0 ;
      RECT  155400.0 185500.0 156000.0 182400.0 ;
      RECT  154300.0 185800.0 155700.0 185200.0 ;
      RECT  152300.0 180100.00000000003 153100.0 179300.0 ;
      RECT  153900.0 185900.0 154700.0 185100.00000000003 ;
      RECT  156100.0 182800.0 155300.0 182000.0 ;
      RECT  155400.0 194400.0 156000.0 195000.0 ;
      RECT  155400.0 188600.00000000003 156000.0 189200.0 ;
      RECT  152700.0 194400.0 155700.0 195000.0 ;
      RECT  155400.0 192000.0 156000.0 194700.0 ;
      RECT  155400.0 188900.0 156000.0 192000.0 ;
      RECT  154300.0 188600.00000000003 155700.0 189200.0 ;
      RECT  152300.0 194300.0 153100.0 195100.00000000003 ;
      RECT  153900.0 188500.0 154700.0 189300.0 ;
      RECT  156100.0 191600.00000000003 155300.0 192400.0 ;
      RECT  155400.0 198400.00000000003 156000.0 197800.0 ;
      RECT  155400.0 204200.0 156000.0 203600.00000000003 ;
      RECT  152700.0 198400.00000000003 155700.0 197800.0 ;
      RECT  155400.0 200800.0 156000.0 198100.00000000003 ;
      RECT  155400.0 203899.99999999997 156000.0 200800.0 ;
      RECT  154300.0 204200.0 155700.0 203600.00000000003 ;
      RECT  152300.0 198500.0 153100.0 197700.0 ;
      RECT  153900.0 204300.0 154700.0 203500.0 ;
      RECT  156100.0 201200.0 155300.0 200399.99999999997 ;
      RECT  155400.0 212800.0 156000.0 213399.99999999997 ;
      RECT  155400.0 207000.0 156000.0 207600.00000000003 ;
      RECT  152700.0 212800.0 155700.0 213399.99999999997 ;
      RECT  155400.0 210399.99999999997 156000.0 213100.00000000003 ;
      RECT  155400.0 207300.0 156000.0 210399.99999999997 ;
      RECT  154300.0 207000.0 155700.0 207600.00000000003 ;
      RECT  152300.0 212700.0 153100.0 213500.0 ;
      RECT  153900.0 206899.99999999997 154700.0 207700.0 ;
      RECT  156100.0 210000.0 155300.0 210800.0 ;
      RECT  155400.0 216800.0 156000.0 216200.0 ;
      RECT  155400.0 222600.00000000003 156000.0 222000.0 ;
      RECT  152700.0 216800.0 155700.0 216200.0 ;
      RECT  155400.0 219200.0 156000.0 216500.0 ;
      RECT  155400.0 222300.0 156000.0 219200.0 ;
      RECT  154300.0 222600.00000000003 155700.0 222000.0 ;
      RECT  152300.0 216899.99999999997 153100.0 216100.00000000003 ;
      RECT  153900.0 222700.0 154700.0 221899.99999999997 ;
      RECT  156100.0 219600.00000000003 155300.0 218800.0 ;
      RECT  155400.0 231200.0 156000.0 231800.0 ;
      RECT  155400.0 225399.99999999997 156000.0 226000.0 ;
      RECT  152700.0 231200.0 155700.0 231800.0 ;
      RECT  155400.0 228800.0 156000.0 231500.0 ;
      RECT  155400.0 225700.0 156000.0 228800.0 ;
      RECT  154300.0 225399.99999999997 155700.0 226000.0 ;
      RECT  152300.0 231100.00000000003 153100.0 231899.99999999997 ;
      RECT  153900.0 225300.0 154700.0 226100.00000000003 ;
      RECT  156100.0 228399.99999999997 155300.0 229200.0 ;
      RECT  155400.0 235200.0 156000.0 234600.00000000003 ;
      RECT  155400.0 241000.0 156000.0 240400.00000000003 ;
      RECT  152700.0 235200.0 155700.0 234600.00000000003 ;
      RECT  155400.0 237600.00000000003 156000.0 234900.00000000003 ;
      RECT  155400.0 240700.0 156000.0 237600.00000000003 ;
      RECT  154300.0 241000.0 155700.0 240400.00000000003 ;
      RECT  152300.0 235300.0 153100.0 234500.0 ;
      RECT  153900.0 241100.00000000003 154700.0 240300.0 ;
      RECT  156100.0 238000.0 155300.0 237200.0 ;
      RECT  155400.0 249600.00000000003 156000.0 250200.0 ;
      RECT  155400.0 243800.0 156000.0 244400.00000000003 ;
      RECT  152700.0 249600.00000000003 155700.0 250200.0 ;
      RECT  155400.0 247200.0 156000.0 249900.00000000003 ;
      RECT  155400.0 244100.00000000003 156000.0 247200.0 ;
      RECT  154300.0 243800.0 155700.0 244400.00000000003 ;
      RECT  152300.0 249500.0 153100.0 250300.0 ;
      RECT  153900.0 243700.0 154700.0 244500.0 ;
      RECT  156100.0 246800.0 155300.0 247600.00000000003 ;
      RECT  155400.0 253600.00000000003 156000.0 253000.0 ;
      RECT  155400.0 259399.99999999997 156000.0 258800.0 ;
      RECT  152700.0 253600.00000000003 155700.0 253000.0 ;
      RECT  155400.0 256000.0 156000.0 253300.0 ;
      RECT  155400.0 259100.00000000003 156000.0 256000.0 ;
      RECT  154300.0 259399.99999999997 155700.0 258800.0 ;
      RECT  152300.0 253700.0 153100.0 252899.99999999997 ;
      RECT  153900.0 259500.0 154700.0 258700.0 ;
      RECT  156100.0 256399.99999999997 155300.0 255600.00000000003 ;
      RECT  155400.0 268000.0 156000.0 268600.0 ;
      RECT  155400.0 262200.0 156000.0 262800.0 ;
      RECT  152700.0 268000.0 155700.0 268600.0 ;
      RECT  155400.0 265600.0 156000.0 268300.0 ;
      RECT  155400.0 262500.0 156000.0 265600.0 ;
      RECT  154300.0 262200.0 155700.0 262800.0 ;
      RECT  152300.0 267900.0 153100.0 268700.0 ;
      RECT  153900.0 262100.00000000003 154700.0 262900.0 ;
      RECT  156100.0 265200.0 155300.0 266000.0 ;
      RECT  155400.0 272000.0 156000.0 271400.00000000006 ;
      RECT  155400.0 277800.0 156000.0 277200.0 ;
      RECT  152700.0 272000.0 155700.0 271400.00000000006 ;
      RECT  155400.0 274400.00000000006 156000.0 271700.0 ;
      RECT  155400.0 277500.0 156000.0 274400.00000000006 ;
      RECT  154300.0 277800.0 155700.0 277200.0 ;
      RECT  152300.0 272100.0 153100.0 271300.0 ;
      RECT  153900.0 277900.00000000006 154700.0 277100.0 ;
      RECT  156100.0 274800.0 155300.0 274000.0 ;
      RECT  155400.0 286400.00000000006 156000.0 287000.0 ;
      RECT  155400.0 280600.0 156000.0 281200.0 ;
      RECT  152700.0 286400.00000000006 155700.0 287000.0 ;
      RECT  155400.0 284000.0 156000.0 286700.0 ;
      RECT  155400.0 280900.00000000006 156000.0 284000.0 ;
      RECT  154300.0 280600.0 155700.0 281200.0 ;
      RECT  152300.0 286300.0 153100.0 287100.0 ;
      RECT  153900.0 280500.0 154700.0 281300.0 ;
      RECT  156100.0 283600.0 155300.0 284400.00000000006 ;
      RECT  155400.0 290400.00000000006 156000.0 289800.0 ;
      RECT  155400.0 296200.0 156000.0 295600.0 ;
      RECT  152700.0 290400.00000000006 155700.0 289800.0 ;
      RECT  155400.0 292800.0 156000.0 290100.0 ;
      RECT  155400.0 295900.00000000006 156000.0 292800.0 ;
      RECT  154300.0 296200.0 155700.0 295600.0 ;
      RECT  152300.0 290500.0 153100.0 289700.0 ;
      RECT  153900.0 296300.0 154700.0 295500.0 ;
      RECT  156100.0 293200.0 155300.0 292400.00000000006 ;
      RECT  155400.0 304800.0 156000.0 305400.00000000006 ;
      RECT  155400.0 299000.0 156000.0 299600.0 ;
      RECT  152700.0 304800.0 155700.0 305400.00000000006 ;
      RECT  155400.0 302400.00000000006 156000.0 305100.0 ;
      RECT  155400.0 299300.0 156000.0 302400.00000000006 ;
      RECT  154300.0 299000.0 155700.0 299600.0 ;
      RECT  152300.0 304700.0 153100.0 305500.0 ;
      RECT  153900.0 298900.00000000006 154700.0 299700.0 ;
      RECT  156100.0 302000.0 155300.0 302800.0 ;
      RECT  155400.0 308800.0 156000.0 308200.0 ;
      RECT  155400.0 314600.0 156000.0 314000.0 ;
      RECT  152700.0 308800.0 155700.0 308200.0 ;
      RECT  155400.0 311200.0 156000.0 308500.0 ;
      RECT  155400.0 314300.0 156000.0 311200.0 ;
      RECT  154300.0 314600.0 155700.0 314000.0 ;
      RECT  152300.0 308900.00000000006 153100.0 308100.0 ;
      RECT  153900.0 314700.0 154700.0 313900.00000000006 ;
      RECT  156100.0 311600.0 155300.0 310800.0 ;
      RECT  147000.0 173200.0 147800.0 174000.0 ;
      RECT  148300.0 171200.0 149100.0 172000.0 ;
      RECT  153100.0 171800.0 152300.0 172600.00000000003 ;
      RECT  147000.0 182000.0 147800.0 182800.0 ;
      RECT  148300.0 184000.0 149100.0 184800.0 ;
      RECT  153100.0 183400.0 152300.0 184200.0 ;
      RECT  147000.0 191600.00000000003 147800.0 192400.0 ;
      RECT  148300.0 189600.00000000003 149100.0 190400.0 ;
      RECT  153100.0 190200.0 152300.0 191000.0 ;
      RECT  147000.0 200399.99999999997 147800.0 201200.0 ;
      RECT  148300.0 202399.99999999997 149100.0 203200.0 ;
      RECT  153100.0 201800.0 152300.0 202600.00000000003 ;
      RECT  147000.0 210000.0 147800.0 210800.0 ;
      RECT  148300.0 208000.0 149100.0 208800.0 ;
      RECT  153100.0 208600.00000000003 152300.0 209399.99999999997 ;
      RECT  147000.0 218800.0 147800.0 219600.00000000003 ;
      RECT  148300.0 220800.0 149100.0 221600.00000000003 ;
      RECT  153100.0 220200.0 152300.0 221000.0 ;
      RECT  147000.0 228399.99999999997 147800.0 229200.0 ;
      RECT  148300.0 226399.99999999997 149100.0 227200.0 ;
      RECT  153100.0 227000.0 152300.0 227800.0 ;
      RECT  147000.0 237200.0 147800.0 238000.0 ;
      RECT  148300.0 239200.0 149100.0 240000.0 ;
      RECT  153100.0 238600.00000000003 152300.0 239399.99999999997 ;
      RECT  147000.0 246800.0 147800.0 247600.00000000003 ;
      RECT  148300.0 244800.0 149100.0 245600.00000000003 ;
      RECT  153100.0 245400.00000000003 152300.0 246200.0 ;
      RECT  147000.0 255600.00000000003 147800.0 256400.00000000003 ;
      RECT  148300.0 257600.00000000003 149100.0 258400.00000000003 ;
      RECT  153100.0 257000.0 152300.0 257800.0 ;
      RECT  147000.0 265200.0 147800.0 266000.0 ;
      RECT  148300.0 263200.0 149100.0 264000.0 ;
      RECT  153100.0 263800.0 152300.0 264600.0 ;
      RECT  147000.0 274000.0 147800.0 274800.0 ;
      RECT  148300.0 276000.0 149100.0 276800.0 ;
      RECT  153100.0 275400.00000000006 152300.0 276200.0 ;
      RECT  147000.0 283600.0 147800.0 284400.00000000006 ;
      RECT  148300.0 281600.0 149100.0 282400.00000000006 ;
      RECT  153100.0 282200.0 152300.0 283000.0 ;
      RECT  147000.0 292400.00000000006 147800.0 293200.0 ;
      RECT  148300.0 294400.00000000006 149100.0 295200.0 ;
      RECT  153100.0 293800.0 152300.0 294600.0 ;
      RECT  147000.0 302000.0 147800.0 302800.0 ;
      RECT  148300.0 300000.0 149100.0 300800.0 ;
      RECT  153100.0 300600.0 152300.0 301400.00000000006 ;
      RECT  147000.0 310800.0 147800.0 311600.0 ;
      RECT  148300.0 312800.0 149100.0 313600.0 ;
      RECT  153100.0 312200.0 152300.0 313000.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 168400.0 158700.0 169200.0 ;
      RECT  159500.0 168400.0 158700.0 169200.0 ;
      RECT  159500.0 168400.0 158700.0 169200.0 ;
      RECT  159500.0 168400.0 158700.0 169200.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 315600.0 158700.0 316400.00000000006 ;
      RECT  159500.0 315600.0 158700.0 316400.00000000006 ;
      RECT  159500.0 315600.0 158700.0 316400.00000000006 ;
      RECT  159500.0 315600.0 158700.0 316400.00000000006 ;
      RECT  147100.0 168800.0 147700.0 316000.0 ;
      RECT  170100.00000000003 154700.0 169300.0 155500.0 ;
      RECT  167300.0 74900.0 166500.0 75700.0 ;
      RECT  168700.0 144500.0 167900.0 145300.0 ;
      RECT  147800.0 164200.0 147000.0 165000.0 ;
      RECT  165900.0 164200.0 165100.00000000003 165000.0 ;
      RECT  172000.0 114800.00000000001 172800.0 117800.00000000001 ;
      RECT  178800.0 114800.00000000001 179600.00000000003 117800.00000000001 ;
      RECT  174400.0 70200.0 175200.0 72200.0 ;
      RECT  181200.0 70200.0 182000.0 72200.0 ;
      RECT  75100.0 168800.0 75700.0 242399.99999999997 ;
      RECT  76500.0 168800.0 77100.0 242399.99999999997 ;
      RECT  77900.0 168800.0 78500.0 242399.99999999997 ;
      RECT  79300.0 168800.0 79900.0 242399.99999999997 ;
      RECT  168000.0 70200.0 168600.00000000003 165600.00000000003 ;
      RECT  169400.0 70200.0 170000.0 165600.00000000003 ;
      RECT  166600.00000000003 70200.0 167200.0 165600.00000000003 ;
      RECT  165200.0 70200.0 165800.0 165600.00000000003 ;
      RECT  36999.99999999999 1400.0000000000057 37599.99999999999 162800.0 ;
      RECT  38399.99999999999 1400.0000000000057 38999.99999999999 162800.0 ;
      RECT  39799.99999999999 1400.0000000000057 40399.99999999999 162800.0 ;
      RECT  41199.99999999999 1400.0000000000057 41800.0 162800.0 ;
      RECT  42599.99999999999 1400.0000000000057 43199.99999999999 162800.0 ;
      RECT  43999.99999999999 1400.0000000000057 44599.99999999999 162800.0 ;
      RECT  43999.99999999999 12400.000000000005 44599.99999999999 82100.00000000001 ;
      RECT  39799.99999999999 30400.000000000007 40399.99999999999 82100.00000000001 ;
      RECT  42599.99999999999 33600.00000000001 43199.99999999999 82100.00000000001 ;
      RECT  5199.999999999992 41400.00000000001 5799.999999999992 44200.0 ;
      RECT  36999.99999999999 72200.0 37599.99999999999 82100.00000000001 ;
      RECT  39799.99999999999 82100.00000000001 40399.99999999999 91000.00000000001 ;
      RECT  36999.99999999999 82100.00000000001 37599.99999999999 116600.00000000001 ;
      RECT  42599.99999999999 82100.00000000001 43199.99999999999 118000.0 ;
      RECT  3999.9999999999914 112200.00000000001 4599.999999999992 170900.0 ;
      RECT  38399.99999999999 82100.00000000001 38999.99999999999 126200.00000000001 ;
      RECT  42599.99999999999 82100.00000000001 43199.99999999999 124800.00000000001 ;
      RECT  11299.999999999993 151800.0 11899.99999999999 166300.0 ;
      RECT  41199.99999999999 10600.000000000007 41800.0 82100.00000000001 ;
      RECT  41199.99999999999 31600.000000000007 41800.0 82100.00000000001 ;
      RECT  43999.99999999999 36600.00000000001 44599.99999999999 82100.00000000001 ;
      RECT  36999.99999999999 32200.000000000004 37599.99999999999 82100.00000000001 ;
      RECT  41199.99999999999 46200.00000000001 41800.0 82100.00000000001 ;
      RECT  43999.99999999999 44800.000000000015 44599.99999999999 82100.00000000003 ;
      RECT  38399.99999999999 50600.00000000001 38999.99999999999 82100.00000000001 ;
      RECT  2399.9999999999914 1400.0000000000057 24199.999999999993 21400.000000000007 ;
      RECT  21199.999999999993 10800.000000000005 21999.999999999993 11600.000000000007 ;
      RECT  25799.999999999993 10600.000000000007 26599.999999999993 11400.000000000007 ;
      RECT  25799.999999999993 10600.000000000007 26599.999999999993 11400.000000000007 ;
      RECT  35199.99999999999 8800.000000000005 35999.99999999999 9600.000000000007 ;
      RECT  29799.999999999993 12000.000000000007 30599.999999999993 12800.000000000007 ;
      RECT  9999.999999999993 10000.000000000005 10799.999999999993 10800.000000000005 ;
      RECT  35299.99999999999 8900.000000000005 35899.99999999999 9500.000000000005 ;
      RECT  29899.999999999993 12100.000000000007 30499.999999999993 12700.000000000007 ;
      RECT  5199.999999999992 8000.000000000007 5999.999999999991 8800.000000000005 ;
      RECT  2399.9999999999914 41400.00000000001 24199.999999999993 21400.000000000007 ;
      RECT  21199.999999999993 32000.000000000007 21999.999999999993 31200.000000000004 ;
      RECT  25799.999999999993 32200.000000000004 26599.999999999993 31400.000000000007 ;
      RECT  25799.999999999993 32200.000000000004 26599.999999999993 31400.000000000007 ;
      RECT  35199.99999999999 34000.00000000001 35999.99999999999 33200.0 ;
      RECT  29799.999999999993 30800.000000000004 30599.999999999993 30000.000000000004 ;
      RECT  9999.999999999993 32800.00000000001 10799.999999999993 32000.000000000007 ;
      RECT  35299.99999999999 33900.00000000001 35899.99999999999 33300.00000000001 ;
      RECT  29899.999999999993 30700.000000000004 30499.999999999993 30100.000000000004 ;
      RECT  5199.999999999992 34800.00000000001 5999.999999999991 34000.00000000001 ;
      RECT  2799.9999999999914 21000.000000000007 1999.9999999999916 21800.000000000007 ;
      RECT  2799.9999999999914 21000.000000000007 1999.9999999999916 21800.000000000007 ;
      RECT  2799.9999999999914 1000.0000000000058 1999.9999999999916 1800.0000000000057 ;
      RECT  2799.9999999999914 1000.0000000000058 1999.9999999999916 1800.0000000000057 ;
      RECT  2799.9999999999914 21000.000000000007 1999.9999999999916 21800.000000000007 ;
      RECT  2799.9999999999914 21000.000000000007 1999.9999999999916 21800.000000000007 ;
      RECT  2799.9999999999914 41000.00000000001 1999.9999999999916 41800.00000000001 ;
      RECT  2799.9999999999914 41000.00000000001 1999.9999999999916 41800.00000000001 ;
      RECT  9999.999999999993 10000.000000000005 10799.999999999993 10800.000000000005 ;
      RECT  9999.999999999993 32000.000000000007 10799.999999999993 32800.000000000015 ;
      RECT  35299.99999999999 8900.000000000005 35899.99999999999 9500.000000000005 ;
      RECT  29899.999999999993 12100.000000000007 30499.999999999993 12700.000000000007 ;
      RECT  35299.99999999999 33300.000000000015 35899.99999999999 33900.00000000001 ;
      RECT  29899.999999999993 30100.000000000007 30499.999999999993 30700.000000000007 ;
      RECT  5199.999999999992 1400.0000000000057 5799.999999999992 41400.00000000001 ;
      RECT  59099.99999999999 23400.000000000007 59699.99999999999 22800.000000000004 ;
      RECT  59099.99999999999 40000.00000000001 59699.99999999999 39400.00000000001 ;
      RECT  56400.0 23400.000000000007 59400.0 22800.000000000004 ;
      RECT  59099.99999999999 36600.00000000001 59699.99999999999 23100.000000000004 ;
      RECT  59099.99999999999 39700.0 59699.99999999999 36600.00000000001 ;
      RECT  58000.0 40000.00000000001 59400.0 39400.00000000001 ;
      RECT  55999.99999999999 23500.000000000004 56800.0 22700.000000000004 ;
      RECT  57599.99999999999 40100.00000000001 58400.0 39300.00000000001 ;
      RECT  59800.0 37000.00000000001 59000.0 36200.0 ;
      RECT  52699.99999999999 59400.00000000001 53300.0 60000.00000000001 ;
      RECT  52699.99999999999 42800.00000000001 53300.0 43400.00000000001 ;
      RECT  50000.0 59400.00000000001 53000.0 60000.00000000001 ;
      RECT  52699.99999999999 46200.0 53300.0 59700.0 ;
      RECT  52699.99999999999 43100.00000000001 53300.0 46200.0 ;
      RECT  51599.99999999999 42800.00000000001 53000.0 43400.00000000001 ;
      RECT  49599.99999999999 59300.000000000015 50400.0 60100.00000000001 ;
      RECT  51199.99999999999 42700.0 52000.0 43500.00000000001 ;
      RECT  53400.0 45800.00000000001 52599.99999999999 46600.00000000001 ;
      RECT  52699.99999999999 103400.0 53300.0 102800.00000000001 ;
      RECT  52699.99999999999 120000.0 53300.0 119400.0 ;
      RECT  50000.0 103400.0 53000.0 102800.00000000001 ;
      RECT  52699.99999999999 116600.00000000001 53300.0 103100.00000000001 ;
      RECT  52699.99999999999 119700.0 53300.0 116600.00000000001 ;
      RECT  51599.99999999999 120000.0 53000.0 119400.0 ;
      RECT  49599.99999999999 103500.0 50400.0 102700.0 ;
      RECT  51199.99999999999 120100.00000000001 52000.0 119300.00000000001 ;
      RECT  53400.0 117000.0 52599.99999999999 116200.0 ;
      RECT  52699.99999999999 139400.0 53300.0 140000.0 ;
      RECT  52699.99999999999 122800.00000000001 53300.0 123400.0 ;
      RECT  50000.0 139400.0 53000.0 140000.0 ;
      RECT  52699.99999999999 126200.0 53300.0 139700.00000000003 ;
      RECT  52699.99999999999 123100.00000000001 53300.0 126200.0 ;
      RECT  51599.99999999999 122800.00000000001 53000.0 123400.0 ;
      RECT  49599.99999999999 139300.0 50400.0 140100.0 ;
      RECT  51199.99999999999 122700.0 52000.0 123500.0 ;
      RECT  53400.0 125800.00000000001 52599.99999999999 126600.00000000001 ;
      RECT  25099.999999999993 173200.00000000003 25699.999999999996 173800.0 ;
      RECT  25099.999999999993 173500.00000000003 25699.999999999996 175500.00000000003 ;
      RECT  19199.999999999993 173200.00000000003 25399.999999999993 173800.0 ;
      RECT  18099.999999999993 164200.00000000003 18699.999999999993 164800.0 ;
      RECT  32099.999999999993 164200.00000000003 32699.999999999996 164800.0 ;
      RECT  18099.999999999993 164500.00000000003 18699.999999999993 171300.0 ;
      RECT  18399.999999999993 164200.00000000003 32399.999999999993 164800.0 ;
      RECT  32099.999999999993 164500.00000000003 32699.999999999996 165900.0 ;
      RECT  5699.999999999992 184400.0 6299.999999999992 185000.00000000003 ;
      RECT  4099.999999999992 184400.0 4699.999999999992 185000.00000000003 ;
      RECT  5699.999999999992 179900.0 6299.999999999992 184700.00000000003 ;
      RECT  4399.999999999992 184400.0 5999.999999999991 185000.00000000003 ;
      RECT  4099.999999999992 184700.00000000003 4699.999999999992 189500.00000000003 ;
      RECT  5699.999999999992 193600.00000000003 6299.999999999992 194200.00000000003 ;
      RECT  4099.999999999992 193600.00000000003 4699.999999999992 194200.00000000003 ;
      RECT  5699.999999999992 189500.00000000003 6299.999999999992 193900.0 ;
      RECT  4399.999999999992 193600.00000000003 5999.999999999991 194200.00000000003 ;
      RECT  4099.999999999992 193900.0 4699.999999999992 198300.00000000003 ;
      RECT  5699.999999999992 202800.0 6299.999999999992 203400.0 ;
      RECT  4099.999999999992 202800.0 4699.999999999992 203400.0 ;
      RECT  5699.999999999992 198300.0 6299.999999999992 203100.00000000003 ;
      RECT  4399.999999999992 202800.0 5999.999999999991 203400.0 ;
      RECT  4099.999999999992 203100.00000000003 4699.999999999992 207900.0 ;
      RECT  25099.999999999993 207600.00000000003 25699.999999999996 208200.00000000003 ;
      RECT  23599.999999999993 207600.00000000003 25399.999999999996 208200.00000000003 ;
      RECT  25099.999999999993 175500.00000000003 25699.999999999996 207900.0 ;
      RECT  10399.99999999999 179500.00000000003 11199.999999999993 180300.0 ;
      RECT  10399.99999999999 179500.00000000003 11199.999999999993 180300.0 ;
      RECT  16799.99999999999 179500.00000000003 17599.999999999993 180300.0 ;
      RECT  16799.99999999999 179500.00000000003 17599.999999999993 180300.0 ;
      RECT  23199.999999999993 179500.00000000003 23999.999999999993 180300.0 ;
      RECT  23199.999999999993 179500.00000000003 23999.999999999993 180300.0 ;
      RECT  3999.9999999999914 179500.00000000003 4799.999999999992 180300.0 ;
      RECT  5599.999999999992 179500.00000000003 6399.999999999992 180300.0 ;
      RECT  5599.999999999992 179500.00000000003 6399.999999999992 180300.0 ;
      RECT  10399.99999999999 189100.00000000003 11199.999999999993 189900.0 ;
      RECT  10399.99999999999 189100.00000000003 11199.999999999993 189900.0 ;
      RECT  16799.99999999999 189100.00000000003 17599.999999999993 189900.0 ;
      RECT  16799.99999999999 189100.00000000003 17599.999999999993 189900.0 ;
      RECT  23199.999999999993 189100.00000000003 23999.999999999993 189900.0 ;
      RECT  23199.999999999993 189100.00000000003 23999.999999999993 189900.0 ;
      RECT  3999.9999999999914 189100.00000000003 4799.999999999992 189900.0 ;
      RECT  5599.999999999992 189100.00000000003 6399.999999999992 189900.0 ;
      RECT  5599.999999999992 189100.00000000003 6399.999999999992 189900.0 ;
      RECT  10399.99999999999 197900.0 11199.999999999993 198700.00000000003 ;
      RECT  10399.99999999999 197900.0 11199.999999999993 198700.00000000003 ;
      RECT  16799.99999999999 197900.0 17599.999999999993 198700.00000000003 ;
      RECT  16799.99999999999 197900.0 17599.999999999993 198700.00000000003 ;
      RECT  23199.999999999993 197900.0 23999.999999999993 198700.00000000003 ;
      RECT  23199.999999999993 197900.0 23999.999999999993 198700.00000000003 ;
      RECT  3999.9999999999914 197900.0 4799.999999999992 198700.00000000003 ;
      RECT  5599.999999999992 197900.0 6399.999999999992 198700.00000000003 ;
      RECT  5599.999999999992 197900.0 6399.999999999992 198700.00000000003 ;
      RECT  10399.99999999999 207500.00000000003 11199.999999999993 208300.0 ;
      RECT  10399.99999999999 207500.00000000003 11199.999999999993 208300.0 ;
      RECT  16799.99999999999 207500.00000000003 17599.999999999993 208300.0 ;
      RECT  16799.99999999999 207500.00000000003 17599.999999999993 208300.0 ;
      RECT  23199.999999999993 207500.00000000003 23999.999999999993 208300.0 ;
      RECT  23199.999999999993 207500.00000000003 23999.999999999993 208300.0 ;
      RECT  3999.9999999999914 207500.00000000003 4799.999999999992 208300.0 ;
      RECT  5599.999999999992 207500.00000000003 6399.999999999992 208300.0 ;
      RECT  5599.999999999992 207500.00000000003 6399.999999999992 208300.0 ;
      RECT  15599.999999999993 184300.0 14799.999999999993 185100.00000000003 ;
      RECT  15599.999999999993 184300.0 14799.999999999993 185100.00000000003 ;
      RECT  15599.999999999993 175100.00000000003 14799.999999999993 175900.0 ;
      RECT  15599.999999999993 175100.00000000003 14799.999999999993 175900.0 ;
      RECT  21999.999999999993 184300.0 21199.999999999993 185100.00000000003 ;
      RECT  21999.999999999993 184300.0 21199.999999999993 185100.00000000003 ;
      RECT  21999.999999999993 175100.00000000003 21199.999999999993 175900.0 ;
      RECT  21999.999999999993 175100.00000000003 21199.999999999993 175900.0 ;
      RECT  15599.999999999993 202700.00000000003 14799.999999999993 203500.00000000003 ;
      RECT  15599.999999999993 202700.00000000003 14799.999999999993 203500.00000000003 ;
      RECT  15599.999999999993 193500.00000000003 14799.999999999993 194300.0 ;
      RECT  15599.999999999993 193500.00000000003 14799.999999999993 194300.0 ;
      RECT  21999.999999999993 202700.00000000003 21199.999999999993 203500.00000000003 ;
      RECT  21999.999999999993 202700.00000000003 21199.999999999993 203500.00000000003 ;
      RECT  21999.999999999993 193500.00000000003 21199.999999999993 194300.0 ;
      RECT  21999.999999999993 193500.00000000003 21199.999999999993 194300.0 ;
      RECT  15599.999999999993 211900.0 14799.999999999993 212700.00000000003 ;
      RECT  15599.999999999993 211900.0 14799.999999999993 212700.00000000003 ;
      RECT  21999.999999999993 211900.0 21199.999999999993 212700.00000000003 ;
      RECT  21999.999999999993 211900.0 21199.999999999993 212700.00000000003 ;
      RECT  3999.9999999999914 179500.00000000003 4799.999999999992 180300.0 ;
      RECT  23199.999999999993 207500.00000000003 23999.999999999993 208300.0 ;
      RECT  3999.9999999999914 175500.00000000003 4599.999999999992 179900.0 ;
      RECT  25099.999999999993 175500.00000000003 25699.999999999993 207900.0 ;
      RECT  30799.999999999993 175500.00000000003 37599.99999999999 166300.0 ;
      RECT  30799.999999999993 175500.00000000003 37599.99999999999 184700.00000000003 ;
      RECT  30799.999999999993 193900.0 37599.99999999999 184700.00000000003 ;
      RECT  30799.999999999993 193900.0 37599.99999999999 203100.00000000003 ;
      RECT  30799.999999999993 212300.00000000003 37599.99999999999 203100.00000000003 ;
      RECT  30799.999999999993 212300.00000000003 37599.99999999999 221500.00000000003 ;
      RECT  30799.999999999993 230700.00000000003 37599.99999999999 221500.00000000003 ;
      RECT  30799.999999999993 230700.00000000003 37599.99999999999 239900.0 ;
      RECT  30799.999999999993 249100.00000000003 37599.99999999999 239900.0 ;
      RECT  33800.0 184300.0 34599.99999999999 185100.00000000003 ;
      RECT  30399.999999999996 179700.00000000003 31199.999999999993 180500.00000000003 ;
      RECT  37199.99999999999 179700.00000000003 37999.99999999999 180500.00000000003 ;
      RECT  33800.0 184300.0 34599.99999999999 185100.00000000003 ;
      RECT  30399.999999999996 188900.0 31199.999999999993 189700.00000000003 ;
      RECT  37199.99999999999 188900.0 37999.99999999999 189700.00000000003 ;
      RECT  33800.0 202700.00000000003 34599.99999999999 203500.00000000003 ;
      RECT  30399.999999999996 198100.00000000003 31199.999999999993 198900.0 ;
      RECT  37199.99999999999 198100.00000000003 37999.99999999999 198900.0 ;
      RECT  33800.0 202700.00000000003 34599.99999999999 203500.00000000003 ;
      RECT  30399.999999999996 207300.0 31199.999999999993 208100.00000000003 ;
      RECT  37199.99999999999 207300.0 37999.99999999999 208100.00000000003 ;
      RECT  33800.0 221100.00000000003 34599.99999999999 221900.0 ;
      RECT  30399.999999999996 216500.00000000003 31199.999999999993 217300.0 ;
      RECT  37199.99999999999 216500.00000000003 37999.99999999999 217300.0 ;
      RECT  33800.0 221100.00000000003 34599.99999999999 221900.0 ;
      RECT  30399.999999999996 225700.00000000003 31199.999999999993 226500.00000000003 ;
      RECT  37199.99999999999 225700.00000000003 37999.99999999999 226500.00000000003 ;
      RECT  33800.0 239500.00000000003 34599.99999999999 240300.0 ;
      RECT  30399.999999999996 234900.0 31199.999999999993 235700.00000000003 ;
      RECT  37199.99999999999 234900.0 37999.99999999999 235700.00000000003 ;
      RECT  33800.0 239500.00000000003 34599.99999999999 240300.0 ;
      RECT  30399.999999999996 244100.00000000003 31199.999999999993 244900.0 ;
      RECT  37199.99999999999 244100.00000000003 37999.99999999999 244900.0 ;
      RECT  31999.999999999993 175100.00000000003 32800.0 250500.00000000003 ;
      RECT  35599.99999999999 175900.0 36399.99999999999 251300.0 ;
      RECT  9199.999999999993 165900.0 8399.99999999999 166700.00000000003 ;
      RECT  9199.999999999993 165900.0 8399.99999999999 166700.00000000003 ;
      RECT  33800.0 165900.0 34599.99999999999 166700.00000000003 ;
      RECT  31199.999999999993 170500.00000000003 30399.999999999993 171300.0 ;
      RECT  31199.999999999993 170500.00000000003 30399.999999999993 171300.0 ;
      RECT  37999.99999999999 170500.00000000003 37199.99999999999 171300.0 ;
      RECT  37999.99999999999 170500.00000000003 37199.99999999999 171300.0 ;
      RECT  40599.99999999999 176500.00000000003 39800.0 177300.0 ;
      RECT  40599.99999999999 176500.00000000003 39800.0 177300.0 ;
      RECT  40599.99999999999 192100.00000000003 39800.0 192900.0 ;
      RECT  40599.99999999999 192100.00000000003 39800.0 192900.0 ;
      RECT  40599.99999999999 194900.0 39800.0 195700.00000000003 ;
      RECT  40599.99999999999 194900.0 39800.0 195700.00000000003 ;
      RECT  40599.99999999999 210500.00000000003 39800.0 211300.0 ;
      RECT  40599.99999999999 210500.00000000003 39800.0 211300.0 ;
      RECT  40599.99999999999 213300.0 39800.0 214100.00000000003 ;
      RECT  40599.99999999999 213300.0 39800.0 214100.00000000003 ;
      RECT  40599.99999999999 228900.0 39800.0 229700.00000000003 ;
      RECT  40599.99999999999 228900.0 39800.0 229700.00000000003 ;
      RECT  40599.99999999999 231700.00000000003 39800.0 232500.00000000003 ;
      RECT  40599.99999999999 231700.00000000003 39800.0 232500.00000000003 ;
      RECT  40599.99999999999 247300.0 39800.0 248100.0 ;
      RECT  40599.99999999999 247300.0 39800.0 248100.0 ;
      RECT  18799.999999999993 173100.00000000003 19599.999999999993 173900.0 ;
      RECT  19599.999999999993 170900.0 20399.999999999996 171700.00000000003 ;
      RECT  19599.999999999993 170900.0 20399.999999999996 171700.00000000003 ;
      RECT  17999.999999999993 170900.0 18799.999999999993 171700.00000000003 ;
      RECT  11199.999999999993 170700.00000000003 11999.999999999993 171500.00000000003 ;
      RECT  3999.9999999999927 166300.0 4599.999999999991 175500.00000000003 ;
      RECT  11299.999999999993 166300.0 11899.99999999999 171100.00000000003 ;
      RECT  44699.99999999999 12000.000000000007 43900.0 12800.000000000007 ;
      RECT  29799.999999999993 12000.000000000007 30599.999999999993 12800.000000000007 ;
      RECT  40499.99999999999 30000.000000000007 39699.99999999999 30800.000000000007 ;
      RECT  29799.999999999993 30000.000000000007 30599.999999999993 30800.000000000007 ;
      RECT  43300.0 33200.0 42500.0 34000.00000000001 ;
      RECT  35199.99999999999 33200.0 35999.99999999999 34000.00000000001 ;
      RECT  5899.999999999992 43800.000000000015 5099.999999999992 44600.00000000001 ;
      RECT  41899.99999999999 43800.000000000015 41099.99999999999 44600.00000000001 ;
      RECT  37699.99999999999 71800.00000000001 36900.0 72600.00000000001 ;
      RECT  40499.99999999999 90600.00000000001 39699.99999999999 91400.0 ;
      RECT  37699.99999999999 116200.00000000001 36900.0 117000.00000000001 ;
      RECT  43300.0 117600.00000000001 42500.0 118400.0 ;
      RECT  4699.999999999992 111800.00000000001 3899.9999999999914 112600.00000000001 ;
      RECT  60399.99999999999 111800.00000000001 59599.99999999999 112600.00000000001 ;
      RECT  60399.99999999999 111800.00000000001 59599.99999999999 112600.00000000001 ;
      RECT  39099.99999999999 125800.00000000001 38300.0 126600.00000000001 ;
      RECT  43300.0 124400.0 42500.0 125200.0 ;
      RECT  11999.999999999993 151400.0 11199.999999999993 152200.00000000003 ;
      RECT  48399.99999999999 10800.000000000005 49199.999999999985 11600.000000000007 ;
      RECT  41899.99999999999 10200.000000000007 41099.99999999999 11000.000000000007 ;
      RECT  56399.99999999999 10200.000000000007 57199.999999999985 11000.000000000007 ;
      RECT  56399.99999999999 10200.000000000007 57199.999999999985 11000.000000000007 ;
      RECT  41899.99999999999 31200.000000000007 41099.99999999999 32000.000000000007 ;
      RECT  44699.99999999999 36200.00000000001 43900.0 37000.00000000001 ;
      RECT  54800.0 36200.00000000001 55599.99999999999 37000.00000000001 ;
      RECT  54800.0 36200.00000000001 55599.99999999999 37000.00000000001 ;
      RECT  37699.99999999999 31800.000000000007 36900.0 32600.000000000007 ;
      RECT  66000.0 31800.000000000007 66800.0 32600.000000000007 ;
      RECT  66000.0 31800.000000000007 66800.0 32600.000000000007 ;
      RECT  41899.99999999999 45800.000000000015 41099.99999999999 46600.00000000001 ;
      RECT  44699.99999999999 44400.00000000001 43900.0 45200.0 ;
      RECT  39099.99999999999 50200.00000000001 38300.0 51000.00000000001 ;
      RECT  59599.99999999999 50200.00000000001 60399.99999999999 51000.00000000001 ;
      RECT  59599.99999999999 50200.00000000001 60399.99999999999 51000.00000000001 ;
      RECT  71199.99999999999 21000.000000000007 70399.99999999999 21800.000000000007 ;
      RECT  71199.99999999999 21000.000000000007 70399.99999999999 21800.000000000007 ;
      RECT  71199.99999999999 1000.0000000000058 70399.99999999999 1800.0000000000057 ;
      RECT  71199.99999999999 1000.0000000000058 70399.99999999999 1800.0000000000057 ;
      RECT  71199.99999999999 21000.000000000007 70399.99999999999 21800.000000000007 ;
      RECT  71199.99999999999 21000.000000000007 70399.99999999999 21800.000000000007 ;
      RECT  71199.99999999999 41000.00000000001 70399.99999999999 41800.00000000001 ;
      RECT  71199.99999999999 41000.00000000001 70399.99999999999 41800.00000000001 ;
      RECT  71199.99999999999 61000.00000000001 70399.99999999999 61800.00000000001 ;
      RECT  71199.99999999999 61000.00000000001 70399.99999999999 61800.00000000001 ;
      RECT  71199.99999999999 41000.00000000001 70399.99999999999 41800.00000000001 ;
      RECT  71199.99999999999 41000.00000000001 70399.99999999999 41800.00000000001 ;
      RECT  71199.99999999999 61000.00000000001 70399.99999999999 61800.00000000001 ;
      RECT  71199.99999999999 61000.00000000001 70399.99999999999 61800.00000000001 ;
      RECT  71199.99999999999 81000.00000000001 70399.99999999999 81800.00000000001 ;
      RECT  71199.99999999999 81000.00000000001 70399.99999999999 81800.00000000001 ;
      RECT  71199.99999999999 101000.00000000001 70399.99999999999 101800.00000000001 ;
      RECT  71199.99999999999 101000.00000000001 70399.99999999999 101800.00000000001 ;
      RECT  71199.99999999999 81000.00000000001 70399.99999999999 81800.00000000001 ;
      RECT  71199.99999999999 81000.00000000001 70399.99999999999 81800.00000000001 ;
      RECT  71199.99999999999 101000.00000000001 70399.99999999999 101800.00000000001 ;
      RECT  71199.99999999999 101000.00000000001 70399.99999999999 101800.00000000001 ;
      RECT  71199.99999999999 121000.00000000001 70399.99999999999 121800.00000000001 ;
      RECT  71199.99999999999 121000.00000000001 70399.99999999999 121800.00000000001 ;
      RECT  71199.99999999999 141000.0 70399.99999999999 141800.0 ;
      RECT  71199.99999999999 141000.0 70399.99999999999 141800.0 ;
      RECT  71199.99999999999 121000.00000000001 70399.99999999999 121800.00000000001 ;
      RECT  71199.99999999999 121000.00000000001 70399.99999999999 121800.00000000001 ;
      RECT  71199.99999999999 141000.0 70399.99999999999 141800.0 ;
      RECT  71199.99999999999 141000.0 70399.99999999999 141800.0 ;
      RECT  71199.99999999999 161000.00000000003 70399.99999999999 161800.00000000003 ;
      RECT  71199.99999999999 161000.00000000003 70399.99999999999 161800.00000000003 ;
      RECT  9999.999999999993 10000.000000000005 10799.999999999993 10800.000000000005 ;
      RECT  9999.999999999993 32000.000000000007 10799.999999999993 32800.000000000015 ;
      RECT  48499.99999999999 1400.0000000000057 49099.99999999999 11200.000000000007 ;
      RECT  53199.99999999999 256100.00000000003 53800.0 336100.0 ;
      RECT  50400.0 256100.00000000003 72200.0 276100.0 ;
      RECT  50400.0 296100.0 72200.0 276100.0 ;
      RECT  50400.0 296100.0 72200.0 316100.0 ;
      RECT  50400.0 336100.0 72200.0 316100.0 ;
      RECT  61700.0 275700.00000000006 60900.0 276500.0 ;
      RECT  61700.0 275700.00000000006 60900.0 276500.0 ;
      RECT  61700.0 255700.00000000003 60900.0 256500.0 ;
      RECT  61700.0 255700.00000000003 60900.0 256500.0 ;
      RECT  61700.0 275700.00000000006 60900.0 276500.0 ;
      RECT  61700.0 275700.00000000006 60900.0 276500.0 ;
      RECT  61700.0 295700.00000000006 60900.0 296500.0 ;
      RECT  61700.0 295700.00000000006 60900.0 296500.0 ;
      RECT  61700.0 315700.00000000006 60900.0 316500.0 ;
      RECT  61700.0 315700.00000000006 60900.0 316500.0 ;
      RECT  61700.0 295700.00000000006 60900.0 296500.0 ;
      RECT  61700.0 295700.00000000006 60900.0 296500.0 ;
      RECT  61700.0 315700.00000000006 60900.0 316500.0 ;
      RECT  61700.0 315700.00000000006 60900.0 316500.0 ;
      RECT  61700.0 335700.00000000006 60900.0 336500.0 ;
      RECT  61700.0 335700.00000000006 60900.0 336500.0 ;
      RECT  53199.99999999999 261100.00000000003 54000.0 261900.00000000003 ;
      RECT  58000.0 264700.00000000006 58800.0 265500.0 ;
      RECT  58000.0 286700.00000000006 58800.0 287500.0 ;
      RECT  58000.0 304700.00000000006 58800.0 305500.0 ;
      RECT  58000.0 326700.00000000006 58800.0 327500.0 ;
      RECT  69200.0 265500.0 70000.0 266300.0 ;
      RECT  69200.0 285900.00000000006 70000.0 286700.00000000006 ;
      RECT  69200.0 305500.0 70000.0 306300.0 ;
      RECT  69200.0 325900.00000000006 70000.0 326700.00000000006 ;
      RECT  174200.00000000003 43200.0 174800.0 63200.0 ;
      RECT  196000.0 43200.0 196600.00000000003 63200.0 ;
      RECT  171400.0 43200.0 193200.00000000003 63200.0 ;
      RECT  193200.00000000003 43200.0 215000.0 63200.0 ;
      RECT  182700.00000000003 62800.00000000001 181900.0 63600.00000000001 ;
      RECT  182700.00000000003 62800.00000000001 181900.0 63600.00000000001 ;
      RECT  182700.00000000003 42800.00000000001 181900.0 43600.0 ;
      RECT  182700.00000000003 42800.00000000001 181900.0 43600.0 ;
      RECT  204500.0 62800.00000000001 203700.00000000003 63600.00000000001 ;
      RECT  204500.0 62800.00000000001 203700.00000000003 63600.00000000001 ;
      RECT  204500.0 42800.00000000001 203700.00000000003 43600.0 ;
      RECT  204500.0 42800.00000000001 203700.00000000003 43600.0 ;
      RECT  174200.00000000003 48200.0 175000.0 49000.0 ;
      RECT  196000.0 48200.0 196800.0 49000.0 ;
      RECT  179000.0 51800.00000000001 179800.0 52600.0 ;
      RECT  200800.0 51800.00000000001 201600.00000000003 52600.0 ;
      RECT  190200.00000000003 52600.0 191000.0 53400.00000000001 ;
      RECT  212000.0 52600.0 212800.0 53400.00000000001 ;
      RECT  74000.0 10200.000000000004 73200.0 11000.000000000004 ;
      RECT  74000.0 261100.00000000003 73200.0 261900.00000000003 ;
      RECT  74000.0 48200.0 73200.0 49000.0 ;
      RECT  168700.0 151800.0 167899.99999999997 152600.00000000003 ;
      RECT  72600.0 151800.0 71800.0 152600.00000000003 ;
      RECT  72600.0 151800.0 71800.0 152600.00000000003 ;
      RECT  167300.0 90200.0 166500.0 91000.0 ;
      RECT  72600.0 90200.0 71800.0 91000.0 ;
      RECT  72600.0 90200.0 71800.0 91000.0 ;
      RECT  170100.00000000003 130199.99999999999 169300.0 131000.0 ;
      RECT  72600.0 130199.99999999999 71800.0 131000.0 ;
      RECT  72600.0 130199.99999999999 71800.0 131000.0 ;
      RECT  165900.0 71800.0 165100.0 72600.0 ;
      RECT  72600.0 71800.0 71800.0 72600.0 ;
      RECT  72600.0 71800.0 71800.0 72600.0 ;
      RECT  75800.0 265500.0 75000.0 266300.0 ;
      RECT  70000.0 265500.0 69200.0 266300.0 ;
      RECT  77200.0 285900.00000000006 76400.0 286700.00000000006 ;
      RECT  70000.0 285900.00000000006 69200.0 286700.00000000006 ;
      RECT  78600.0 305500.0 77800.0 306300.0 ;
      RECT  70000.0 305500.0 69200.0 306300.0 ;
      RECT  80000.0 325900.00000000006 79200.0 326700.00000000006 ;
      RECT  70000.0 325900.00000000006 69200.0 326700.00000000006 ;
      RECT  174400.0 65600.00000000001 175200.00000000003 66400.0 ;
      RECT  190200.0 65600.00000000001 191000.0 66400.0 ;
      RECT  181200.0 67000.0 182000.0 67800.0 ;
      RECT  212000.0 67000.0 212800.0 67800.0 ;
   LAYER  metal3 ;
      RECT  72200.0 261200.0 73600.00000000001 261800.0 ;
      RECT  73600.0 48300.0 193200.0 48900.0 ;
      RECT  72200.0 151900.0 168300.0 152500.0 ;
      RECT  72200.0 90300.00000000001 166900.0 90900.0 ;
      RECT  72200.0 130300.00000000001 169700.0 130900.0 ;
      RECT  72200.0 71900.0 165500.0 72500.0 ;
      RECT  69600.0 265600.0 75399.99999999999 266200.00000000006 ;
      RECT  69600.0 286000.0 76800.0 286600.0 ;
      RECT  69600.0 305600.0 78199.99999999999 306200.00000000006 ;
      RECT  69600.0 326000.0 79600.0 326600.0 ;
      RECT  0.0 19200.000000000004 3600.0 22800.000000000004 ;
      RECT  7200.000000000003 165600.00000000003 10800.000000000002 166800.0 ;
      RECT  14399.999999999998 201600.00000000003 18000.0 205200.00000000003 ;
      RECT  16799.999999999996 182400.0 17999.999999999996 186000.0 ;
      RECT  14399.999999999998 184800.0 18000.0 186000.0 ;
      RECT  14799.999999999996 184300.0 17400.0 185100.00000000003 ;
      RECT  19199.999999999996 170400.0 22799.999999999996 171600.0 ;
      RECT  21599.999999999993 172800.0 22799.999999999993 174000.0 ;
      RECT  19199.999999999996 182400.0 22799.999999999996 186000.0 ;
      RECT  19199.999999999996 201600.00000000003 22799.999999999996 205200.00000000003 ;
      RECT  33599.99999999999 182400.0 34800.0 186000.0 ;
      RECT  33599.99999999999 201600.00000000003 34800.0 205200.00000000003 ;
      RECT  33599.99999999999 220800.0 34800.0 222000.0 ;
      RECT  33599.99999999999 237600.00000000003 34800.0 241200.00000000003 ;
      RECT  33599.99999999999 165600.00000000003 34800.0 166800.0 ;
      RECT  60000.0 273600.0 63600.0 277200.00000000006 ;
      RECT  60000.0 314400.00000000006 63600.0 318000.00000000006 ;
      RECT  69600.0 100800.00000000001 73199.99999999999 102000.00000000001 ;
      RECT  69600.0 19200.000000000004 73199.99999999999 22800.000000000004 ;
      RECT  69600.0 139200.0 73199.99999999999 142799.99999999997 ;
      RECT  69600.0 60000.0 73199.99999999999 63600.0 ;
      RECT  88800.0 230400.00000000003 92399.99999999999 231600.00000000003 ;
      RECT  91200.0 230400.00000000003 92400.0 234000.00000000003 ;
      RECT  90900.0 231000.0 91700.0 233600.0 ;
      RECT  91200.0 175200.0 92400.0 178799.99999999997 ;
      RECT  88800.0 175200.0 92399.99999999999 176399.99999999997 ;
      RECT  90900.0 175800.0 91700.0 178400.0 ;
      RECT  88800.0 213600.00000000003 92399.99999999999 217200.00000000003 ;
      RECT  88800.0 194400.0 92399.99999999999 198000.0 ;
      RECT  108000.0 230400.00000000003 109200.0 234000.00000000003 ;
      RECT  108000.0 194400.0 109200.0 198000.0 ;
      RECT  108000.0 175200.0 109200.0 178799.99999999997 ;
      RECT  108000.0 213600.00000000003 109200.0 217200.00000000003 ;
      RECT  129600.0 213600.00000000003 133200.0 217200.00000000003 ;
      RECT  129600.0 268800.0 133200.0 272400.00000000006 ;
      RECT  129600.0 249600.00000000003 133200.0 253200.00000000003 ;
      RECT  129600.0 230400.00000000003 133200.0 234000.00000000003 ;
      RECT  129600.0 175200.0 133200.0 178799.99999999997 ;
      RECT  129600.0 285600.0 133200.0 289200.00000000006 ;
      RECT  129600.0 194400.0 133200.0 198000.0 ;
      RECT  129600.0 304800.0 133200.0 308400.00000000006 ;
      RECT  158400.0 249600.00000000003 159600.0 253200.00000000003 ;
      RECT  158400.0 213600.00000000003 159600.0 217200.00000000003 ;
      RECT  158400.0 175200.0 159600.0 178799.99999999997 ;
      RECT  158400.0 194400.0 159600.0 198000.0 ;
      RECT  158400.0 230400.00000000003 159600.0 234000.00000000003 ;
      RECT  158400.0 304800.0 159600.0 308400.00000000006 ;
      RECT  158400.0 268800.0 159600.0 272400.00000000006 ;
      RECT  158400.0 285600.0 159600.0 289200.00000000006 ;
      RECT  172800.0 156000.0 176400.0 159600.0 ;
      RECT  172800.0 285600.0 176400.0 289200.00000000006 ;
      RECT  172800.0 194400.0 176400.0 198000.0 ;
      RECT  172800.0 213600.00000000003 176400.0 217200.00000000003 ;
      RECT  172800.0 304800.0 176400.0 308400.00000000006 ;
      RECT  172800.0 268800.0 176400.0 272400.00000000006 ;
      RECT  172800.0 175200.0 176400.0 178799.99999999997 ;
      RECT  172800.0 230400.00000000003 176400.0 234000.00000000003 ;
      RECT  172800.0 249600.00000000003 176400.0 253200.00000000003 ;
      RECT  172800.0 93600.00000000001 176400.0 94800.00000000001 ;
      RECT  172800.0 74400.0 176400.0 78000.0 ;
      RECT  175200.0 127200.0 178799.99999999997 130800.00000000001 ;
      RECT  180000.0 156000.0 183600.0 159600.0 ;
      RECT  180000.0 230400.00000000003 183600.0 234000.00000000003 ;
      RECT  180000.0 285600.0 183600.0 289200.00000000006 ;
      RECT  180000.0 268800.0 183600.0 272400.00000000006 ;
      RECT  180000.0 175200.0 183600.0 178799.99999999997 ;
      RECT  180000.0 249600.00000000003 183600.0 253200.00000000003 ;
      RECT  180000.0 304800.0 183600.0 308400.00000000006 ;
      RECT  180000.0 213600.00000000003 183600.0 217200.00000000003 ;
      RECT  180000.0 194400.0 183600.0 198000.0 ;
      RECT  180000.0 93600.00000000001 183600.0 94800.00000000001 ;
      RECT  180000.0 64800.0 183600.0 66000.0 ;
      RECT  182400.0 62400.00000000001 183600.0 66000.0 ;
      RECT  181900.0 62800.00000000001 182700.00000000003 65400.00000000001 ;
      RECT  180000.0 74400.0 183600.0 78000.0 ;
      RECT  182400.0 127200.0 186000.0 130800.00000000001 ;
      RECT  201600.00000000003 64800.0 205200.00000000003 66000.0 ;
      RECT  204000.0 62400.00000000001 205200.0 66000.0 ;
      RECT  203700.00000000003 62800.00000000001 204500.00000000003 65400.00000000001 ;
      RECT  0.0 40800.0 3600.0 42000.0 ;
      RECT  0.0 0.0 3600.0 3600.0 ;
      RECT  14399.999999999998 192000.0 18000.0 195600.0 ;
      RECT  16799.999999999996 172800.0 17999.999999999996 176400.0 ;
      RECT  14399.999999999998 175200.0 18000.0 176399.99999999997 ;
      RECT  14799.999999999996 175100.00000000003 17400.0 175900.00000000003 ;
      RECT  16799.999999999996 211200.0 17999.999999999996 214799.99999999997 ;
      RECT  14399.999999999998 211200.0 18000.0 212399.99999999997 ;
      RECT  14799.999999999996 211900.00000000003 17400.0 212700.00000000006 ;
      RECT  19199.999999999996 172800.0 20399.999999999996 176400.0 ;
      RECT  19199.999999999996 175200.0 22799.999999999996 176399.99999999997 ;
      RECT  19799.999999999996 175100.00000000003 21999.999999999996 175900.00000000003 ;
      RECT  19199.999999999996 211200.0 22799.999999999996 214799.99999999997 ;
      RECT  19199.999999999996 192000.0 22799.999999999996 195600.0 ;
      RECT  28799.999999999996 170400.0 32400.0 171600.0 ;
      RECT  28799.999999999996 225600.00000000003 32400.0 226800.0 ;
      RECT  28799.999999999996 206400.00000000003 32400.0 210000.00000000003 ;
      RECT  28799.999999999996 177600.00000000003 32400.0 181200.00000000003 ;
      RECT  28799.999999999996 196800.0 32400.0 200400.0 ;
      RECT  28799.999999999996 232800.0 32400.0 236400.0 ;
      RECT  28799.999999999996 216000.0 32400.0 219600.0 ;
      RECT  28799.999999999996 187200.0 32400.0 190799.99999999997 ;
      RECT  28799.999999999996 242400.00000000003 32400.0 246000.00000000003 ;
      RECT  36000.0 242400.00000000003 39600.0 246000.00000000003 ;
      RECT  36000.0 170400.0 39600.0 171600.0 ;
      RECT  36000.0 232800.0 39600.0 236400.0 ;
      RECT  36000.0 216000.0 39600.0 219600.0 ;
      RECT  36000.0 225600.00000000003 39600.0 226800.0 ;
      RECT  36000.0 196800.0 39600.0 200400.0 ;
      RECT  36000.0 206400.00000000003 39600.0 210000.00000000003 ;
      RECT  36000.0 187200.0 39600.0 190799.99999999997 ;
      RECT  36000.0 177600.00000000003 39600.0 181200.00000000003 ;
      RECT  38400.0 230400.00000000003 42000.0 234000.00000000003 ;
      RECT  38400.0 194400.0 42000.0 198000.0 ;
      RECT  38400.0 192000.0 42000.0 193200.0 ;
      RECT  38400.0 211200.0 42000.0 214799.99999999997 ;
      RECT  38400.0 247200.0 42000.0 248399.99999999997 ;
      RECT  38400.0 175200.0 42000.0 178799.99999999997 ;
      RECT  38400.0 208800.0 42000.0 212400.0 ;
      RECT  38400.0 228000.0 42000.0 231600.0 ;
      RECT  60000.0 295200.0 63600.0 298800.0 ;
      RECT  60000.0 254400.00000000003 63600.0 258000.00000000006 ;
      RECT  60000.0 333600.0 63600.0 337200.00000000006 ;
      RECT  69600.0 0.0 73199.99999999999 3600.0 ;
      RECT  69600.0 120000.0 73199.99999999999 123600.0 ;
      RECT  69600.0 40800.0 73199.99999999999 42000.0 ;
      RECT  69600.0 160800.0 73199.99999999999 162000.0 ;
      RECT  69600.0 79200.0 73199.99999999999 82800.0 ;
      RECT  88800.0 170400.0 92399.99999999999 171600.0 ;
      RECT  91200.0 168000.0 92400.0 171600.0 ;
      RECT  90900.0 168400.0 91700.0 171000.0 ;
      RECT  88800.0 225600.00000000003 92399.99999999999 226800.0 ;
      RECT  91200.0 223200.0 92400.0 226799.99999999997 ;
      RECT  90900.0 223600.00000000003 91700.0 226200.00000000003 ;
      RECT  88800.0 240000.0 92399.99999999999 243600.0 ;
      RECT  88800.0 184800.0 92399.99999999999 188400.0 ;
      RECT  88800.0 204000.0 92399.99999999999 207600.0 ;
      RECT  108000.0 184800.0 109200.0 188400.0 ;
      RECT  108000.0 223200.0 109200.0 226799.99999999997 ;
      RECT  108000.0 204000.0 109200.0 207600.0 ;
      RECT  108000.0 240000.0 109200.0 243600.0 ;
      RECT  108000.0 168000.0 109200.0 171600.0 ;
      RECT  129600.0 240000.0 133200.0 243600.0 ;
      RECT  129600.0 314400.00000000006 133200.0 318000.00000000006 ;
      RECT  129600.0 259200.0 133200.0 262800.0 ;
      RECT  129600.0 184800.0 133200.0 188400.0 ;
      RECT  129600.0 295200.0 133200.0 298800.0 ;
      RECT  129600.0 168000.0 133200.0 171600.0 ;
      RECT  129600.0 223200.0 133200.0 226799.99999999997 ;
      RECT  129600.0 278400.00000000006 133200.0 282000.00000000006 ;
      RECT  129600.0 204000.0 133200.0 207600.0 ;
      RECT  158400.0 295200.0 159600.0 298800.0 ;
      RECT  158400.0 240000.0 159600.0 243600.0 ;
      RECT  158400.0 223200.0 159600.0 226799.99999999997 ;
      RECT  158400.0 314400.00000000006 159600.0 318000.00000000006 ;
      RECT  158400.0 168000.0 159600.0 171600.0 ;
      RECT  158400.0 184800.0 159600.0 188400.0 ;
      RECT  158400.0 278400.00000000006 159600.0 282000.00000000006 ;
      RECT  158400.0 204000.0 159600.0 207600.0 ;
      RECT  158400.0 259200.0 159600.0 262800.0 ;
      RECT  170400.0 189600.00000000003 174000.0 193200.00000000003 ;
      RECT  170400.0 235200.0 174000.0 238799.99999999997 ;
      RECT  170400.0 180000.0 174000.0 183600.0 ;
      RECT  170400.0 280800.0 174000.0 284400.00000000006 ;
      RECT  170400.0 170400.0 174000.0 174000.0 ;
      RECT  170400.0 309600.0 174000.0 313200.00000000006 ;
      RECT  170400.0 208800.0 174000.0 212400.0 ;
      RECT  170400.0 244800.0 174000.0 248400.0 ;
      RECT  170400.0 225600.00000000003 174000.0 229200.00000000003 ;
      RECT  170400.0 300000.0 174000.0 303600.0 ;
      RECT  170400.0 273600.0 174000.0 274800.0 ;
      RECT  170400.0 199200.0 174000.0 202799.99999999997 ;
      RECT  170400.0 254400.00000000003 174000.0 258000.00000000006 ;
      RECT  170400.0 218400.00000000003 174000.0 219600.00000000003 ;
      RECT  170400.0 264000.0 174000.0 267600.0 ;
      RECT  170400.0 290400.00000000006 174000.0 294000.00000000006 ;
      RECT  172800.0 81600.00000000001 176400.0 85200.0 ;
      RECT  175200.0 98400.0 178799.99999999997 102000.0 ;
      RECT  175200.0 86400.0 178799.99999999997 90000.0 ;
      RECT  177600.00000000003 235200.0 178800.0 238799.99999999997 ;
      RECT  177600.00000000003 280800.0 178800.0 284400.00000000006 ;
      RECT  177600.00000000003 139200.0 178800.0 142799.99999999997 ;
      RECT  177600.00000000003 189600.00000000003 178800.0 193200.00000000003 ;
      RECT  177600.00000000003 199200.0 178800.0 202799.99999999997 ;
      RECT  177600.00000000003 300000.0 178800.0 303600.0 ;
      RECT  177600.00000000003 218400.00000000003 178800.0 219600.00000000003 ;
      RECT  177600.00000000003 170400.0 178800.0 174000.0 ;
      RECT  177600.00000000003 273600.0 178800.0 274800.0 ;
      RECT  177600.00000000003 208800.0 178800.0 212400.0 ;
      RECT  177600.00000000003 309600.0 178800.0 313200.00000000006 ;
      RECT  177600.00000000003 290400.00000000006 178800.0 294000.00000000006 ;
      RECT  177600.00000000003 180000.0 178800.0 183600.0 ;
      RECT  177600.00000000003 225600.00000000003 178800.0 229200.00000000003 ;
      RECT  177600.00000000003 254400.00000000003 178800.0 258000.00000000006 ;
      RECT  177600.00000000003 264000.0 178800.0 267600.0 ;
      RECT  177600.00000000003 244800.0 178800.0 248400.0 ;
      RECT  180000.0 40800.0 183600.0 44400.0 ;
      RECT  180000.0 81600.00000000001 183600.0 85200.0 ;
      RECT  182400.0 100800.00000000001 183600.0 102000.00000000001 ;
      RECT  182400.0 86400.0 186000.0 90000.0 ;
      RECT  182400.0 244800.0 186000.0 248400.0 ;
      RECT  182400.0 235200.0 186000.0 238799.99999999997 ;
      RECT  182400.0 208800.0 186000.0 212400.0 ;
      RECT  182400.0 290400.00000000006 186000.0 294000.00000000006 ;
      RECT  182400.0 264000.0 186000.0 267600.0 ;
      RECT  182400.0 139200.0 186000.0 142799.99999999997 ;
      RECT  182400.0 280800.0 186000.0 284400.00000000006 ;
      RECT  182400.0 170400.0 186000.0 174000.0 ;
      RECT  182400.0 189600.00000000003 186000.0 193200.00000000003 ;
      RECT  182400.0 180000.0 186000.0 183600.0 ;
      RECT  182400.0 300000.0 186000.0 303600.0 ;
      RECT  182400.0 199200.0 186000.0 202799.99999999997 ;
      RECT  182400.0 225600.00000000003 186000.0 229200.00000000003 ;
      RECT  182400.0 309600.0 186000.0 313200.00000000006 ;
      RECT  182400.0 218400.00000000003 186000.0 219600.00000000003 ;
      RECT  182400.0 273600.0 186000.0 274800.0 ;
      RECT  182400.0 254400.00000000003 186000.0 258000.00000000006 ;
      RECT  201600.00000000003 40800.0 205200.00000000003 44400.0 ;
      RECT  19199.999999999996 170400.0 20399.999999999996 171600.0 ;
      RECT  33599.99999999999 223200.0 34800.0 224399.99999999997 ;
      RECT  33599.99999999999 221400.00000000003 34800.0 223800.00000000003 ;
      RECT  33599.99999999999 220800.0 34800.0 222000.0 ;
      RECT  33599.99999999999 223200.0 34800.0 224399.99999999997 ;
      RECT  72000.0 103200.0 73200.0 104400.0 ;
      RECT  72000.0 101400.0 73200.0 103800.00000000001 ;
      RECT  72000.0 100800.00000000001 73200.0 102000.00000000001 ;
      RECT  72000.0 103200.0 73200.0 104400.0 ;
      RECT  91200.0 213600.00000000003 92400.0 214800.0 ;
      RECT  108000.0 218400.00000000003 109200.0 219600.00000000003 ;
      RECT  108000.0 216600.00000000003 109200.0 219000.00000000003 ;
      RECT  108000.0 216000.0 109200.0 217200.0 ;
      RECT  108000.0 218400.00000000003 109200.0 219600.00000000003 ;
      RECT  2399.9999999999914 43200.0 3599.999999999992 44400.00000000001 ;
      RECT  2399.9999999999914 41400.00000000001 3599.999999999992 43800.00000000001 ;
      RECT  2399.9999999999914 40800.0 3599.999999999992 42000.0 ;
      RECT  2399.9999999999914 43200.0 3599.999999999992 44400.00000000001 ;
      RECT  2399.9999999999914 4799.999999999997 3599.999999999992 5999.999999999997 ;
      RECT  2399.9999999999914 3000.0 3599.999999999992 5400.0 ;
      RECT  2399.9999999999914 2400.0000000000055 3599.999999999992 3600.000000000006 ;
      RECT  2399.9999999999914 4799.999999999997 3599.999999999992 5999.999999999997 ;
      RECT  16799.999999999996 172800.0 17999.999999999996 174000.0 ;
      RECT  21599.999999999993 175200.0 22799.999999999993 176399.99999999997 ;
      RECT  31199.999999999996 172800.0 32400.0 174000.0 ;
      RECT  31199.999999999996 171000.0 32400.0 173400.0 ;
      RECT  31199.999999999996 170400.0 32400.0 171600.0 ;
      RECT  31199.999999999996 172800.0 32400.0 174000.0 ;
      RECT  36000.0 172800.0 37200.0 174000.0 ;
      RECT  36000.0 171000.0 37200.0 173400.0 ;
      RECT  36000.0 170400.0 37200.0 171600.0 ;
      RECT  36000.0 172800.0 37200.0 174000.0 ;
      RECT  40800.0 249600.00000000003 42000.0 250800.0 ;
      RECT  40800.0 247800.0 42000.0 250200.00000000003 ;
      RECT  40800.0 247200.0 42000.0 248399.99999999997 ;
      RECT  40800.0 249600.00000000003 42000.0 250800.0 ;
      RECT  60000.0 331200.0 61200.0 332400.0 ;
      RECT  60000.0 331800.0 61200.0 334200.0 ;
      RECT  60000.0 333600.0 61200.0 334800.0 ;
      RECT  60000.0 331200.0 61200.0 332400.0 ;
      RECT  69600.0 0.0 70800.0 1200.0000000000002 ;
      RECT  69600.0 43200.0 70800.0 44400.00000000001 ;
      RECT  69600.0 41400.00000000001 70800.0 43800.00000000001 ;
      RECT  69600.0 40800.0 70800.0 42000.0 ;
      RECT  69600.0 43200.0 70800.0 44400.00000000001 ;
      RECT  69600.0 163200.0 70800.0 164399.99999999997 ;
      RECT  69600.0 161400.0 70800.0 163800.0 ;
      RECT  69600.0 160800.0 70800.0 162000.0 ;
      RECT  69600.0 163200.0 70800.0 164399.99999999997 ;
      RECT  88800.0 187200.0 90000.0 188399.99999999997 ;
      RECT  108000.0 187200.0 109200.0 188399.99999999997 ;
      RECT  170400.0 220800.0 171600.0 222000.0 ;
      RECT  170400.0 219000.0 171600.0 221400.0 ;
      RECT  170400.0 218400.00000000003 171600.0 219600.00000000003 ;
      RECT  170400.0 220800.0 171600.0 222000.0 ;
      RECT  177600.00000000003 220800.0 178800.0 222000.0 ;
      RECT  177600.00000000003 219000.0 178800.0 221400.0 ;
      RECT  177600.00000000003 218400.00000000003 178800.0 219600.00000000003 ;
      RECT  177600.00000000003 220800.0 178800.0 222000.0 ;
      RECT  184800.0 220800.0 186000.0 222000.0 ;
      RECT  184800.0 219000.0 186000.0 221400.0 ;
      RECT  184800.0 218400.00000000003 186000.0 219600.00000000003 ;
      RECT  184800.0 220800.0 186000.0 222000.0 ;
      RECT  174400.0 177200.0 175200.0 178000.0 ;
      RECT  171000.0 172600.00000000003 171800.0 173400.0 ;
      RECT  177800.0 172600.00000000003 178600.00000000003 173400.0 ;
      RECT  181200.0 177200.0 182000.0 178000.0 ;
      RECT  177800.0 172600.00000000003 178600.00000000003 173400.0 ;
      RECT  184600.00000000003 172600.00000000003 185400.0 173400.0 ;
      RECT  174400.0 177200.0 175200.0 178000.0 ;
      RECT  171000.0 181800.0 171800.0 182600.00000000003 ;
      RECT  177800.0 181800.0 178600.00000000003 182600.00000000003 ;
      RECT  181200.0 177200.0 182000.0 178000.0 ;
      RECT  177800.0 181800.0 178600.00000000003 182600.00000000003 ;
      RECT  184600.00000000003 181800.0 185400.0 182600.00000000003 ;
      RECT  174400.0 195600.00000000003 175200.0 196400.0 ;
      RECT  171000.0 191000.0 171800.0 191800.0 ;
      RECT  177800.0 191000.0 178600.00000000003 191800.0 ;
      RECT  181200.0 195600.00000000003 182000.0 196400.0 ;
      RECT  177800.0 191000.0 178600.00000000003 191800.0 ;
      RECT  184600.00000000003 191000.0 185400.0 191800.0 ;
      RECT  174400.0 195600.00000000003 175200.0 196400.0 ;
      RECT  171000.0 200200.0 171800.0 201000.0 ;
      RECT  177800.0 200200.0 178600.00000000003 201000.0 ;
      RECT  181200.0 195600.00000000003 182000.0 196400.0 ;
      RECT  177800.0 200200.0 178600.00000000003 201000.0 ;
      RECT  184600.00000000003 200200.0 185400.0 201000.0 ;
      RECT  174400.0 214000.0 175200.0 214800.0 ;
      RECT  171000.0 209399.99999999997 171800.0 210200.0 ;
      RECT  177800.0 209399.99999999997 178600.00000000003 210200.0 ;
      RECT  181200.0 214000.0 182000.0 214800.0 ;
      RECT  177800.0 209399.99999999997 178600.00000000003 210200.0 ;
      RECT  184600.00000000003 209399.99999999997 185400.0 210200.0 ;
      RECT  174400.0 214000.0 175200.0 214800.0 ;
      RECT  171000.0 218600.00000000003 171800.0 219399.99999999997 ;
      RECT  177800.0 218600.00000000003 178600.00000000003 219399.99999999997 ;
      RECT  181200.0 214000.0 182000.0 214800.0 ;
      RECT  177800.0 218600.00000000003 178600.00000000003 219399.99999999997 ;
      RECT  184600.00000000003 218600.00000000003 185400.0 219399.99999999997 ;
      RECT  174400.0 232399.99999999997 175200.0 233200.0 ;
      RECT  171000.0 227800.0 171800.0 228600.00000000003 ;
      RECT  177800.0 227800.0 178600.00000000003 228600.00000000003 ;
      RECT  181200.0 232399.99999999997 182000.0 233200.0 ;
      RECT  177800.0 227800.0 178600.00000000003 228600.00000000003 ;
      RECT  184600.00000000003 227800.0 185400.0 228600.00000000003 ;
      RECT  174400.0 232399.99999999997 175200.0 233200.0 ;
      RECT  171000.0 237000.0 171800.0 237800.0 ;
      RECT  177800.0 237000.0 178600.00000000003 237800.0 ;
      RECT  181200.0 232399.99999999997 182000.0 233200.0 ;
      RECT  177800.0 237000.0 178600.00000000003 237800.0 ;
      RECT  184600.00000000003 237000.0 185400.0 237800.0 ;
      RECT  174400.0 250800.0 175200.0 251600.00000000003 ;
      RECT  171000.0 246200.0 171800.0 247000.0 ;
      RECT  177800.0 246200.0 178600.00000000003 247000.0 ;
      RECT  181200.0 250800.0 182000.0 251600.00000000003 ;
      RECT  177800.0 246200.0 178600.00000000003 247000.0 ;
      RECT  184600.00000000003 246200.0 185400.0 247000.0 ;
      RECT  174400.0 250800.0 175200.0 251600.00000000003 ;
      RECT  171000.0 255399.99999999997 171800.0 256200.0 ;
      RECT  177800.0 255399.99999999997 178600.00000000003 256200.0 ;
      RECT  181200.0 250800.0 182000.0 251600.00000000003 ;
      RECT  177800.0 255399.99999999997 178600.00000000003 256200.0 ;
      RECT  184600.00000000003 255399.99999999997 185400.0 256200.0 ;
      RECT  174400.0 269200.0 175200.0 270000.0 ;
      RECT  171000.0 264600.0 171800.0 265400.0 ;
      RECT  177800.0 264600.0 178600.00000000003 265400.0 ;
      RECT  181200.0 269200.0 182000.0 270000.0 ;
      RECT  177800.0 264600.0 178600.00000000003 265400.0 ;
      RECT  184600.00000000003 264600.0 185400.0 265400.0 ;
      RECT  174400.0 269200.0 175200.0 270000.0 ;
      RECT  171000.0 273800.0 171800.0 274600.0 ;
      RECT  177800.0 273800.0 178600.00000000003 274600.0 ;
      RECT  181200.0 269200.0 182000.0 270000.0 ;
      RECT  177800.0 273800.0 178600.00000000003 274600.0 ;
      RECT  184600.00000000003 273800.0 185400.0 274600.0 ;
      RECT  174400.0 287600.0 175200.0 288400.0 ;
      RECT  171000.0 283000.0 171800.0 283800.0 ;
      RECT  177800.0 283000.0 178600.00000000003 283800.0 ;
      RECT  181200.0 287600.0 182000.0 288400.0 ;
      RECT  177800.0 283000.0 178600.00000000003 283800.0 ;
      RECT  184600.00000000003 283000.0 185400.0 283800.0 ;
      RECT  174400.0 287600.0 175200.0 288400.0 ;
      RECT  171000.0 292200.0 171800.0 293000.0 ;
      RECT  177800.0 292200.0 178600.00000000003 293000.0 ;
      RECT  181200.0 287600.0 182000.0 288400.0 ;
      RECT  177800.0 292200.0 178600.00000000003 293000.0 ;
      RECT  184600.00000000003 292200.0 185400.0 293000.0 ;
      RECT  174400.0 306000.0 175200.0 306800.0 ;
      RECT  171000.0 301400.0 171800.0 302200.0 ;
      RECT  177800.0 301400.0 178600.00000000003 302200.0 ;
      RECT  181200.0 306000.0 182000.0 306800.0 ;
      RECT  177800.0 301400.0 178600.00000000003 302200.0 ;
      RECT  184600.00000000003 301400.0 185400.0 302200.0 ;
      RECT  174400.0 306000.0 175200.0 306800.0 ;
      RECT  171000.0 310600.0 171800.0 311400.00000000006 ;
      RECT  177800.0 310600.0 178600.00000000003 311400.00000000006 ;
      RECT  181200.0 306000.0 182000.0 306800.0 ;
      RECT  177800.0 310600.0 178600.00000000003 311400.00000000006 ;
      RECT  184600.00000000003 310600.0 185400.0 311400.00000000006 ;
      RECT  174400.0 177200.0 175200.0 178000.0 ;
      RECT  181200.0 177200.0 182000.0 178000.0 ;
      RECT  174400.0 195600.00000000003 175200.0 196400.0 ;
      RECT  181200.0 195600.00000000003 182000.0 196400.0 ;
      RECT  174400.0 214000.0 175200.0 214800.0 ;
      RECT  181200.0 214000.0 182000.0 214800.0 ;
      RECT  174400.0 232399.99999999997 175200.0 233200.0 ;
      RECT  181200.0 232399.99999999997 182000.0 233200.0 ;
      RECT  174400.0 250800.0 175200.0 251600.00000000003 ;
      RECT  181200.0 250800.0 182000.0 251600.00000000003 ;
      RECT  174400.0 269200.0 175200.0 270000.0 ;
      RECT  181200.0 269200.0 182000.0 270000.0 ;
      RECT  174400.0 287600.0 175200.0 288400.0 ;
      RECT  181200.0 287600.0 182000.0 288400.0 ;
      RECT  174400.0 306000.0 175200.0 306800.0 ;
      RECT  181200.0 306000.0 182000.0 306800.0 ;
      RECT  171000.0 172600.00000000003 171800.0 173400.0 ;
      RECT  177800.0 172600.00000000003 178600.00000000003 173400.0 ;
      RECT  184600.00000000003 172600.00000000003 185400.0 173400.0 ;
      RECT  171000.0 181800.0 171800.0 182600.00000000003 ;
      RECT  177800.0 181800.0 178600.00000000003 182600.00000000003 ;
      RECT  184600.00000000003 181800.0 185400.0 182600.00000000003 ;
      RECT  171000.0 191000.0 171800.0 191800.0 ;
      RECT  177800.0 191000.0 178600.00000000003 191800.0 ;
      RECT  184600.00000000003 191000.0 185400.0 191800.0 ;
      RECT  171000.0 200200.0 171800.0 201000.0 ;
      RECT  177800.0 200200.0 178600.00000000003 201000.0 ;
      RECT  184600.00000000003 200200.0 185400.0 201000.0 ;
      RECT  171000.0 209399.99999999997 171800.0 210200.0 ;
      RECT  177800.0 209399.99999999997 178600.00000000003 210200.0 ;
      RECT  184600.00000000003 209399.99999999997 185400.0 210200.0 ;
      RECT  171000.0 218600.00000000003 171800.0 219399.99999999997 ;
      RECT  177800.0 218600.00000000003 178600.00000000003 219399.99999999997 ;
      RECT  184600.00000000003 218600.00000000003 185400.0 219399.99999999997 ;
      RECT  171000.0 227800.0 171800.0 228600.00000000003 ;
      RECT  177800.0 227800.0 178600.00000000003 228600.00000000003 ;
      RECT  184600.00000000003 227800.0 185400.0 228600.00000000003 ;
      RECT  171000.0 237000.0 171800.0 237800.0 ;
      RECT  177800.0 237000.0 178600.00000000003 237800.0 ;
      RECT  184600.00000000003 237000.0 185400.0 237800.0 ;
      RECT  171000.0 246200.0 171800.0 247000.0 ;
      RECT  177800.0 246200.0 178600.00000000003 247000.0 ;
      RECT  184600.00000000003 246200.0 185400.0 247000.0 ;
      RECT  171000.0 255399.99999999997 171800.0 256200.0 ;
      RECT  177800.0 255399.99999999997 178600.00000000003 256200.0 ;
      RECT  184600.00000000003 255399.99999999997 185400.0 256200.0 ;
      RECT  171000.0 264600.0 171800.0 265400.0 ;
      RECT  177800.0 264600.0 178600.00000000003 265400.0 ;
      RECT  184600.00000000003 264600.0 185400.0 265400.0 ;
      RECT  171000.0 273800.0 171800.0 274600.0 ;
      RECT  177800.0 273800.0 178600.00000000003 274600.0 ;
      RECT  184600.00000000003 273800.0 185400.0 274600.0 ;
      RECT  171000.0 283000.0 171800.0 283800.0 ;
      RECT  177800.0 283000.0 178600.00000000003 283800.0 ;
      RECT  184600.00000000003 283000.0 185400.0 283800.0 ;
      RECT  171000.0 292200.0 171800.0 293000.0 ;
      RECT  177800.0 292200.0 178600.00000000003 293000.0 ;
      RECT  184600.00000000003 292200.0 185400.0 293000.0 ;
      RECT  171000.0 301400.0 171800.0 302200.0 ;
      RECT  177800.0 301400.0 178600.00000000003 302200.0 ;
      RECT  184600.00000000003 301400.0 185400.0 302200.0 ;
      RECT  171000.0 310600.0 171800.0 311400.0 ;
      RECT  177800.0 310600.0 178600.00000000003 311400.0 ;
      RECT  184600.00000000003 310600.0 185400.0 311400.0 ;
      RECT  174200.0 158000.0 175000.0 158800.0 ;
      RECT  174200.0 158000.0 175000.0 158800.0 ;
      RECT  181000.0 158000.0 181800.0 158800.0 ;
      RECT  181000.0 158000.0 181800.0 158800.0 ;
      RECT  174200.0 158000.0 175000.0 158800.0 ;
      RECT  181000.0 158000.0 181800.0 158800.0 ;
      RECT  177800.0 141000.0 178600.00000000003 141800.0 ;
      RECT  176800.0 127600.00000000001 177600.00000000003 128400.0 ;
      RECT  184600.00000000003 141000.0 185400.0 141800.0 ;
      RECT  183600.00000000003 127600.00000000001 184400.0 128400.0 ;
      RECT  176900.0 127700.0 177500.0 128300.00000000001 ;
      RECT  183700.0 127700.0 184300.0 128300.00000000001 ;
      RECT  177900.0 141100.00000000003 178500.0 141700.0 ;
      RECT  184700.0 141100.00000000003 185300.0 141700.0 ;
      RECT  175200.0 76400.0 176000.0 77200.0 ;
      RECT  174600.00000000003 93800.00000000001 175400.0 94600.00000000001 ;
      RECT  175200.0 83000.0 176000.0 83800.00000000001 ;
      RECT  176600.00000000003 87400.0 177400.0 88200.0 ;
      RECT  176000.0 100800.00000000001 176800.0 101600.00000000001 ;
      RECT  182000.0 76400.0 182800.0 77200.0 ;
      RECT  181400.0 93800.00000000001 182200.0 94600.00000000001 ;
      RECT  182000.0 83000.0 182800.0 83800.00000000001 ;
      RECT  183400.0 87400.0 184200.0 88200.0 ;
      RECT  182800.0 100800.00000000001 183600.00000000003 101600.00000000001 ;
      RECT  175300.0 76500.0 175900.0 77100.00000000001 ;
      RECT  174700.0 93900.0 175300.0 94500.0 ;
      RECT  182100.00000000003 76500.0 182700.0 77100.00000000001 ;
      RECT  181500.0 93900.0 182100.00000000003 94500.0 ;
      RECT  175300.0 83100.00000000001 175900.0 83700.0 ;
      RECT  176700.0 87500.0 177300.0 88100.00000000001 ;
      RECT  176100.00000000003 100900.0 176700.0 101500.0 ;
      RECT  182100.00000000003 83100.00000000001 182700.0 83700.0 ;
      RECT  183500.0 87500.0 184100.00000000003 88100.00000000001 ;
      RECT  182900.0 100900.0 183500.0 101500.0 ;
      RECT  75400.0 178900.0 82700.0 179500.0 ;
      RECT  76800.0 188100.00000000003 84100.0 188700.0 ;
      RECT  78200.0 215700.0 82700.0 216300.0 ;
      RECT  79600.0 224899.99999999997 84100.0 225500.0 ;
      RECT  112900.0 177500.0 116300.00000000001 178100.00000000003 ;
      RECT  112900.0 187100.00000000003 117700.0 187700.0 ;
      RECT  112900.0 195900.0 119100.00000000001 196500.0 ;
      RECT  112900.0 205500.0 120500.0 206100.00000000003 ;
      RECT  112900.0 214300.0 121900.0 214899.99999999997 ;
      RECT  112900.0 223899.99999999997 123300.00000000001 224500.0 ;
      RECT  112900.0 232700.0 124700.0 233300.0 ;
      RECT  112900.0 242300.0 126100.00000000001 242899.99999999997 ;
      RECT  91700.0 177600.00000000003 90900.0 178400.0 ;
      RECT  109100.0 177600.00000000003 108300.0 178400.0 ;
      RECT  91700.0 168400.0 90900.0 169200.0 ;
      RECT  109100.0 168400.0 108300.0 169200.0 ;
      RECT  91700.0 177600.00000000003 90900.0 178400.0 ;
      RECT  109100.0 177600.00000000003 108300.0 178400.0 ;
      RECT  91700.0 186800.0 90900.0 187600.00000000003 ;
      RECT  109100.0 186800.0 108300.0 187600.00000000003 ;
      RECT  91700.0 196000.0 90900.0 196800.0 ;
      RECT  109100.0 196000.0 108300.0 196800.0 ;
      RECT  91700.0 186800.0 90900.0 187600.00000000003 ;
      RECT  109100.0 186800.0 108300.0 187600.00000000003 ;
      RECT  91700.0 196000.0 90900.0 196800.0 ;
      RECT  109100.0 196000.0 108300.0 196800.0 ;
      RECT  91700.0 205200.0 90900.0 206000.0 ;
      RECT  109100.0 205200.0 108300.0 206000.0 ;
      RECT  90900.0 177600.00000000003 91700.0 178400.0 ;
      RECT  108300.00000000001 177600.00000000003 109100.0 178400.0 ;
      RECT  90900.0 196000.0 91700.0 196800.0 ;
      RECT  108300.00000000001 196000.0 109100.0 196800.0 ;
      RECT  90900.0 168400.0 91700.0 169200.0 ;
      RECT  108300.00000000001 168400.0 109100.0 169200.0 ;
      RECT  90900.0 186800.0 91700.0 187600.00000000003 ;
      RECT  108300.00000000001 186800.0 109100.0 187600.00000000003 ;
      RECT  90900.0 205200.0 91700.0 206000.0 ;
      RECT  108300.00000000001 205200.0 109100.0 206000.0 ;
      RECT  91700.0 214399.99999999997 90900.0 215200.0 ;
      RECT  109100.0 214399.99999999997 108300.0 215200.0 ;
      RECT  91700.0 205200.0 90900.0 206000.0 ;
      RECT  109100.0 205200.0 108300.0 206000.0 ;
      RECT  91700.0 214399.99999999997 90900.0 215200.0 ;
      RECT  109100.0 214399.99999999997 108300.0 215200.0 ;
      RECT  91700.0 223600.00000000003 90900.0 224399.99999999997 ;
      RECT  109100.0 223600.00000000003 108300.0 224399.99999999997 ;
      RECT  91700.0 232800.0 90900.0 233600.00000000003 ;
      RECT  109100.0 232800.0 108300.0 233600.00000000003 ;
      RECT  91700.0 223600.00000000003 90900.0 224399.99999999997 ;
      RECT  109100.0 223600.00000000003 108300.0 224399.99999999997 ;
      RECT  91700.0 232800.0 90900.0 233600.00000000003 ;
      RECT  109100.0 232800.0 108300.0 233600.00000000003 ;
      RECT  91700.0 242000.0 90900.0 242800.0 ;
      RECT  109100.0 242000.0 108300.0 242800.0 ;
      RECT  90900.0 214399.99999999997 91700.0 215200.0 ;
      RECT  108300.00000000001 214399.99999999997 109100.0 215200.0 ;
      RECT  90900.0 232800.0 91700.0 233600.00000000003 ;
      RECT  108300.00000000001 232800.0 109100.0 233600.00000000003 ;
      RECT  90900.0 205200.0 91700.0 206000.0 ;
      RECT  108300.00000000001 205200.0 109100.0 206000.0 ;
      RECT  90900.0 223600.00000000003 91700.0 224399.99999999997 ;
      RECT  108300.00000000001 223600.00000000003 109100.0 224399.99999999997 ;
      RECT  90900.0 242000.0 91700.0 242800.0 ;
      RECT  108300.00000000001 242000.0 109100.0 242800.0 ;
      RECT  83100.0 178800.0 82300.0 179600.00000000003 ;
      RECT  75800.0 178800.0 75000.0 179600.00000000003 ;
      RECT  84500.0 188000.0 83700.0 188800.0 ;
      RECT  77200.0 188000.0 76400.0 188800.0 ;
      RECT  83100.0 215600.00000000003 82300.0 216399.99999999997 ;
      RECT  78600.0 215600.00000000003 77800.0 216399.99999999997 ;
      RECT  84500.0 224800.0 83700.0 225600.00000000003 ;
      RECT  80000.0 224800.0 79200.0 225600.00000000003 ;
      RECT  113300.00000000001 177400.0 112500.0 178200.0 ;
      RECT  116700.0 177400.0 115900.0 178200.0 ;
      RECT  113300.00000000001 187000.0 112500.0 187800.0 ;
      RECT  118100.0 187000.0 117300.00000000001 187800.0 ;
      RECT  113300.00000000001 195800.0 112500.0 196600.00000000003 ;
      RECT  119500.0 195800.0 118700.0 196600.00000000003 ;
      RECT  113300.00000000001 205399.99999999997 112500.0 206200.0 ;
      RECT  120900.0 205399.99999999997 120100.00000000001 206200.0 ;
      RECT  113300.00000000001 214200.0 112500.0 215000.0 ;
      RECT  122300.00000000001 214200.0 121500.0 215000.0 ;
      RECT  113300.00000000001 223800.0 112500.0 224600.00000000003 ;
      RECT  123700.0 223800.0 122900.0 224600.00000000003 ;
      RECT  113300.00000000001 232600.00000000003 112500.0 233399.99999999997 ;
      RECT  125100.0 232600.00000000003 124300.00000000001 233399.99999999997 ;
      RECT  113300.00000000001 242200.0 112500.0 243000.0 ;
      RECT  126500.0 242200.0 125700.0 243000.0 ;
      RECT  132100.00000000003 177600.00000000003 131300.0 178400.0 ;
      RECT  132100.00000000003 168400.0 131300.0 169200.0 ;
      RECT  132100.00000000003 177600.00000000003 131300.0 178400.0 ;
      RECT  132100.00000000003 186800.0 131300.0 187600.00000000003 ;
      RECT  132100.00000000003 196000.0 131300.0 196800.0 ;
      RECT  132100.00000000003 186800.0 131300.0 187600.00000000003 ;
      RECT  132100.00000000003 196000.0 131300.0 196800.0 ;
      RECT  132100.00000000003 205200.0 131300.0 206000.0 ;
      RECT  132100.00000000003 214399.99999999997 131300.0 215200.0 ;
      RECT  132100.00000000003 205200.0 131300.0 206000.0 ;
      RECT  132100.00000000003 214399.99999999997 131300.0 215200.0 ;
      RECT  132100.00000000003 223600.00000000003 131300.0 224399.99999999997 ;
      RECT  132100.00000000003 232800.0 131300.0 233600.00000000003 ;
      RECT  132100.00000000003 223600.00000000003 131300.0 224399.99999999997 ;
      RECT  132100.00000000003 232800.0 131300.0 233600.00000000003 ;
      RECT  132100.00000000003 242000.0 131300.0 242800.0 ;
      RECT  132100.00000000003 251200.0 131300.0 252000.0 ;
      RECT  132100.00000000003 242000.0 131300.0 242800.0 ;
      RECT  132100.00000000003 251200.0 131300.0 252000.0 ;
      RECT  132100.00000000003 260400.00000000003 131300.0 261200.0 ;
      RECT  132100.00000000003 269600.0 131300.0 270400.00000000006 ;
      RECT  132100.00000000003 260400.00000000003 131300.0 261200.0 ;
      RECT  132100.00000000003 269600.0 131300.0 270400.00000000006 ;
      RECT  132100.00000000003 278800.0 131300.0 279600.0 ;
      RECT  132100.00000000003 288000.0 131300.0 288800.0 ;
      RECT  132100.00000000003 278800.0 131300.0 279600.0 ;
      RECT  132100.00000000003 288000.0 131300.0 288800.0 ;
      RECT  132100.00000000003 297200.0 131300.0 298000.0 ;
      RECT  132100.00000000003 306400.0 131300.0 307200.0 ;
      RECT  132100.00000000003 297200.0 131300.0 298000.0 ;
      RECT  132100.00000000003 306400.0 131300.0 307200.0 ;
      RECT  132100.00000000003 315600.0 131300.0 316400.00000000006 ;
      RECT  131300.0 177600.00000000003 132100.00000000003 178400.0 ;
      RECT  131300.0 196000.0 132100.00000000003 196800.0 ;
      RECT  131300.0 214399.99999999997 132100.00000000003 215200.0 ;
      RECT  131300.0 232800.0 132100.00000000003 233600.00000000003 ;
      RECT  131300.0 251200.0 132100.00000000003 252000.0 ;
      RECT  131300.0 269600.0 132100.00000000003 270400.00000000006 ;
      RECT  131300.0 288000.0 132100.00000000003 288800.0 ;
      RECT  131300.0 306400.0 132100.00000000003 307200.0 ;
      RECT  90900.0 177600.00000000003 91700.0 178400.0 ;
      RECT  108300.00000000001 177600.00000000003 109100.0 178400.0 ;
      RECT  90900.0 196000.0 91700.0 196800.0 ;
      RECT  108300.00000000001 196000.0 109100.0 196800.0 ;
      RECT  90900.0 214399.99999999997 91700.0 215200.0 ;
      RECT  108300.00000000001 214399.99999999997 109100.0 215200.0 ;
      RECT  90900.0 232800.0 91700.0 233600.00000000003 ;
      RECT  108300.00000000001 232800.0 109100.0 233600.00000000003 ;
      RECT  131300.0 168400.0 132100.00000000003 169200.0 ;
      RECT  131300.0 186800.0 132100.00000000003 187600.00000000003 ;
      RECT  131300.0 205200.0 132100.00000000003 206000.0 ;
      RECT  131300.0 223600.00000000003 132100.00000000003 224399.99999999997 ;
      RECT  131300.0 242000.0 132100.00000000003 242800.0 ;
      RECT  131300.0 260400.00000000003 132100.00000000003 261200.0 ;
      RECT  131300.0 278800.0 132100.00000000003 279600.0 ;
      RECT  131300.0 297200.0 132100.00000000003 298000.0 ;
      RECT  131300.0 315600.0 132100.00000000003 316400.0 ;
      RECT  90900.0 168400.0 91700.0 169200.0 ;
      RECT  108300.00000000001 168400.0 109100.0 169200.0 ;
      RECT  90900.0 186800.0 91700.0 187600.00000000003 ;
      RECT  108300.00000000001 186800.0 109100.0 187600.00000000003 ;
      RECT  90900.0 205200.0 91700.0 206000.0 ;
      RECT  108300.00000000001 205200.0 109100.0 206000.0 ;
      RECT  90900.0 223600.00000000003 91700.0 224399.99999999997 ;
      RECT  108300.00000000001 223600.00000000003 109100.0 224399.99999999997 ;
      RECT  90900.0 242000.0 91700.0 242800.0 ;
      RECT  108300.00000000001 242000.0 109100.0 242800.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 168400.0 158700.0 169200.0 ;
      RECT  159500.0 168400.0 158700.0 169200.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 177600.00000000003 158700.0 178400.0 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 186800.0 158700.0 187600.00000000003 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 196000.0 158700.0 196800.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 205200.0 158700.0 206000.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 214399.99999999997 158700.0 215200.0 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 223600.00000000003 158700.0 224399.99999999997 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 232800.0 158700.0 233600.00000000003 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 242000.0 158700.0 242800.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 251200.0 158700.0 252000.0 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 260400.00000000003 158700.0 261200.0 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 269600.0 158700.0 270400.00000000006 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 278800.0 158700.0 279600.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 288000.0 158700.0 288800.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 297200.0 158700.0 298000.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 306400.0 158700.0 307200.0 ;
      RECT  159500.0 315600.0 158700.0 316400.00000000006 ;
      RECT  159500.0 315600.0 158700.0 316400.00000000006 ;
      RECT  158800.0 177700.0 159400.0 178300.0 ;
      RECT  158800.0 196100.00000000003 159400.0 196700.0 ;
      RECT  158800.0 214500.0 159400.0 215100.00000000003 ;
      RECT  158800.0 232900.00000000003 159400.0 233500.0 ;
      RECT  158800.0 251300.0 159400.0 251900.00000000003 ;
      RECT  158800.0 269700.0 159400.0 270300.0 ;
      RECT  158800.0 288100.0 159400.0 288700.0 ;
      RECT  158800.0 306500.0 159400.0 307100.0 ;
      RECT  158800.0 168500.0 159400.0 169100.00000000003 ;
      RECT  158800.0 186900.0 159400.0 187500.0 ;
      RECT  158800.0 205300.0 159400.0 205899.99999999997 ;
      RECT  158800.0 223700.0 159400.0 224300.0 ;
      RECT  158800.0 242100.00000000003 159400.0 242700.0 ;
      RECT  158800.0 260500.0 159400.0 261100.00000000003 ;
      RECT  158800.0 278900.00000000006 159400.0 279500.0 ;
      RECT  158800.0 297300.0 159400.0 297900.0 ;
      RECT  158800.0 315700.0 159400.0 316300.0 ;
      RECT  174400.0 177200.0 175200.0 178000.0 ;
      RECT  181200.0 177200.0 182000.0 178000.0 ;
      RECT  174400.0 195600.00000000003 175200.0 196400.0 ;
      RECT  181200.0 195600.00000000003 182000.0 196400.0 ;
      RECT  174400.0 214000.0 175200.0 214800.0 ;
      RECT  181200.0 214000.0 182000.0 214800.0 ;
      RECT  174400.0 232399.99999999997 175200.0 233200.0 ;
      RECT  181200.0 232399.99999999997 182000.0 233200.0 ;
      RECT  174400.0 250800.0 175200.0 251600.00000000003 ;
      RECT  181200.0 250800.0 182000.0 251600.00000000003 ;
      RECT  174400.0 269200.0 175200.0 270000.0 ;
      RECT  181200.0 269200.0 182000.0 270000.0 ;
      RECT  174400.0 287600.0 175200.0 288400.0 ;
      RECT  181200.0 287600.0 182000.0 288400.0 ;
      RECT  174400.0 306000.0 175200.0 306800.0 ;
      RECT  181200.0 306000.0 182000.0 306800.0 ;
      RECT  174200.0 158000.0 175000.0 158800.0 ;
      RECT  181000.0 158000.0 181800.0 158800.0 ;
      RECT  176900.0 127700.0 177500.0 128300.00000000001 ;
      RECT  183700.0 127700.0 184300.0 128300.00000000001 ;
      RECT  175300.0 76500.0 175900.0 77100.0 ;
      RECT  174700.0 93900.0 175300.0 94500.0 ;
      RECT  182100.00000000003 76500.0 182700.0 77100.0 ;
      RECT  181500.0 93900.0 182100.00000000003 94500.0 ;
      RECT  131300.0 177600.00000000003 132100.0 178400.0 ;
      RECT  131300.0 196000.0 132100.0 196800.0 ;
      RECT  131300.0 214399.99999999997 132100.0 215200.0 ;
      RECT  131300.0 232800.0 132100.0 233600.00000000003 ;
      RECT  131300.0 251200.0 132100.0 252000.0 ;
      RECT  131300.0 269600.0 132100.0 270400.0 ;
      RECT  131300.0 288000.0 132100.0 288800.0 ;
      RECT  131300.0 306400.0 132100.0 307200.0 ;
      RECT  90900.0 177600.00000000003 91700.0 178400.0 ;
      RECT  108300.00000000001 177600.00000000003 109100.0 178400.0 ;
      RECT  90900.0 196000.0 91700.0 196800.0 ;
      RECT  108300.00000000001 196000.0 109100.0 196800.0 ;
      RECT  90900.0 214399.99999999997 91700.0 215200.0 ;
      RECT  108300.00000000001 214399.99999999997 109100.0 215200.0 ;
      RECT  90900.0 232800.0 91700.0 233600.00000000003 ;
      RECT  108300.00000000001 232800.0 109100.0 233600.00000000003 ;
      RECT  158800.0 177700.0 159400.0 178300.0 ;
      RECT  158800.0 196100.00000000003 159400.0 196700.0 ;
      RECT  158800.0 214500.0 159400.0 215100.00000000003 ;
      RECT  158800.0 232899.99999999997 159400.0 233500.0 ;
      RECT  158800.0 251300.0 159400.0 251899.99999999997 ;
      RECT  158800.0 269700.0 159400.0 270300.0 ;
      RECT  158800.0 288100.0 159400.0 288700.0 ;
      RECT  158800.0 306500.0 159400.0 307100.0 ;
      RECT  171000.0 172600.00000000003 171800.0 173400.0 ;
      RECT  177800.0 172600.00000000003 178600.00000000003 173400.0 ;
      RECT  184600.00000000003 172600.00000000003 185400.0 173400.0 ;
      RECT  171000.0 181800.0 171800.0 182600.00000000003 ;
      RECT  177800.0 181800.0 178600.00000000003 182600.00000000003 ;
      RECT  184600.00000000003 181800.0 185400.0 182600.00000000003 ;
      RECT  171000.0 191000.0 171800.0 191800.0 ;
      RECT  177800.0 191000.0 178600.00000000003 191800.0 ;
      RECT  184600.00000000003 191000.0 185400.0 191800.0 ;
      RECT  171000.0 200200.0 171800.0 201000.0 ;
      RECT  177800.0 200200.0 178600.00000000003 201000.0 ;
      RECT  184600.00000000003 200200.0 185400.0 201000.0 ;
      RECT  171000.0 209399.99999999997 171800.0 210200.0 ;
      RECT  177800.0 209399.99999999997 178600.00000000003 210200.0 ;
      RECT  184600.00000000003 209399.99999999997 185400.0 210200.0 ;
      RECT  171000.0 218600.00000000003 171800.0 219399.99999999997 ;
      RECT  177800.0 218600.00000000003 178600.00000000003 219399.99999999997 ;
      RECT  184600.00000000003 218600.00000000003 185400.0 219399.99999999997 ;
      RECT  171000.0 227800.0 171800.0 228600.00000000003 ;
      RECT  177800.0 227800.0 178600.00000000003 228600.00000000003 ;
      RECT  184600.00000000003 227800.0 185400.0 228600.00000000003 ;
      RECT  171000.0 237000.0 171800.0 237800.0 ;
      RECT  177800.0 237000.0 178600.00000000003 237800.0 ;
      RECT  184600.00000000003 237000.0 185400.0 237800.0 ;
      RECT  171000.0 246200.0 171800.0 247000.0 ;
      RECT  177800.0 246200.0 178600.00000000003 247000.0 ;
      RECT  184600.00000000003 246200.0 185400.0 247000.0 ;
      RECT  171000.0 255399.99999999997 171800.0 256200.0 ;
      RECT  177800.0 255399.99999999997 178600.00000000003 256200.0 ;
      RECT  184600.00000000003 255399.99999999997 185400.0 256200.0 ;
      RECT  171000.0 264600.0 171800.0 265400.0 ;
      RECT  177800.0 264600.0 178600.00000000003 265400.0 ;
      RECT  184600.00000000003 264600.0 185400.0 265400.0 ;
      RECT  171000.0 273800.0 171800.0 274600.0 ;
      RECT  177800.0 273800.0 178600.00000000003 274600.0 ;
      RECT  184600.00000000003 273800.0 185400.0 274600.0 ;
      RECT  171000.0 283000.0 171800.0 283800.0 ;
      RECT  177800.0 283000.0 178600.00000000003 283800.0 ;
      RECT  184600.00000000003 283000.0 185400.0 283800.0 ;
      RECT  171000.0 292200.0 171800.0 293000.0 ;
      RECT  177800.0 292200.0 178600.00000000003 293000.0 ;
      RECT  184600.00000000003 292200.0 185400.0 293000.0 ;
      RECT  171000.0 301400.0 171800.0 302200.0 ;
      RECT  177800.0 301400.0 178600.00000000003 302200.0 ;
      RECT  184600.00000000003 301400.0 185400.0 302200.0 ;
      RECT  171000.0 310600.0 171800.0 311400.0 ;
      RECT  177800.0 310600.0 178600.00000000003 311400.0 ;
      RECT  184600.00000000003 310600.0 185400.0 311400.0 ;
      RECT  177900.0 141100.00000000003 178500.0 141700.0 ;
      RECT  184700.0 141100.00000000003 185300.0 141700.0 ;
      RECT  175300.0 83100.0 175900.0 83700.0 ;
      RECT  176700.0 87500.0 177300.0 88100.0 ;
      RECT  176100.00000000003 100900.0 176700.0 101500.0 ;
      RECT  182100.00000000003 83100.0 182700.0 83700.0 ;
      RECT  183500.0 87500.0 184100.00000000003 88100.0 ;
      RECT  182900.0 100900.0 183500.0 101500.0 ;
      RECT  131300.0 168400.0 132100.0 169200.0 ;
      RECT  131300.0 186800.0 132100.0 187600.00000000003 ;
      RECT  131300.0 205200.0 132100.0 206000.0 ;
      RECT  131300.0 223600.00000000003 132100.0 224399.99999999997 ;
      RECT  131300.0 242000.0 132100.0 242800.0 ;
      RECT  131300.0 260399.99999999997 132100.0 261200.0 ;
      RECT  131300.0 278800.0 132100.0 279600.0 ;
      RECT  131300.0 297200.0 132100.0 298000.0 ;
      RECT  131300.0 315600.0 132100.0 316400.0 ;
      RECT  90900.0 168400.0 91700.0 169200.0 ;
      RECT  108300.00000000001 168400.0 109100.0 169200.0 ;
      RECT  90900.0 186800.0 91700.0 187600.00000000003 ;
      RECT  108300.00000000001 186800.0 109100.0 187600.00000000003 ;
      RECT  90900.0 205200.0 91700.0 206000.0 ;
      RECT  108300.00000000001 205200.0 109100.0 206000.0 ;
      RECT  90900.0 223600.00000000003 91700.0 224399.99999999997 ;
      RECT  108300.00000000001 223600.00000000003 109100.0 224399.99999999997 ;
      RECT  90900.0 242000.0 91700.0 242800.0 ;
      RECT  108300.00000000001 242000.0 109100.0 242800.0 ;
      RECT  158800.0 168500.0 159400.0 169100.00000000003 ;
      RECT  158800.0 186900.0 159400.0 187500.0 ;
      RECT  158800.0 205300.0 159400.0 205899.99999999997 ;
      RECT  158800.0 223700.0 159400.0 224300.0 ;
      RECT  158800.0 242100.00000000003 159400.0 242700.0 ;
      RECT  158800.0 260500.0 159400.0 261100.00000000003 ;
      RECT  158800.0 278900.0 159400.0 279500.0 ;
      RECT  158800.0 297300.0 159400.0 297900.0 ;
      RECT  158800.0 315700.0 159400.0 316300.0 ;
      RECT  30199.999999999993 12100.000000000007 44300.0 12700.000000000007 ;
      RECT  30199.999999999993 30100.000000000007 40099.99999999999 30700.00000000001 ;
      RECT  35599.99999999999 33300.000000000015 42899.99999999999 33900.00000000001 ;
      RECT  4299.999999999992 111900.0 59999.99999999999 112500.0 ;
      RECT  41499.99999999999 10300.000000000005 56800.0 10900.000000000005 ;
      RECT  44300.0 36300.00000000001 55199.99999999999 36900.00000000001 ;
      RECT  37299.99999999999 31900.000000000007 66399.99999999999 32500.000000000007 ;
      RECT  38699.99999999999 50300.000000000015 60000.0 50900.000000000015 ;
      RECT  23599.999999999993 10900.000000000005 24199.999999999996 11500.000000000005 ;
      RECT  23599.999999999993 10700.000000000007 24199.999999999996 11300.000000000005 ;
      RECT  21599.999999999993 10900.000000000005 23899.999999999996 11500.000000000005 ;
      RECT  23599.999999999993 11000.000000000007 24199.999999999996 11200.000000000007 ;
      RECT  23899.999999999993 10700.000000000007 26199.999999999993 11300.000000000005 ;
      RECT  21199.999999999993 10800.000000000005 21999.999999999993 11600.000000000007 ;
      RECT  25799.999999999993 10600.000000000007 26599.999999999993 11400.000000000007 ;
      RECT  23599.999999999993 31900.000000000007 24199.999999999996 31300.000000000004 ;
      RECT  23599.999999999993 32100.000000000007 24199.999999999996 31500.000000000007 ;
      RECT  21599.999999999993 31900.000000000007 23899.999999999996 31300.000000000004 ;
      RECT  23599.999999999993 31800.000000000004 24199.999999999996 31600.000000000004 ;
      RECT  23899.999999999993 32100.000000000007 26199.999999999993 31500.000000000007 ;
      RECT  21199.999999999993 32000.000000000007 21999.999999999993 31200.000000000004 ;
      RECT  25799.999999999993 32200.000000000004 26599.999999999993 31400.000000000007 ;
      RECT  2799.9999999999914 21000.000000000007 1999.9999999999916 21800.000000000007 ;
      RECT  2799.9999999999914 1000.0000000000058 1999.9999999999916 1800.0000000000057 ;
      RECT  2799.9999999999914 21000.000000000007 1999.9999999999916 21800.000000000007 ;
      RECT  2799.9999999999914 41000.00000000001 1999.9999999999916 41800.00000000001 ;
      RECT  1999.9999999999916 21000.000000000007 2799.9999999999914 21800.000000000007 ;
      RECT  1999.9999999999916 1000.0000000000058 2799.9999999999914 1800.0000000000057 ;
      RECT  1999.9999999999916 41000.00000000001 2799.9999999999914 41800.000000000015 ;
      RECT  5999.999999999991 179600.00000000003 23599.999999999993 180200.00000000003 ;
      RECT  5999.999999999991 189200.00000000003 23599.999999999993 189800.0 ;
      RECT  5999.999999999991 198000.00000000003 23599.999999999993 198600.00000000003 ;
      RECT  5999.999999999991 207600.00000000003 23599.999999999993 208200.00000000003 ;
      RECT  10399.99999999999 179500.00000000003 11199.999999999993 180300.0 ;
      RECT  16799.99999999999 179500.00000000003 17599.999999999993 180300.0 ;
      RECT  23199.999999999993 179500.00000000003 23999.999999999993 180300.0 ;
      RECT  5599.999999999992 179500.00000000003 6399.999999999992 180300.0 ;
      RECT  10399.99999999999 189100.00000000003 11199.999999999993 189900.0 ;
      RECT  16799.99999999999 189100.00000000003 17599.999999999993 189900.0 ;
      RECT  23199.999999999993 189100.00000000003 23999.999999999993 189900.0 ;
      RECT  5599.999999999992 189100.00000000003 6399.999999999992 189900.0 ;
      RECT  10399.99999999999 197900.0 11199.999999999993 198700.00000000003 ;
      RECT  16799.99999999999 197900.0 17599.999999999993 198700.00000000003 ;
      RECT  23199.999999999993 197900.0 23999.999999999993 198700.00000000003 ;
      RECT  5599.999999999992 197900.0 6399.999999999992 198700.00000000003 ;
      RECT  10399.99999999999 207500.00000000003 11199.999999999993 208300.0 ;
      RECT  16799.99999999999 207500.00000000003 17599.999999999993 208300.0 ;
      RECT  23199.999999999993 207500.00000000003 23999.999999999993 208300.0 ;
      RECT  5599.999999999992 207500.00000000003 6399.999999999992 208300.0 ;
      RECT  15599.999999999993 184300.0 14799.999999999993 185100.00000000003 ;
      RECT  15599.999999999993 175100.00000000003 14799.999999999993 175900.0 ;
      RECT  21999.999999999993 184300.0 21199.999999999993 185100.00000000003 ;
      RECT  21999.999999999993 175100.00000000003 21199.999999999993 175900.0 ;
      RECT  15599.999999999993 202700.00000000003 14799.999999999993 203500.00000000003 ;
      RECT  15599.999999999993 193500.00000000003 14799.999999999993 194300.0 ;
      RECT  21999.999999999993 202700.00000000003 21199.999999999993 203500.00000000003 ;
      RECT  21999.999999999993 193500.00000000003 21199.999999999993 194300.0 ;
      RECT  15599.999999999993 211900.0 14799.999999999993 212700.00000000003 ;
      RECT  21999.999999999993 211900.0 21199.999999999993 212700.00000000003 ;
      RECT  14799.999999999993 184300.0 15599.999999999993 185100.00000000003 ;
      RECT  21199.999999999993 184300.0 21999.999999999993 185100.00000000003 ;
      RECT  14799.999999999993 202700.00000000003 15599.999999999993 203500.00000000003 ;
      RECT  21199.999999999993 202700.00000000003 21999.999999999993 203500.00000000003 ;
      RECT  14799.999999999993 175100.00000000003 15599.999999999993 175900.0 ;
      RECT  21199.999999999993 175100.00000000003 21999.999999999993 175900.0 ;
      RECT  14799.999999999993 193500.00000000003 15599.999999999993 194300.0 ;
      RECT  21199.999999999993 193500.00000000003 21999.999999999993 194300.0 ;
      RECT  14799.999999999993 211900.0 15599.999999999993 212700.00000000003 ;
      RECT  21199.999999999993 211900.0 21999.999999999993 212700.00000000003 ;
      RECT  33800.0 184300.0 34599.99999999999 185100.00000000003 ;
      RECT  30399.999999999996 179700.00000000003 31199.999999999993 180500.00000000003 ;
      RECT  37199.99999999999 179700.00000000003 37999.99999999999 180500.00000000003 ;
      RECT  33800.0 184300.0 34599.99999999999 185100.00000000003 ;
      RECT  30399.999999999996 188900.0 31199.999999999993 189700.00000000003 ;
      RECT  37199.99999999999 188900.0 37999.99999999999 189700.00000000003 ;
      RECT  33800.0 202700.00000000003 34599.99999999999 203500.00000000003 ;
      RECT  30399.999999999996 198100.00000000003 31199.999999999993 198900.0 ;
      RECT  37199.99999999999 198100.00000000003 37999.99999999999 198900.0 ;
      RECT  33800.0 202700.00000000003 34599.99999999999 203500.00000000003 ;
      RECT  30399.999999999996 207300.0 31199.999999999993 208100.00000000003 ;
      RECT  37199.99999999999 207300.0 37999.99999999999 208100.00000000003 ;
      RECT  33800.0 221100.00000000003 34599.99999999999 221900.0 ;
      RECT  30399.999999999996 216500.00000000003 31199.999999999993 217300.0 ;
      RECT  37199.99999999999 216500.00000000003 37999.99999999999 217300.0 ;
      RECT  33800.0 221100.00000000003 34599.99999999999 221900.0 ;
      RECT  30399.999999999996 225700.00000000003 31199.999999999993 226500.00000000003 ;
      RECT  37199.99999999999 225700.00000000003 37999.99999999999 226500.00000000003 ;
      RECT  33800.0 239500.00000000003 34599.99999999999 240300.0 ;
      RECT  30399.999999999996 234900.0 31199.999999999993 235700.00000000003 ;
      RECT  37199.99999999999 234900.0 37999.99999999999 235700.00000000003 ;
      RECT  33800.0 239500.00000000003 34599.99999999999 240300.0 ;
      RECT  30399.999999999996 244100.00000000003 31199.999999999993 244900.0 ;
      RECT  37199.99999999999 244100.00000000003 37999.99999999999 244900.0 ;
      RECT  33800.0 184300.0 34599.99999999999 185100.00000000003 ;
      RECT  33800.0 202700.00000000003 34599.99999999999 203500.00000000003 ;
      RECT  33800.0 221100.00000000003 34599.99999999999 221900.0 ;
      RECT  33800.0 239500.00000000003 34599.99999999999 240300.0 ;
      RECT  30399.999999999996 179700.00000000003 31199.999999999993 180500.00000000003 ;
      RECT  37199.99999999999 179700.00000000003 37999.99999999999 180500.00000000003 ;
      RECT  30399.999999999996 188900.0 31199.999999999993 189700.00000000003 ;
      RECT  37199.99999999999 188900.0 37999.99999999999 189700.00000000003 ;
      RECT  30399.999999999996 198100.00000000003 31199.999999999993 198900.0 ;
      RECT  37199.99999999999 198100.00000000003 37999.99999999999 198900.0 ;
      RECT  30399.999999999996 207300.0 31199.999999999993 208100.00000000003 ;
      RECT  37199.99999999999 207300.0 37999.99999999999 208100.00000000003 ;
      RECT  30399.999999999996 216500.00000000003 31199.999999999993 217300.00000000003 ;
      RECT  37199.99999999999 216500.00000000003 37999.99999999999 217300.00000000003 ;
      RECT  30399.999999999996 225700.00000000003 31199.999999999993 226500.00000000003 ;
      RECT  37199.99999999999 225700.00000000003 37999.99999999999 226500.00000000003 ;
      RECT  30399.999999999996 234900.0 31199.999999999993 235700.00000000003 ;
      RECT  37199.99999999999 234900.0 37999.99999999999 235700.00000000003 ;
      RECT  30399.999999999996 244100.00000000003 31199.999999999993 244900.0 ;
      RECT  37199.99999999999 244100.00000000003 37999.99999999999 244900.0 ;
      RECT  9199.999999999993 165900.0 8399.99999999999 166700.00000000003 ;
      RECT  33800.0 165900.0 34599.99999999999 166700.00000000003 ;
      RECT  31199.999999999993 170500.00000000003 30399.999999999993 171300.0 ;
      RECT  37999.99999999999 170500.00000000003 37199.99999999999 171300.0 ;
      RECT  40599.99999999999 176500.00000000003 39800.0 177300.0 ;
      RECT  40599.99999999999 192100.00000000003 39800.0 192900.0 ;
      RECT  40599.99999999999 194900.0 39800.0 195700.00000000003 ;
      RECT  40599.99999999999 210500.00000000003 39800.0 211300.0 ;
      RECT  40599.99999999999 213300.0 39800.0 214100.00000000003 ;
      RECT  40599.99999999999 228900.0 39800.0 229700.00000000003 ;
      RECT  40599.99999999999 231700.00000000003 39800.0 232500.00000000003 ;
      RECT  40599.99999999999 247300.0 39800.0 248100.0 ;
      RECT  19599.999999999993 170900.0 20399.999999999996 171700.00000000003 ;
      RECT  33800.0 184300.0 34599.99999999999 185100.00000000003 ;
      RECT  33800.0 202700.00000000003 34599.99999999999 203500.00000000003 ;
      RECT  33800.0 221100.00000000003 34599.99999999999 221900.0 ;
      RECT  33800.0 239500.00000000003 34599.99999999999 240300.0 ;
      RECT  14799.999999999993 184300.0 15599.999999999993 185100.00000000003 ;
      RECT  21199.999999999993 184300.0 21999.999999999993 185100.00000000003 ;
      RECT  14799.999999999993 202700.00000000003 15599.999999999993 203500.00000000003 ;
      RECT  21199.999999999993 202700.00000000003 21999.999999999993 203500.00000000003 ;
      RECT  8399.99999999999 165900.0 9199.999999999993 166700.00000000003 ;
      RECT  33800.0 165900.0 34599.99999999999 166700.00000000003 ;
      RECT  19599.999999999993 170900.0 20399.999999999993 171700.00000000003 ;
      RECT  30399.999999999996 179700.00000000003 31199.999999999993 180500.00000000003 ;
      RECT  37199.99999999999 179700.00000000003 37999.99999999999 180500.00000000003 ;
      RECT  30399.999999999996 188900.0 31199.999999999993 189700.00000000003 ;
      RECT  37199.99999999999 188900.0 37999.99999999999 189700.00000000003 ;
      RECT  30399.999999999996 198100.00000000003 31199.999999999993 198900.0 ;
      RECT  37199.99999999999 198100.00000000003 37999.99999999999 198900.0 ;
      RECT  30399.999999999996 207300.0 31199.999999999993 208100.00000000003 ;
      RECT  37199.99999999999 207300.0 37999.99999999999 208100.00000000003 ;
      RECT  30399.999999999996 216500.00000000003 31199.999999999993 217300.0 ;
      RECT  37199.99999999999 216500.00000000003 37999.99999999999 217300.0 ;
      RECT  30399.999999999996 225700.00000000003 31199.999999999993 226500.00000000003 ;
      RECT  37199.99999999999 225700.00000000003 37999.99999999999 226500.00000000003 ;
      RECT  30399.999999999996 234900.0 31199.999999999993 235700.00000000003 ;
      RECT  37199.99999999999 234900.0 37999.99999999999 235700.00000000003 ;
      RECT  30399.999999999996 244100.00000000003 31199.999999999993 244900.0 ;
      RECT  37199.99999999999 244100.00000000003 37999.99999999999 244900.0 ;
      RECT  14799.999999999993 175100.00000000003 15599.999999999993 175900.0 ;
      RECT  21199.999999999993 175100.00000000003 21999.999999999993 175900.0 ;
      RECT  14799.999999999993 193500.00000000003 15599.999999999993 194300.0 ;
      RECT  21199.999999999993 193500.00000000003 21999.999999999993 194300.0 ;
      RECT  14799.999999999993 211900.0 15599.999999999993 212700.00000000003 ;
      RECT  21199.999999999993 211900.0 21999.999999999993 212700.00000000003 ;
      RECT  30399.999999999996 170500.00000000003 31199.999999999993 171300.0 ;
      RECT  37199.99999999999 170500.00000000003 37999.99999999999 171300.0 ;
      RECT  39800.0 176500.00000000003 40599.99999999999 177300.0 ;
      RECT  39800.0 192100.00000000003 40599.99999999999 192900.0 ;
      RECT  39800.0 194900.0 40599.99999999999 195700.00000000003 ;
      RECT  39800.0 210500.00000000003 40599.99999999999 211300.0 ;
      RECT  39800.0 213300.0 40599.99999999999 214100.00000000003 ;
      RECT  39800.0 228900.0 40599.99999999999 229700.00000000003 ;
      RECT  39800.0 231700.00000000003 40599.99999999999 232500.00000000003 ;
      RECT  39800.0 247300.0 40599.99999999999 248100.00000000003 ;
      RECT  44699.99999999999 12000.000000000007 43900.0 12800.000000000007 ;
      RECT  29799.999999999993 12000.000000000007 30599.999999999993 12800.000000000007 ;
      RECT  40499.99999999999 30000.000000000007 39699.99999999999 30800.000000000007 ;
      RECT  29799.999999999993 30000.000000000007 30599.999999999993 30800.000000000007 ;
      RECT  43300.0 33200.0 42500.0 34000.00000000001 ;
      RECT  35199.99999999999 33200.0 35999.99999999999 34000.00000000001 ;
      RECT  4699.999999999992 111800.00000000001 3899.9999999999914 112600.00000000001 ;
      RECT  60399.99999999999 111800.00000000001 59599.99999999999 112600.00000000001 ;
      RECT  41899.99999999999 10200.000000000007 41099.99999999999 11000.000000000007 ;
      RECT  56399.99999999999 10200.000000000007 57199.999999999985 11000.000000000007 ;
      RECT  44699.99999999999 36200.00000000001 43900.0 37000.00000000001 ;
      RECT  54800.0 36200.00000000001 55599.99999999999 37000.00000000001 ;
      RECT  37699.99999999999 31800.000000000007 36900.0 32600.000000000007 ;
      RECT  66000.0 31800.000000000007 66800.0 32600.000000000007 ;
      RECT  39099.99999999999 50200.00000000001 38300.0 51000.00000000001 ;
      RECT  59599.99999999999 50200.00000000001 60399.99999999999 51000.00000000001 ;
      RECT  71199.99999999999 21000.000000000007 70399.99999999999 21800.000000000007 ;
      RECT  71199.99999999999 1000.0000000000058 70399.99999999999 1800.0000000000057 ;
      RECT  71199.99999999999 21000.000000000007 70399.99999999999 21800.000000000007 ;
      RECT  71199.99999999999 41000.00000000001 70399.99999999999 41800.00000000001 ;
      RECT  71199.99999999999 61000.00000000001 70399.99999999999 61800.00000000001 ;
      RECT  71199.99999999999 41000.00000000001 70399.99999999999 41800.00000000001 ;
      RECT  71199.99999999999 61000.00000000001 70399.99999999999 61800.00000000001 ;
      RECT  71199.99999999999 81000.00000000001 70399.99999999999 81800.00000000001 ;
      RECT  71199.99999999999 101000.00000000001 70399.99999999999 101800.00000000001 ;
      RECT  71199.99999999999 81000.00000000001 70399.99999999999 81800.00000000001 ;
      RECT  71199.99999999999 101000.00000000001 70399.99999999999 101800.00000000001 ;
      RECT  71199.99999999999 121000.00000000001 70399.99999999999 121800.00000000001 ;
      RECT  71199.99999999999 141000.0 70399.99999999999 141800.0 ;
      RECT  71199.99999999999 121000.00000000001 70399.99999999999 121800.00000000001 ;
      RECT  71199.99999999999 141000.0 70399.99999999999 141800.0 ;
      RECT  71199.99999999999 161000.00000000003 70399.99999999999 161800.00000000003 ;
      RECT  70399.99999999999 21000.000000000007 71199.99999999999 21800.000000000007 ;
      RECT  70399.99999999999 61000.00000000001 71199.99999999999 61800.000000000015 ;
      RECT  70399.99999999999 101000.00000000001 71199.99999999999 101800.00000000001 ;
      RECT  70399.99999999999 141000.0 71199.99999999999 141800.0 ;
      RECT  33800.0 184300.0 34599.99999999999 185100.00000000003 ;
      RECT  33800.0 202700.00000000003 34599.99999999999 203500.00000000003 ;
      RECT  33800.0 221100.00000000003 34599.99999999999 221900.0 ;
      RECT  33800.0 239500.00000000003 34599.99999999999 240300.0 ;
      RECT  14799.999999999993 184300.0 15599.999999999993 185100.00000000003 ;
      RECT  21199.999999999993 184300.0 21999.999999999993 185100.00000000003 ;
      RECT  14799.999999999993 202700.00000000003 15599.999999999993 203500.00000000003 ;
      RECT  21199.999999999993 202700.00000000003 21999.999999999993 203500.00000000003 ;
      RECT  8399.99999999999 165900.0 9199.999999999993 166700.00000000003 ;
      RECT  33800.0 165900.0 34599.99999999999 166700.00000000003 ;
      RECT  19599.99999999999 170900.0 20399.999999999993 171700.00000000003 ;
      RECT  1999.9999999999916 21000.000000000007 2799.9999999999914 21800.000000000007 ;
      RECT  70399.99999999999 1000.0000000000058 71199.99999999999 1800.0000000000057 ;
      RECT  70399.99999999999 41000.00000000001 71199.99999999999 41800.000000000015 ;
      RECT  70399.99999999999 81000.00000000001 71199.99999999999 81800.00000000001 ;
      RECT  70399.99999999999 121000.00000000001 71199.99999999999 121800.00000000001 ;
      RECT  70399.99999999999 161000.00000000003 71199.99999999999 161800.0 ;
      RECT  30399.999999999993 179700.00000000003 31199.999999999993 180500.00000000003 ;
      RECT  37199.99999999999 179700.00000000003 37999.99999999999 180500.00000000003 ;
      RECT  30399.999999999993 188900.0 31199.999999999993 189700.00000000003 ;
      RECT  37199.99999999999 188900.0 37999.99999999999 189700.00000000003 ;
      RECT  30399.999999999993 198100.00000000003 31199.999999999993 198900.0 ;
      RECT  37199.99999999999 198100.00000000003 37999.99999999999 198900.0 ;
      RECT  30399.999999999993 207300.0 31199.999999999993 208100.00000000003 ;
      RECT  37199.99999999999 207300.0 37999.99999999999 208100.00000000003 ;
      RECT  30399.999999999993 216500.00000000003 31199.999999999993 217300.0 ;
      RECT  37199.99999999999 216500.00000000003 37999.99999999999 217300.0 ;
      RECT  30399.999999999993 225700.00000000003 31199.999999999993 226500.00000000003 ;
      RECT  37199.99999999999 225700.00000000003 37999.99999999999 226500.00000000003 ;
      RECT  30399.999999999993 234900.0 31199.999999999993 235700.00000000003 ;
      RECT  37199.99999999999 234900.0 37999.99999999999 235700.00000000003 ;
      RECT  30399.999999999993 244100.00000000003 31199.999999999993 244900.0 ;
      RECT  37199.99999999999 244100.00000000003 37999.99999999999 244900.0 ;
      RECT  14799.999999999993 175100.00000000003 15599.999999999993 175900.0 ;
      RECT  21199.999999999993 175100.00000000003 21999.999999999993 175900.0 ;
      RECT  14799.999999999993 193500.00000000003 15599.999999999993 194300.0 ;
      RECT  21199.999999999993 193500.00000000003 21999.999999999993 194300.0 ;
      RECT  14799.999999999993 211900.0 15599.999999999993 212700.00000000003 ;
      RECT  21199.999999999993 211900.0 21999.999999999993 212700.00000000003 ;
      RECT  30399.999999999993 170500.00000000003 31199.999999999993 171300.0 ;
      RECT  37199.99999999999 170500.00000000003 37999.99999999999 171300.0 ;
      RECT  39799.99999999999 176500.00000000003 40599.99999999999 177300.0 ;
      RECT  39799.99999999999 192100.00000000003 40599.99999999999 192900.0 ;
      RECT  39799.99999999999 194900.0 40599.99999999999 195700.00000000003 ;
      RECT  39799.99999999999 210500.00000000003 40599.99999999999 211300.0 ;
      RECT  39799.99999999999 213300.0 40599.99999999999 214100.00000000003 ;
      RECT  39799.99999999999 228900.0 40599.99999999999 229700.00000000003 ;
      RECT  39799.99999999999 231700.00000000003 40599.99999999999 232500.00000000003 ;
      RECT  39799.99999999999 247300.0 40599.99999999999 248100.00000000003 ;
      RECT  1999.9999999999916 1000.0000000000058 2799.9999999999914 1800.0000000000057 ;
      RECT  1999.9999999999916 41000.00000000001 2799.9999999999914 41800.000000000015 ;
      RECT  61700.0 275700.00000000006 60900.0 276500.0 ;
      RECT  61700.0 255700.00000000003 60900.0 256500.0 ;
      RECT  61700.0 275700.00000000006 60900.0 276500.0 ;
      RECT  61700.0 295700.00000000006 60900.0 296500.0 ;
      RECT  61700.0 315700.00000000006 60900.0 316500.0 ;
      RECT  61700.0 295700.00000000006 60900.0 296500.0 ;
      RECT  61700.0 315700.00000000006 60900.0 316500.0 ;
      RECT  61700.0 335700.00000000006 60900.0 336500.0 ;
      RECT  53199.99999999999 261100.00000000003 54000.0 261900.00000000003 ;
      RECT  50400.0 261200.00000000006 72200.0 261800.0 ;
      RECT  60900.0 275700.00000000006 61700.0 276500.0 ;
      RECT  60900.0 315700.00000000006 61700.0 316500.0 ;
      RECT  60900.0 255700.00000000003 61700.0 256500.0 ;
      RECT  60900.0 295700.00000000006 61700.0 296500.0 ;
      RECT  60900.0 335700.00000000006 61700.0 336500.0 ;
      RECT  182700.00000000003 62800.00000000001 181900.0 63600.00000000001 ;
      RECT  182700.00000000003 42800.00000000001 181900.0 43600.0 ;
      RECT  204500.0 62800.00000000001 203700.00000000003 63600.00000000001 ;
      RECT  204500.0 42800.00000000001 203700.00000000003 43600.0 ;
      RECT  174200.00000000003 48200.0 175000.0 49000.0 ;
      RECT  196000.0 48200.0 196800.0 49000.0 ;
      RECT  171400.0 48300.00000000001 215000.0 48900.00000000001 ;
      RECT  181900.0 62800.00000000001 182700.00000000003 63600.00000000001 ;
      RECT  203700.00000000003 62800.00000000001 204500.0 63600.00000000001 ;
      RECT  181900.0 42800.00000000001 182700.00000000003 43600.0 ;
      RECT  203700.00000000003 42800.00000000001 204500.0 43600.0 ;
      RECT  74000.0 261100.00000000003 73200.0 261900.00000000003 ;
      RECT  74000.0 48200.0 73200.0 49000.0 ;
      RECT  168700.0 151800.0 167899.99999999997 152600.00000000003 ;
      RECT  72600.0 151800.0 71800.0 152600.00000000003 ;
      RECT  167300.0 90200.0 166500.0 91000.0 ;
      RECT  72600.0 90200.0 71800.0 91000.0 ;
      RECT  170100.00000000003 130199.99999999999 169300.0 131000.0 ;
      RECT  72600.0 130199.99999999999 71800.0 131000.0 ;
      RECT  165900.0 71800.0 165100.0 72600.0 ;
      RECT  72600.0 71800.0 71800.0 72600.0 ;
      RECT  75800.0 265500.0 75000.0 266300.0 ;
      RECT  70000.0 265500.0 69200.0 266300.0 ;
      RECT  77200.0 285900.00000000006 76400.0 286700.00000000006 ;
      RECT  70000.0 285900.00000000006 69200.0 286700.00000000006 ;
      RECT  78600.0 305500.0 77800.0 306300.0 ;
      RECT  70000.0 305500.0 69200.0 306300.0 ;
      RECT  80000.0 325900.00000000006 79200.0 326700.00000000006 ;
      RECT  70000.0 325900.00000000006 69200.0 326700.00000000006 ;
      RECT  7400.000000000003 4999.999999999997 8200.000000000004 5799.999999999997 ;
      RECT  12200.0 4999.999999999997 13000.0 5799.999999999997 ;
      RECT  16999.999999999996 4999.999999999997 17799.999999999996 5799.999999999997 ;
      RECT  21799.999999999993 4999.999999999997 22599.999999999993 5799.999999999997 ;
      RECT  26599.999999999996 4999.999999999997 27400.0 5799.999999999997 ;
      RECT  31399.999999999996 4999.999999999997 32199.999999999996 5799.999999999997 ;
      RECT  36200.0 4999.999999999997 37000.0 5799.999999999997 ;
      RECT  41000.0 4999.999999999997 41800.0 5799.999999999997 ;
      RECT  45800.0 4999.999999999997 46599.99999999999 5799.999999999997 ;
      RECT  50600.0 4999.999999999997 51400.0 5799.999999999997 ;
      RECT  55400.00000000001 4999.999999999997 56200.0 5799.999999999997 ;
      RECT  60200.0 4999.999999999997 61000.0 5799.999999999997 ;
      RECT  65000.0 4999.999999999997 65800.0 5799.999999999997 ;
      RECT  69800.0 4999.999999999997 70600.0 5799.999999999997 ;
      RECT  74600.00000000001 4999.999999999997 75400.0 5799.999999999997 ;
      RECT  79400.0 4999.999999999997 80200.0 5799.999999999997 ;
      RECT  84200.0 4999.999999999997 85000.0 5799.999999999997 ;
      RECT  89000.0 4999.999999999997 89800.0 5799.999999999997 ;
      RECT  93800.0 4999.999999999997 94600.0 5799.999999999997 ;
      RECT  98600.00000000001 4999.999999999997 99400.0 5799.999999999997 ;
      RECT  103400.0 4999.999999999997 104200.0 5799.999999999997 ;
      RECT  108200.0 4999.999999999997 109000.0 5799.999999999997 ;
      RECT  113000.00000000001 4999.999999999997 113800.00000000001 5799.999999999997 ;
      RECT  117800.0 4999.999999999997 118600.0 5799.999999999997 ;
      RECT  122600.00000000001 4999.999999999997 123400.0 5799.999999999997 ;
      RECT  127400.0 4999.999999999997 128199.99999999999 5799.999999999997 ;
      RECT  132200.0 4999.999999999997 133000.0 5799.999999999997 ;
      RECT  137000.0 4999.999999999997 137800.0 5799.999999999997 ;
      RECT  141800.0 4999.999999999997 142600.00000000003 5799.999999999997 ;
      RECT  146600.0 4999.999999999997 147400.0 5799.999999999997 ;
      RECT  151399.99999999997 4999.999999999997 152200.0 5799.999999999997 ;
      RECT  156200.0 4999.999999999997 157000.0 5799.999999999997 ;
      RECT  161000.0 4999.999999999997 161800.0 5799.999999999997 ;
      RECT  165800.0 4999.999999999997 166600.00000000003 5799.999999999997 ;
      RECT  170600.0 4999.999999999997 171400.0 5799.999999999997 ;
      RECT  175399.99999999997 4999.999999999997 176200.0 5799.999999999997 ;
      RECT  180200.0 4999.999999999997 181000.0 5799.999999999997 ;
      RECT  185000.0 4999.999999999997 185800.0 5799.999999999997 ;
      RECT  189800.0 4999.999999999997 190600.00000000003 5799.999999999997 ;
      RECT  194600.0 4999.999999999997 195400.0 5799.999999999997 ;
      RECT  199399.99999999997 4999.999999999997 200200.0 5799.999999999997 ;
      RECT  204200.0 4999.999999999997 205000.0 5799.999999999997 ;
      RECT  209000.0 4999.999999999997 209800.0 5799.999999999997 ;
      RECT  65000.0 9800.0 65800.0 10600.000000000002 ;
      RECT  69800.0 9800.0 70600.0 10600.000000000002 ;
      RECT  74600.00000000001 9800.0 75400.0 10600.000000000002 ;
      RECT  79400.0 9800.0 80200.0 10600.000000000002 ;
      RECT  84200.0 9800.0 85000.0 10600.000000000002 ;
      RECT  89000.0 9800.0 89800.0 10600.000000000002 ;
      RECT  93800.0 9800.0 94600.0 10600.000000000002 ;
      RECT  98600.00000000001 9800.0 99400.0 10600.000000000002 ;
      RECT  103400.0 9800.0 104200.0 10600.000000000002 ;
      RECT  108200.0 9800.0 109000.0 10600.000000000002 ;
      RECT  113000.00000000001 9800.0 113800.00000000001 10600.000000000002 ;
      RECT  117800.0 9800.0 118600.0 10600.000000000002 ;
      RECT  122600.00000000001 9800.0 123400.0 10600.000000000002 ;
      RECT  127400.0 9800.0 128199.99999999999 10600.000000000002 ;
      RECT  132200.0 9800.0 133000.0 10600.000000000002 ;
      RECT  137000.0 9800.0 137800.0 10600.000000000002 ;
      RECT  141800.0 9800.0 142600.00000000003 10600.000000000002 ;
      RECT  146600.0 9800.0 147400.0 10600.000000000002 ;
      RECT  151399.99999999997 9800.0 152200.0 10600.000000000002 ;
      RECT  156200.0 9800.0 157000.0 10600.000000000002 ;
      RECT  161000.0 9800.0 161800.0 10600.000000000002 ;
      RECT  165800.0 9800.0 166600.00000000003 10600.000000000002 ;
      RECT  170600.0 9800.0 171400.0 10600.000000000002 ;
      RECT  175399.99999999997 9800.0 176200.0 10600.000000000002 ;
      RECT  180200.0 9800.0 181000.0 10600.000000000002 ;
      RECT  185000.0 9800.0 185800.0 10600.000000000002 ;
      RECT  189800.0 9800.0 190600.00000000003 10600.000000000002 ;
      RECT  194600.0 9800.0 195400.0 10600.000000000002 ;
      RECT  199399.99999999997 9800.0 200200.0 10600.000000000002 ;
      RECT  204200.0 9800.0 205000.0 10600.000000000002 ;
      RECT  209000.0 9800.0 209800.0 10600.000000000002 ;
      RECT  7400.000000000003 14599.999999999998 8200.000000000004 15399.999999999998 ;
      RECT  12200.0 14599.999999999998 13000.0 15399.999999999998 ;
      RECT  16999.999999999996 14599.999999999998 17799.999999999996 15399.999999999998 ;
      RECT  21799.999999999993 14599.999999999998 22599.999999999993 15399.999999999998 ;
      RECT  26599.999999999996 14599.999999999998 27400.0 15399.999999999998 ;
      RECT  31399.999999999996 14599.999999999998 32199.999999999996 15399.999999999998 ;
      RECT  36200.0 14599.999999999998 37000.0 15399.999999999998 ;
      RECT  41000.0 14599.999999999998 41800.0 15399.999999999998 ;
      RECT  45800.0 14599.999999999998 46599.99999999999 15399.999999999998 ;
      RECT  50600.0 14599.999999999998 51400.0 15399.999999999998 ;
      RECT  55400.00000000001 14599.999999999998 56200.0 15399.999999999998 ;
      RECT  60200.0 14599.999999999998 61000.0 15399.999999999998 ;
      RECT  65000.0 14599.999999999998 65800.0 15399.999999999998 ;
      RECT  69800.0 14599.999999999998 70600.0 15399.999999999998 ;
      RECT  74600.00000000001 14599.999999999998 75400.0 15399.999999999998 ;
      RECT  79400.0 14599.999999999998 80200.0 15399.999999999998 ;
      RECT  84200.0 14599.999999999998 85000.0 15399.999999999998 ;
      RECT  89000.0 14599.999999999998 89800.0 15399.999999999998 ;
      RECT  93800.0 14599.999999999998 94600.0 15399.999999999998 ;
      RECT  98600.00000000001 14599.999999999998 99400.0 15399.999999999998 ;
      RECT  103400.0 14599.999999999998 104200.0 15399.999999999998 ;
      RECT  108200.0 14599.999999999998 109000.0 15399.999999999998 ;
      RECT  113000.00000000001 14599.999999999998 113800.00000000001 15399.999999999998 ;
      RECT  117800.0 14599.999999999998 118600.0 15399.999999999998 ;
      RECT  122600.00000000001 14599.999999999998 123400.0 15399.999999999998 ;
      RECT  127400.0 14599.999999999998 128199.99999999999 15399.999999999998 ;
      RECT  132200.0 14599.999999999998 133000.0 15399.999999999998 ;
      RECT  137000.0 14599.999999999998 137800.0 15399.999999999998 ;
      RECT  141800.0 14599.999999999998 142600.00000000003 15399.999999999998 ;
      RECT  146600.0 14599.999999999998 147400.0 15399.999999999998 ;
      RECT  151399.99999999997 14599.999999999998 152200.0 15399.999999999998 ;
      RECT  156200.0 14599.999999999998 157000.0 15399.999999999998 ;
      RECT  161000.0 14599.999999999998 161800.0 15399.999999999998 ;
      RECT  165800.0 14599.999999999998 166600.00000000003 15399.999999999998 ;
      RECT  170600.0 14599.999999999998 171400.0 15399.999999999998 ;
      RECT  175399.99999999997 14599.999999999998 176200.0 15399.999999999998 ;
      RECT  180200.0 14599.999999999998 181000.0 15399.999999999998 ;
      RECT  185000.0 14599.999999999998 185800.0 15399.999999999998 ;
      RECT  189800.0 14599.999999999998 190600.00000000003 15399.999999999998 ;
      RECT  194600.0 14599.999999999998 195400.0 15399.999999999998 ;
      RECT  199399.99999999997 14599.999999999998 200200.0 15399.999999999998 ;
      RECT  204200.0 14599.999999999998 205000.0 15399.999999999998 ;
      RECT  209000.0 14599.999999999998 209800.0 15399.999999999998 ;
      RECT  7400.000000000003 19400.000000000004 8200.000000000004 20200.000000000004 ;
      RECT  12200.0 19400.000000000004 13000.0 20200.000000000004 ;
      RECT  16999.999999999996 19400.000000000004 17799.999999999996 20200.000000000004 ;
      RECT  21799.999999999993 19400.000000000004 22599.999999999993 20200.000000000004 ;
      RECT  26599.999999999996 19400.000000000004 27400.0 20200.000000000004 ;
      RECT  31399.999999999996 19400.000000000004 32199.999999999996 20200.000000000004 ;
      RECT  36200.0 19400.000000000004 37000.0 20200.000000000004 ;
      RECT  41000.0 19400.000000000004 41800.0 20200.000000000004 ;
      RECT  45800.0 19400.000000000004 46599.99999999999 20200.000000000004 ;
      RECT  50600.0 19400.000000000004 51400.0 20200.000000000004 ;
      RECT  55400.00000000001 19400.000000000004 56200.0 20200.000000000004 ;
      RECT  60200.0 19400.000000000004 61000.0 20200.000000000004 ;
      RECT  79400.0 19400.000000000004 80200.0 20200.000000000004 ;
      RECT  84200.0 19400.000000000004 85000.0 20200.000000000004 ;
      RECT  89000.0 19400.000000000004 89800.0 20200.000000000004 ;
      RECT  93800.0 19400.000000000004 94600.0 20200.000000000004 ;
      RECT  98600.00000000001 19400.000000000004 99400.0 20200.000000000004 ;
      RECT  103400.0 19400.000000000004 104200.0 20200.000000000004 ;
      RECT  108200.0 19400.000000000004 109000.0 20200.000000000004 ;
      RECT  113000.00000000001 19400.000000000004 113800.00000000001 20200.000000000004 ;
      RECT  117800.0 19400.000000000004 118600.0 20200.000000000004 ;
      RECT  122600.00000000001 19400.000000000004 123400.0 20200.000000000004 ;
      RECT  127400.0 19400.000000000004 128199.99999999999 20200.000000000004 ;
      RECT  132200.0 19400.000000000004 133000.0 20200.000000000004 ;
      RECT  137000.0 19400.000000000004 137800.0 20200.000000000004 ;
      RECT  141800.0 19400.000000000004 142600.00000000003 20200.000000000004 ;
      RECT  146600.0 19400.000000000004 147400.0 20200.000000000004 ;
      RECT  151399.99999999997 19400.000000000004 152200.0 20200.000000000004 ;
      RECT  156200.0 19400.000000000004 157000.0 20200.000000000004 ;
      RECT  161000.0 19400.000000000004 161800.0 20200.000000000004 ;
      RECT  165800.0 19400.000000000004 166600.00000000003 20200.000000000004 ;
      RECT  170600.0 19400.000000000004 171400.0 20200.000000000004 ;
      RECT  175399.99999999997 19400.000000000004 176200.0 20200.000000000004 ;
      RECT  180200.0 19400.000000000004 181000.0 20200.000000000004 ;
      RECT  185000.0 19400.000000000004 185800.0 20200.000000000004 ;
      RECT  189800.0 19400.000000000004 190600.00000000003 20200.000000000004 ;
      RECT  194600.0 19400.000000000004 195400.0 20200.000000000004 ;
      RECT  199399.99999999997 19400.000000000004 200200.0 20200.000000000004 ;
      RECT  204200.0 19400.000000000004 205000.0 20200.000000000004 ;
      RECT  209000.0 19400.000000000004 209800.0 20200.000000000004 ;
      RECT  7400.000000000003 24200.0 8200.000000000004 25000.0 ;
      RECT  12200.0 24200.0 13000.0 25000.0 ;
      RECT  16999.999999999996 24200.0 17799.999999999996 25000.0 ;
      RECT  21799.999999999993 24200.0 22599.999999999993 25000.0 ;
      RECT  26599.999999999996 24200.0 27400.0 25000.0 ;
      RECT  31399.999999999996 24200.0 32199.999999999996 25000.0 ;
      RECT  36200.0 24200.0 37000.0 25000.0 ;
      RECT  41000.0 24200.0 41800.0 25000.0 ;
      RECT  45800.0 24200.0 46599.99999999999 25000.0 ;
      RECT  50600.0 24200.0 51400.0 25000.0 ;
      RECT  55400.00000000001 24200.0 56200.0 25000.0 ;
      RECT  60200.0 24200.0 61000.0 25000.0 ;
      RECT  65000.0 24200.0 65800.0 25000.0 ;
      RECT  69800.0 24200.0 70600.0 25000.0 ;
      RECT  74600.00000000001 24200.0 75400.0 25000.0 ;
      RECT  79400.0 24200.0 80200.0 25000.0 ;
      RECT  84200.0 24200.0 85000.0 25000.0 ;
      RECT  89000.0 24200.0 89800.0 25000.0 ;
      RECT  93800.0 24200.0 94600.0 25000.0 ;
      RECT  98600.00000000001 24200.0 99400.0 25000.0 ;
      RECT  103400.0 24200.0 104200.0 25000.0 ;
      RECT  108200.0 24200.0 109000.0 25000.0 ;
      RECT  113000.00000000001 24200.0 113800.00000000001 25000.0 ;
      RECT  117800.0 24200.0 118600.0 25000.0 ;
      RECT  122600.00000000001 24200.0 123400.0 25000.0 ;
      RECT  127400.0 24200.0 128199.99999999999 25000.0 ;
      RECT  132200.0 24200.0 133000.0 25000.0 ;
      RECT  137000.0 24200.0 137800.0 25000.0 ;
      RECT  141800.0 24200.0 142600.00000000003 25000.0 ;
      RECT  146600.0 24200.0 147400.0 25000.0 ;
      RECT  151399.99999999997 24200.0 152200.0 25000.0 ;
      RECT  156200.0 24200.0 157000.0 25000.0 ;
      RECT  161000.0 24200.0 161800.0 25000.0 ;
      RECT  165800.0 24200.0 166600.00000000003 25000.0 ;
      RECT  170600.0 24200.0 171400.0 25000.0 ;
      RECT  175399.99999999997 24200.0 176200.0 25000.0 ;
      RECT  180200.0 24200.0 181000.0 25000.0 ;
      RECT  185000.0 24200.0 185800.0 25000.0 ;
      RECT  189800.0 24200.0 190600.00000000003 25000.0 ;
      RECT  194600.0 24200.0 195400.0 25000.0 ;
      RECT  199399.99999999997 24200.0 200200.0 25000.0 ;
      RECT  204200.0 24200.0 205000.0 25000.0 ;
      RECT  209000.0 24200.0 209800.0 25000.0 ;
      RECT  45800.0 28999.999999999996 46599.99999999999 29799.999999999996 ;
      RECT  50600.0 28999.999999999996 51400.0 29799.999999999996 ;
      RECT  55400.00000000001 28999.999999999996 56200.0 29799.999999999996 ;
      RECT  60200.0 28999.999999999996 61000.0 29799.999999999996 ;
      RECT  65000.0 28999.999999999996 65800.0 29799.999999999996 ;
      RECT  69800.0 28999.999999999996 70600.0 29799.999999999996 ;
      RECT  74600.00000000001 28999.999999999996 75400.0 29799.999999999996 ;
      RECT  79400.0 28999.999999999996 80200.0 29799.999999999996 ;
      RECT  84200.0 28999.999999999996 85000.0 29799.999999999996 ;
      RECT  89000.0 28999.999999999996 89800.0 29799.999999999996 ;
      RECT  93800.0 28999.999999999996 94600.0 29799.999999999996 ;
      RECT  98600.00000000001 28999.999999999996 99400.0 29799.999999999996 ;
      RECT  103400.0 28999.999999999996 104200.0 29799.999999999996 ;
      RECT  108200.0 28999.999999999996 109000.0 29799.999999999996 ;
      RECT  113000.00000000001 28999.999999999996 113800.00000000001 29799.999999999996 ;
      RECT  117800.0 28999.999999999996 118600.0 29799.999999999996 ;
      RECT  122600.00000000001 28999.999999999996 123400.0 29799.999999999996 ;
      RECT  127400.0 28999.999999999996 128199.99999999999 29799.999999999996 ;
      RECT  132200.0 28999.999999999996 133000.0 29799.999999999996 ;
      RECT  137000.0 28999.999999999996 137800.0 29799.999999999996 ;
      RECT  141800.0 28999.999999999996 142600.00000000003 29799.999999999996 ;
      RECT  146600.0 28999.999999999996 147400.0 29799.999999999996 ;
      RECT  151399.99999999997 28999.999999999996 152200.0 29799.999999999996 ;
      RECT  156200.0 28999.999999999996 157000.0 29799.999999999996 ;
      RECT  161000.0 28999.999999999996 161800.0 29799.999999999996 ;
      RECT  165800.0 28999.999999999996 166600.00000000003 29799.999999999996 ;
      RECT  170600.0 28999.999999999996 171400.0 29799.999999999996 ;
      RECT  175399.99999999997 28999.999999999996 176200.0 29799.999999999996 ;
      RECT  180200.0 28999.999999999996 181000.0 29799.999999999996 ;
      RECT  185000.0 28999.999999999996 185800.0 29799.999999999996 ;
      RECT  189800.0 28999.999999999996 190600.00000000003 29799.999999999996 ;
      RECT  194600.0 28999.999999999996 195400.0 29799.999999999996 ;
      RECT  199399.99999999997 28999.999999999996 200200.0 29799.999999999996 ;
      RECT  204200.0 28999.999999999996 205000.0 29799.999999999996 ;
      RECT  209000.0 28999.999999999996 209800.0 29799.999999999996 ;
      RECT  7400.000000000003 33800.00000000001 8200.000000000004 34600.0 ;
      RECT  12200.0 33800.00000000001 13000.0 34600.0 ;
      RECT  16999.999999999996 33800.00000000001 17799.999999999996 34600.0 ;
      RECT  21799.999999999993 33800.00000000001 22599.999999999993 34600.0 ;
      RECT  26599.999999999996 33800.00000000001 27400.0 34600.0 ;
      RECT  50600.0 33800.00000000001 51400.0 34600.0 ;
      RECT  55400.00000000001 33800.00000000001 56200.0 34600.0 ;
      RECT  60200.0 33800.00000000001 61000.0 34600.0 ;
      RECT  65000.0 33800.00000000001 65800.0 34600.0 ;
      RECT  69800.0 33800.00000000001 70600.0 34600.0 ;
      RECT  74600.00000000001 33800.00000000001 75400.0 34600.0 ;
      RECT  79400.0 33800.00000000001 80200.0 34600.0 ;
      RECT  84200.0 33800.00000000001 85000.0 34600.0 ;
      RECT  89000.0 33800.00000000001 89800.0 34600.0 ;
      RECT  93800.0 33800.00000000001 94600.0 34600.0 ;
      RECT  98600.00000000001 33800.00000000001 99400.0 34600.0 ;
      RECT  103400.0 33800.00000000001 104200.0 34600.0 ;
      RECT  108200.0 33800.00000000001 109000.0 34600.0 ;
      RECT  113000.00000000001 33800.00000000001 113800.00000000001 34600.0 ;
      RECT  117800.0 33800.00000000001 118600.0 34600.0 ;
      RECT  122600.00000000001 33800.00000000001 123400.0 34600.0 ;
      RECT  127400.0 33800.00000000001 128199.99999999999 34600.0 ;
      RECT  132200.0 33800.00000000001 133000.0 34600.0 ;
      RECT  137000.0 33800.00000000001 137800.0 34600.0 ;
      RECT  141800.0 33800.00000000001 142600.00000000003 34600.0 ;
      RECT  146600.0 33800.00000000001 147400.0 34600.0 ;
      RECT  151399.99999999997 33800.00000000001 152200.0 34600.0 ;
      RECT  156200.0 33800.00000000001 157000.0 34600.0 ;
      RECT  161000.0 33800.00000000001 161800.0 34600.0 ;
      RECT  165800.0 33800.00000000001 166600.00000000003 34600.0 ;
      RECT  170600.0 33800.00000000001 171400.0 34600.0 ;
      RECT  175399.99999999997 33800.00000000001 176200.0 34600.0 ;
      RECT  180200.0 33800.00000000001 181000.0 34600.0 ;
      RECT  185000.0 33800.00000000001 185800.0 34600.0 ;
      RECT  189800.0 33800.00000000001 190600.00000000003 34600.0 ;
      RECT  194600.0 33800.00000000001 195400.0 34600.0 ;
      RECT  199399.99999999997 33800.00000000001 200200.0 34600.0 ;
      RECT  204200.0 33800.00000000001 205000.0 34600.0 ;
      RECT  209000.0 33800.00000000001 209800.0 34600.0 ;
      RECT  7400.000000000003 38600.00000000001 8200.000000000004 39400.00000000001 ;
      RECT  12200.0 38600.00000000001 13000.0 39400.00000000001 ;
      RECT  16999.999999999996 38600.00000000001 17799.999999999996 39400.00000000001 ;
      RECT  21799.999999999993 38600.00000000001 22599.999999999993 39400.00000000001 ;
      RECT  26599.999999999996 38600.00000000001 27400.0 39400.00000000001 ;
      RECT  31399.999999999996 38600.00000000001 32199.999999999996 39400.00000000001 ;
      RECT  36200.0 38600.00000000001 37000.0 39400.00000000001 ;
      RECT  41000.0 38600.00000000001 41800.0 39400.00000000001 ;
      RECT  45800.0 38600.00000000001 46599.99999999999 39400.00000000001 ;
      RECT  50600.0 38600.00000000001 51400.0 39400.00000000001 ;
      RECT  55400.00000000001 38600.00000000001 56200.0 39400.00000000001 ;
      RECT  60200.0 38600.00000000001 61000.0 39400.00000000001 ;
      RECT  65000.0 38600.00000000001 65800.0 39400.00000000001 ;
      RECT  69800.0 38600.00000000001 70600.0 39400.00000000001 ;
      RECT  74600.00000000001 38600.00000000001 75400.0 39400.00000000001 ;
      RECT  79400.0 38600.00000000001 80200.0 39400.00000000001 ;
      RECT  84200.0 38600.00000000001 85000.0 39400.00000000001 ;
      RECT  89000.0 38600.00000000001 89800.0 39400.00000000001 ;
      RECT  93800.0 38600.00000000001 94600.0 39400.00000000001 ;
      RECT  98600.00000000001 38600.00000000001 99400.0 39400.00000000001 ;
      RECT  103400.0 38600.00000000001 104200.0 39400.00000000001 ;
      RECT  108200.0 38600.00000000001 109000.0 39400.00000000001 ;
      RECT  113000.00000000001 38600.00000000001 113800.00000000001 39400.00000000001 ;
      RECT  117800.0 38600.00000000001 118600.0 39400.00000000001 ;
      RECT  122600.00000000001 38600.00000000001 123400.0 39400.00000000001 ;
      RECT  127400.0 38600.00000000001 128199.99999999999 39400.00000000001 ;
      RECT  132200.0 38600.00000000001 133000.0 39400.00000000001 ;
      RECT  137000.0 38600.00000000001 137800.0 39400.00000000001 ;
      RECT  141800.0 38600.00000000001 142600.00000000003 39400.00000000001 ;
      RECT  146600.0 38600.00000000001 147400.0 39400.00000000001 ;
      RECT  151399.99999999997 38600.00000000001 152200.0 39400.00000000001 ;
      RECT  156200.0 38600.00000000001 157000.0 39400.00000000001 ;
      RECT  161000.0 38600.00000000001 161800.0 39400.00000000001 ;
      RECT  165800.0 38600.00000000001 166600.00000000003 39400.00000000001 ;
      RECT  170600.0 38600.00000000001 171400.0 39400.00000000001 ;
      RECT  175399.99999999997 38600.00000000001 176200.0 39400.00000000001 ;
      RECT  180200.0 38600.00000000001 181000.0 39400.00000000001 ;
      RECT  185000.0 38600.00000000001 185800.0 39400.00000000001 ;
      RECT  189800.0 38600.00000000001 190600.00000000003 39400.00000000001 ;
      RECT  194600.0 38600.00000000001 195400.0 39400.00000000001 ;
      RECT  199399.99999999997 38600.00000000001 200200.0 39400.00000000001 ;
      RECT  204200.0 38600.00000000001 205000.0 39400.00000000001 ;
      RECT  209000.0 38600.00000000001 209800.0 39400.00000000001 ;
      RECT  7400.000000000003 43400.00000000001 8200.000000000004 44200.0 ;
      RECT  12200.0 43400.00000000001 13000.0 44200.0 ;
      RECT  16999.999999999996 43400.00000000001 17799.999999999996 44200.0 ;
      RECT  21799.999999999993 43400.00000000001 22599.999999999993 44200.0 ;
      RECT  26599.999999999996 43400.00000000001 27400.0 44200.0 ;
      RECT  31399.999999999996 43400.00000000001 32199.999999999996 44200.0 ;
      RECT  36200.0 43400.00000000001 37000.0 44200.0 ;
      RECT  41000.0 43400.00000000001 41800.0 44200.0 ;
      RECT  45800.0 43400.00000000001 46599.99999999999 44200.0 ;
      RECT  50600.0 43400.00000000001 51400.0 44200.0 ;
      RECT  55400.00000000001 43400.00000000001 56200.0 44200.0 ;
      RECT  60200.0 43400.00000000001 61000.0 44200.0 ;
      RECT  65000.0 43400.00000000001 65800.0 44200.0 ;
      RECT  69800.0 43400.00000000001 70600.0 44200.0 ;
      RECT  74600.00000000001 43400.00000000001 75400.0 44200.0 ;
      RECT  79400.0 43400.00000000001 80200.0 44200.0 ;
      RECT  84200.0 43400.00000000001 85000.0 44200.0 ;
      RECT  89000.0 43400.00000000001 89800.0 44200.0 ;
      RECT  93800.0 43400.00000000001 94600.0 44200.0 ;
      RECT  98600.00000000001 43400.00000000001 99400.0 44200.0 ;
      RECT  103400.0 43400.00000000001 104200.0 44200.0 ;
      RECT  108200.0 43400.00000000001 109000.0 44200.0 ;
      RECT  113000.00000000001 43400.00000000001 113800.00000000001 44200.0 ;
      RECT  117800.0 43400.00000000001 118600.0 44200.0 ;
      RECT  122600.00000000001 43400.00000000001 123400.0 44200.0 ;
      RECT  127400.0 43400.00000000001 128199.99999999999 44200.0 ;
      RECT  132200.0 43400.00000000001 133000.0 44200.0 ;
      RECT  137000.0 43400.00000000001 137800.0 44200.0 ;
      RECT  141800.0 43400.00000000001 142600.00000000003 44200.0 ;
      RECT  146600.0 43400.00000000001 147400.0 44200.0 ;
      RECT  151399.99999999997 43400.00000000001 152200.0 44200.0 ;
      RECT  156200.0 43400.00000000001 157000.0 44200.0 ;
      RECT  161000.0 43400.00000000001 161800.0 44200.0 ;
      RECT  165800.0 43400.00000000001 166600.00000000003 44200.0 ;
      RECT  170600.0 43400.00000000001 171400.0 44200.0 ;
      RECT  175399.99999999997 43400.00000000001 176200.0 44200.0 ;
      RECT  180200.0 43400.00000000001 181000.0 44200.0 ;
      RECT  185000.0 43400.00000000001 185800.0 44200.0 ;
      RECT  189800.0 43400.00000000001 190600.00000000003 44200.0 ;
      RECT  194600.0 43400.00000000001 195400.0 44200.0 ;
      RECT  199399.99999999997 43400.00000000001 200200.0 44200.0 ;
      RECT  204200.0 43400.00000000001 205000.0 44200.0 ;
      RECT  209000.0 43400.00000000001 209800.0 44200.0 ;
      RECT  7400.000000000003 48200.0 8200.000000000004 49000.0 ;
      RECT  12200.0 48200.0 13000.0 49000.0 ;
      RECT  16999.999999999996 48200.0 17799.999999999996 49000.0 ;
      RECT  21799.999999999993 48200.0 22599.999999999993 49000.0 ;
      RECT  26599.999999999996 48200.0 27400.0 49000.0 ;
      RECT  31399.999999999996 48200.0 32199.999999999996 49000.0 ;
      RECT  36200.0 48200.0 37000.0 49000.0 ;
      RECT  41000.0 48200.0 41800.0 49000.0 ;
      RECT  45800.0 48200.0 46599.99999999999 49000.0 ;
      RECT  50600.0 48200.0 51400.0 49000.0 ;
      RECT  55400.00000000001 48200.0 56200.0 49000.0 ;
      RECT  60200.0 48200.0 61000.0 49000.0 ;
      RECT  65000.0 48200.0 65800.0 49000.0 ;
      RECT  7400.000000000003 53000.0 8200.000000000004 53800.0 ;
      RECT  12200.0 53000.0 13000.0 53800.0 ;
      RECT  16999.999999999996 53000.0 17799.999999999996 53800.0 ;
      RECT  21799.999999999993 53000.0 22599.999999999993 53800.0 ;
      RECT  26599.999999999996 53000.0 27400.0 53800.0 ;
      RECT  31399.999999999996 53000.0 32199.999999999996 53800.0 ;
      RECT  36200.0 53000.0 37000.0 53800.0 ;
      RECT  41000.0 53000.0 41800.0 53800.0 ;
      RECT  45800.0 53000.0 46599.99999999999 53800.0 ;
      RECT  50600.0 53000.0 51400.0 53800.0 ;
      RECT  55400.00000000001 53000.0 56200.0 53800.0 ;
      RECT  60200.0 53000.0 61000.0 53800.0 ;
      RECT  65000.0 53000.0 65800.0 53800.0 ;
      RECT  69800.0 53000.0 70600.0 53800.0 ;
      RECT  74600.00000000001 53000.0 75400.0 53800.0 ;
      RECT  79400.0 53000.0 80200.0 53800.0 ;
      RECT  84200.0 53000.0 85000.0 53800.0 ;
      RECT  89000.0 53000.0 89800.0 53800.0 ;
      RECT  93800.0 53000.0 94600.0 53800.0 ;
      RECT  98600.00000000001 53000.0 99400.0 53800.0 ;
      RECT  103400.0 53000.0 104200.0 53800.0 ;
      RECT  108200.0 53000.0 109000.0 53800.0 ;
      RECT  113000.00000000001 53000.0 113800.00000000001 53800.0 ;
      RECT  117800.0 53000.0 118600.0 53800.0 ;
      RECT  122600.00000000001 53000.0 123400.0 53800.0 ;
      RECT  127400.0 53000.0 128199.99999999999 53800.0 ;
      RECT  132200.0 53000.0 133000.0 53800.0 ;
      RECT  137000.0 53000.0 137800.0 53800.0 ;
      RECT  141800.0 53000.0 142600.00000000003 53800.0 ;
      RECT  146600.0 53000.0 147400.0 53800.0 ;
      RECT  151399.99999999997 53000.0 152200.0 53800.0 ;
      RECT  156200.0 53000.0 157000.0 53800.0 ;
      RECT  161000.0 53000.0 161800.0 53800.0 ;
      RECT  165800.0 53000.0 166600.00000000003 53800.0 ;
      RECT  170600.0 53000.0 171400.0 53800.0 ;
      RECT  175399.99999999997 53000.0 176200.0 53800.0 ;
      RECT  180200.0 53000.0 181000.0 53800.0 ;
      RECT  185000.0 53000.0 185800.0 53800.0 ;
      RECT  189800.0 53000.0 190600.00000000003 53800.0 ;
      RECT  194600.0 53000.0 195400.0 53800.0 ;
      RECT  199399.99999999997 53000.0 200200.0 53800.0 ;
      RECT  204200.0 53000.0 205000.0 53800.0 ;
      RECT  209000.0 53000.0 209800.0 53800.0 ;
      RECT  7400.000000000003 57800.00000000001 8200.000000000004 58600.0 ;
      RECT  12200.0 57800.00000000001 13000.0 58600.0 ;
      RECT  16999.999999999996 57800.00000000001 17799.999999999996 58600.0 ;
      RECT  21799.999999999993 57800.00000000001 22599.999999999993 58600.0 ;
      RECT  26599.999999999996 57800.00000000001 27400.0 58600.0 ;
      RECT  31399.999999999996 57800.00000000001 32199.999999999996 58600.0 ;
      RECT  36200.0 57800.00000000001 37000.0 58600.0 ;
      RECT  41000.0 57800.00000000001 41800.0 58600.0 ;
      RECT  45800.0 57800.00000000001 46599.99999999999 58600.0 ;
      RECT  50600.0 57800.00000000001 51400.0 58600.0 ;
      RECT  55400.00000000001 57800.00000000001 56200.0 58600.0 ;
      RECT  60200.0 57800.00000000001 61000.0 58600.0 ;
      RECT  65000.0 57800.00000000001 65800.0 58600.0 ;
      RECT  69800.0 57800.00000000001 70600.0 58600.0 ;
      RECT  74600.00000000001 57800.00000000001 75400.0 58600.0 ;
      RECT  79400.0 57800.00000000001 80200.0 58600.0 ;
      RECT  84200.0 57800.00000000001 85000.0 58600.0 ;
      RECT  89000.0 57800.00000000001 89800.0 58600.0 ;
      RECT  93800.0 57800.00000000001 94600.0 58600.0 ;
      RECT  98600.00000000001 57800.00000000001 99400.0 58600.0 ;
      RECT  103400.0 57800.00000000001 104200.0 58600.0 ;
      RECT  108200.0 57800.00000000001 109000.0 58600.0 ;
      RECT  113000.00000000001 57800.00000000001 113800.00000000001 58600.0 ;
      RECT  117800.0 57800.00000000001 118600.0 58600.0 ;
      RECT  122600.00000000001 57800.00000000001 123400.0 58600.0 ;
      RECT  127400.0 57800.00000000001 128199.99999999999 58600.0 ;
      RECT  132200.0 57800.00000000001 133000.0 58600.0 ;
      RECT  137000.0 57800.00000000001 137800.0 58600.0 ;
      RECT  141800.0 57800.00000000001 142600.00000000003 58600.0 ;
      RECT  146600.0 57800.00000000001 147400.0 58600.0 ;
      RECT  151399.99999999997 57800.00000000001 152200.0 58600.0 ;
      RECT  156200.0 57800.00000000001 157000.0 58600.0 ;
      RECT  161000.0 57800.00000000001 161800.0 58600.0 ;
      RECT  165800.0 57800.00000000001 166600.00000000003 58600.0 ;
      RECT  170600.0 57800.00000000001 171400.0 58600.0 ;
      RECT  175399.99999999997 57800.00000000001 176200.0 58600.0 ;
      RECT  180200.0 57800.00000000001 181000.0 58600.0 ;
      RECT  185000.0 57800.00000000001 185800.0 58600.0 ;
      RECT  189800.0 57800.00000000001 190600.00000000003 58600.0 ;
      RECT  194600.0 57800.00000000001 195400.0 58600.0 ;
      RECT  199399.99999999997 57800.00000000001 200200.0 58600.0 ;
      RECT  204200.0 57800.00000000001 205000.0 58600.0 ;
      RECT  209000.0 57800.00000000001 209800.0 58600.0 ;
      RECT  7400.000000000003 62600.00000000001 8200.000000000004 63400.00000000001 ;
      RECT  12200.0 62600.00000000001 13000.0 63400.00000000001 ;
      RECT  16999.999999999996 62600.00000000001 17799.999999999996 63400.00000000001 ;
      RECT  21799.999999999993 62600.00000000001 22599.999999999993 63400.00000000001 ;
      RECT  26599.999999999996 62600.00000000001 27400.0 63400.00000000001 ;
      RECT  31399.999999999996 62600.00000000001 32199.999999999996 63400.00000000001 ;
      RECT  36200.0 62600.00000000001 37000.0 63400.00000000001 ;
      RECT  41000.0 62600.00000000001 41800.0 63400.00000000001 ;
      RECT  45800.0 62600.00000000001 46599.99999999999 63400.00000000001 ;
      RECT  50600.0 62600.00000000001 51400.0 63400.00000000001 ;
      RECT  55400.00000000001 62600.00000000001 56200.0 63400.00000000001 ;
      RECT  60200.0 62600.00000000001 61000.0 63400.00000000001 ;
      RECT  79400.0 62600.00000000001 80200.0 63400.00000000001 ;
      RECT  84200.0 62600.00000000001 85000.0 63400.00000000001 ;
      RECT  89000.0 62600.00000000001 89800.0 63400.00000000001 ;
      RECT  93800.0 62600.00000000001 94600.0 63400.00000000001 ;
      RECT  98600.00000000001 62600.00000000001 99400.0 63400.00000000001 ;
      RECT  103400.0 62600.00000000001 104200.0 63400.00000000001 ;
      RECT  108200.0 62600.00000000001 109000.0 63400.00000000001 ;
      RECT  113000.00000000001 62600.00000000001 113800.00000000001 63400.00000000001 ;
      RECT  117800.0 62600.00000000001 118600.0 63400.00000000001 ;
      RECT  122600.00000000001 62600.00000000001 123400.0 63400.00000000001 ;
      RECT  127400.0 62600.00000000001 128199.99999999999 63400.00000000001 ;
      RECT  132200.0 62600.00000000001 133000.0 63400.00000000001 ;
      RECT  137000.0 62600.00000000001 137800.0 63400.00000000001 ;
      RECT  141800.0 62600.00000000001 142600.00000000003 63400.00000000001 ;
      RECT  146600.0 62600.00000000001 147400.0 63400.00000000001 ;
      RECT  151399.99999999997 62600.00000000001 152200.0 63400.00000000001 ;
      RECT  156200.0 62600.00000000001 157000.0 63400.00000000001 ;
      RECT  161000.0 62600.00000000001 161800.0 63400.00000000001 ;
      RECT  165800.0 62600.00000000001 166600.00000000003 63400.00000000001 ;
      RECT  170600.0 62600.00000000001 171400.0 63400.00000000001 ;
      RECT  175399.99999999997 62600.00000000001 176200.0 63400.00000000001 ;
      RECT  7400.000000000003 67400.0 8200.000000000004 68200.0 ;
      RECT  12200.0 67400.0 13000.0 68200.0 ;
      RECT  16999.999999999996 67400.0 17799.999999999996 68200.0 ;
      RECT  21799.999999999993 67400.0 22599.999999999993 68200.0 ;
      RECT  26599.999999999996 67400.0 27400.0 68200.0 ;
      RECT  31399.999999999996 67400.0 32199.999999999996 68200.0 ;
      RECT  36200.0 67400.0 37000.0 68200.0 ;
      RECT  41000.0 67400.0 41800.0 68200.0 ;
      RECT  45800.0 67400.0 46599.99999999999 68200.0 ;
      RECT  50600.0 67400.0 51400.0 68200.0 ;
      RECT  55400.00000000001 67400.0 56200.0 68200.0 ;
      RECT  60200.0 67400.0 61000.0 68200.0 ;
      RECT  65000.0 67400.0 65800.0 68200.0 ;
      RECT  69800.0 67400.0 70600.0 68200.0 ;
      RECT  74600.00000000001 67400.0 75400.0 68200.0 ;
      RECT  79400.0 67400.0 80200.0 68200.0 ;
      RECT  84200.0 67400.0 85000.0 68200.0 ;
      RECT  89000.0 67400.0 89800.0 68200.0 ;
      RECT  93800.0 67400.0 94600.0 68200.0 ;
      RECT  98600.00000000001 67400.0 99400.0 68200.0 ;
      RECT  103400.0 67400.0 104200.0 68200.0 ;
      RECT  108200.0 67400.0 109000.0 68200.0 ;
      RECT  113000.00000000001 67400.0 113800.00000000001 68200.0 ;
      RECT  117800.0 67400.0 118600.0 68200.0 ;
      RECT  122600.00000000001 67400.0 123400.0 68200.0 ;
      RECT  127400.0 67400.0 128199.99999999999 68200.0 ;
      RECT  132200.0 67400.0 133000.0 68200.0 ;
      RECT  137000.0 67400.0 137800.0 68200.0 ;
      RECT  141800.0 67400.0 142600.00000000003 68200.0 ;
      RECT  146600.0 67400.0 147400.0 68200.0 ;
      RECT  151399.99999999997 67400.0 152200.0 68200.0 ;
      RECT  156200.0 67400.0 157000.0 68200.0 ;
      RECT  161000.0 67400.0 161800.0 68200.0 ;
      RECT  165800.0 67400.0 166600.00000000003 68200.0 ;
      RECT  170600.0 67400.0 171400.0 68200.0 ;
      RECT  175399.99999999997 67400.0 176200.0 68200.0 ;
      RECT  180200.0 67400.0 181000.0 68200.0 ;
      RECT  185000.0 67400.0 185800.0 68200.0 ;
      RECT  189800.0 67400.0 190600.00000000003 68200.0 ;
      RECT  194600.0 67400.0 195400.0 68200.0 ;
      RECT  199399.99999999997 67400.0 200200.0 68200.0 ;
      RECT  204200.0 67400.0 205000.0 68200.0 ;
      RECT  209000.0 67400.0 209800.0 68200.0 ;
      RECT  7400.000000000003 72200.0 8200.000000000004 73000.0 ;
      RECT  12200.0 72200.0 13000.0 73000.0 ;
      RECT  16999.999999999996 72200.0 17799.999999999996 73000.0 ;
      RECT  21799.999999999993 72200.0 22599.999999999993 73000.0 ;
      RECT  26599.999999999996 72200.0 27400.0 73000.0 ;
      RECT  31399.999999999996 72200.0 32199.999999999996 73000.0 ;
      RECT  36200.0 72200.0 37000.0 73000.0 ;
      RECT  41000.0 72200.0 41800.0 73000.0 ;
      RECT  45800.0 72200.0 46599.99999999999 73000.0 ;
      RECT  50600.0 72200.0 51400.0 73000.0 ;
      RECT  55400.00000000001 72200.0 56200.0 73000.0 ;
      RECT  60200.0 72200.0 61000.0 73000.0 ;
      RECT  65000.0 72200.0 65800.0 73000.0 ;
      RECT  175399.99999999997 72200.0 176200.0 73000.0 ;
      RECT  180200.0 72200.0 181000.0 73000.0 ;
      RECT  185000.0 72200.0 185800.0 73000.0 ;
      RECT  189800.0 72200.0 190600.00000000003 73000.0 ;
      RECT  194600.0 72200.0 195400.0 73000.0 ;
      RECT  199399.99999999997 72200.0 200200.0 73000.0 ;
      RECT  204200.0 72200.0 205000.0 73000.0 ;
      RECT  209000.0 72200.0 209800.0 73000.0 ;
      RECT  7400.000000000003 77000.0 8200.000000000004 77800.0 ;
      RECT  12200.0 77000.0 13000.0 77800.0 ;
      RECT  16999.999999999996 77000.0 17799.999999999996 77800.0 ;
      RECT  21799.999999999993 77000.0 22599.999999999993 77800.0 ;
      RECT  26599.999999999996 77000.0 27400.0 77800.0 ;
      RECT  31399.999999999996 77000.0 32199.999999999996 77800.0 ;
      RECT  36200.0 77000.0 37000.0 77800.0 ;
      RECT  41000.0 77000.0 41800.0 77800.0 ;
      RECT  45800.0 77000.0 46599.99999999999 77800.0 ;
      RECT  50600.0 77000.0 51400.0 77800.0 ;
      RECT  55400.00000000001 77000.0 56200.0 77800.0 ;
      RECT  60200.0 77000.0 61000.0 77800.0 ;
      RECT  65000.0 77000.0 65800.0 77800.0 ;
      RECT  69800.0 77000.0 70600.0 77800.0 ;
      RECT  74600.00000000001 77000.0 75400.0 77800.0 ;
      RECT  79400.0 77000.0 80200.0 77800.0 ;
      RECT  84200.0 77000.0 85000.0 77800.0 ;
      RECT  89000.0 77000.0 89800.0 77800.0 ;
      RECT  93800.0 77000.0 94600.0 77800.0 ;
      RECT  98600.00000000001 77000.0 99400.0 77800.0 ;
      RECT  103400.0 77000.0 104200.0 77800.0 ;
      RECT  108200.0 77000.0 109000.0 77800.0 ;
      RECT  113000.00000000001 77000.0 113800.00000000001 77800.0 ;
      RECT  117800.0 77000.0 118600.0 77800.0 ;
      RECT  122600.00000000001 77000.0 123400.0 77800.0 ;
      RECT  127400.0 77000.0 128199.99999999999 77800.0 ;
      RECT  132200.0 77000.0 133000.0 77800.0 ;
      RECT  137000.0 77000.0 137800.0 77800.0 ;
      RECT  141800.0 77000.0 142600.00000000003 77800.0 ;
      RECT  146600.0 77000.0 147400.0 77800.0 ;
      RECT  151399.99999999997 77000.0 152200.0 77800.0 ;
      RECT  156200.0 77000.0 157000.0 77800.0 ;
      RECT  161000.0 77000.0 161800.0 77800.0 ;
      RECT  165800.0 77000.0 166600.00000000003 77800.0 ;
      RECT  7400.000000000003 81800.00000000001 8200.000000000004 82600.00000000001 ;
      RECT  12200.0 81800.00000000001 13000.0 82600.00000000001 ;
      RECT  16999.999999999996 81800.00000000001 17799.999999999996 82600.00000000001 ;
      RECT  21799.999999999993 81800.00000000001 22599.999999999993 82600.00000000001 ;
      RECT  26599.999999999996 81800.00000000001 27400.0 82600.00000000001 ;
      RECT  31399.999999999996 81800.00000000001 32199.999999999996 82600.00000000001 ;
      RECT  36200.0 81800.00000000001 37000.0 82600.00000000001 ;
      RECT  41000.0 81800.00000000001 41800.0 82600.00000000001 ;
      RECT  45800.0 81800.00000000001 46599.99999999999 82600.00000000001 ;
      RECT  50600.0 81800.00000000001 51400.0 82600.00000000001 ;
      RECT  55400.00000000001 81800.00000000001 56200.0 82600.00000000001 ;
      RECT  60200.0 81800.00000000001 61000.0 82600.00000000001 ;
      RECT  65000.0 81800.00000000001 65800.0 82600.00000000001 ;
      RECT  69800.0 81800.00000000001 70600.0 82600.00000000001 ;
      RECT  74600.00000000001 81800.00000000001 75400.0 82600.00000000001 ;
      RECT  79400.0 81800.00000000001 80200.0 82600.00000000001 ;
      RECT  84200.0 81800.00000000001 85000.0 82600.00000000001 ;
      RECT  89000.0 81800.00000000001 89800.0 82600.00000000001 ;
      RECT  93800.0 81800.00000000001 94600.0 82600.00000000001 ;
      RECT  98600.00000000001 81800.00000000001 99400.0 82600.00000000001 ;
      RECT  103400.0 81800.00000000001 104200.0 82600.00000000001 ;
      RECT  108200.0 81800.00000000001 109000.0 82600.00000000001 ;
      RECT  113000.00000000001 81800.00000000001 113800.00000000001 82600.00000000001 ;
      RECT  117800.0 81800.00000000001 118600.0 82600.00000000001 ;
      RECT  122600.00000000001 81800.00000000001 123400.0 82600.00000000001 ;
      RECT  127400.0 81800.00000000001 128199.99999999999 82600.00000000001 ;
      RECT  132200.0 81800.00000000001 133000.0 82600.00000000001 ;
      RECT  137000.0 81800.00000000001 137800.0 82600.00000000001 ;
      RECT  141800.0 81800.00000000001 142600.00000000003 82600.00000000001 ;
      RECT  146600.0 81800.00000000001 147400.0 82600.00000000001 ;
      RECT  151399.99999999997 81800.00000000001 152200.0 82600.00000000001 ;
      RECT  156200.0 81800.00000000001 157000.0 82600.00000000001 ;
      RECT  161000.0 81800.00000000001 161800.0 82600.00000000001 ;
      RECT  165800.0 81800.00000000001 166600.00000000003 82600.00000000001 ;
      RECT  170600.0 81800.00000000001 171400.0 82600.00000000001 ;
      RECT  175399.99999999997 81800.00000000001 176200.0 82600.00000000001 ;
      RECT  180200.0 81800.00000000001 181000.0 82600.00000000001 ;
      RECT  185000.0 81800.00000000001 185800.0 82600.00000000001 ;
      RECT  189800.0 81800.00000000001 190600.00000000003 82600.00000000001 ;
      RECT  194600.0 81800.00000000001 195400.0 82600.00000000001 ;
      RECT  199399.99999999997 81800.00000000001 200200.0 82600.00000000001 ;
      RECT  204200.0 81800.00000000001 205000.0 82600.00000000001 ;
      RECT  209000.0 81800.00000000001 209800.0 82600.00000000001 ;
      RECT  7400.000000000003 86600.00000000001 8200.000000000004 87400.0 ;
      RECT  12200.0 86600.00000000001 13000.0 87400.0 ;
      RECT  16999.999999999996 86600.00000000001 17799.999999999996 87400.0 ;
      RECT  21799.999999999993 86600.00000000001 22599.999999999993 87400.0 ;
      RECT  26599.999999999996 86600.00000000001 27400.0 87400.0 ;
      RECT  31399.999999999996 86600.00000000001 32199.999999999996 87400.0 ;
      RECT  36200.0 86600.00000000001 37000.0 87400.0 ;
      RECT  41000.0 86600.00000000001 41800.0 87400.0 ;
      RECT  45800.0 86600.00000000001 46599.99999999999 87400.0 ;
      RECT  50600.0 86600.00000000001 51400.0 87400.0 ;
      RECT  55400.00000000001 86600.00000000001 56200.0 87400.0 ;
      RECT  60200.0 86600.00000000001 61000.0 87400.0 ;
      RECT  65000.0 86600.00000000001 65800.0 87400.0 ;
      RECT  69800.0 86600.00000000001 70600.0 87400.0 ;
      RECT  74600.00000000001 86600.00000000001 75400.0 87400.0 ;
      RECT  79400.0 86600.00000000001 80200.0 87400.0 ;
      RECT  84200.0 86600.00000000001 85000.0 87400.0 ;
      RECT  89000.0 86600.00000000001 89800.0 87400.0 ;
      RECT  93800.0 86600.00000000001 94600.0 87400.0 ;
      RECT  98600.00000000001 86600.00000000001 99400.0 87400.0 ;
      RECT  103400.0 86600.00000000001 104200.0 87400.0 ;
      RECT  108200.0 86600.00000000001 109000.0 87400.0 ;
      RECT  113000.00000000001 86600.00000000001 113800.00000000001 87400.0 ;
      RECT  117800.0 86600.00000000001 118600.0 87400.0 ;
      RECT  122600.00000000001 86600.00000000001 123400.0 87400.0 ;
      RECT  127400.0 86600.00000000001 128199.99999999999 87400.0 ;
      RECT  132200.0 86600.00000000001 133000.0 87400.0 ;
      RECT  137000.0 86600.00000000001 137800.0 87400.0 ;
      RECT  141800.0 86600.00000000001 142600.00000000003 87400.0 ;
      RECT  146600.0 86600.00000000001 147400.0 87400.0 ;
      RECT  151399.99999999997 86600.00000000001 152200.0 87400.0 ;
      RECT  156200.0 86600.00000000001 157000.0 87400.0 ;
      RECT  161000.0 86600.00000000001 161800.0 87400.0 ;
      RECT  165800.0 86600.00000000001 166600.00000000003 87400.0 ;
      RECT  170600.0 86600.00000000001 171400.0 87400.0 ;
      RECT  175399.99999999997 86600.00000000001 176200.0 87400.0 ;
      RECT  180200.0 86600.00000000001 181000.0 87400.0 ;
      RECT  185000.0 86600.00000000001 185800.0 87400.0 ;
      RECT  189800.0 86600.00000000001 190600.00000000003 87400.0 ;
      RECT  194600.0 86600.00000000001 195400.0 87400.0 ;
      RECT  199399.99999999997 86600.00000000001 200200.0 87400.0 ;
      RECT  204200.0 86600.00000000001 205000.0 87400.0 ;
      RECT  209000.0 86600.00000000001 209800.0 87400.0 ;
      RECT  7400.000000000003 91400.0 8200.000000000004 92200.0 ;
      RECT  12200.0 91400.0 13000.0 92200.0 ;
      RECT  16999.999999999996 91400.0 17799.999999999996 92200.0 ;
      RECT  21799.999999999993 91400.0 22599.999999999993 92200.0 ;
      RECT  26599.999999999996 91400.0 27400.0 92200.0 ;
      RECT  31399.999999999996 91400.0 32199.999999999996 92200.0 ;
      RECT  36200.0 91400.0 37000.0 92200.0 ;
      RECT  41000.0 91400.0 41800.0 92200.0 ;
      RECT  45800.0 91400.0 46599.99999999999 92200.0 ;
      RECT  50600.0 91400.0 51400.0 92200.0 ;
      RECT  55400.00000000001 91400.0 56200.0 92200.0 ;
      RECT  60200.0 91400.0 61000.0 92200.0 ;
      RECT  65000.0 91400.0 65800.0 92200.0 ;
      RECT  175399.99999999997 91400.0 176200.0 92200.0 ;
      RECT  180200.0 91400.0 181000.0 92200.0 ;
      RECT  185000.0 91400.0 185800.0 92200.0 ;
      RECT  189800.0 91400.0 190600.00000000003 92200.0 ;
      RECT  194600.0 91400.0 195400.0 92200.0 ;
      RECT  199399.99999999997 91400.0 200200.0 92200.0 ;
      RECT  204200.0 91400.0 205000.0 92200.0 ;
      RECT  209000.0 91400.0 209800.0 92200.0 ;
      RECT  7400.000000000003 96200.0 8200.000000000004 97000.0 ;
      RECT  12200.0 96200.0 13000.0 97000.0 ;
      RECT  16999.999999999996 96200.0 17799.999999999996 97000.0 ;
      RECT  21799.999999999993 96200.0 22599.999999999993 97000.0 ;
      RECT  26599.999999999996 96200.0 27400.0 97000.0 ;
      RECT  31399.999999999996 96200.0 32199.999999999996 97000.0 ;
      RECT  36200.0 96200.0 37000.0 97000.0 ;
      RECT  41000.0 96200.0 41800.0 97000.0 ;
      RECT  45800.0 96200.0 46599.99999999999 97000.0 ;
      RECT  50600.0 96200.0 51400.0 97000.0 ;
      RECT  55400.00000000001 96200.0 56200.0 97000.0 ;
      RECT  60200.0 96200.0 61000.0 97000.0 ;
      RECT  65000.0 96200.0 65800.0 97000.0 ;
      RECT  69800.0 96200.0 70600.0 97000.0 ;
      RECT  74600.00000000001 96200.0 75400.0 97000.0 ;
      RECT  79400.0 96200.0 80200.0 97000.0 ;
      RECT  84200.0 96200.0 85000.0 97000.0 ;
      RECT  89000.0 96200.0 89800.0 97000.0 ;
      RECT  93800.0 96200.0 94600.0 97000.0 ;
      RECT  98600.00000000001 96200.0 99400.0 97000.0 ;
      RECT  103400.0 96200.0 104200.0 97000.0 ;
      RECT  108200.0 96200.0 109000.0 97000.0 ;
      RECT  113000.00000000001 96200.0 113800.00000000001 97000.0 ;
      RECT  117800.0 96200.0 118600.0 97000.0 ;
      RECT  122600.00000000001 96200.0 123400.0 97000.0 ;
      RECT  127400.0 96200.0 128199.99999999999 97000.0 ;
      RECT  132200.0 96200.0 133000.0 97000.0 ;
      RECT  137000.0 96200.0 137800.0 97000.0 ;
      RECT  141800.0 96200.0 142600.00000000003 97000.0 ;
      RECT  146600.0 96200.0 147400.0 97000.0 ;
      RECT  151399.99999999997 96200.0 152200.0 97000.0 ;
      RECT  156200.0 96200.0 157000.0 97000.0 ;
      RECT  161000.0 96200.0 161800.0 97000.0 ;
      RECT  165800.0 96200.0 166600.00000000003 97000.0 ;
      RECT  170600.0 96200.0 171400.0 97000.0 ;
      RECT  175399.99999999997 96200.0 176200.0 97000.0 ;
      RECT  180200.0 96200.0 181000.0 97000.0 ;
      RECT  185000.0 96200.0 185800.0 97000.0 ;
      RECT  189800.0 96200.0 190600.00000000003 97000.0 ;
      RECT  194600.0 96200.0 195400.0 97000.0 ;
      RECT  199399.99999999997 96200.0 200200.0 97000.0 ;
      RECT  204200.0 96200.0 205000.0 97000.0 ;
      RECT  209000.0 96200.0 209800.0 97000.0 ;
      RECT  7400.000000000003 101000.00000000001 8200.000000000004 101800.00000000001 ;
      RECT  12200.0 101000.00000000001 13000.0 101800.00000000001 ;
      RECT  16999.999999999996 101000.00000000001 17799.999999999996 101800.00000000001 ;
      RECT  21799.999999999993 101000.00000000001 22599.999999999993 101800.00000000001 ;
      RECT  26599.999999999996 101000.00000000001 27400.0 101800.00000000001 ;
      RECT  31399.999999999996 101000.00000000001 32199.999999999996 101800.00000000001 ;
      RECT  36200.0 101000.00000000001 37000.0 101800.00000000001 ;
      RECT  41000.0 101000.00000000001 41800.0 101800.00000000001 ;
      RECT  45800.0 101000.00000000001 46599.99999999999 101800.00000000001 ;
      RECT  50600.0 101000.00000000001 51400.0 101800.00000000001 ;
      RECT  55400.00000000001 101000.00000000001 56200.0 101800.00000000001 ;
      RECT  60200.0 101000.00000000001 61000.0 101800.00000000001 ;
      RECT  79400.0 101000.00000000001 80200.0 101800.00000000001 ;
      RECT  84200.0 101000.00000000001 85000.0 101800.00000000001 ;
      RECT  89000.0 101000.00000000001 89800.0 101800.00000000001 ;
      RECT  93800.0 101000.00000000001 94600.0 101800.00000000001 ;
      RECT  98600.00000000001 101000.00000000001 99400.0 101800.00000000001 ;
      RECT  103400.0 101000.00000000001 104200.0 101800.00000000001 ;
      RECT  108200.0 101000.00000000001 109000.0 101800.00000000001 ;
      RECT  113000.00000000001 101000.00000000001 113800.00000000001 101800.00000000001 ;
      RECT  117800.0 101000.00000000001 118600.0 101800.00000000001 ;
      RECT  122600.00000000001 101000.00000000001 123400.0 101800.00000000001 ;
      RECT  127400.0 101000.00000000001 128199.99999999999 101800.00000000001 ;
      RECT  132200.0 101000.00000000001 133000.0 101800.00000000001 ;
      RECT  137000.0 101000.00000000001 137800.0 101800.00000000001 ;
      RECT  141800.0 101000.00000000001 142600.00000000003 101800.00000000001 ;
      RECT  146600.0 101000.00000000001 147400.0 101800.00000000001 ;
      RECT  151399.99999999997 101000.00000000001 152200.0 101800.00000000001 ;
      RECT  156200.0 101000.00000000001 157000.0 101800.00000000001 ;
      RECT  161000.0 101000.00000000001 161800.0 101800.00000000001 ;
      RECT  165800.0 101000.00000000001 166600.00000000003 101800.00000000001 ;
      RECT  170600.0 101000.00000000001 171400.0 101800.00000000001 ;
      RECT  175399.99999999997 101000.00000000001 176200.0 101800.00000000001 ;
      RECT  180200.0 101000.00000000001 181000.0 101800.00000000001 ;
      RECT  185000.0 101000.00000000001 185800.0 101800.00000000001 ;
      RECT  189800.0 101000.00000000001 190600.00000000003 101800.00000000001 ;
      RECT  194600.0 101000.00000000001 195400.0 101800.00000000001 ;
      RECT  199399.99999999997 101000.00000000001 200200.0 101800.00000000001 ;
      RECT  204200.0 101000.00000000001 205000.0 101800.00000000001 ;
      RECT  209000.0 101000.00000000001 209800.0 101800.00000000001 ;
      RECT  7400.000000000003 105800.0 8200.000000000004 106600.0 ;
      RECT  12200.0 105800.0 13000.0 106600.0 ;
      RECT  16999.999999999996 105800.0 17799.999999999996 106600.0 ;
      RECT  21799.999999999993 105800.0 22599.999999999993 106600.0 ;
      RECT  26599.999999999996 105800.0 27400.0 106600.0 ;
      RECT  31399.999999999996 105800.0 32199.999999999996 106600.0 ;
      RECT  36200.0 105800.0 37000.0 106600.0 ;
      RECT  41000.0 105800.0 41800.0 106600.0 ;
      RECT  45800.0 105800.0 46599.99999999999 106600.0 ;
      RECT  50600.0 105800.0 51400.0 106600.0 ;
      RECT  55400.00000000001 105800.0 56200.0 106600.0 ;
      RECT  60200.0 105800.0 61000.0 106600.0 ;
      RECT  65000.0 105800.0 65800.0 106600.0 ;
      RECT  69800.0 105800.0 70600.0 106600.0 ;
      RECT  74600.00000000001 105800.0 75400.0 106600.0 ;
      RECT  79400.0 105800.0 80200.0 106600.0 ;
      RECT  84200.0 105800.0 85000.0 106600.0 ;
      RECT  89000.0 105800.0 89800.0 106600.0 ;
      RECT  93800.0 105800.0 94600.0 106600.0 ;
      RECT  98600.00000000001 105800.0 99400.0 106600.0 ;
      RECT  103400.0 105800.0 104200.0 106600.0 ;
      RECT  108200.0 105800.0 109000.0 106600.0 ;
      RECT  113000.00000000001 105800.0 113800.00000000001 106600.0 ;
      RECT  117800.0 105800.0 118600.0 106600.0 ;
      RECT  122600.00000000001 105800.0 123400.0 106600.0 ;
      RECT  127400.0 105800.0 128199.99999999999 106600.0 ;
      RECT  132200.0 105800.0 133000.0 106600.0 ;
      RECT  137000.0 105800.0 137800.0 106600.0 ;
      RECT  141800.0 105800.0 142600.00000000003 106600.0 ;
      RECT  146600.0 105800.0 147400.0 106600.0 ;
      RECT  151399.99999999997 105800.0 152200.0 106600.0 ;
      RECT  156200.0 105800.0 157000.0 106600.0 ;
      RECT  161000.0 105800.0 161800.0 106600.0 ;
      RECT  165800.0 105800.0 166600.00000000003 106600.0 ;
      RECT  170600.0 105800.0 171400.0 106600.0 ;
      RECT  175399.99999999997 105800.0 176200.0 106600.0 ;
      RECT  180200.0 105800.0 181000.0 106600.0 ;
      RECT  185000.0 105800.0 185800.0 106600.0 ;
      RECT  189800.0 105800.0 190600.00000000003 106600.0 ;
      RECT  194600.0 105800.0 195400.0 106600.0 ;
      RECT  199399.99999999997 105800.0 200200.0 106600.0 ;
      RECT  204200.0 105800.0 205000.0 106600.0 ;
      RECT  209000.0 105800.0 209800.0 106600.0 ;
      RECT  65000.0 110600.00000000001 65800.0 111400.0 ;
      RECT  69800.0 110600.00000000001 70600.0 111400.0 ;
      RECT  74600.00000000001 110600.00000000001 75400.0 111400.0 ;
      RECT  79400.0 110600.00000000001 80200.0 111400.0 ;
      RECT  84200.0 110600.00000000001 85000.0 111400.0 ;
      RECT  89000.0 110600.00000000001 89800.0 111400.0 ;
      RECT  93800.0 110600.00000000001 94600.0 111400.0 ;
      RECT  98600.00000000001 110600.00000000001 99400.0 111400.0 ;
      RECT  103400.0 110600.00000000001 104200.0 111400.0 ;
      RECT  108200.0 110600.00000000001 109000.0 111400.0 ;
      RECT  113000.00000000001 110600.00000000001 113800.00000000001 111400.0 ;
      RECT  117800.0 110600.00000000001 118600.0 111400.0 ;
      RECT  122600.00000000001 110600.00000000001 123400.0 111400.0 ;
      RECT  127400.0 110600.00000000001 128199.99999999999 111400.0 ;
      RECT  132200.0 110600.00000000001 133000.0 111400.0 ;
      RECT  137000.0 110600.00000000001 137800.0 111400.0 ;
      RECT  141800.0 110600.00000000001 142600.00000000003 111400.0 ;
      RECT  146600.0 110600.00000000001 147400.0 111400.0 ;
      RECT  151399.99999999997 110600.00000000001 152200.0 111400.0 ;
      RECT  156200.0 110600.00000000001 157000.0 111400.0 ;
      RECT  161000.0 110600.00000000001 161800.0 111400.0 ;
      RECT  165800.0 110600.00000000001 166600.00000000003 111400.0 ;
      RECT  170600.0 110600.00000000001 171400.0 111400.0 ;
      RECT  175399.99999999997 110600.00000000001 176200.0 111400.0 ;
      RECT  180200.0 110600.00000000001 181000.0 111400.0 ;
      RECT  185000.0 110600.00000000001 185800.0 111400.0 ;
      RECT  189800.0 110600.00000000001 190600.00000000003 111400.0 ;
      RECT  194600.0 110600.00000000001 195400.0 111400.0 ;
      RECT  199399.99999999997 110600.00000000001 200200.0 111400.0 ;
      RECT  204200.0 110600.00000000001 205000.0 111400.0 ;
      RECT  209000.0 110600.00000000001 209800.0 111400.0 ;
      RECT  7400.000000000003 115400.0 8200.000000000004 116200.0 ;
      RECT  12200.0 115400.0 13000.0 116200.0 ;
      RECT  16999.999999999996 115400.0 17799.999999999996 116200.0 ;
      RECT  21799.999999999993 115400.0 22599.999999999993 116200.0 ;
      RECT  26599.999999999996 115400.0 27400.0 116200.0 ;
      RECT  31399.999999999996 115400.0 32199.999999999996 116200.0 ;
      RECT  36200.0 115400.0 37000.0 116200.0 ;
      RECT  41000.0 115400.0 41800.0 116200.0 ;
      RECT  45800.0 115400.0 46599.99999999999 116200.0 ;
      RECT  50600.0 115400.0 51400.0 116200.0 ;
      RECT  55400.00000000001 115400.0 56200.0 116200.0 ;
      RECT  60200.0 115400.0 61000.0 116200.0 ;
      RECT  65000.0 115400.0 65800.0 116200.0 ;
      RECT  69800.0 115400.0 70600.0 116200.0 ;
      RECT  74600.00000000001 115400.0 75400.0 116200.0 ;
      RECT  79400.0 115400.0 80200.0 116200.0 ;
      RECT  84200.0 115400.0 85000.0 116200.0 ;
      RECT  89000.0 115400.0 89800.0 116200.0 ;
      RECT  93800.0 115400.0 94600.0 116200.0 ;
      RECT  98600.00000000001 115400.0 99400.0 116200.0 ;
      RECT  103400.0 115400.0 104200.0 116200.0 ;
      RECT  108200.0 115400.0 109000.0 116200.0 ;
      RECT  113000.00000000001 115400.0 113800.00000000001 116200.0 ;
      RECT  117800.0 115400.0 118600.0 116200.0 ;
      RECT  122600.00000000001 115400.0 123400.0 116200.0 ;
      RECT  127400.0 115400.0 128199.99999999999 116200.0 ;
      RECT  132200.0 115400.0 133000.0 116200.0 ;
      RECT  137000.0 115400.0 137800.0 116200.0 ;
      RECT  141800.0 115400.0 142600.00000000003 116200.0 ;
      RECT  146600.0 115400.0 147400.0 116200.0 ;
      RECT  151399.99999999997 115400.0 152200.0 116200.0 ;
      RECT  156200.0 115400.0 157000.0 116200.0 ;
      RECT  161000.0 115400.0 161800.0 116200.0 ;
      RECT  165800.0 115400.0 166600.00000000003 116200.0 ;
      RECT  170600.0 115400.0 171400.0 116200.0 ;
      RECT  175399.99999999997 115400.0 176200.0 116200.0 ;
      RECT  180200.0 115400.0 181000.0 116200.0 ;
      RECT  185000.0 115400.0 185800.0 116200.0 ;
      RECT  189800.0 115400.0 190600.00000000003 116200.0 ;
      RECT  194600.0 115400.0 195400.0 116200.0 ;
      RECT  199399.99999999997 115400.0 200200.0 116200.0 ;
      RECT  204200.0 115400.0 205000.0 116200.0 ;
      RECT  209000.0 115400.0 209800.0 116200.0 ;
      RECT  7400.000000000003 120200.0 8200.000000000004 121000.0 ;
      RECT  12200.0 120200.0 13000.0 121000.0 ;
      RECT  16999.999999999996 120200.0 17799.999999999996 121000.0 ;
      RECT  21799.999999999993 120200.0 22599.999999999993 121000.0 ;
      RECT  26599.999999999996 120200.0 27400.0 121000.0 ;
      RECT  31399.999999999996 120200.0 32199.999999999996 121000.0 ;
      RECT  36200.0 120200.0 37000.0 121000.0 ;
      RECT  41000.0 120200.0 41800.0 121000.0 ;
      RECT  45800.0 120200.0 46599.99999999999 121000.0 ;
      RECT  50600.0 120200.0 51400.0 121000.0 ;
      RECT  55400.00000000001 120200.0 56200.0 121000.0 ;
      RECT  60200.0 120200.0 61000.0 121000.0 ;
      RECT  65000.0 120200.0 65800.0 121000.0 ;
      RECT  69800.0 120200.0 70600.0 121000.0 ;
      RECT  74600.00000000001 120200.0 75400.0 121000.0 ;
      RECT  79400.0 120200.0 80200.0 121000.0 ;
      RECT  84200.0 120200.0 85000.0 121000.0 ;
      RECT  89000.0 120200.0 89800.0 121000.0 ;
      RECT  93800.0 120200.0 94600.0 121000.0 ;
      RECT  98600.00000000001 120200.0 99400.0 121000.0 ;
      RECT  103400.0 120200.0 104200.0 121000.0 ;
      RECT  108200.0 120200.0 109000.0 121000.0 ;
      RECT  113000.00000000001 120200.0 113800.00000000001 121000.0 ;
      RECT  117800.0 120200.0 118600.0 121000.0 ;
      RECT  122600.00000000001 120200.0 123400.0 121000.0 ;
      RECT  127400.0 120200.0 128199.99999999999 121000.0 ;
      RECT  132200.0 120200.0 133000.0 121000.0 ;
      RECT  137000.0 120200.0 137800.0 121000.0 ;
      RECT  141800.0 120200.0 142600.00000000003 121000.0 ;
      RECT  146600.0 120200.0 147400.0 121000.0 ;
      RECT  151399.99999999997 120200.0 152200.0 121000.0 ;
      RECT  156200.0 120200.0 157000.0 121000.0 ;
      RECT  161000.0 120200.0 161800.0 121000.0 ;
      RECT  165800.0 120200.0 166600.00000000003 121000.0 ;
      RECT  170600.0 120200.0 171400.0 121000.0 ;
      RECT  175399.99999999997 120200.0 176200.0 121000.0 ;
      RECT  180200.0 120200.0 181000.0 121000.0 ;
      RECT  185000.0 120200.0 185800.0 121000.0 ;
      RECT  189800.0 120200.0 190600.00000000003 121000.0 ;
      RECT  194600.0 120200.0 195400.0 121000.0 ;
      RECT  199399.99999999997 120200.0 200200.0 121000.0 ;
      RECT  204200.0 120200.0 205000.0 121000.0 ;
      RECT  209000.0 120200.0 209800.0 121000.0 ;
      RECT  7400.000000000003 125000.00000000001 8200.000000000004 125800.00000000001 ;
      RECT  12200.0 125000.00000000001 13000.0 125800.00000000001 ;
      RECT  16999.999999999996 125000.00000000001 17799.999999999996 125800.00000000001 ;
      RECT  21799.999999999993 125000.00000000001 22599.999999999993 125800.00000000001 ;
      RECT  26599.999999999996 125000.00000000001 27400.0 125800.00000000001 ;
      RECT  31399.999999999996 125000.00000000001 32199.999999999996 125800.00000000001 ;
      RECT  36200.0 125000.00000000001 37000.0 125800.00000000001 ;
      RECT  41000.0 125000.00000000001 41800.0 125800.00000000001 ;
      RECT  45800.0 125000.00000000001 46599.99999999999 125800.00000000001 ;
      RECT  50600.0 125000.00000000001 51400.0 125800.00000000001 ;
      RECT  55400.00000000001 125000.00000000001 56200.0 125800.00000000001 ;
      RECT  60200.0 125000.00000000001 61000.0 125800.00000000001 ;
      RECT  65000.0 125000.00000000001 65800.0 125800.00000000001 ;
      RECT  69800.0 125000.00000000001 70600.0 125800.00000000001 ;
      RECT  74600.00000000001 125000.00000000001 75400.0 125800.00000000001 ;
      RECT  79400.0 125000.00000000001 80200.0 125800.00000000001 ;
      RECT  84200.0 125000.00000000001 85000.0 125800.00000000001 ;
      RECT  89000.0 125000.00000000001 89800.0 125800.00000000001 ;
      RECT  93800.0 125000.00000000001 94600.0 125800.00000000001 ;
      RECT  98600.00000000001 125000.00000000001 99400.0 125800.00000000001 ;
      RECT  103400.0 125000.00000000001 104200.0 125800.00000000001 ;
      RECT  108200.0 125000.00000000001 109000.0 125800.00000000001 ;
      RECT  113000.00000000001 125000.00000000001 113800.00000000001 125800.00000000001 ;
      RECT  117800.0 125000.00000000001 118600.0 125800.00000000001 ;
      RECT  122600.00000000001 125000.00000000001 123400.0 125800.00000000001 ;
      RECT  127400.0 125000.00000000001 128199.99999999999 125800.00000000001 ;
      RECT  132200.0 125000.00000000001 133000.0 125800.00000000001 ;
      RECT  137000.0 125000.00000000001 137800.0 125800.00000000001 ;
      RECT  141800.0 125000.00000000001 142600.00000000003 125800.00000000001 ;
      RECT  146600.0 125000.00000000001 147400.0 125800.00000000001 ;
      RECT  151399.99999999997 125000.00000000001 152200.0 125800.00000000001 ;
      RECT  156200.0 125000.00000000001 157000.0 125800.00000000001 ;
      RECT  161000.0 125000.00000000001 161800.0 125800.00000000001 ;
      RECT  165800.0 125000.00000000001 166600.00000000003 125800.00000000001 ;
      RECT  170600.0 125000.00000000001 171400.0 125800.00000000001 ;
      RECT  175399.99999999997 125000.00000000001 176200.0 125800.00000000001 ;
      RECT  180200.0 125000.00000000001 181000.0 125800.00000000001 ;
      RECT  185000.0 125000.00000000001 185800.0 125800.00000000001 ;
      RECT  189800.0 125000.00000000001 190600.00000000003 125800.00000000001 ;
      RECT  194600.0 125000.00000000001 195400.0 125800.00000000001 ;
      RECT  199399.99999999997 125000.00000000001 200200.0 125800.00000000001 ;
      RECT  204200.0 125000.00000000001 205000.0 125800.00000000001 ;
      RECT  209000.0 125000.00000000001 209800.0 125800.00000000001 ;
      RECT  7400.000000000003 129800.00000000001 8200.000000000004 130600.00000000003 ;
      RECT  12200.0 129800.00000000001 13000.0 130600.00000000003 ;
      RECT  16999.999999999996 129800.00000000001 17799.999999999996 130600.00000000003 ;
      RECT  21799.999999999993 129800.00000000001 22599.999999999993 130600.00000000003 ;
      RECT  26599.999999999996 129800.00000000001 27400.0 130600.00000000003 ;
      RECT  31399.999999999996 129800.00000000001 32199.999999999996 130600.00000000003 ;
      RECT  36200.0 129800.00000000001 37000.0 130600.00000000003 ;
      RECT  41000.0 129800.00000000001 41800.0 130600.00000000003 ;
      RECT  45800.0 129800.00000000001 46599.99999999999 130600.00000000003 ;
      RECT  50600.0 129800.00000000001 51400.0 130600.00000000003 ;
      RECT  55400.00000000001 129800.00000000001 56200.0 130600.00000000003 ;
      RECT  60200.0 129800.00000000001 61000.0 130600.00000000003 ;
      RECT  65000.0 129800.00000000001 65800.0 130600.00000000003 ;
      RECT  7400.000000000003 134600.0 8200.000000000004 135400.0 ;
      RECT  12200.0 134600.0 13000.0 135400.0 ;
      RECT  16999.999999999996 134600.0 17799.999999999996 135400.0 ;
      RECT  21799.999999999993 134600.0 22599.999999999993 135400.0 ;
      RECT  26599.999999999996 134600.0 27400.0 135400.0 ;
      RECT  31399.999999999996 134600.0 32199.999999999996 135400.0 ;
      RECT  36200.0 134600.0 37000.0 135400.0 ;
      RECT  41000.0 134600.0 41800.0 135400.0 ;
      RECT  45800.0 134600.0 46599.99999999999 135400.0 ;
      RECT  50600.0 134600.0 51400.0 135400.0 ;
      RECT  55400.00000000001 134600.0 56200.0 135400.0 ;
      RECT  60200.0 134600.0 61000.0 135400.0 ;
      RECT  65000.0 134600.0 65800.0 135400.0 ;
      RECT  69800.0 134600.0 70600.0 135400.0 ;
      RECT  74600.00000000001 134600.0 75400.0 135400.0 ;
      RECT  79400.0 134600.0 80200.0 135400.0 ;
      RECT  84200.0 134600.0 85000.0 135400.0 ;
      RECT  89000.0 134600.0 89800.0 135400.0 ;
      RECT  93800.0 134600.0 94600.0 135400.0 ;
      RECT  98600.00000000001 134600.0 99400.0 135400.0 ;
      RECT  103400.0 134600.0 104200.0 135400.0 ;
      RECT  108200.0 134600.0 109000.0 135400.0 ;
      RECT  113000.00000000001 134600.0 113800.00000000001 135400.0 ;
      RECT  117800.0 134600.0 118600.0 135400.0 ;
      RECT  122600.00000000001 134600.0 123400.0 135400.0 ;
      RECT  127400.0 134600.0 128199.99999999999 135400.0 ;
      RECT  132200.0 134600.0 133000.0 135400.0 ;
      RECT  137000.0 134600.0 137800.0 135400.0 ;
      RECT  141800.0 134600.0 142600.00000000003 135400.0 ;
      RECT  146600.0 134600.0 147400.0 135400.0 ;
      RECT  151399.99999999997 134600.0 152200.0 135400.0 ;
      RECT  156200.0 134600.0 157000.0 135400.0 ;
      RECT  161000.0 134600.0 161800.0 135400.0 ;
      RECT  165800.0 134600.0 166600.00000000003 135400.0 ;
      RECT  170600.0 134600.0 171400.0 135400.0 ;
      RECT  175399.99999999997 134600.0 176200.0 135400.0 ;
      RECT  180200.0 134600.0 181000.0 135400.0 ;
      RECT  185000.0 134600.0 185800.0 135400.0 ;
      RECT  189800.0 134600.0 190600.00000000003 135400.0 ;
      RECT  194600.0 134600.0 195400.0 135400.0 ;
      RECT  199399.99999999997 134600.0 200200.0 135400.0 ;
      RECT  204200.0 134600.0 205000.0 135400.0 ;
      RECT  209000.0 134600.0 209800.0 135400.0 ;
      RECT  7400.000000000003 139399.99999999997 8200.000000000004 140200.0 ;
      RECT  12200.0 139399.99999999997 13000.0 140200.0 ;
      RECT  16999.999999999996 139399.99999999997 17799.999999999996 140200.0 ;
      RECT  21799.999999999993 139399.99999999997 22599.999999999993 140200.0 ;
      RECT  26599.999999999996 139399.99999999997 27400.0 140200.0 ;
      RECT  31399.999999999996 139399.99999999997 32199.999999999996 140200.0 ;
      RECT  36200.0 139399.99999999997 37000.0 140200.0 ;
      RECT  41000.0 139399.99999999997 41800.0 140200.0 ;
      RECT  45800.0 139399.99999999997 46599.99999999999 140200.0 ;
      RECT  50600.0 139399.99999999997 51400.0 140200.0 ;
      RECT  55400.00000000001 139399.99999999997 56200.0 140200.0 ;
      RECT  60200.0 139399.99999999997 61000.0 140200.0 ;
      RECT  79400.0 139399.99999999997 80200.0 140200.0 ;
      RECT  84200.0 139399.99999999997 85000.0 140200.0 ;
      RECT  89000.0 139399.99999999997 89800.0 140200.0 ;
      RECT  93800.0 139399.99999999997 94600.0 140200.0 ;
      RECT  98600.00000000001 139399.99999999997 99400.0 140200.0 ;
      RECT  103400.0 139399.99999999997 104200.0 140200.0 ;
      RECT  108200.0 139399.99999999997 109000.0 140200.0 ;
      RECT  113000.00000000001 139399.99999999997 113800.00000000001 140200.0 ;
      RECT  117800.0 139399.99999999997 118600.0 140200.0 ;
      RECT  122600.00000000001 139399.99999999997 123400.0 140200.0 ;
      RECT  127400.0 139399.99999999997 128199.99999999999 140200.0 ;
      RECT  132200.0 139399.99999999997 133000.0 140200.0 ;
      RECT  137000.0 139399.99999999997 137800.0 140200.0 ;
      RECT  141800.0 139399.99999999997 142600.00000000003 140200.0 ;
      RECT  146600.0 139399.99999999997 147400.0 140200.0 ;
      RECT  151399.99999999997 139399.99999999997 152200.0 140200.0 ;
      RECT  156200.0 139399.99999999997 157000.0 140200.0 ;
      RECT  161000.0 139399.99999999997 161800.0 140200.0 ;
      RECT  165800.0 139399.99999999997 166600.00000000003 140200.0 ;
      RECT  170600.0 139399.99999999997 171400.0 140200.0 ;
      RECT  175399.99999999997 139399.99999999997 176200.0 140200.0 ;
      RECT  180200.0 139399.99999999997 181000.0 140200.0 ;
      RECT  185000.0 139399.99999999997 185800.0 140200.0 ;
      RECT  189800.0 139399.99999999997 190600.00000000003 140200.0 ;
      RECT  194600.0 139399.99999999997 195400.0 140200.0 ;
      RECT  199399.99999999997 139399.99999999997 200200.0 140200.0 ;
      RECT  204200.0 139399.99999999997 205000.0 140200.0 ;
      RECT  209000.0 139399.99999999997 209800.0 140200.0 ;
      RECT  7400.000000000003 144200.0 8200.000000000004 145000.0 ;
      RECT  12200.0 144200.0 13000.0 145000.0 ;
      RECT  16999.999999999996 144200.0 17799.999999999996 145000.0 ;
      RECT  21799.999999999993 144200.0 22599.999999999993 145000.0 ;
      RECT  26599.999999999996 144200.0 27400.0 145000.0 ;
      RECT  31399.999999999996 144200.0 32199.999999999996 145000.0 ;
      RECT  36200.0 144200.0 37000.0 145000.0 ;
      RECT  41000.0 144200.0 41800.0 145000.0 ;
      RECT  45800.0 144200.0 46599.99999999999 145000.0 ;
      RECT  50600.0 144200.0 51400.0 145000.0 ;
      RECT  55400.00000000001 144200.0 56200.0 145000.0 ;
      RECT  60200.0 144200.0 61000.0 145000.0 ;
      RECT  65000.0 144200.0 65800.0 145000.0 ;
      RECT  69800.0 144200.0 70600.0 145000.0 ;
      RECT  74600.00000000001 144200.0 75400.0 145000.0 ;
      RECT  79400.0 144200.0 80200.0 145000.0 ;
      RECT  84200.0 144200.0 85000.0 145000.0 ;
      RECT  89000.0 144200.0 89800.0 145000.0 ;
      RECT  93800.0 144200.0 94600.0 145000.0 ;
      RECT  98600.00000000001 144200.0 99400.0 145000.0 ;
      RECT  103400.0 144200.0 104200.0 145000.0 ;
      RECT  108200.0 144200.0 109000.0 145000.0 ;
      RECT  113000.00000000001 144200.0 113800.00000000001 145000.0 ;
      RECT  117800.0 144200.0 118600.0 145000.0 ;
      RECT  122600.00000000001 144200.0 123400.0 145000.0 ;
      RECT  127400.0 144200.0 128199.99999999999 145000.0 ;
      RECT  132200.0 144200.0 133000.0 145000.0 ;
      RECT  137000.0 144200.0 137800.0 145000.0 ;
      RECT  141800.0 144200.0 142600.00000000003 145000.0 ;
      RECT  146600.0 144200.0 147400.0 145000.0 ;
      RECT  151399.99999999997 144200.0 152200.0 145000.0 ;
      RECT  156200.0 144200.0 157000.0 145000.0 ;
      RECT  161000.0 144200.0 161800.0 145000.0 ;
      RECT  165800.0 144200.0 166600.00000000003 145000.0 ;
      RECT  170600.0 144200.0 171400.0 145000.0 ;
      RECT  175399.99999999997 144200.0 176200.0 145000.0 ;
      RECT  180200.0 144200.0 181000.0 145000.0 ;
      RECT  185000.0 144200.0 185800.0 145000.0 ;
      RECT  189800.0 144200.0 190600.00000000003 145000.0 ;
      RECT  194600.0 144200.0 195400.0 145000.0 ;
      RECT  199399.99999999997 144200.0 200200.0 145000.0 ;
      RECT  204200.0 144200.0 205000.0 145000.0 ;
      RECT  209000.0 144200.0 209800.0 145000.0 ;
      RECT  7400.000000000003 149000.0 8200.000000000004 149800.0 ;
      RECT  12200.0 149000.0 13000.0 149800.0 ;
      RECT  16999.999999999996 149000.0 17799.999999999996 149800.0 ;
      RECT  21799.999999999993 149000.0 22599.999999999993 149800.0 ;
      RECT  26599.999999999996 149000.0 27400.0 149800.0 ;
      RECT  31399.999999999996 149000.0 32199.999999999996 149800.0 ;
      RECT  36200.0 149000.0 37000.0 149800.0 ;
      RECT  41000.0 149000.0 41800.0 149800.0 ;
      RECT  45800.0 149000.0 46599.99999999999 149800.0 ;
      RECT  50600.0 149000.0 51400.0 149800.0 ;
      RECT  55400.00000000001 149000.0 56200.0 149800.0 ;
      RECT  60200.0 149000.0 61000.0 149800.0 ;
      RECT  65000.0 149000.0 65800.0 149800.0 ;
      RECT  69800.0 149000.0 70600.0 149800.0 ;
      RECT  74600.00000000001 149000.0 75400.0 149800.0 ;
      RECT  79400.0 149000.0 80200.0 149800.0 ;
      RECT  84200.0 149000.0 85000.0 149800.0 ;
      RECT  89000.0 149000.0 89800.0 149800.0 ;
      RECT  93800.0 149000.0 94600.0 149800.0 ;
      RECT  98600.00000000001 149000.0 99400.0 149800.0 ;
      RECT  103400.0 149000.0 104200.0 149800.0 ;
      RECT  108200.0 149000.0 109000.0 149800.0 ;
      RECT  113000.00000000001 149000.0 113800.00000000001 149800.0 ;
      RECT  117800.0 149000.0 118600.0 149800.0 ;
      RECT  122600.00000000001 149000.0 123400.0 149800.0 ;
      RECT  127400.0 149000.0 128199.99999999999 149800.0 ;
      RECT  132200.0 149000.0 133000.0 149800.0 ;
      RECT  137000.0 149000.0 137800.0 149800.0 ;
      RECT  141800.0 149000.0 142600.00000000003 149800.0 ;
      RECT  146600.0 149000.0 147400.0 149800.0 ;
      RECT  151399.99999999997 149000.0 152200.0 149800.0 ;
      RECT  156200.0 149000.0 157000.0 149800.0 ;
      RECT  161000.0 149000.0 161800.0 149800.0 ;
      RECT  165800.0 149000.0 166600.00000000003 149800.0 ;
      RECT  170600.0 149000.0 171400.0 149800.0 ;
      RECT  175399.99999999997 149000.0 176200.0 149800.0 ;
      RECT  180200.0 149000.0 181000.0 149800.0 ;
      RECT  185000.0 149000.0 185800.0 149800.0 ;
      RECT  189800.0 149000.0 190600.00000000003 149800.0 ;
      RECT  194600.0 149000.0 195400.0 149800.0 ;
      RECT  199399.99999999997 149000.0 200200.0 149800.0 ;
      RECT  204200.0 149000.0 205000.0 149800.0 ;
      RECT  209000.0 149000.0 209800.0 149800.0 ;
      RECT  7400.000000000003 153800.0 8200.000000000004 154600.00000000003 ;
      RECT  12200.0 153800.0 13000.0 154600.00000000003 ;
      RECT  16999.999999999996 153800.0 17799.999999999996 154600.00000000003 ;
      RECT  21799.999999999993 153800.0 22599.999999999993 154600.00000000003 ;
      RECT  26599.999999999996 153800.0 27400.0 154600.00000000003 ;
      RECT  31399.999999999996 153800.0 32199.999999999996 154600.00000000003 ;
      RECT  36200.0 153800.0 37000.0 154600.00000000003 ;
      RECT  41000.0 153800.0 41800.0 154600.00000000003 ;
      RECT  45800.0 153800.0 46599.99999999999 154600.00000000003 ;
      RECT  50600.0 153800.0 51400.0 154600.00000000003 ;
      RECT  55400.00000000001 153800.0 56200.0 154600.00000000003 ;
      RECT  60200.0 153800.0 61000.0 154600.00000000003 ;
      RECT  65000.0 153800.0 65800.0 154600.00000000003 ;
      RECT  69800.0 153800.0 70600.0 154600.00000000003 ;
      RECT  74600.00000000001 153800.0 75400.0 154600.00000000003 ;
      RECT  79400.0 153800.0 80200.0 154600.00000000003 ;
      RECT  84200.0 153800.0 85000.0 154600.00000000003 ;
      RECT  89000.0 153800.0 89800.0 154600.00000000003 ;
      RECT  93800.0 153800.0 94600.0 154600.00000000003 ;
      RECT  98600.00000000001 153800.0 99400.0 154600.00000000003 ;
      RECT  103400.0 153800.0 104200.0 154600.00000000003 ;
      RECT  108200.0 153800.0 109000.0 154600.00000000003 ;
      RECT  113000.00000000001 153800.0 113800.00000000001 154600.00000000003 ;
      RECT  117800.0 153800.0 118600.0 154600.00000000003 ;
      RECT  122600.00000000001 153800.0 123400.0 154600.00000000003 ;
      RECT  127400.0 153800.0 128199.99999999999 154600.00000000003 ;
      RECT  132200.0 153800.0 133000.0 154600.00000000003 ;
      RECT  137000.0 153800.0 137800.0 154600.00000000003 ;
      RECT  141800.0 153800.0 142600.00000000003 154600.00000000003 ;
      RECT  146600.0 153800.0 147400.0 154600.00000000003 ;
      RECT  151399.99999999997 153800.0 152200.0 154600.00000000003 ;
      RECT  156200.0 153800.0 157000.0 154600.00000000003 ;
      RECT  161000.0 153800.0 161800.0 154600.00000000003 ;
      RECT  165800.0 153800.0 166600.00000000003 154600.00000000003 ;
      RECT  170600.0 153800.0 171400.0 154600.00000000003 ;
      RECT  175399.99999999997 153800.0 176200.0 154600.00000000003 ;
      RECT  180200.0 153800.0 181000.0 154600.00000000003 ;
      RECT  185000.0 153800.0 185800.0 154600.00000000003 ;
      RECT  189800.0 153800.0 190600.00000000003 154600.00000000003 ;
      RECT  194600.0 153800.0 195400.0 154600.00000000003 ;
      RECT  199399.99999999997 153800.0 200200.0 154600.00000000003 ;
      RECT  204200.0 153800.0 205000.0 154600.00000000003 ;
      RECT  209000.0 153800.0 209800.0 154600.00000000003 ;
      RECT  7400.000000000003 158600.0 8200.000000000004 159400.0 ;
      RECT  12200.0 158600.0 13000.0 159400.0 ;
      RECT  16999.999999999996 158600.0 17799.999999999996 159400.0 ;
      RECT  21799.999999999993 158600.0 22599.999999999993 159400.0 ;
      RECT  26599.999999999996 158600.0 27400.0 159400.0 ;
      RECT  31399.999999999996 158600.0 32199.999999999996 159400.0 ;
      RECT  36200.0 158600.0 37000.0 159400.0 ;
      RECT  41000.0 158600.0 41800.0 159400.0 ;
      RECT  45800.0 158600.0 46599.99999999999 159400.0 ;
      RECT  50600.0 158600.0 51400.0 159400.0 ;
      RECT  55400.00000000001 158600.0 56200.0 159400.0 ;
      RECT  60200.0 158600.0 61000.0 159400.0 ;
      RECT  65000.0 158600.0 65800.0 159400.0 ;
      RECT  69800.0 158600.0 70600.0 159400.0 ;
      RECT  74600.00000000001 158600.0 75400.0 159400.0 ;
      RECT  79400.0 158600.0 80200.0 159400.0 ;
      RECT  84200.0 158600.0 85000.0 159400.0 ;
      RECT  89000.0 158600.0 89800.0 159400.0 ;
      RECT  93800.0 158600.0 94600.0 159400.0 ;
      RECT  98600.00000000001 158600.0 99400.0 159400.0 ;
      RECT  103400.0 158600.0 104200.0 159400.0 ;
      RECT  108200.0 158600.0 109000.0 159400.0 ;
      RECT  113000.00000000001 158600.0 113800.00000000001 159400.0 ;
      RECT  117800.0 158600.0 118600.0 159400.0 ;
      RECT  122600.00000000001 158600.0 123400.0 159400.0 ;
      RECT  127400.0 158600.0 128199.99999999999 159400.0 ;
      RECT  132200.0 158600.0 133000.0 159400.0 ;
      RECT  137000.0 158600.0 137800.0 159400.0 ;
      RECT  141800.0 158600.0 142600.00000000003 159400.0 ;
      RECT  146600.0 158600.0 147400.0 159400.0 ;
      RECT  151399.99999999997 158600.0 152200.0 159400.0 ;
      RECT  156200.0 158600.0 157000.0 159400.0 ;
      RECT  161000.0 158600.0 161800.0 159400.0 ;
      RECT  165800.0 158600.0 166600.00000000003 159400.0 ;
      RECT  7400.000000000003 163399.99999999997 8200.000000000004 164200.0 ;
      RECT  12200.0 163399.99999999997 13000.0 164200.0 ;
      RECT  16999.999999999996 163399.99999999997 17799.999999999996 164200.0 ;
      RECT  21799.999999999993 163399.99999999997 22599.999999999993 164200.0 ;
      RECT  26599.999999999996 163399.99999999997 27400.0 164200.0 ;
      RECT  31399.999999999996 163399.99999999997 32199.999999999996 164200.0 ;
      RECT  36200.0 163399.99999999997 37000.0 164200.0 ;
      RECT  41000.0 163399.99999999997 41800.0 164200.0 ;
      RECT  45800.0 163399.99999999997 46599.99999999999 164200.0 ;
      RECT  50600.0 163399.99999999997 51400.0 164200.0 ;
      RECT  55400.00000000001 163399.99999999997 56200.0 164200.0 ;
      RECT  60200.0 163399.99999999997 61000.0 164200.0 ;
      RECT  65000.0 163399.99999999997 65800.0 164200.0 ;
      RECT  69800.0 163399.99999999997 70600.0 164200.0 ;
      RECT  74600.00000000001 163399.99999999997 75400.0 164200.0 ;
      RECT  79400.0 163399.99999999997 80200.0 164200.0 ;
      RECT  84200.0 163399.99999999997 85000.0 164200.0 ;
      RECT  89000.0 163399.99999999997 89800.0 164200.0 ;
      RECT  93800.0 163399.99999999997 94600.0 164200.0 ;
      RECT  98600.00000000001 163399.99999999997 99400.0 164200.0 ;
      RECT  103400.0 163399.99999999997 104200.0 164200.0 ;
      RECT  108200.0 163399.99999999997 109000.0 164200.0 ;
      RECT  113000.00000000001 163399.99999999997 113800.00000000001 164200.0 ;
      RECT  117800.0 163399.99999999997 118600.0 164200.0 ;
      RECT  122600.00000000001 163399.99999999997 123400.0 164200.0 ;
      RECT  127400.0 163399.99999999997 128199.99999999999 164200.0 ;
      RECT  132200.0 163399.99999999997 133000.0 164200.0 ;
      RECT  137000.0 163399.99999999997 137800.0 164200.0 ;
      RECT  141800.0 163399.99999999997 142600.00000000003 164200.0 ;
      RECT  146600.0 163399.99999999997 147400.0 164200.0 ;
      RECT  151399.99999999997 163399.99999999997 152200.0 164200.0 ;
      RECT  156200.0 163399.99999999997 157000.0 164200.0 ;
      RECT  161000.0 163399.99999999997 161800.0 164200.0 ;
      RECT  165800.0 163399.99999999997 166600.00000000003 164200.0 ;
      RECT  170600.0 163399.99999999997 171400.0 164200.0 ;
      RECT  175399.99999999997 163399.99999999997 176200.0 164200.0 ;
      RECT  180200.0 163399.99999999997 181000.0 164200.0 ;
      RECT  185000.0 163399.99999999997 185800.0 164200.0 ;
      RECT  189800.0 163399.99999999997 190600.00000000003 164200.0 ;
      RECT  194600.0 163399.99999999997 195400.0 164200.0 ;
      RECT  199399.99999999997 163399.99999999997 200200.0 164200.0 ;
      RECT  204200.0 163399.99999999997 205000.0 164200.0 ;
      RECT  209000.0 163399.99999999997 209800.0 164200.0 ;
      RECT  7400.000000000003 168200.0 8200.000000000004 169000.0 ;
      RECT  12200.0 168200.0 13000.0 169000.0 ;
      RECT  16999.999999999996 168200.0 17799.999999999996 169000.0 ;
      RECT  21799.999999999993 168200.0 22599.999999999993 169000.0 ;
      RECT  26599.999999999996 168200.0 27400.0 169000.0 ;
      RECT  31399.999999999996 168200.0 32199.999999999996 169000.0 ;
      RECT  36200.0 168200.0 37000.0 169000.0 ;
      RECT  41000.0 168200.0 41800.0 169000.0 ;
      RECT  45800.0 168200.0 46599.99999999999 169000.0 ;
      RECT  50600.0 168200.0 51400.0 169000.0 ;
      RECT  55400.00000000001 168200.0 56200.0 169000.0 ;
      RECT  60200.0 168200.0 61000.0 169000.0 ;
      RECT  65000.0 168200.0 65800.0 169000.0 ;
      RECT  69800.0 168200.0 70600.0 169000.0 ;
      RECT  74600.00000000001 168200.0 75400.0 169000.0 ;
      RECT  79400.0 168200.0 80200.0 169000.0 ;
      RECT  84200.0 168200.0 85000.0 169000.0 ;
      RECT  89000.0 168200.0 89800.0 169000.0 ;
      RECT  93800.0 168200.0 94600.0 169000.0 ;
      RECT  98600.00000000001 168200.0 99400.0 169000.0 ;
      RECT  103400.0 168200.0 104200.0 169000.0 ;
      RECT  108200.0 168200.0 109000.0 169000.0 ;
      RECT  113000.00000000001 168200.0 113800.00000000001 169000.0 ;
      RECT  117800.0 168200.0 118600.0 169000.0 ;
      RECT  122600.00000000001 168200.0 123400.0 169000.0 ;
      RECT  127400.0 168200.0 128199.99999999999 169000.0 ;
      RECT  132200.0 168200.0 133000.0 169000.0 ;
      RECT  137000.0 168200.0 137800.0 169000.0 ;
      RECT  141800.0 168200.0 142600.00000000003 169000.0 ;
      RECT  146600.0 168200.0 147400.0 169000.0 ;
      RECT  151399.99999999997 168200.0 152200.0 169000.0 ;
      RECT  156200.0 168200.0 157000.0 169000.0 ;
      RECT  161000.0 168200.0 161800.0 169000.0 ;
      RECT  165800.0 168200.0 166600.00000000003 169000.0 ;
      RECT  170600.0 168200.0 171400.0 169000.0 ;
      RECT  175399.99999999997 168200.0 176200.0 169000.0 ;
      RECT  180200.0 168200.0 181000.0 169000.0 ;
      RECT  185000.0 168200.0 185800.0 169000.0 ;
      RECT  189800.0 168200.0 190600.00000000003 169000.0 ;
      RECT  194600.0 168200.0 195400.0 169000.0 ;
      RECT  199399.99999999997 168200.0 200200.0 169000.0 ;
      RECT  204200.0 168200.0 205000.0 169000.0 ;
      RECT  209000.0 168200.0 209800.0 169000.0 ;
      RECT  26599.999999999996 173000.0 27400.0 173800.0 ;
      RECT  31399.999999999996 173000.0 32199.999999999996 173800.0 ;
      RECT  36200.0 173000.0 37000.0 173800.0 ;
      RECT  41000.0 173000.0 41800.0 173800.0 ;
      RECT  45800.0 173000.0 46599.99999999999 173800.0 ;
      RECT  50600.0 173000.0 51400.0 173800.0 ;
      RECT  55400.00000000001 173000.0 56200.0 173800.0 ;
      RECT  60200.0 173000.0 61000.0 173800.0 ;
      RECT  65000.0 173000.0 65800.0 173800.0 ;
      RECT  69800.0 173000.0 70600.0 173800.0 ;
      RECT  74600.00000000001 173000.0 75400.0 173800.0 ;
      RECT  79400.0 173000.0 80200.0 173800.0 ;
      RECT  84200.0 173000.0 85000.0 173800.0 ;
      RECT  89000.0 173000.0 89800.0 173800.0 ;
      RECT  93800.0 173000.0 94600.0 173800.0 ;
      RECT  98600.00000000001 173000.0 99400.0 173800.0 ;
      RECT  103400.0 173000.0 104200.0 173800.0 ;
      RECT  108200.0 173000.0 109000.0 173800.0 ;
      RECT  113000.00000000001 173000.0 113800.00000000001 173800.0 ;
      RECT  117800.0 173000.0 118600.0 173800.0 ;
      RECT  122600.00000000001 173000.0 123400.0 173800.0 ;
      RECT  127400.0 173000.0 128199.99999999999 173800.0 ;
      RECT  132200.0 173000.0 133000.0 173800.0 ;
      RECT  137000.0 173000.0 137800.0 173800.0 ;
      RECT  141800.0 173000.0 142600.00000000003 173800.0 ;
      RECT  146600.0 173000.0 147400.0 173800.0 ;
      RECT  151399.99999999997 173000.0 152200.0 173800.0 ;
      RECT  156200.0 173000.0 157000.0 173800.0 ;
      RECT  161000.0 173000.0 161800.0 173800.0 ;
      RECT  165800.0 173000.0 166600.00000000003 173800.0 ;
      RECT  170600.0 173000.0 171400.0 173800.0 ;
      RECT  175399.99999999997 173000.0 176200.0 173800.0 ;
      RECT  180200.0 173000.0 181000.0 173800.0 ;
      RECT  185000.0 173000.0 185800.0 173800.0 ;
      RECT  189800.0 173000.0 190600.00000000003 173800.0 ;
      RECT  194600.0 173000.0 195400.0 173800.0 ;
      RECT  199399.99999999997 173000.0 200200.0 173800.0 ;
      RECT  204200.0 173000.0 205000.0 173800.0 ;
      RECT  209000.0 173000.0 209800.0 173800.0 ;
      RECT  31399.999999999996 177800.0 32199.999999999996 178600.00000000003 ;
      RECT  36200.0 177800.0 37000.0 178600.00000000003 ;
      RECT  41000.0 177800.0 41800.0 178600.00000000003 ;
      RECT  45800.0 177800.0 46599.99999999999 178600.00000000003 ;
      RECT  50600.0 177800.0 51400.0 178600.00000000003 ;
      RECT  55400.00000000001 177800.0 56200.0 178600.00000000003 ;
      RECT  60200.0 177800.0 61000.0 178600.00000000003 ;
      RECT  65000.0 177800.0 65800.0 178600.00000000003 ;
      RECT  41000.0 182600.0 41800.0 183400.0 ;
      RECT  45800.0 182600.0 46599.99999999999 183400.0 ;
      RECT  50600.0 182600.0 51400.0 183400.0 ;
      RECT  55400.00000000001 182600.0 56200.0 183400.0 ;
      RECT  60200.0 182600.0 61000.0 183400.0 ;
      RECT  65000.0 182600.0 65800.0 183400.0 ;
      RECT  69800.0 182600.0 70600.0 183400.0 ;
      RECT  74600.00000000001 182600.0 75400.0 183400.0 ;
      RECT  79400.0 182600.0 80200.0 183400.0 ;
      RECT  84200.0 182600.0 85000.0 183400.0 ;
      RECT  89000.0 182600.0 89800.0 183400.0 ;
      RECT  93800.0 182600.0 94600.0 183400.0 ;
      RECT  98600.00000000001 182600.0 99400.0 183400.0 ;
      RECT  103400.0 182600.0 104200.0 183400.0 ;
      RECT  108200.0 182600.0 109000.0 183400.0 ;
      RECT  113000.00000000001 182600.0 113800.00000000001 183400.0 ;
      RECT  117800.0 182600.0 118600.0 183400.0 ;
      RECT  122600.00000000001 182600.0 123400.0 183400.0 ;
      RECT  127400.0 182600.0 128199.99999999999 183400.0 ;
      RECT  132200.0 182600.0 133000.0 183400.0 ;
      RECT  137000.0 182600.0 137800.0 183400.0 ;
      RECT  141800.0 182600.0 142600.00000000003 183400.0 ;
      RECT  146600.0 182600.0 147400.0 183400.0 ;
      RECT  151399.99999999997 182600.0 152200.0 183400.0 ;
      RECT  156200.0 182600.0 157000.0 183400.0 ;
      RECT  161000.0 182600.0 161800.0 183400.0 ;
      RECT  165800.0 182600.0 166600.00000000003 183400.0 ;
      RECT  170600.0 182600.0 171400.0 183400.0 ;
      RECT  175399.99999999997 182600.0 176200.0 183400.0 ;
      RECT  180200.0 182600.0 181000.0 183400.0 ;
      RECT  185000.0 182600.0 185800.0 183400.0 ;
      RECT  189800.0 182600.0 190600.00000000003 183400.0 ;
      RECT  194600.0 182600.0 195400.0 183400.0 ;
      RECT  199399.99999999997 182600.0 200200.0 183400.0 ;
      RECT  204200.0 182600.0 205000.0 183400.0 ;
      RECT  209000.0 182600.0 209800.0 183400.0 ;
      RECT  31399.999999999996 187399.99999999997 32199.999999999996 188200.0 ;
      RECT  36200.0 187399.99999999997 37000.0 188200.0 ;
      RECT  41000.0 187399.99999999997 41800.0 188200.0 ;
      RECT  45800.0 187399.99999999997 46599.99999999999 188200.0 ;
      RECT  50600.0 187399.99999999997 51400.0 188200.0 ;
      RECT  55400.00000000001 187399.99999999997 56200.0 188200.0 ;
      RECT  60200.0 187399.99999999997 61000.0 188200.0 ;
      RECT  65000.0 187399.99999999997 65800.0 188200.0 ;
      RECT  127400.0 187399.99999999997 128199.99999999999 188200.0 ;
      RECT  132200.0 187399.99999999997 133000.0 188200.0 ;
      RECT  137000.0 187399.99999999997 137800.0 188200.0 ;
      RECT  141800.0 187399.99999999997 142600.00000000003 188200.0 ;
      RECT  146600.0 187399.99999999997 147400.0 188200.0 ;
      RECT  151399.99999999997 187399.99999999997 152200.0 188200.0 ;
      RECT  156200.0 187399.99999999997 157000.0 188200.0 ;
      RECT  161000.0 187399.99999999997 161800.0 188200.0 ;
      RECT  165800.0 187399.99999999997 166600.00000000003 188200.0 ;
      RECT  170600.0 187399.99999999997 171400.0 188200.0 ;
      RECT  175399.99999999997 187399.99999999997 176200.0 188200.0 ;
      RECT  180200.0 187399.99999999997 181000.0 188200.0 ;
      RECT  185000.0 187399.99999999997 185800.0 188200.0 ;
      RECT  189800.0 187399.99999999997 190600.00000000003 188200.0 ;
      RECT  194600.0 187399.99999999997 195400.0 188200.0 ;
      RECT  199399.99999999997 187399.99999999997 200200.0 188200.0 ;
      RECT  204200.0 187399.99999999997 205000.0 188200.0 ;
      RECT  209000.0 187399.99999999997 209800.0 188200.0 ;
      RECT  7400.000000000003 192200.0 8200.000000000004 193000.0 ;
      RECT  12200.0 192200.0 13000.0 193000.0 ;
      RECT  16999.999999999996 192200.0 17799.999999999996 193000.0 ;
      RECT  21799.999999999993 192200.0 22599.999999999993 193000.0 ;
      RECT  26599.999999999996 192200.0 27400.0 193000.0 ;
      RECT  31399.999999999996 192200.0 32199.999999999996 193000.0 ;
      RECT  36200.0 192200.0 37000.0 193000.0 ;
      RECT  41000.0 192200.0 41800.0 193000.0 ;
      RECT  45800.0 192200.0 46599.99999999999 193000.0 ;
      RECT  50600.0 192200.0 51400.0 193000.0 ;
      RECT  55400.00000000001 192200.0 56200.0 193000.0 ;
      RECT  60200.0 192200.0 61000.0 193000.0 ;
      RECT  65000.0 192200.0 65800.0 193000.0 ;
      RECT  69800.0 192200.0 70600.0 193000.0 ;
      RECT  74600.00000000001 192200.0 75400.0 193000.0 ;
      RECT  79400.0 192200.0 80200.0 193000.0 ;
      RECT  84200.0 192200.0 85000.0 193000.0 ;
      RECT  89000.0 192200.0 89800.0 193000.0 ;
      RECT  93800.0 192200.0 94600.0 193000.0 ;
      RECT  98600.00000000001 192200.0 99400.0 193000.0 ;
      RECT  103400.0 192200.0 104200.0 193000.0 ;
      RECT  108200.0 192200.0 109000.0 193000.0 ;
      RECT  113000.00000000001 192200.0 113800.00000000001 193000.0 ;
      RECT  117800.0 192200.0 118600.0 193000.0 ;
      RECT  122600.00000000001 192200.0 123400.0 193000.0 ;
      RECT  127400.0 192200.0 128199.99999999999 193000.0 ;
      RECT  132200.0 192200.0 133000.0 193000.0 ;
      RECT  137000.0 192200.0 137800.0 193000.0 ;
      RECT  141800.0 192200.0 142600.00000000003 193000.0 ;
      RECT  146600.0 192200.0 147400.0 193000.0 ;
      RECT  151399.99999999997 192200.0 152200.0 193000.0 ;
      RECT  156200.0 192200.0 157000.0 193000.0 ;
      RECT  161000.0 192200.0 161800.0 193000.0 ;
      RECT  165800.0 192200.0 166600.00000000003 193000.0 ;
      RECT  170600.0 192200.0 171400.0 193000.0 ;
      RECT  175399.99999999997 192200.0 176200.0 193000.0 ;
      RECT  180200.0 192200.0 181000.0 193000.0 ;
      RECT  185000.0 192200.0 185800.0 193000.0 ;
      RECT  189800.0 192200.0 190600.00000000003 193000.0 ;
      RECT  194600.0 192200.0 195400.0 193000.0 ;
      RECT  199399.99999999997 192200.0 200200.0 193000.0 ;
      RECT  204200.0 192200.0 205000.0 193000.0 ;
      RECT  209000.0 192200.0 209800.0 193000.0 ;
      RECT  31399.999999999996 197000.0 32199.999999999996 197800.0 ;
      RECT  36200.0 197000.0 37000.0 197800.0 ;
      RECT  41000.0 197000.0 41800.0 197800.0 ;
      RECT  45800.0 197000.0 46599.99999999999 197800.0 ;
      RECT  50600.0 197000.0 51400.0 197800.0 ;
      RECT  55400.00000000001 197000.0 56200.0 197800.0 ;
      RECT  60200.0 197000.0 61000.0 197800.0 ;
      RECT  65000.0 197000.0 65800.0 197800.0 ;
      RECT  69800.0 197000.0 70600.0 197800.0 ;
      RECT  74600.00000000001 197000.0 75400.0 197800.0 ;
      RECT  79400.0 197000.0 80200.0 197800.0 ;
      RECT  41000.0 201800.0 41800.0 202600.00000000003 ;
      RECT  45800.0 201800.0 46599.99999999999 202600.00000000003 ;
      RECT  50600.0 201800.0 51400.0 202600.00000000003 ;
      RECT  55400.00000000001 201800.0 56200.0 202600.00000000003 ;
      RECT  60200.0 201800.0 61000.0 202600.00000000003 ;
      RECT  65000.0 201800.0 65800.0 202600.00000000003 ;
      RECT  69800.0 201800.0 70600.0 202600.00000000003 ;
      RECT  74600.00000000001 201800.0 75400.0 202600.00000000003 ;
      RECT  79400.0 201800.0 80200.0 202600.00000000003 ;
      RECT  84200.0 201800.0 85000.0 202600.00000000003 ;
      RECT  89000.0 201800.0 89800.0 202600.00000000003 ;
      RECT  93800.0 201800.0 94600.0 202600.00000000003 ;
      RECT  98600.00000000001 201800.0 99400.0 202600.00000000003 ;
      RECT  103400.0 201800.0 104200.0 202600.00000000003 ;
      RECT  108200.0 201800.0 109000.0 202600.00000000003 ;
      RECT  113000.00000000001 201800.0 113800.00000000001 202600.00000000003 ;
      RECT  117800.0 201800.0 118600.0 202600.00000000003 ;
      RECT  122600.00000000001 201800.0 123400.0 202600.00000000003 ;
      RECT  127400.0 201800.0 128199.99999999999 202600.00000000003 ;
      RECT  132200.0 201800.0 133000.0 202600.00000000003 ;
      RECT  137000.0 201800.0 137800.0 202600.00000000003 ;
      RECT  141800.0 201800.0 142600.00000000003 202600.00000000003 ;
      RECT  146600.0 201800.0 147400.0 202600.00000000003 ;
      RECT  151399.99999999997 201800.0 152200.0 202600.00000000003 ;
      RECT  156200.0 201800.0 157000.0 202600.00000000003 ;
      RECT  161000.0 201800.0 161800.0 202600.00000000003 ;
      RECT  165800.0 201800.0 166600.00000000003 202600.00000000003 ;
      RECT  170600.0 201800.0 171400.0 202600.00000000003 ;
      RECT  175399.99999999997 201800.0 176200.0 202600.00000000003 ;
      RECT  180200.0 201800.0 181000.0 202600.00000000003 ;
      RECT  185000.0 201800.0 185800.0 202600.00000000003 ;
      RECT  189800.0 201800.0 190600.00000000003 202600.00000000003 ;
      RECT  194600.0 201800.0 195400.0 202600.00000000003 ;
      RECT  199399.99999999997 201800.0 200200.0 202600.00000000003 ;
      RECT  204200.0 201800.0 205000.0 202600.00000000003 ;
      RECT  209000.0 201800.0 209800.0 202600.00000000003 ;
      RECT  31399.999999999996 206600.00000000003 32199.999999999996 207400.00000000003 ;
      RECT  36200.0 206600.00000000003 37000.0 207400.00000000003 ;
      RECT  41000.0 206600.00000000003 41800.0 207400.00000000003 ;
      RECT  45800.0 206600.00000000003 46599.99999999999 207400.00000000003 ;
      RECT  50600.0 206600.00000000003 51400.0 207400.00000000003 ;
      RECT  55400.00000000001 206600.00000000003 56200.0 207400.00000000003 ;
      RECT  60200.0 206600.00000000003 61000.0 207400.00000000003 ;
      RECT  65000.0 206600.00000000003 65800.0 207400.00000000003 ;
      RECT  69800.0 206600.00000000003 70600.0 207400.00000000003 ;
      RECT  74600.00000000001 206600.00000000003 75400.0 207400.00000000003 ;
      RECT  79400.0 206600.00000000003 80200.0 207400.00000000003 ;
      RECT  84200.0 206600.00000000003 85000.0 207400.00000000003 ;
      RECT  89000.0 206600.00000000003 89800.0 207400.00000000003 ;
      RECT  93800.0 206600.00000000003 94600.0 207400.00000000003 ;
      RECT  98600.00000000001 206600.00000000003 99400.0 207400.00000000003 ;
      RECT  103400.0 206600.00000000003 104200.0 207400.00000000003 ;
      RECT  127400.0 206600.00000000003 128199.99999999999 207400.00000000003 ;
      RECT  132200.0 206600.00000000003 133000.0 207400.00000000003 ;
      RECT  137000.0 206600.00000000003 137800.0 207400.00000000003 ;
      RECT  141800.0 206600.00000000003 142600.00000000003 207400.00000000003 ;
      RECT  146600.0 206600.00000000003 147400.0 207400.00000000003 ;
      RECT  151399.99999999997 206600.00000000003 152200.0 207400.00000000003 ;
      RECT  156200.0 206600.00000000003 157000.0 207400.00000000003 ;
      RECT  161000.0 206600.00000000003 161800.0 207400.00000000003 ;
      RECT  165800.0 206600.00000000003 166600.00000000003 207400.00000000003 ;
      RECT  170600.0 206600.00000000003 171400.0 207400.00000000003 ;
      RECT  175399.99999999997 206600.00000000003 176200.0 207400.00000000003 ;
      RECT  180200.0 206600.00000000003 181000.0 207400.00000000003 ;
      RECT  185000.0 206600.00000000003 185800.0 207400.00000000003 ;
      RECT  189800.0 206600.00000000003 190600.00000000003 207400.00000000003 ;
      RECT  194600.0 206600.00000000003 195400.0 207400.00000000003 ;
      RECT  199399.99999999997 206600.00000000003 200200.0 207400.00000000003 ;
      RECT  204200.0 206600.00000000003 205000.0 207400.00000000003 ;
      RECT  209000.0 206600.00000000003 209800.0 207400.00000000003 ;
      RECT  7400.000000000003 211399.99999999997 8200.000000000004 212200.0 ;
      RECT  12200.0 211399.99999999997 13000.0 212200.0 ;
      RECT  16999.999999999996 211399.99999999997 17799.999999999996 212200.0 ;
      RECT  21799.999999999993 211399.99999999997 22599.999999999993 212200.0 ;
      RECT  26599.999999999996 211399.99999999997 27400.0 212200.0 ;
      RECT  31399.999999999996 211399.99999999997 32199.999999999996 212200.0 ;
      RECT  36200.0 211399.99999999997 37000.0 212200.0 ;
      RECT  41000.0 211399.99999999997 41800.0 212200.0 ;
      RECT  45800.0 211399.99999999997 46599.99999999999 212200.0 ;
      RECT  50600.0 211399.99999999997 51400.0 212200.0 ;
      RECT  55400.00000000001 211399.99999999997 56200.0 212200.0 ;
      RECT  60200.0 211399.99999999997 61000.0 212200.0 ;
      RECT  65000.0 211399.99999999997 65800.0 212200.0 ;
      RECT  69800.0 211399.99999999997 70600.0 212200.0 ;
      RECT  74600.00000000001 211399.99999999997 75400.0 212200.0 ;
      RECT  79400.0 211399.99999999997 80200.0 212200.0 ;
      RECT  84200.0 211399.99999999997 85000.0 212200.0 ;
      RECT  89000.0 211399.99999999997 89800.0 212200.0 ;
      RECT  93800.0 211399.99999999997 94600.0 212200.0 ;
      RECT  98600.00000000001 211399.99999999997 99400.0 212200.0 ;
      RECT  103400.0 211399.99999999997 104200.0 212200.0 ;
      RECT  108200.0 211399.99999999997 109000.0 212200.0 ;
      RECT  113000.00000000001 211399.99999999997 113800.00000000001 212200.0 ;
      RECT  117800.0 211399.99999999997 118600.0 212200.0 ;
      RECT  122600.00000000001 211399.99999999997 123400.0 212200.0 ;
      RECT  127400.0 211399.99999999997 128199.99999999999 212200.0 ;
      RECT  132200.0 211399.99999999997 133000.0 212200.0 ;
      RECT  137000.0 211399.99999999997 137800.0 212200.0 ;
      RECT  141800.0 211399.99999999997 142600.00000000003 212200.0 ;
      RECT  146600.0 211399.99999999997 147400.0 212200.0 ;
      RECT  151399.99999999997 211399.99999999997 152200.0 212200.0 ;
      RECT  156200.0 211399.99999999997 157000.0 212200.0 ;
      RECT  161000.0 211399.99999999997 161800.0 212200.0 ;
      RECT  165800.0 211399.99999999997 166600.00000000003 212200.0 ;
      RECT  170600.0 211399.99999999997 171400.0 212200.0 ;
      RECT  175399.99999999997 211399.99999999997 176200.0 212200.0 ;
      RECT  180200.0 211399.99999999997 181000.0 212200.0 ;
      RECT  185000.0 211399.99999999997 185800.0 212200.0 ;
      RECT  189800.0 211399.99999999997 190600.00000000003 212200.0 ;
      RECT  194600.0 211399.99999999997 195400.0 212200.0 ;
      RECT  199399.99999999997 211399.99999999997 200200.0 212200.0 ;
      RECT  204200.0 211399.99999999997 205000.0 212200.0 ;
      RECT  209000.0 211399.99999999997 209800.0 212200.0 ;
      RECT  7400.000000000003 216200.0 8200.000000000004 217000.0 ;
      RECT  12200.0 216200.0 13000.0 217000.0 ;
      RECT  16999.999999999996 216200.0 17799.999999999996 217000.0 ;
      RECT  21799.999999999993 216200.0 22599.999999999993 217000.0 ;
      RECT  26599.999999999996 216200.0 27400.0 217000.0 ;
      RECT  31399.999999999996 216200.0 32199.999999999996 217000.0 ;
      RECT  36200.0 216200.0 37000.0 217000.0 ;
      RECT  41000.0 216200.0 41800.0 217000.0 ;
      RECT  45800.0 216200.0 46599.99999999999 217000.0 ;
      RECT  50600.0 216200.0 51400.0 217000.0 ;
      RECT  55400.00000000001 216200.0 56200.0 217000.0 ;
      RECT  60200.0 216200.0 61000.0 217000.0 ;
      RECT  65000.0 216200.0 65800.0 217000.0 ;
      RECT  69800.0 216200.0 70600.0 217000.0 ;
      RECT  7400.000000000003 221000.0 8200.000000000004 221800.0 ;
      RECT  12200.0 221000.0 13000.0 221800.0 ;
      RECT  16999.999999999996 221000.0 17799.999999999996 221800.0 ;
      RECT  21799.999999999993 221000.0 22599.999999999993 221800.0 ;
      RECT  26599.999999999996 221000.0 27400.0 221800.0 ;
      RECT  41000.0 221000.0 41800.0 221800.0 ;
      RECT  45800.0 221000.0 46599.99999999999 221800.0 ;
      RECT  50600.0 221000.0 51400.0 221800.0 ;
      RECT  55400.00000000001 221000.0 56200.0 221800.0 ;
      RECT  60200.0 221000.0 61000.0 221800.0 ;
      RECT  65000.0 221000.0 65800.0 221800.0 ;
      RECT  69800.0 221000.0 70600.0 221800.0 ;
      RECT  74600.00000000001 221000.0 75400.0 221800.0 ;
      RECT  79400.0 221000.0 80200.0 221800.0 ;
      RECT  84200.0 221000.0 85000.0 221800.0 ;
      RECT  89000.0 221000.0 89800.0 221800.0 ;
      RECT  93800.0 221000.0 94600.0 221800.0 ;
      RECT  98600.00000000001 221000.0 99400.0 221800.0 ;
      RECT  103400.0 221000.0 104200.0 221800.0 ;
      RECT  108200.0 221000.0 109000.0 221800.0 ;
      RECT  113000.00000000001 221000.0 113800.00000000001 221800.0 ;
      RECT  117800.0 221000.0 118600.0 221800.0 ;
      RECT  122600.00000000001 221000.0 123400.0 221800.0 ;
      RECT  127400.0 221000.0 128199.99999999999 221800.0 ;
      RECT  132200.0 221000.0 133000.0 221800.0 ;
      RECT  137000.0 221000.0 137800.0 221800.0 ;
      RECT  141800.0 221000.0 142600.00000000003 221800.0 ;
      RECT  146600.0 221000.0 147400.0 221800.0 ;
      RECT  151399.99999999997 221000.0 152200.0 221800.0 ;
      RECT  156200.0 221000.0 157000.0 221800.0 ;
      RECT  161000.0 221000.0 161800.0 221800.0 ;
      RECT  165800.0 221000.0 166600.00000000003 221800.0 ;
      RECT  170600.0 221000.0 171400.0 221800.0 ;
      RECT  175399.99999999997 221000.0 176200.0 221800.0 ;
      RECT  180200.0 221000.0 181000.0 221800.0 ;
      RECT  185000.0 221000.0 185800.0 221800.0 ;
      RECT  189800.0 221000.0 190600.00000000003 221800.0 ;
      RECT  194600.0 221000.0 195400.0 221800.0 ;
      RECT  199399.99999999997 221000.0 200200.0 221800.0 ;
      RECT  204200.0 221000.0 205000.0 221800.0 ;
      RECT  209000.0 221000.0 209800.0 221800.0 ;
      RECT  7400.000000000003 225800.0 8200.000000000004 226600.00000000003 ;
      RECT  12200.0 225800.0 13000.0 226600.00000000003 ;
      RECT  16999.999999999996 225800.0 17799.999999999996 226600.00000000003 ;
      RECT  21799.999999999993 225800.0 22599.999999999993 226600.00000000003 ;
      RECT  26599.999999999996 225800.0 27400.0 226600.00000000003 ;
      RECT  31399.999999999996 225800.0 32199.999999999996 226600.00000000003 ;
      RECT  36200.0 225800.0 37000.0 226600.00000000003 ;
      RECT  41000.0 225800.0 41800.0 226600.00000000003 ;
      RECT  45800.0 225800.0 46599.99999999999 226600.00000000003 ;
      RECT  50600.0 225800.0 51400.0 226600.00000000003 ;
      RECT  55400.00000000001 225800.0 56200.0 226600.00000000003 ;
      RECT  60200.0 225800.0 61000.0 226600.00000000003 ;
      RECT  65000.0 225800.0 65800.0 226600.00000000003 ;
      RECT  69800.0 225800.0 70600.0 226600.00000000003 ;
      RECT  93800.0 225800.0 94600.0 226600.00000000003 ;
      RECT  98600.00000000001 225800.0 99400.0 226600.00000000003 ;
      RECT  103400.0 225800.0 104200.0 226600.00000000003 ;
      RECT  108200.0 225800.0 109000.0 226600.00000000003 ;
      RECT  113000.00000000001 225800.0 113800.00000000001 226600.00000000003 ;
      RECT  117800.0 225800.0 118600.0 226600.00000000003 ;
      RECT  122600.00000000001 225800.0 123400.0 226600.00000000003 ;
      RECT  127400.0 225800.0 128199.99999999999 226600.00000000003 ;
      RECT  132200.0 225800.0 133000.0 226600.00000000003 ;
      RECT  137000.0 225800.0 137800.0 226600.00000000003 ;
      RECT  141800.0 225800.0 142600.00000000003 226600.00000000003 ;
      RECT  146600.0 225800.0 147400.0 226600.00000000003 ;
      RECT  151399.99999999997 225800.0 152200.0 226600.00000000003 ;
      RECT  156200.0 225800.0 157000.0 226600.00000000003 ;
      RECT  161000.0 225800.0 161800.0 226600.00000000003 ;
      RECT  165800.0 225800.0 166600.00000000003 226600.00000000003 ;
      RECT  170600.0 225800.0 171400.0 226600.00000000003 ;
      RECT  175399.99999999997 225800.0 176200.0 226600.00000000003 ;
      RECT  180200.0 225800.0 181000.0 226600.00000000003 ;
      RECT  185000.0 225800.0 185800.0 226600.00000000003 ;
      RECT  189800.0 225800.0 190600.00000000003 226600.00000000003 ;
      RECT  194600.0 225800.0 195400.0 226600.00000000003 ;
      RECT  199399.99999999997 225800.0 200200.0 226600.00000000003 ;
      RECT  204200.0 225800.0 205000.0 226600.00000000003 ;
      RECT  209000.0 225800.0 209800.0 226600.00000000003 ;
      RECT  7400.000000000003 230600.00000000003 8200.000000000004 231400.00000000003 ;
      RECT  12200.0 230600.00000000003 13000.0 231400.00000000003 ;
      RECT  16999.999999999996 230600.00000000003 17799.999999999996 231400.00000000003 ;
      RECT  21799.999999999993 230600.00000000003 22599.999999999993 231400.00000000003 ;
      RECT  26599.999999999996 230600.00000000003 27400.0 231400.00000000003 ;
      RECT  31399.999999999996 230600.00000000003 32199.999999999996 231400.00000000003 ;
      RECT  36200.0 230600.00000000003 37000.0 231400.00000000003 ;
      RECT  41000.0 230600.00000000003 41800.0 231400.00000000003 ;
      RECT  45800.0 230600.00000000003 46599.99999999999 231400.00000000003 ;
      RECT  50600.0 230600.00000000003 51400.0 231400.00000000003 ;
      RECT  55400.00000000001 230600.00000000003 56200.0 231400.00000000003 ;
      RECT  60200.0 230600.00000000003 61000.0 231400.00000000003 ;
      RECT  65000.0 230600.00000000003 65800.0 231400.00000000003 ;
      RECT  69800.0 230600.00000000003 70600.0 231400.00000000003 ;
      RECT  74600.00000000001 230600.00000000003 75400.0 231400.00000000003 ;
      RECT  79400.0 230600.00000000003 80200.0 231400.00000000003 ;
      RECT  7400.000000000003 235399.99999999997 8200.000000000004 236200.0 ;
      RECT  12200.0 235399.99999999997 13000.0 236200.0 ;
      RECT  16999.999999999996 235399.99999999997 17799.999999999996 236200.0 ;
      RECT  21799.999999999993 235399.99999999997 22599.999999999993 236200.0 ;
      RECT  26599.999999999996 235399.99999999997 27400.0 236200.0 ;
      RECT  31399.999999999996 235399.99999999997 32199.999999999996 236200.0 ;
      RECT  36200.0 235399.99999999997 37000.0 236200.0 ;
      RECT  41000.0 235399.99999999997 41800.0 236200.0 ;
      RECT  45800.0 235399.99999999997 46599.99999999999 236200.0 ;
      RECT  50600.0 235399.99999999997 51400.0 236200.0 ;
      RECT  55400.00000000001 235399.99999999997 56200.0 236200.0 ;
      RECT  60200.0 235399.99999999997 61000.0 236200.0 ;
      RECT  65000.0 235399.99999999997 65800.0 236200.0 ;
      RECT  69800.0 235399.99999999997 70600.0 236200.0 ;
      RECT  74600.00000000001 235399.99999999997 75400.0 236200.0 ;
      RECT  79400.0 235399.99999999997 80200.0 236200.0 ;
      RECT  84200.0 235399.99999999997 85000.0 236200.0 ;
      RECT  89000.0 235399.99999999997 89800.0 236200.0 ;
      RECT  93800.0 235399.99999999997 94600.0 236200.0 ;
      RECT  98600.00000000001 235399.99999999997 99400.0 236200.0 ;
      RECT  103400.0 235399.99999999997 104200.0 236200.0 ;
      RECT  108200.0 235399.99999999997 109000.0 236200.0 ;
      RECT  113000.00000000001 235399.99999999997 113800.00000000001 236200.0 ;
      RECT  117800.0 235399.99999999997 118600.0 236200.0 ;
      RECT  122600.00000000001 235399.99999999997 123400.0 236200.0 ;
      RECT  127400.0 235399.99999999997 128199.99999999999 236200.0 ;
      RECT  132200.0 235399.99999999997 133000.0 236200.0 ;
      RECT  137000.0 235399.99999999997 137800.0 236200.0 ;
      RECT  141800.0 235399.99999999997 142600.00000000003 236200.0 ;
      RECT  146600.0 235399.99999999997 147400.0 236200.0 ;
      RECT  151399.99999999997 235399.99999999997 152200.0 236200.0 ;
      RECT  156200.0 235399.99999999997 157000.0 236200.0 ;
      RECT  161000.0 235399.99999999997 161800.0 236200.0 ;
      RECT  165800.0 235399.99999999997 166600.00000000003 236200.0 ;
      RECT  170600.0 235399.99999999997 171400.0 236200.0 ;
      RECT  175399.99999999997 235399.99999999997 176200.0 236200.0 ;
      RECT  180200.0 235399.99999999997 181000.0 236200.0 ;
      RECT  185000.0 235399.99999999997 185800.0 236200.0 ;
      RECT  189800.0 235399.99999999997 190600.00000000003 236200.0 ;
      RECT  194600.0 235399.99999999997 195400.0 236200.0 ;
      RECT  199399.99999999997 235399.99999999997 200200.0 236200.0 ;
      RECT  204200.0 235399.99999999997 205000.0 236200.0 ;
      RECT  209000.0 235399.99999999997 209800.0 236200.0 ;
      RECT  7400.000000000003 240200.0 8200.000000000004 241000.0 ;
      RECT  12200.0 240200.0 13000.0 241000.0 ;
      RECT  16999.999999999996 240200.0 17799.999999999996 241000.0 ;
      RECT  21799.999999999993 240200.0 22599.999999999993 241000.0 ;
      RECT  26599.999999999996 240200.0 27400.0 241000.0 ;
      RECT  41000.0 240200.0 41800.0 241000.0 ;
      RECT  45800.0 240200.0 46599.99999999999 241000.0 ;
      RECT  50600.0 240200.0 51400.0 241000.0 ;
      RECT  55400.00000000001 240200.0 56200.0 241000.0 ;
      RECT  60200.0 240200.0 61000.0 241000.0 ;
      RECT  65000.0 240200.0 65800.0 241000.0 ;
      RECT  69800.0 240200.0 70600.0 241000.0 ;
      RECT  74600.00000000001 240200.0 75400.0 241000.0 ;
      RECT  79400.0 240200.0 80200.0 241000.0 ;
      RECT  84200.0 240200.0 85000.0 241000.0 ;
      RECT  89000.0 240200.0 89800.0 241000.0 ;
      RECT  93800.0 240200.0 94600.0 241000.0 ;
      RECT  98600.00000000001 240200.0 99400.0 241000.0 ;
      RECT  103400.0 240200.0 104200.0 241000.0 ;
      RECT  108200.0 240200.0 109000.0 241000.0 ;
      RECT  113000.00000000001 240200.0 113800.00000000001 241000.0 ;
      RECT  117800.0 240200.0 118600.0 241000.0 ;
      RECT  122600.00000000001 240200.0 123400.0 241000.0 ;
      RECT  127400.0 240200.0 128199.99999999999 241000.0 ;
      RECT  132200.0 240200.0 133000.0 241000.0 ;
      RECT  137000.0 240200.0 137800.0 241000.0 ;
      RECT  141800.0 240200.0 142600.00000000003 241000.0 ;
      RECT  146600.0 240200.0 147400.0 241000.0 ;
      RECT  151399.99999999997 240200.0 152200.0 241000.0 ;
      RECT  156200.0 240200.0 157000.0 241000.0 ;
      RECT  161000.0 240200.0 161800.0 241000.0 ;
      RECT  165800.0 240200.0 166600.00000000003 241000.0 ;
      RECT  170600.0 240200.0 171400.0 241000.0 ;
      RECT  175399.99999999997 240200.0 176200.0 241000.0 ;
      RECT  180200.0 240200.0 181000.0 241000.0 ;
      RECT  185000.0 240200.0 185800.0 241000.0 ;
      RECT  189800.0 240200.0 190600.00000000003 241000.0 ;
      RECT  194600.0 240200.0 195400.0 241000.0 ;
      RECT  199399.99999999997 240200.0 200200.0 241000.0 ;
      RECT  204200.0 240200.0 205000.0 241000.0 ;
      RECT  209000.0 240200.0 209800.0 241000.0 ;
      RECT  7400.000000000003 245000.0 8200.000000000004 245800.0 ;
      RECT  12200.0 245000.0 13000.0 245800.0 ;
      RECT  16999.999999999996 245000.0 17799.999999999996 245800.0 ;
      RECT  21799.999999999993 245000.0 22599.999999999993 245800.0 ;
      RECT  26599.999999999996 245000.0 27400.0 245800.0 ;
      RECT  31399.999999999996 245000.0 32199.999999999996 245800.0 ;
      RECT  36200.0 245000.0 37000.0 245800.0 ;
      RECT  41000.0 245000.0 41800.0 245800.0 ;
      RECT  45800.0 245000.0 46599.99999999999 245800.0 ;
      RECT  50600.0 245000.0 51400.0 245800.0 ;
      RECT  55400.00000000001 245000.0 56200.0 245800.0 ;
      RECT  60200.0 245000.0 61000.0 245800.0 ;
      RECT  65000.0 245000.0 65800.0 245800.0 ;
      RECT  69800.0 245000.0 70600.0 245800.0 ;
      RECT  74600.00000000001 245000.0 75400.0 245800.0 ;
      RECT  79400.0 245000.0 80200.0 245800.0 ;
      RECT  84200.0 245000.0 85000.0 245800.0 ;
      RECT  89000.0 245000.0 89800.0 245800.0 ;
      RECT  93800.0 245000.0 94600.0 245800.0 ;
      RECT  98600.00000000001 245000.0 99400.0 245800.0 ;
      RECT  103400.0 245000.0 104200.0 245800.0 ;
      RECT  108200.0 245000.0 109000.0 245800.0 ;
      RECT  113000.00000000001 245000.0 113800.00000000001 245800.0 ;
      RECT  117800.0 245000.0 118600.0 245800.0 ;
      RECT  122600.00000000001 245000.0 123400.0 245800.0 ;
      RECT  127400.0 245000.0 128199.99999999999 245800.0 ;
      RECT  132200.0 245000.0 133000.0 245800.0 ;
      RECT  137000.0 245000.0 137800.0 245800.0 ;
      RECT  141800.0 245000.0 142600.00000000003 245800.0 ;
      RECT  146600.0 245000.0 147400.0 245800.0 ;
      RECT  151399.99999999997 245000.0 152200.0 245800.0 ;
      RECT  156200.0 245000.0 157000.0 245800.0 ;
      RECT  161000.0 245000.0 161800.0 245800.0 ;
      RECT  165800.0 245000.0 166600.00000000003 245800.0 ;
      RECT  170600.0 245000.0 171400.0 245800.0 ;
      RECT  175399.99999999997 245000.0 176200.0 245800.0 ;
      RECT  180200.0 245000.0 181000.0 245800.0 ;
      RECT  185000.0 245000.0 185800.0 245800.0 ;
      RECT  189800.0 245000.0 190600.00000000003 245800.0 ;
      RECT  194600.0 245000.0 195400.0 245800.0 ;
      RECT  199399.99999999997 245000.0 200200.0 245800.0 ;
      RECT  204200.0 245000.0 205000.0 245800.0 ;
      RECT  209000.0 245000.0 209800.0 245800.0 ;
      RECT  7400.000000000003 249800.0 8200.000000000004 250600.00000000003 ;
      RECT  12200.0 249800.0 13000.0 250600.00000000003 ;
      RECT  16999.999999999996 249800.0 17799.999999999996 250600.00000000003 ;
      RECT  21799.999999999993 249800.0 22599.999999999993 250600.00000000003 ;
      RECT  26599.999999999996 249800.0 27400.0 250600.00000000003 ;
      RECT  31399.999999999996 249800.0 32199.999999999996 250600.00000000003 ;
      RECT  36200.0 249800.0 37000.0 250600.00000000003 ;
      RECT  41000.0 249800.0 41800.0 250600.00000000003 ;
      RECT  45800.0 249800.0 46599.99999999999 250600.00000000003 ;
      RECT  50600.0 249800.0 51400.0 250600.00000000003 ;
      RECT  55400.00000000001 249800.0 56200.0 250600.00000000003 ;
      RECT  60200.0 249800.0 61000.0 250600.00000000003 ;
      RECT  65000.0 249800.0 65800.0 250600.00000000003 ;
      RECT  69800.0 249800.0 70600.0 250600.00000000003 ;
      RECT  74600.00000000001 249800.0 75400.0 250600.00000000003 ;
      RECT  79400.0 249800.0 80200.0 250600.00000000003 ;
      RECT  84200.0 249800.0 85000.0 250600.00000000003 ;
      RECT  89000.0 249800.0 89800.0 250600.00000000003 ;
      RECT  93800.0 249800.0 94600.0 250600.00000000003 ;
      RECT  98600.00000000001 249800.0 99400.0 250600.00000000003 ;
      RECT  103400.0 249800.0 104200.0 250600.00000000003 ;
      RECT  108200.0 249800.0 109000.0 250600.00000000003 ;
      RECT  113000.00000000001 249800.0 113800.00000000001 250600.00000000003 ;
      RECT  117800.0 249800.0 118600.0 250600.00000000003 ;
      RECT  122600.00000000001 249800.0 123400.0 250600.00000000003 ;
      RECT  7400.000000000003 254600.00000000003 8200.000000000004 255400.00000000003 ;
      RECT  12200.0 254600.00000000003 13000.0 255400.00000000003 ;
      RECT  16999.999999999996 254600.00000000003 17799.999999999996 255400.00000000003 ;
      RECT  21799.999999999993 254600.00000000003 22599.999999999993 255400.00000000003 ;
      RECT  26599.999999999996 254600.00000000003 27400.0 255400.00000000003 ;
      RECT  31399.999999999996 254600.00000000003 32199.999999999996 255400.00000000003 ;
      RECT  36200.0 254600.00000000003 37000.0 255400.00000000003 ;
      RECT  41000.0 254600.00000000003 41800.0 255400.00000000003 ;
      RECT  45800.0 254600.00000000003 46599.99999999999 255400.00000000003 ;
      RECT  50600.0 254600.00000000003 51400.0 255400.00000000003 ;
      RECT  55400.00000000001 254600.00000000003 56200.0 255400.00000000003 ;
      RECT  60200.0 254600.00000000003 61000.0 255400.00000000003 ;
      RECT  65000.0 254600.00000000003 65800.0 255400.00000000003 ;
      RECT  69800.0 254600.00000000003 70600.0 255400.00000000003 ;
      RECT  74600.00000000001 254600.00000000003 75400.0 255400.00000000003 ;
      RECT  79400.0 254600.00000000003 80200.0 255400.00000000003 ;
      RECT  84200.0 254600.00000000003 85000.0 255400.00000000003 ;
      RECT  89000.0 254600.00000000003 89800.0 255400.00000000003 ;
      RECT  93800.0 254600.00000000003 94600.0 255400.00000000003 ;
      RECT  98600.00000000001 254600.00000000003 99400.0 255400.00000000003 ;
      RECT  103400.0 254600.00000000003 104200.0 255400.00000000003 ;
      RECT  108200.0 254600.00000000003 109000.0 255400.00000000003 ;
      RECT  113000.00000000001 254600.00000000003 113800.00000000001 255400.00000000003 ;
      RECT  117800.0 254600.00000000003 118600.0 255400.00000000003 ;
      RECT  122600.00000000001 254600.00000000003 123400.0 255400.00000000003 ;
      RECT  127400.0 254600.00000000003 128199.99999999999 255400.00000000003 ;
      RECT  132200.0 254600.00000000003 133000.0 255400.00000000003 ;
      RECT  137000.0 254600.00000000003 137800.0 255400.00000000003 ;
      RECT  141800.0 254600.00000000003 142600.00000000003 255400.00000000003 ;
      RECT  146600.0 254600.00000000003 147400.0 255400.00000000003 ;
      RECT  151399.99999999997 254600.00000000003 152200.0 255400.00000000003 ;
      RECT  156200.0 254600.00000000003 157000.0 255400.00000000003 ;
      RECT  161000.0 254600.00000000003 161800.0 255400.00000000003 ;
      RECT  165800.0 254600.00000000003 166600.00000000003 255400.00000000003 ;
      RECT  170600.0 254600.00000000003 171400.0 255400.00000000003 ;
      RECT  175399.99999999997 254600.00000000003 176200.0 255400.00000000003 ;
      RECT  180200.0 254600.00000000003 181000.0 255400.00000000003 ;
      RECT  185000.0 254600.00000000003 185800.0 255400.00000000003 ;
      RECT  189800.0 254600.00000000003 190600.00000000003 255400.00000000003 ;
      RECT  194600.0 254600.00000000003 195400.0 255400.00000000003 ;
      RECT  199399.99999999997 254600.00000000003 200200.0 255400.00000000003 ;
      RECT  204200.0 254600.00000000003 205000.0 255400.00000000003 ;
      RECT  209000.0 254600.00000000003 209800.0 255400.00000000003 ;
      RECT  7400.000000000003 259399.99999999997 8200.000000000004 260200.0 ;
      RECT  12200.0 259399.99999999997 13000.0 260200.0 ;
      RECT  16999.999999999996 259399.99999999997 17799.999999999996 260200.0 ;
      RECT  21799.999999999993 259399.99999999997 22599.999999999993 260200.0 ;
      RECT  26599.999999999996 259399.99999999997 27400.0 260200.0 ;
      RECT  31399.999999999996 259399.99999999997 32199.999999999996 260200.0 ;
      RECT  36200.0 259399.99999999997 37000.0 260200.0 ;
      RECT  41000.0 259399.99999999997 41800.0 260200.0 ;
      RECT  84200.0 259399.99999999997 85000.0 260200.0 ;
      RECT  89000.0 259399.99999999997 89800.0 260200.0 ;
      RECT  93800.0 259399.99999999997 94600.0 260200.0 ;
      RECT  98600.00000000001 259399.99999999997 99400.0 260200.0 ;
      RECT  103400.0 259399.99999999997 104200.0 260200.0 ;
      RECT  108200.0 259399.99999999997 109000.0 260200.0 ;
      RECT  113000.00000000001 259399.99999999997 113800.00000000001 260200.0 ;
      RECT  117800.0 259399.99999999997 118600.0 260200.0 ;
      RECT  122600.00000000001 259399.99999999997 123400.0 260200.0 ;
      RECT  127400.0 259399.99999999997 128199.99999999999 260200.0 ;
      RECT  132200.0 259399.99999999997 133000.0 260200.0 ;
      RECT  137000.0 259399.99999999997 137800.0 260200.0 ;
      RECT  141800.0 259399.99999999997 142600.00000000003 260200.0 ;
      RECT  146600.0 259399.99999999997 147400.0 260200.0 ;
      RECT  151399.99999999997 259399.99999999997 152200.0 260200.0 ;
      RECT  156200.0 259399.99999999997 157000.0 260200.0 ;
      RECT  161000.0 259399.99999999997 161800.0 260200.0 ;
      RECT  165800.0 259399.99999999997 166600.00000000003 260200.0 ;
      RECT  170600.0 259399.99999999997 171400.0 260200.0 ;
      RECT  175399.99999999997 259399.99999999997 176200.0 260200.0 ;
      RECT  180200.0 259399.99999999997 181000.0 260200.0 ;
      RECT  185000.0 259399.99999999997 185800.0 260200.0 ;
      RECT  189800.0 259399.99999999997 190600.00000000003 260200.0 ;
      RECT  194600.0 259399.99999999997 195400.0 260200.0 ;
      RECT  199399.99999999997 259399.99999999997 200200.0 260200.0 ;
      RECT  204200.0 259399.99999999997 205000.0 260200.0 ;
      RECT  209000.0 259399.99999999997 209800.0 260200.0 ;
      RECT  7400.000000000003 264200.0 8200.000000000004 265000.0 ;
      RECT  12200.0 264200.0 13000.0 265000.0 ;
      RECT  16999.999999999996 264200.0 17799.999999999996 265000.0 ;
      RECT  21799.999999999993 264200.0 22599.999999999993 265000.0 ;
      RECT  26599.999999999996 264200.0 27400.0 265000.0 ;
      RECT  31399.999999999996 264200.0 32199.999999999996 265000.0 ;
      RECT  36200.0 264200.0 37000.0 265000.0 ;
      RECT  41000.0 264200.0 41800.0 265000.0 ;
      RECT  45800.0 264200.0 46599.99999999999 265000.0 ;
      RECT  50600.0 264200.0 51400.0 265000.0 ;
      RECT  55400.00000000001 264200.0 56200.0 265000.0 ;
      RECT  60200.0 264200.0 61000.0 265000.0 ;
      RECT  84200.0 264200.0 85000.0 265000.0 ;
      RECT  89000.0 264200.0 89800.0 265000.0 ;
      RECT  93800.0 264200.0 94600.0 265000.0 ;
      RECT  98600.00000000001 264200.0 99400.0 265000.0 ;
      RECT  103400.0 264200.0 104200.0 265000.0 ;
      RECT  108200.0 264200.0 109000.0 265000.0 ;
      RECT  113000.00000000001 264200.0 113800.00000000001 265000.0 ;
      RECT  117800.0 264200.0 118600.0 265000.0 ;
      RECT  122600.00000000001 264200.0 123400.0 265000.0 ;
      RECT  127400.0 264200.0 128199.99999999999 265000.0 ;
      RECT  132200.0 264200.0 133000.0 265000.0 ;
      RECT  137000.0 264200.0 137800.0 265000.0 ;
      RECT  141800.0 264200.0 142600.00000000003 265000.0 ;
      RECT  146600.0 264200.0 147400.0 265000.0 ;
      RECT  151399.99999999997 264200.0 152200.0 265000.0 ;
      RECT  156200.0 264200.0 157000.0 265000.0 ;
      RECT  161000.0 264200.0 161800.0 265000.0 ;
      RECT  165800.0 264200.0 166600.00000000003 265000.0 ;
      RECT  170600.0 264200.0 171400.0 265000.0 ;
      RECT  175399.99999999997 264200.0 176200.0 265000.0 ;
      RECT  180200.0 264200.0 181000.0 265000.0 ;
      RECT  185000.0 264200.0 185800.0 265000.0 ;
      RECT  189800.0 264200.0 190600.00000000003 265000.0 ;
      RECT  194600.0 264200.0 195400.0 265000.0 ;
      RECT  199399.99999999997 264200.0 200200.0 265000.0 ;
      RECT  204200.0 264200.0 205000.0 265000.0 ;
      RECT  209000.0 264200.0 209800.0 265000.0 ;
      RECT  7400.000000000003 269000.0 8200.000000000004 269800.0 ;
      RECT  12200.0 269000.0 13000.0 269800.0 ;
      RECT  16999.999999999996 269000.0 17799.999999999996 269800.0 ;
      RECT  21799.999999999993 269000.0 22599.999999999993 269800.0 ;
      RECT  26599.999999999996 269000.0 27400.0 269800.0 ;
      RECT  31399.999999999996 269000.0 32199.999999999996 269800.0 ;
      RECT  36200.0 269000.0 37000.0 269800.0 ;
      RECT  41000.0 269000.0 41800.0 269800.0 ;
      RECT  45800.0 269000.0 46599.99999999999 269800.0 ;
      RECT  50600.0 269000.0 51400.0 269800.0 ;
      RECT  55400.00000000001 269000.0 56200.0 269800.0 ;
      RECT  60200.0 269000.0 61000.0 269800.0 ;
      RECT  65000.0 269000.0 65800.0 269800.0 ;
      RECT  69800.0 269000.0 70600.0 269800.0 ;
      RECT  74600.00000000001 269000.0 75400.0 269800.0 ;
      RECT  79400.0 269000.0 80200.0 269800.0 ;
      RECT  84200.0 269000.0 85000.0 269800.0 ;
      RECT  89000.0 269000.0 89800.0 269800.0 ;
      RECT  93800.0 269000.0 94600.0 269800.0 ;
      RECT  98600.00000000001 269000.0 99400.0 269800.0 ;
      RECT  103400.0 269000.0 104200.0 269800.0 ;
      RECT  108200.0 269000.0 109000.0 269800.0 ;
      RECT  113000.00000000001 269000.0 113800.00000000001 269800.0 ;
      RECT  117800.0 269000.0 118600.0 269800.0 ;
      RECT  122600.00000000001 269000.0 123400.0 269800.0 ;
      RECT  7400.000000000003 273800.0 8200.000000000004 274600.0 ;
      RECT  12200.0 273800.0 13000.0 274600.0 ;
      RECT  16999.999999999996 273800.0 17799.999999999996 274600.0 ;
      RECT  21799.999999999993 273800.0 22599.999999999993 274600.0 ;
      RECT  26599.999999999996 273800.0 27400.0 274600.0 ;
      RECT  31399.999999999996 273800.0 32199.999999999996 274600.0 ;
      RECT  36200.0 273800.0 37000.0 274600.0 ;
      RECT  41000.0 273800.0 41800.0 274600.0 ;
      RECT  45800.0 273800.0 46599.99999999999 274600.0 ;
      RECT  50600.0 273800.0 51400.0 274600.0 ;
      RECT  69800.0 273800.0 70600.0 274600.0 ;
      RECT  74600.00000000001 273800.0 75400.0 274600.0 ;
      RECT  79400.0 273800.0 80200.0 274600.0 ;
      RECT  84200.0 273800.0 85000.0 274600.0 ;
      RECT  89000.0 273800.0 89800.0 274600.0 ;
      RECT  93800.0 273800.0 94600.0 274600.0 ;
      RECT  98600.00000000001 273800.0 99400.0 274600.0 ;
      RECT  103400.0 273800.0 104200.0 274600.0 ;
      RECT  108200.0 273800.0 109000.0 274600.0 ;
      RECT  113000.00000000001 273800.0 113800.00000000001 274600.0 ;
      RECT  117800.0 273800.0 118600.0 274600.0 ;
      RECT  122600.00000000001 273800.0 123400.0 274600.0 ;
      RECT  127400.0 273800.0 128199.99999999999 274600.0 ;
      RECT  132200.0 273800.0 133000.0 274600.0 ;
      RECT  137000.0 273800.0 137800.0 274600.0 ;
      RECT  141800.0 273800.0 142600.00000000003 274600.0 ;
      RECT  146600.0 273800.0 147400.0 274600.0 ;
      RECT  151399.99999999997 273800.0 152200.0 274600.0 ;
      RECT  156200.0 273800.0 157000.0 274600.0 ;
      RECT  161000.0 273800.0 161800.0 274600.0 ;
      RECT  165800.0 273800.0 166600.00000000003 274600.0 ;
      RECT  170600.0 273800.0 171400.0 274600.0 ;
      RECT  175399.99999999997 273800.0 176200.0 274600.0 ;
      RECT  180200.0 273800.0 181000.0 274600.0 ;
      RECT  185000.0 273800.0 185800.0 274600.0 ;
      RECT  189800.0 273800.0 190600.00000000003 274600.0 ;
      RECT  194600.0 273800.0 195400.0 274600.0 ;
      RECT  199399.99999999997 273800.0 200200.0 274600.0 ;
      RECT  204200.0 273800.0 205000.0 274600.0 ;
      RECT  209000.0 273800.0 209800.0 274600.0 ;
      RECT  7400.000000000003 278600.0 8200.000000000004 279400.00000000006 ;
      RECT  12200.0 278600.0 13000.0 279400.00000000006 ;
      RECT  16999.999999999996 278600.0 17799.999999999996 279400.00000000006 ;
      RECT  21799.999999999993 278600.0 22599.999999999993 279400.00000000006 ;
      RECT  26599.999999999996 278600.0 27400.0 279400.00000000006 ;
      RECT  31399.999999999996 278600.0 32199.999999999996 279400.00000000006 ;
      RECT  36200.0 278600.0 37000.0 279400.00000000006 ;
      RECT  41000.0 278600.0 41800.0 279400.00000000006 ;
      RECT  45800.0 278600.0 46599.99999999999 279400.00000000006 ;
      RECT  50600.0 278600.0 51400.0 279400.00000000006 ;
      RECT  55400.00000000001 278600.0 56200.0 279400.00000000006 ;
      RECT  60200.0 278600.0 61000.0 279400.00000000006 ;
      RECT  65000.0 278600.0 65800.0 279400.00000000006 ;
      RECT  69800.0 278600.0 70600.0 279400.00000000006 ;
      RECT  74600.00000000001 278600.0 75400.0 279400.00000000006 ;
      RECT  79400.0 278600.0 80200.0 279400.00000000006 ;
      RECT  84200.0 278600.0 85000.0 279400.00000000006 ;
      RECT  89000.0 278600.0 89800.0 279400.00000000006 ;
      RECT  93800.0 278600.0 94600.0 279400.00000000006 ;
      RECT  98600.00000000001 278600.0 99400.0 279400.00000000006 ;
      RECT  103400.0 278600.0 104200.0 279400.00000000006 ;
      RECT  108200.0 278600.0 109000.0 279400.00000000006 ;
      RECT  113000.00000000001 278600.0 113800.00000000001 279400.00000000006 ;
      RECT  117800.0 278600.0 118600.0 279400.00000000006 ;
      RECT  122600.00000000001 278600.0 123400.0 279400.00000000006 ;
      RECT  127400.0 278600.0 128199.99999999999 279400.00000000006 ;
      RECT  132200.0 278600.0 133000.0 279400.00000000006 ;
      RECT  137000.0 278600.0 137800.0 279400.00000000006 ;
      RECT  141800.0 278600.0 142600.00000000003 279400.00000000006 ;
      RECT  146600.0 278600.0 147400.0 279400.00000000006 ;
      RECT  151399.99999999997 278600.0 152200.0 279400.00000000006 ;
      RECT  156200.0 278600.0 157000.0 279400.00000000006 ;
      RECT  161000.0 278600.0 161800.0 279400.00000000006 ;
      RECT  165800.0 278600.0 166600.00000000003 279400.00000000006 ;
      RECT  170600.0 278600.0 171400.0 279400.00000000006 ;
      RECT  175399.99999999997 278600.0 176200.0 279400.00000000006 ;
      RECT  180200.0 278600.0 181000.0 279400.00000000006 ;
      RECT  185000.0 278600.0 185800.0 279400.00000000006 ;
      RECT  189800.0 278600.0 190600.00000000003 279400.00000000006 ;
      RECT  194600.0 278600.0 195400.0 279400.00000000006 ;
      RECT  199399.99999999997 278600.0 200200.0 279400.00000000006 ;
      RECT  204200.0 278600.0 205000.0 279400.00000000006 ;
      RECT  209000.0 278600.0 209800.0 279400.00000000006 ;
      RECT  7400.000000000003 283400.0 8200.000000000004 284200.0 ;
      RECT  12200.0 283400.0 13000.0 284200.0 ;
      RECT  16999.999999999996 283400.0 17799.999999999996 284200.0 ;
      RECT  21799.999999999993 283400.0 22599.999999999993 284200.0 ;
      RECT  26599.999999999996 283400.0 27400.0 284200.0 ;
      RECT  31399.999999999996 283400.0 32199.999999999996 284200.0 ;
      RECT  36200.0 283400.0 37000.0 284200.0 ;
      RECT  41000.0 283400.0 41800.0 284200.0 ;
      RECT  45800.0 283400.0 46599.99999999999 284200.0 ;
      RECT  50600.0 283400.0 51400.0 284200.0 ;
      RECT  55400.00000000001 283400.0 56200.0 284200.0 ;
      RECT  60200.0 283400.0 61000.0 284200.0 ;
      RECT  65000.0 283400.0 65800.0 284200.0 ;
      RECT  69800.0 283400.0 70600.0 284200.0 ;
      RECT  74600.00000000001 283400.0 75400.0 284200.0 ;
      RECT  79400.0 283400.0 80200.0 284200.0 ;
      RECT  84200.0 283400.0 85000.0 284200.0 ;
      RECT  89000.0 283400.0 89800.0 284200.0 ;
      RECT  93800.0 283400.0 94600.0 284200.0 ;
      RECT  98600.00000000001 283400.0 99400.0 284200.0 ;
      RECT  103400.0 283400.0 104200.0 284200.0 ;
      RECT  108200.0 283400.0 109000.0 284200.0 ;
      RECT  113000.00000000001 283400.0 113800.00000000001 284200.0 ;
      RECT  117800.0 283400.0 118600.0 284200.0 ;
      RECT  122600.00000000001 283400.0 123400.0 284200.0 ;
      RECT  127400.0 283400.0 128199.99999999999 284200.0 ;
      RECT  132200.0 283400.0 133000.0 284200.0 ;
      RECT  137000.0 283400.0 137800.0 284200.0 ;
      RECT  141800.0 283400.0 142600.00000000003 284200.0 ;
      RECT  146600.0 283400.0 147400.0 284200.0 ;
      RECT  151399.99999999997 283400.0 152200.0 284200.0 ;
      RECT  156200.0 283400.0 157000.0 284200.0 ;
      RECT  161000.0 283400.0 161800.0 284200.0 ;
      RECT  165800.0 283400.0 166600.00000000003 284200.0 ;
      RECT  170600.0 283400.0 171400.0 284200.0 ;
      RECT  175399.99999999997 283400.0 176200.0 284200.0 ;
      RECT  180200.0 283400.0 181000.0 284200.0 ;
      RECT  185000.0 283400.0 185800.0 284200.0 ;
      RECT  189800.0 283400.0 190600.00000000003 284200.0 ;
      RECT  194600.0 283400.0 195400.0 284200.0 ;
      RECT  199399.99999999997 283400.0 200200.0 284200.0 ;
      RECT  204200.0 283400.0 205000.0 284200.0 ;
      RECT  209000.0 283400.0 209800.0 284200.0 ;
      RECT  7400.000000000003 288200.0 8200.000000000004 289000.0 ;
      RECT  12200.0 288200.0 13000.0 289000.0 ;
      RECT  16999.999999999996 288200.0 17799.999999999996 289000.0 ;
      RECT  21799.999999999993 288200.0 22599.999999999993 289000.0 ;
      RECT  26599.999999999996 288200.0 27400.0 289000.0 ;
      RECT  31399.999999999996 288200.0 32199.999999999996 289000.0 ;
      RECT  36200.0 288200.0 37000.0 289000.0 ;
      RECT  41000.0 288200.0 41800.0 289000.0 ;
      RECT  45800.0 288200.0 46599.99999999999 289000.0 ;
      RECT  50600.0 288200.0 51400.0 289000.0 ;
      RECT  55400.00000000001 288200.0 56200.0 289000.0 ;
      RECT  60200.0 288200.0 61000.0 289000.0 ;
      RECT  65000.0 288200.0 65800.0 289000.0 ;
      RECT  69800.0 288200.0 70600.0 289000.0 ;
      RECT  74600.00000000001 288200.0 75400.0 289000.0 ;
      RECT  79400.0 288200.0 80200.0 289000.0 ;
      RECT  84200.0 288200.0 85000.0 289000.0 ;
      RECT  89000.0 288200.0 89800.0 289000.0 ;
      RECT  93800.0 288200.0 94600.0 289000.0 ;
      RECT  98600.00000000001 288200.0 99400.0 289000.0 ;
      RECT  103400.0 288200.0 104200.0 289000.0 ;
      RECT  108200.0 288200.0 109000.0 289000.0 ;
      RECT  113000.00000000001 288200.0 113800.00000000001 289000.0 ;
      RECT  117800.0 288200.0 118600.0 289000.0 ;
      RECT  122600.00000000001 288200.0 123400.0 289000.0 ;
      RECT  7400.000000000003 293000.0 8200.000000000004 293800.0 ;
      RECT  12200.0 293000.0 13000.0 293800.0 ;
      RECT  16999.999999999996 293000.0 17799.999999999996 293800.0 ;
      RECT  21799.999999999993 293000.0 22599.999999999993 293800.0 ;
      RECT  26599.999999999996 293000.0 27400.0 293800.0 ;
      RECT  31399.999999999996 293000.0 32199.999999999996 293800.0 ;
      RECT  36200.0 293000.0 37000.0 293800.0 ;
      RECT  41000.0 293000.0 41800.0 293800.0 ;
      RECT  45800.0 293000.0 46599.99999999999 293800.0 ;
      RECT  50600.0 293000.0 51400.0 293800.0 ;
      RECT  55400.00000000001 293000.0 56200.0 293800.0 ;
      RECT  60200.0 293000.0 61000.0 293800.0 ;
      RECT  65000.0 293000.0 65800.0 293800.0 ;
      RECT  69800.0 293000.0 70600.0 293800.0 ;
      RECT  74600.00000000001 293000.0 75400.0 293800.0 ;
      RECT  79400.0 293000.0 80200.0 293800.0 ;
      RECT  84200.0 293000.0 85000.0 293800.0 ;
      RECT  89000.0 293000.0 89800.0 293800.0 ;
      RECT  93800.0 293000.0 94600.0 293800.0 ;
      RECT  98600.00000000001 293000.0 99400.0 293800.0 ;
      RECT  103400.0 293000.0 104200.0 293800.0 ;
      RECT  108200.0 293000.0 109000.0 293800.0 ;
      RECT  113000.00000000001 293000.0 113800.00000000001 293800.0 ;
      RECT  117800.0 293000.0 118600.0 293800.0 ;
      RECT  122600.00000000001 293000.0 123400.0 293800.0 ;
      RECT  127400.0 293000.0 128199.99999999999 293800.0 ;
      RECT  132200.0 293000.0 133000.0 293800.0 ;
      RECT  137000.0 293000.0 137800.0 293800.0 ;
      RECT  141800.0 293000.0 142600.00000000003 293800.0 ;
      RECT  146600.0 293000.0 147400.0 293800.0 ;
      RECT  151399.99999999997 293000.0 152200.0 293800.0 ;
      RECT  156200.0 293000.0 157000.0 293800.0 ;
      RECT  161000.0 293000.0 161800.0 293800.0 ;
      RECT  165800.0 293000.0 166600.00000000003 293800.0 ;
      RECT  170600.0 293000.0 171400.0 293800.0 ;
      RECT  175399.99999999997 293000.0 176200.0 293800.0 ;
      RECT  180200.0 293000.0 181000.0 293800.0 ;
      RECT  185000.0 293000.0 185800.0 293800.0 ;
      RECT  189800.0 293000.0 190600.00000000003 293800.0 ;
      RECT  194600.0 293000.0 195400.0 293800.0 ;
      RECT  199399.99999999997 293000.0 200200.0 293800.0 ;
      RECT  204200.0 293000.0 205000.0 293800.0 ;
      RECT  209000.0 293000.0 209800.0 293800.0 ;
      RECT  7400.000000000003 297800.0 8200.000000000004 298600.0 ;
      RECT  12200.0 297800.0 13000.0 298600.0 ;
      RECT  16999.999999999996 297800.0 17799.999999999996 298600.0 ;
      RECT  21799.999999999993 297800.0 22599.999999999993 298600.0 ;
      RECT  26599.999999999996 297800.0 27400.0 298600.0 ;
      RECT  31399.999999999996 297800.0 32199.999999999996 298600.0 ;
      RECT  36200.0 297800.0 37000.0 298600.0 ;
      RECT  41000.0 297800.0 41800.0 298600.0 ;
      RECT  45800.0 297800.0 46599.99999999999 298600.0 ;
      RECT  50600.0 297800.0 51400.0 298600.0 ;
      RECT  55400.00000000001 297800.0 56200.0 298600.0 ;
      RECT  60200.0 297800.0 61000.0 298600.0 ;
      RECT  65000.0 297800.0 65800.0 298600.0 ;
      RECT  69800.0 297800.0 70600.0 298600.0 ;
      RECT  74600.00000000001 297800.0 75400.0 298600.0 ;
      RECT  79400.0 297800.0 80200.0 298600.0 ;
      RECT  84200.0 297800.0 85000.0 298600.0 ;
      RECT  89000.0 297800.0 89800.0 298600.0 ;
      RECT  93800.0 297800.0 94600.0 298600.0 ;
      RECT  98600.00000000001 297800.0 99400.0 298600.0 ;
      RECT  103400.0 297800.0 104200.0 298600.0 ;
      RECT  108200.0 297800.0 109000.0 298600.0 ;
      RECT  113000.00000000001 297800.0 113800.00000000001 298600.0 ;
      RECT  117800.0 297800.0 118600.0 298600.0 ;
      RECT  122600.00000000001 297800.0 123400.0 298600.0 ;
      RECT  127400.0 297800.0 128199.99999999999 298600.0 ;
      RECT  132200.0 297800.0 133000.0 298600.0 ;
      RECT  137000.0 297800.0 137800.0 298600.0 ;
      RECT  141800.0 297800.0 142600.00000000003 298600.0 ;
      RECT  146600.0 297800.0 147400.0 298600.0 ;
      RECT  151399.99999999997 297800.0 152200.0 298600.0 ;
      RECT  156200.0 297800.0 157000.0 298600.0 ;
      RECT  161000.0 297800.0 161800.0 298600.0 ;
      RECT  165800.0 297800.0 166600.00000000003 298600.0 ;
      RECT  170600.0 297800.0 171400.0 298600.0 ;
      RECT  175399.99999999997 297800.0 176200.0 298600.0 ;
      RECT  180200.0 297800.0 181000.0 298600.0 ;
      RECT  185000.0 297800.0 185800.0 298600.0 ;
      RECT  189800.0 297800.0 190600.00000000003 298600.0 ;
      RECT  194600.0 297800.0 195400.0 298600.0 ;
      RECT  199399.99999999997 297800.0 200200.0 298600.0 ;
      RECT  204200.0 297800.0 205000.0 298600.0 ;
      RECT  209000.0 297800.0 209800.0 298600.0 ;
      RECT  7400.000000000003 302600.0 8200.000000000004 303400.00000000006 ;
      RECT  12200.0 302600.0 13000.0 303400.00000000006 ;
      RECT  16999.999999999996 302600.0 17799.999999999996 303400.00000000006 ;
      RECT  21799.999999999993 302600.0 22599.999999999993 303400.00000000006 ;
      RECT  26599.999999999996 302600.0 27400.0 303400.00000000006 ;
      RECT  31399.999999999996 302600.0 32199.999999999996 303400.00000000006 ;
      RECT  36200.0 302600.0 37000.0 303400.00000000006 ;
      RECT  41000.0 302600.0 41800.0 303400.00000000006 ;
      RECT  45800.0 302600.0 46599.99999999999 303400.00000000006 ;
      RECT  50600.0 302600.0 51400.0 303400.00000000006 ;
      RECT  55400.00000000001 302600.0 56200.0 303400.00000000006 ;
      RECT  60200.0 302600.0 61000.0 303400.00000000006 ;
      RECT  65000.0 302600.0 65800.0 303400.00000000006 ;
      RECT  69800.0 302600.0 70600.0 303400.00000000006 ;
      RECT  74600.00000000001 302600.0 75400.0 303400.00000000006 ;
      RECT  79400.0 302600.0 80200.0 303400.00000000006 ;
      RECT  84200.0 302600.0 85000.0 303400.00000000006 ;
      RECT  89000.0 302600.0 89800.0 303400.00000000006 ;
      RECT  93800.0 302600.0 94600.0 303400.00000000006 ;
      RECT  98600.00000000001 302600.0 99400.0 303400.00000000006 ;
      RECT  103400.0 302600.0 104200.0 303400.00000000006 ;
      RECT  108200.0 302600.0 109000.0 303400.00000000006 ;
      RECT  113000.00000000001 302600.0 113800.00000000001 303400.00000000006 ;
      RECT  117800.0 302600.0 118600.0 303400.00000000006 ;
      RECT  122600.00000000001 302600.0 123400.0 303400.00000000006 ;
      RECT  127400.0 302600.0 128199.99999999999 303400.00000000006 ;
      RECT  132200.0 302600.0 133000.0 303400.00000000006 ;
      RECT  137000.0 302600.0 137800.0 303400.00000000006 ;
      RECT  141800.0 302600.0 142600.00000000003 303400.00000000006 ;
      RECT  146600.0 302600.0 147400.0 303400.00000000006 ;
      RECT  151399.99999999997 302600.0 152200.0 303400.00000000006 ;
      RECT  156200.0 302600.0 157000.0 303400.00000000006 ;
      RECT  161000.0 302600.0 161800.0 303400.00000000006 ;
      RECT  165800.0 302600.0 166600.00000000003 303400.00000000006 ;
      RECT  170600.0 302600.0 171400.0 303400.00000000006 ;
      RECT  175399.99999999997 302600.0 176200.0 303400.00000000006 ;
      RECT  180200.0 302600.0 181000.0 303400.00000000006 ;
      RECT  185000.0 302600.0 185800.0 303400.00000000006 ;
      RECT  189800.0 302600.0 190600.00000000003 303400.00000000006 ;
      RECT  194600.0 302600.0 195400.0 303400.00000000006 ;
      RECT  199399.99999999997 302600.0 200200.0 303400.00000000006 ;
      RECT  204200.0 302600.0 205000.0 303400.00000000006 ;
      RECT  209000.0 302600.0 209800.0 303400.00000000006 ;
      RECT  7400.000000000003 307400.0 8200.000000000004 308200.0 ;
      RECT  12200.0 307400.0 13000.0 308200.0 ;
      RECT  16999.999999999996 307400.0 17799.999999999996 308200.0 ;
      RECT  21799.999999999993 307400.0 22599.999999999993 308200.0 ;
      RECT  26599.999999999996 307400.0 27400.0 308200.0 ;
      RECT  31399.999999999996 307400.0 32199.999999999996 308200.0 ;
      RECT  36200.0 307400.0 37000.0 308200.0 ;
      RECT  41000.0 307400.0 41800.0 308200.0 ;
      RECT  45800.0 307400.0 46599.99999999999 308200.0 ;
      RECT  50600.0 307400.0 51400.0 308200.0 ;
      RECT  55400.00000000001 307400.0 56200.0 308200.0 ;
      RECT  60200.0 307400.0 61000.0 308200.0 ;
      RECT  65000.0 307400.0 65800.0 308200.0 ;
      RECT  69800.0 307400.0 70600.0 308200.0 ;
      RECT  74600.00000000001 307400.0 75400.0 308200.0 ;
      RECT  79400.0 307400.0 80200.0 308200.0 ;
      RECT  84200.0 307400.0 85000.0 308200.0 ;
      RECT  89000.0 307400.0 89800.0 308200.0 ;
      RECT  93800.0 307400.0 94600.0 308200.0 ;
      RECT  98600.00000000001 307400.0 99400.0 308200.0 ;
      RECT  103400.0 307400.0 104200.0 308200.0 ;
      RECT  108200.0 307400.0 109000.0 308200.0 ;
      RECT  113000.00000000001 307400.0 113800.00000000001 308200.0 ;
      RECT  117800.0 307400.0 118600.0 308200.0 ;
      RECT  122600.00000000001 307400.0 123400.0 308200.0 ;
      RECT  7400.000000000003 312200.0 8200.000000000004 313000.0 ;
      RECT  12200.0 312200.0 13000.0 313000.0 ;
      RECT  16999.999999999996 312200.0 17799.999999999996 313000.0 ;
      RECT  21799.999999999993 312200.0 22599.999999999993 313000.0 ;
      RECT  26599.999999999996 312200.0 27400.0 313000.0 ;
      RECT  31399.999999999996 312200.0 32199.999999999996 313000.0 ;
      RECT  36200.0 312200.0 37000.0 313000.0 ;
      RECT  41000.0 312200.0 41800.0 313000.0 ;
      RECT  45800.0 312200.0 46599.99999999999 313000.0 ;
      RECT  50600.0 312200.0 51400.0 313000.0 ;
      RECT  55400.00000000001 312200.0 56200.0 313000.0 ;
      RECT  60200.0 312200.0 61000.0 313000.0 ;
      RECT  65000.0 312200.0 65800.0 313000.0 ;
      RECT  69800.0 312200.0 70600.0 313000.0 ;
      RECT  74600.00000000001 312200.0 75400.0 313000.0 ;
      RECT  79400.0 312200.0 80200.0 313000.0 ;
      RECT  84200.0 312200.0 85000.0 313000.0 ;
      RECT  89000.0 312200.0 89800.0 313000.0 ;
      RECT  93800.0 312200.0 94600.0 313000.0 ;
      RECT  98600.00000000001 312200.0 99400.0 313000.0 ;
      RECT  103400.0 312200.0 104200.0 313000.0 ;
      RECT  108200.0 312200.0 109000.0 313000.0 ;
      RECT  113000.00000000001 312200.0 113800.00000000001 313000.0 ;
      RECT  117800.0 312200.0 118600.0 313000.0 ;
      RECT  122600.00000000001 312200.0 123400.0 313000.0 ;
      RECT  127400.0 312200.0 128199.99999999999 313000.0 ;
      RECT  132200.0 312200.0 133000.0 313000.0 ;
      RECT  137000.0 312200.0 137800.0 313000.0 ;
      RECT  141800.0 312200.0 142600.00000000003 313000.0 ;
      RECT  146600.0 312200.0 147400.0 313000.0 ;
      RECT  151399.99999999997 312200.0 152200.0 313000.0 ;
      RECT  156200.0 312200.0 157000.0 313000.0 ;
      RECT  161000.0 312200.0 161800.0 313000.0 ;
      RECT  165800.0 312200.0 166600.00000000003 313000.0 ;
      RECT  170600.0 312200.0 171400.0 313000.0 ;
      RECT  175399.99999999997 312200.0 176200.0 313000.0 ;
      RECT  180200.0 312200.0 181000.0 313000.0 ;
      RECT  185000.0 312200.0 185800.0 313000.0 ;
      RECT  189800.0 312200.0 190600.00000000003 313000.0 ;
      RECT  194600.0 312200.0 195400.0 313000.0 ;
      RECT  199399.99999999997 312200.0 200200.0 313000.0 ;
      RECT  204200.0 312200.0 205000.0 313000.0 ;
      RECT  209000.0 312200.0 209800.0 313000.0 ;
      RECT  7400.000000000003 317000.0 8200.000000000004 317800.0 ;
      RECT  12200.0 317000.0 13000.0 317800.0 ;
      RECT  16999.999999999996 317000.0 17799.999999999996 317800.0 ;
      RECT  21799.999999999993 317000.0 22599.999999999993 317800.0 ;
      RECT  26599.999999999996 317000.0 27400.0 317800.0 ;
      RECT  31399.999999999996 317000.0 32199.999999999996 317800.0 ;
      RECT  36200.0 317000.0 37000.0 317800.0 ;
      RECT  41000.0 317000.0 41800.0 317800.0 ;
      RECT  45800.0 317000.0 46599.99999999999 317800.0 ;
      RECT  50600.0 317000.0 51400.0 317800.0 ;
      RECT  69800.0 317000.0 70600.0 317800.0 ;
      RECT  74600.00000000001 317000.0 75400.0 317800.0 ;
      RECT  79400.0 317000.0 80200.0 317800.0 ;
      RECT  84200.0 317000.0 85000.0 317800.0 ;
      RECT  89000.0 317000.0 89800.0 317800.0 ;
      RECT  93800.0 317000.0 94600.0 317800.0 ;
      RECT  98600.00000000001 317000.0 99400.0 317800.0 ;
      RECT  103400.0 317000.0 104200.0 317800.0 ;
      RECT  108200.0 317000.0 109000.0 317800.0 ;
      RECT  113000.00000000001 317000.0 113800.00000000001 317800.0 ;
      RECT  117800.0 317000.0 118600.0 317800.0 ;
      RECT  122600.00000000001 317000.0 123400.0 317800.0 ;
      RECT  127400.0 317000.0 128199.99999999999 317800.0 ;
      RECT  132200.0 317000.0 133000.0 317800.0 ;
      RECT  137000.0 317000.0 137800.0 317800.0 ;
      RECT  141800.0 317000.0 142600.00000000003 317800.0 ;
      RECT  146600.0 317000.0 147400.0 317800.0 ;
      RECT  151399.99999999997 317000.0 152200.0 317800.0 ;
      RECT  156200.0 317000.0 157000.0 317800.0 ;
      RECT  161000.0 317000.0 161800.0 317800.0 ;
      RECT  165800.0 317000.0 166600.00000000003 317800.0 ;
      RECT  170600.0 317000.0 171400.0 317800.0 ;
      RECT  175399.99999999997 317000.0 176200.0 317800.0 ;
      RECT  180200.0 317000.0 181000.0 317800.0 ;
      RECT  185000.0 317000.0 185800.0 317800.0 ;
      RECT  189800.0 317000.0 190600.00000000003 317800.0 ;
      RECT  194600.0 317000.0 195400.0 317800.0 ;
      RECT  199399.99999999997 317000.0 200200.0 317800.0 ;
      RECT  204200.0 317000.0 205000.0 317800.0 ;
      RECT  209000.0 317000.0 209800.0 317800.0 ;
      RECT  7400.000000000003 321800.0 8200.000000000004 322600.0 ;
      RECT  12200.0 321800.0 13000.0 322600.0 ;
      RECT  16999.999999999996 321800.0 17799.999999999996 322600.0 ;
      RECT  21799.999999999993 321800.0 22599.999999999993 322600.0 ;
      RECT  26599.999999999996 321800.0 27400.0 322600.0 ;
      RECT  31399.999999999996 321800.0 32199.999999999996 322600.0 ;
      RECT  36200.0 321800.0 37000.0 322600.0 ;
      RECT  41000.0 321800.0 41800.0 322600.0 ;
      RECT  45800.0 321800.0 46599.99999999999 322600.0 ;
      RECT  50600.0 321800.0 51400.0 322600.0 ;
      RECT  55400.00000000001 321800.0 56200.0 322600.0 ;
      RECT  60200.0 321800.0 61000.0 322600.0 ;
      RECT  65000.0 321800.0 65800.0 322600.0 ;
      RECT  69800.0 321800.0 70600.0 322600.0 ;
      RECT  74600.00000000001 321800.0 75400.0 322600.0 ;
      RECT  79400.0 321800.0 80200.0 322600.0 ;
      RECT  84200.0 321800.0 85000.0 322600.0 ;
      RECT  89000.0 321800.0 89800.0 322600.0 ;
      RECT  93800.0 321800.0 94600.0 322600.0 ;
      RECT  98600.00000000001 321800.0 99400.0 322600.0 ;
      RECT  103400.0 321800.0 104200.0 322600.0 ;
      RECT  108200.0 321800.0 109000.0 322600.0 ;
      RECT  113000.00000000001 321800.0 113800.00000000001 322600.0 ;
      RECT  117800.0 321800.0 118600.0 322600.0 ;
      RECT  122600.00000000001 321800.0 123400.0 322600.0 ;
      RECT  127400.0 321800.0 128199.99999999999 322600.0 ;
      RECT  132200.0 321800.0 133000.0 322600.0 ;
      RECT  137000.0 321800.0 137800.0 322600.0 ;
      RECT  141800.0 321800.0 142600.00000000003 322600.0 ;
      RECT  146600.0 321800.0 147400.0 322600.0 ;
      RECT  151399.99999999997 321800.0 152200.0 322600.0 ;
      RECT  156200.0 321800.0 157000.0 322600.0 ;
      RECT  161000.0 321800.0 161800.0 322600.0 ;
      RECT  165800.0 321800.0 166600.00000000003 322600.0 ;
      RECT  170600.0 321800.0 171400.0 322600.0 ;
      RECT  175399.99999999997 321800.0 176200.0 322600.0 ;
      RECT  180200.0 321800.0 181000.0 322600.0 ;
      RECT  185000.0 321800.0 185800.0 322600.0 ;
      RECT  189800.0 321800.0 190600.00000000003 322600.0 ;
      RECT  194600.0 321800.0 195400.0 322600.0 ;
      RECT  199399.99999999997 321800.0 200200.0 322600.0 ;
      RECT  204200.0 321800.0 205000.0 322600.0 ;
      RECT  209000.0 321800.0 209800.0 322600.0 ;
      RECT  7400.000000000003 326599.99999999994 8200.000000000004 327400.0 ;
      RECT  12200.0 326599.99999999994 13000.0 327400.0 ;
      RECT  16999.999999999996 326599.99999999994 17799.999999999996 327400.0 ;
      RECT  21799.999999999993 326599.99999999994 22599.999999999993 327400.0 ;
      RECT  26599.999999999996 326599.99999999994 27400.0 327400.0 ;
      RECT  31399.999999999996 326599.99999999994 32199.999999999996 327400.0 ;
      RECT  36200.0 326599.99999999994 37000.0 327400.0 ;
      RECT  41000.0 326599.99999999994 41800.0 327400.0 ;
      RECT  45800.0 326599.99999999994 46599.99999999999 327400.0 ;
      RECT  50600.0 326599.99999999994 51400.0 327400.0 ;
      RECT  55400.00000000001 326599.99999999994 56200.0 327400.0 ;
      RECT  60200.0 326599.99999999994 61000.0 327400.0 ;
      RECT  89000.0 326599.99999999994 89800.0 327400.0 ;
      RECT  93800.0 326599.99999999994 94600.0 327400.0 ;
      RECT  98600.00000000001 326599.99999999994 99400.0 327400.0 ;
      RECT  103400.0 326599.99999999994 104200.0 327400.0 ;
      RECT  108200.0 326599.99999999994 109000.0 327400.0 ;
      RECT  113000.00000000001 326599.99999999994 113800.00000000001 327400.0 ;
      RECT  117800.0 326599.99999999994 118600.0 327400.0 ;
      RECT  122600.00000000001 326599.99999999994 123400.0 327400.0 ;
      RECT  127400.0 326599.99999999994 128199.99999999999 327400.0 ;
      RECT  132200.0 326599.99999999994 133000.0 327400.0 ;
      RECT  137000.0 326599.99999999994 137800.0 327400.0 ;
      RECT  141800.0 326599.99999999994 142600.00000000003 327400.0 ;
      RECT  146600.0 326599.99999999994 147400.0 327400.0 ;
      RECT  151399.99999999997 326599.99999999994 152200.0 327400.0 ;
      RECT  156200.0 326599.99999999994 157000.0 327400.0 ;
      RECT  161000.0 326599.99999999994 161800.0 327400.0 ;
      RECT  165800.0 326599.99999999994 166600.00000000003 327400.0 ;
      RECT  170600.0 326599.99999999994 171400.0 327400.0 ;
      RECT  175399.99999999997 326599.99999999994 176200.0 327400.0 ;
      RECT  180200.0 326599.99999999994 181000.0 327400.0 ;
      RECT  185000.0 326599.99999999994 185800.0 327400.0 ;
      RECT  189800.0 326599.99999999994 190600.00000000003 327400.0 ;
      RECT  194600.0 326599.99999999994 195400.0 327400.0 ;
      RECT  199399.99999999997 326599.99999999994 200200.0 327400.0 ;
      RECT  204200.0 326599.99999999994 205000.0 327400.0 ;
      RECT  209000.0 326599.99999999994 209800.0 327400.0 ;
      RECT  7400.000000000003 331400.0 8200.000000000004 332200.0 ;
      RECT  12200.0 331400.0 13000.0 332200.0 ;
      RECT  16999.999999999996 331400.0 17799.999999999996 332200.0 ;
      RECT  21799.999999999993 331400.0 22599.999999999993 332200.0 ;
      RECT  26599.999999999996 331400.0 27400.0 332200.0 ;
      RECT  31399.999999999996 331400.0 32199.999999999996 332200.0 ;
      RECT  36200.0 331400.0 37000.0 332200.0 ;
      RECT  41000.0 331400.0 41800.0 332200.0 ;
      RECT  45800.0 331400.0 46599.99999999999 332200.0 ;
      RECT  50600.0 331400.0 51400.0 332200.0 ;
      RECT  55400.00000000001 331400.0 56200.0 332200.0 ;
      RECT  60200.0 331400.0 61000.0 332200.0 ;
      RECT  65000.0 331400.0 65800.0 332200.0 ;
      RECT  69800.0 331400.0 70600.0 332200.0 ;
      RECT  74600.00000000001 331400.0 75400.0 332200.0 ;
      RECT  79400.0 331400.0 80200.0 332200.0 ;
      RECT  84200.0 331400.0 85000.0 332200.0 ;
      RECT  89000.0 331400.0 89800.0 332200.0 ;
      RECT  93800.0 331400.0 94600.0 332200.0 ;
      RECT  98600.00000000001 331400.0 99400.0 332200.0 ;
      RECT  103400.0 331400.0 104200.0 332200.0 ;
      RECT  108200.0 331400.0 109000.0 332200.0 ;
      RECT  113000.00000000001 331400.0 113800.00000000001 332200.0 ;
      RECT  117800.0 331400.0 118600.0 332200.0 ;
      RECT  122600.00000000001 331400.0 123400.0 332200.0 ;
      RECT  127400.0 331400.0 128199.99999999999 332200.0 ;
      RECT  132200.0 331400.0 133000.0 332200.0 ;
      RECT  137000.0 331400.0 137800.0 332200.0 ;
      RECT  141800.0 331400.0 142600.00000000003 332200.0 ;
      RECT  146600.0 331400.0 147400.0 332200.0 ;
      RECT  151399.99999999997 331400.0 152200.0 332200.0 ;
      RECT  156200.0 331400.0 157000.0 332200.0 ;
      RECT  161000.0 331400.0 161800.0 332200.0 ;
      RECT  165800.0 331400.0 166600.00000000003 332200.0 ;
      RECT  170600.0 331400.0 171400.0 332200.0 ;
      RECT  175399.99999999997 331400.0 176200.0 332200.0 ;
      RECT  180200.0 331400.0 181000.0 332200.0 ;
      RECT  185000.0 331400.0 185800.0 332200.0 ;
      RECT  189800.0 331400.0 190600.00000000003 332200.0 ;
      RECT  194600.0 331400.0 195400.0 332200.0 ;
      RECT  199399.99999999997 331400.0 200200.0 332200.0 ;
      RECT  204200.0 331400.0 205000.0 332200.0 ;
      RECT  209000.0 331400.0 209800.0 332200.0 ;
      RECT  9799.999999999993 2600.000000000006 10599.999999999995 3400.0000000000055 ;
      RECT  14599.999999999998 2600.000000000006 15399.999999999998 3400.0000000000055 ;
      RECT  19399.999999999996 2600.000000000006 20199.999999999996 3400.0000000000055 ;
      RECT  24200.0 2600.000000000006 25000.0 3400.0000000000055 ;
      RECT  28999.999999999996 2600.000000000006 29799.999999999996 3400.0000000000055 ;
      RECT  33800.0 2600.000000000006 34599.99999999999 3400.0000000000055 ;
      RECT  38600.0 2600.000000000006 39400.0 3400.0000000000055 ;
      RECT  43400.00000000001 2600.000000000006 44200.0 3400.0000000000055 ;
      RECT  48200.0 2600.000000000006 49000.0 3400.0000000000055 ;
      RECT  53000.0 2600.000000000006 53800.0 3400.0000000000055 ;
      RECT  57800.0 2600.000000000006 58599.99999999999 3400.0000000000055 ;
      RECT  62600.0 2600.000000000006 63400.0 3400.0000000000055 ;
      RECT  77000.0 2600.000000000006 77800.0 3400.0000000000055 ;
      RECT  81800.0 2600.000000000006 82600.0 3400.0000000000055 ;
      RECT  86600.00000000001 2600.000000000006 87400.0 3400.0000000000055 ;
      RECT  91400.0 2600.000000000006 92200.0 3400.0000000000055 ;
      RECT  96200.0 2600.000000000006 97000.0 3400.0000000000055 ;
      RECT  101000.0 2600.000000000006 101800.0 3400.0000000000055 ;
      RECT  105800.0 2600.000000000006 106600.0 3400.0000000000055 ;
      RECT  110600.00000000001 2600.000000000006 111400.0 3400.0000000000055 ;
      RECT  115400.0 2600.000000000006 116200.0 3400.0000000000055 ;
      RECT  120200.0 2600.000000000006 121000.0 3400.0000000000055 ;
      RECT  125000.00000000001 2600.000000000006 125800.00000000001 3400.0000000000055 ;
      RECT  129799.99999999999 2600.000000000006 130600.0 3400.0000000000055 ;
      RECT  134600.0 2600.000000000006 135400.0 3400.0000000000055 ;
      RECT  139399.99999999997 2600.000000000006 140200.0 3400.0000000000055 ;
      RECT  144200.0 2600.000000000006 145000.0 3400.0000000000055 ;
      RECT  149000.0 2600.000000000006 149800.0 3400.0000000000055 ;
      RECT  153800.0 2600.000000000006 154600.00000000003 3400.0000000000055 ;
      RECT  158600.0 2600.000000000006 159400.0 3400.0000000000055 ;
      RECT  163399.99999999997 2600.000000000006 164200.0 3400.0000000000055 ;
      RECT  168200.0 2600.000000000006 169000.0 3400.0000000000055 ;
      RECT  173000.0 2600.000000000006 173800.0 3400.0000000000055 ;
      RECT  177800.0 2600.000000000006 178600.00000000003 3400.0000000000055 ;
      RECT  182600.0 2600.000000000006 183400.0 3400.0000000000055 ;
      RECT  187399.99999999997 2600.000000000006 188200.0 3400.0000000000055 ;
      RECT  192200.0 2600.000000000006 193000.0 3400.0000000000055 ;
      RECT  197000.0 2600.000000000006 197800.0 3400.0000000000055 ;
      RECT  201800.0 2600.000000000006 202600.00000000003 3400.0000000000055 ;
      RECT  206600.0 2600.000000000006 207400.0 3400.0000000000055 ;
      RECT  4999.999999999997 7400.000000000003 5799.999999999997 8200.000000000004 ;
      RECT  9799.999999999993 7400.000000000003 10599.999999999995 8200.000000000004 ;
      RECT  14599.999999999998 7400.000000000003 15399.999999999998 8200.000000000004 ;
      RECT  19399.999999999996 7400.000000000003 20199.999999999996 8200.000000000004 ;
      RECT  24200.0 7400.000000000003 25000.0 8200.000000000004 ;
      RECT  28999.999999999996 7400.000000000003 29799.999999999996 8200.000000000004 ;
      RECT  33800.0 7400.000000000003 34599.99999999999 8200.000000000004 ;
      RECT  38600.0 7400.000000000003 39400.0 8200.000000000004 ;
      RECT  43400.00000000001 7400.000000000003 44200.0 8200.000000000004 ;
      RECT  48200.0 7400.000000000003 49000.0 8200.000000000004 ;
      RECT  53000.0 7400.000000000003 53800.0 8200.000000000004 ;
      RECT  57800.0 7400.000000000003 58599.99999999999 8200.000000000004 ;
      RECT  62600.0 7400.000000000003 63400.0 8200.000000000004 ;
      RECT  67400.0 7400.000000000003 68200.0 8200.000000000004 ;
      RECT  72200.0 7400.000000000003 73000.0 8200.000000000004 ;
      RECT  77000.0 7400.000000000003 77800.0 8200.000000000004 ;
      RECT  81800.0 7400.000000000003 82600.0 8200.000000000004 ;
      RECT  86600.00000000001 7400.000000000003 87400.0 8200.000000000004 ;
      RECT  91400.0 7400.000000000003 92200.0 8200.000000000004 ;
      RECT  96200.0 7400.000000000003 97000.0 8200.000000000004 ;
      RECT  101000.0 7400.000000000003 101800.0 8200.000000000004 ;
      RECT  105800.0 7400.000000000003 106600.0 8200.000000000004 ;
      RECT  110600.00000000001 7400.000000000003 111400.0 8200.000000000004 ;
      RECT  115400.0 7400.000000000003 116200.0 8200.000000000004 ;
      RECT  120200.0 7400.000000000003 121000.0 8200.000000000004 ;
      RECT  125000.00000000001 7400.000000000003 125800.00000000001 8200.000000000004 ;
      RECT  129799.99999999999 7400.000000000003 130600.0 8200.000000000004 ;
      RECT  134600.0 7400.000000000003 135400.0 8200.000000000004 ;
      RECT  139399.99999999997 7400.000000000003 140200.0 8200.000000000004 ;
      RECT  144200.0 7400.000000000003 145000.0 8200.000000000004 ;
      RECT  149000.0 7400.000000000003 149800.0 8200.000000000004 ;
      RECT  153800.0 7400.000000000003 154600.00000000003 8200.000000000004 ;
      RECT  158600.0 7400.000000000003 159400.0 8200.000000000004 ;
      RECT  163399.99999999997 7400.000000000003 164200.0 8200.000000000004 ;
      RECT  168200.0 7400.000000000003 169000.0 8200.000000000004 ;
      RECT  173000.0 7400.000000000003 173800.0 8200.000000000004 ;
      RECT  177800.0 7400.000000000003 178600.00000000003 8200.000000000004 ;
      RECT  182600.0 7400.000000000003 183400.0 8200.000000000004 ;
      RECT  187399.99999999997 7400.000000000003 188200.0 8200.000000000004 ;
      RECT  192200.0 7400.000000000003 193000.0 8200.000000000004 ;
      RECT  197000.0 7400.000000000003 197800.0 8200.000000000004 ;
      RECT  201800.0 7400.000000000003 202600.00000000003 8200.000000000004 ;
      RECT  206600.0 7400.000000000003 207400.0 8200.000000000004 ;
      RECT  53000.0 12200.0 53800.0 13000.0 ;
      RECT  57800.0 12200.0 58599.99999999999 13000.0 ;
      RECT  62600.0 12200.0 63400.0 13000.0 ;
      RECT  67400.0 12200.0 68200.0 13000.0 ;
      RECT  72200.0 12200.0 73000.0 13000.0 ;
      RECT  77000.0 12200.0 77800.0 13000.0 ;
      RECT  81800.0 12200.0 82600.0 13000.0 ;
      RECT  86600.00000000001 12200.0 87400.0 13000.0 ;
      RECT  91400.0 12200.0 92200.0 13000.0 ;
      RECT  96200.0 12200.0 97000.0 13000.0 ;
      RECT  101000.0 12200.0 101800.0 13000.0 ;
      RECT  105800.0 12200.0 106600.0 13000.0 ;
      RECT  110600.00000000001 12200.0 111400.0 13000.0 ;
      RECT  115400.0 12200.0 116200.0 13000.0 ;
      RECT  120200.0 12200.0 121000.0 13000.0 ;
      RECT  125000.00000000001 12200.0 125800.00000000001 13000.0 ;
      RECT  129799.99999999999 12200.0 130600.0 13000.0 ;
      RECT  134600.0 12200.0 135400.0 13000.0 ;
      RECT  139399.99999999997 12200.0 140200.0 13000.0 ;
      RECT  144200.0 12200.0 145000.0 13000.0 ;
      RECT  149000.0 12200.0 149800.0 13000.0 ;
      RECT  153800.0 12200.0 154600.00000000003 13000.0 ;
      RECT  158600.0 12200.0 159400.0 13000.0 ;
      RECT  163399.99999999997 12200.0 164200.0 13000.0 ;
      RECT  168200.0 12200.0 169000.0 13000.0 ;
      RECT  173000.0 12200.0 173800.0 13000.0 ;
      RECT  177800.0 12200.0 178600.00000000003 13000.0 ;
      RECT  182600.0 12200.0 183400.0 13000.0 ;
      RECT  187399.99999999997 12200.0 188200.0 13000.0 ;
      RECT  192200.0 12200.0 193000.0 13000.0 ;
      RECT  197000.0 12200.0 197800.0 13000.0 ;
      RECT  201800.0 12200.0 202600.00000000003 13000.0 ;
      RECT  206600.0 12200.0 207400.0 13000.0 ;
      RECT  4999.999999999997 16999.999999999996 5799.999999999997 17799.999999999996 ;
      RECT  9799.999999999993 16999.999999999996 10599.999999999995 17799.999999999996 ;
      RECT  14599.999999999998 16999.999999999996 15399.999999999998 17799.999999999996 ;
      RECT  19399.999999999996 16999.999999999996 20199.999999999996 17799.999999999996 ;
      RECT  24200.0 16999.999999999996 25000.0 17799.999999999996 ;
      RECT  28999.999999999996 16999.999999999996 29799.999999999996 17799.999999999996 ;
      RECT  33800.0 16999.999999999996 34599.99999999999 17799.999999999996 ;
      RECT  38600.0 16999.999999999996 39400.0 17799.999999999996 ;
      RECT  43400.00000000001 16999.999999999996 44200.0 17799.999999999996 ;
      RECT  48200.0 16999.999999999996 49000.0 17799.999999999996 ;
      RECT  53000.0 16999.999999999996 53800.0 17799.999999999996 ;
      RECT  57800.0 16999.999999999996 58599.99999999999 17799.999999999996 ;
      RECT  62600.0 16999.999999999996 63400.0 17799.999999999996 ;
      RECT  67400.0 16999.999999999996 68200.0 17799.999999999996 ;
      RECT  72200.0 16999.999999999996 73000.0 17799.999999999996 ;
      RECT  77000.0 16999.999999999996 77800.0 17799.999999999996 ;
      RECT  81800.0 16999.999999999996 82600.0 17799.999999999996 ;
      RECT  86600.00000000001 16999.999999999996 87400.0 17799.999999999996 ;
      RECT  91400.0 16999.999999999996 92200.0 17799.999999999996 ;
      RECT  96200.0 16999.999999999996 97000.0 17799.999999999996 ;
      RECT  101000.0 16999.999999999996 101800.0 17799.999999999996 ;
      RECT  105800.0 16999.999999999996 106600.0 17799.999999999996 ;
      RECT  110600.00000000001 16999.999999999996 111400.0 17799.999999999996 ;
      RECT  115400.0 16999.999999999996 116200.0 17799.999999999996 ;
      RECT  120200.0 16999.999999999996 121000.0 17799.999999999996 ;
      RECT  125000.00000000001 16999.999999999996 125800.00000000001 17799.999999999996 ;
      RECT  129799.99999999999 16999.999999999996 130600.0 17799.999999999996 ;
      RECT  134600.0 16999.999999999996 135400.0 17799.999999999996 ;
      RECT  139399.99999999997 16999.999999999996 140200.0 17799.999999999996 ;
      RECT  144200.0 16999.999999999996 145000.0 17799.999999999996 ;
      RECT  149000.0 16999.999999999996 149800.0 17799.999999999996 ;
      RECT  153800.0 16999.999999999996 154600.00000000003 17799.999999999996 ;
      RECT  158600.0 16999.999999999996 159400.0 17799.999999999996 ;
      RECT  163399.99999999997 16999.999999999996 164200.0 17799.999999999996 ;
      RECT  168200.0 16999.999999999996 169000.0 17799.999999999996 ;
      RECT  173000.0 16999.999999999996 173800.0 17799.999999999996 ;
      RECT  177800.0 16999.999999999996 178600.00000000003 17799.999999999996 ;
      RECT  182600.0 16999.999999999996 183400.0 17799.999999999996 ;
      RECT  187399.99999999997 16999.999999999996 188200.0 17799.999999999996 ;
      RECT  192200.0 16999.999999999996 193000.0 17799.999999999996 ;
      RECT  197000.0 16999.999999999996 197800.0 17799.999999999996 ;
      RECT  201800.0 16999.999999999996 202600.00000000003 17799.999999999996 ;
      RECT  206600.0 16999.999999999996 207400.0 17799.999999999996 ;
      RECT  4999.999999999997 21800.0 5799.999999999997 22600.0 ;
      RECT  9799.999999999993 21800.0 10599.999999999995 22600.0 ;
      RECT  14599.999999999998 21800.0 15399.999999999998 22600.0 ;
      RECT  19399.999999999996 21800.0 20199.999999999996 22600.0 ;
      RECT  24200.0 21800.0 25000.0 22600.0 ;
      RECT  28999.999999999996 21800.0 29799.999999999996 22600.0 ;
      RECT  33800.0 21800.0 34599.99999999999 22600.0 ;
      RECT  38600.0 21800.0 39400.0 22600.0 ;
      RECT  43400.00000000001 21800.0 44200.0 22600.0 ;
      RECT  48200.0 21800.0 49000.0 22600.0 ;
      RECT  53000.0 21800.0 53800.0 22600.0 ;
      RECT  57800.0 21800.0 58599.99999999999 22600.0 ;
      RECT  62600.0 21800.0 63400.0 22600.0 ;
      RECT  67400.0 21800.0 68200.0 22600.0 ;
      RECT  72200.0 21800.0 73000.0 22600.0 ;
      RECT  77000.0 21800.0 77800.0 22600.0 ;
      RECT  81800.0 21800.0 82600.0 22600.0 ;
      RECT  86600.00000000001 21800.0 87400.0 22600.0 ;
      RECT  91400.0 21800.0 92200.0 22600.0 ;
      RECT  96200.0 21800.0 97000.0 22600.0 ;
      RECT  101000.0 21800.0 101800.0 22600.0 ;
      RECT  105800.0 21800.0 106600.0 22600.0 ;
      RECT  110600.00000000001 21800.0 111400.0 22600.0 ;
      RECT  115400.0 21800.0 116200.0 22600.0 ;
      RECT  120200.0 21800.0 121000.0 22600.0 ;
      RECT  125000.00000000001 21800.0 125800.00000000001 22600.0 ;
      RECT  129799.99999999999 21800.0 130600.0 22600.0 ;
      RECT  134600.0 21800.0 135400.0 22600.0 ;
      RECT  139399.99999999997 21800.0 140200.0 22600.0 ;
      RECT  144200.0 21800.0 145000.0 22600.0 ;
      RECT  149000.0 21800.0 149800.0 22600.0 ;
      RECT  153800.0 21800.0 154600.00000000003 22600.0 ;
      RECT  158600.0 21800.0 159400.0 22600.0 ;
      RECT  163399.99999999997 21800.0 164200.0 22600.0 ;
      RECT  168200.0 21800.0 169000.0 22600.0 ;
      RECT  173000.0 21800.0 173800.0 22600.0 ;
      RECT  177800.0 21800.0 178600.00000000003 22600.0 ;
      RECT  182600.0 21800.0 183400.0 22600.0 ;
      RECT  187399.99999999997 21800.0 188200.0 22600.0 ;
      RECT  192200.0 21800.0 193000.0 22600.0 ;
      RECT  197000.0 21800.0 197800.0 22600.0 ;
      RECT  201800.0 21800.0 202600.00000000003 22600.0 ;
      RECT  206600.0 21800.0 207400.0 22600.0 ;
      RECT  4999.999999999997 26599.999999999996 5799.999999999997 27400.0 ;
      RECT  9799.999999999993 26599.999999999996 10599.999999999995 27400.0 ;
      RECT  14599.999999999998 26599.999999999996 15399.999999999998 27400.0 ;
      RECT  19399.999999999996 26599.999999999996 20199.999999999996 27400.0 ;
      RECT  24200.0 26599.999999999996 25000.0 27400.0 ;
      RECT  28999.999999999996 26599.999999999996 29799.999999999996 27400.0 ;
      RECT  33800.0 26599.999999999996 34599.99999999999 27400.0 ;
      RECT  38600.0 26599.999999999996 39400.0 27400.0 ;
      RECT  43400.00000000001 26599.999999999996 44200.0 27400.0 ;
      RECT  48200.0 26599.999999999996 49000.0 27400.0 ;
      RECT  53000.0 26599.999999999996 53800.0 27400.0 ;
      RECT  57800.0 26599.999999999996 58599.99999999999 27400.0 ;
      RECT  62600.0 26599.999999999996 63400.0 27400.0 ;
      RECT  67400.0 26599.999999999996 68200.0 27400.0 ;
      RECT  72200.0 26599.999999999996 73000.0 27400.0 ;
      RECT  77000.0 26599.999999999996 77800.0 27400.0 ;
      RECT  81800.0 26599.999999999996 82600.0 27400.0 ;
      RECT  86600.00000000001 26599.999999999996 87400.0 27400.0 ;
      RECT  91400.0 26599.999999999996 92200.0 27400.0 ;
      RECT  96200.0 26599.999999999996 97000.0 27400.0 ;
      RECT  101000.0 26599.999999999996 101800.0 27400.0 ;
      RECT  105800.0 26599.999999999996 106600.0 27400.0 ;
      RECT  110600.00000000001 26599.999999999996 111400.0 27400.0 ;
      RECT  115400.0 26599.999999999996 116200.0 27400.0 ;
      RECT  120200.0 26599.999999999996 121000.0 27400.0 ;
      RECT  125000.00000000001 26599.999999999996 125800.00000000001 27400.0 ;
      RECT  129799.99999999999 26599.999999999996 130600.0 27400.0 ;
      RECT  134600.0 26599.999999999996 135400.0 27400.0 ;
      RECT  139399.99999999997 26599.999999999996 140200.0 27400.0 ;
      RECT  144200.0 26599.999999999996 145000.0 27400.0 ;
      RECT  149000.0 26599.999999999996 149800.0 27400.0 ;
      RECT  153800.0 26599.999999999996 154600.00000000003 27400.0 ;
      RECT  158600.0 26599.999999999996 159400.0 27400.0 ;
      RECT  163399.99999999997 26599.999999999996 164200.0 27400.0 ;
      RECT  168200.0 26599.999999999996 169000.0 27400.0 ;
      RECT  173000.0 26599.999999999996 173800.0 27400.0 ;
      RECT  177800.0 26599.999999999996 178600.00000000003 27400.0 ;
      RECT  182600.0 26599.999999999996 183400.0 27400.0 ;
      RECT  187399.99999999997 26599.999999999996 188200.0 27400.0 ;
      RECT  192200.0 26599.999999999996 193000.0 27400.0 ;
      RECT  197000.0 26599.999999999996 197800.0 27400.0 ;
      RECT  201800.0 26599.999999999996 202600.00000000003 27400.0 ;
      RECT  206600.0 26599.999999999996 207400.0 27400.0 ;
      RECT  72200.0 31400.000000000004 73000.0 32200.000000000004 ;
      RECT  77000.0 31400.000000000004 77800.0 32200.000000000004 ;
      RECT  81800.0 31400.000000000004 82600.0 32200.000000000004 ;
      RECT  86600.00000000001 31400.000000000004 87400.0 32200.000000000004 ;
      RECT  91400.0 31400.000000000004 92200.0 32200.000000000004 ;
      RECT  96200.0 31400.000000000004 97000.0 32200.000000000004 ;
      RECT  101000.0 31400.000000000004 101800.0 32200.000000000004 ;
      RECT  105800.0 31400.000000000004 106600.0 32200.000000000004 ;
      RECT  110600.00000000001 31400.000000000004 111400.0 32200.000000000004 ;
      RECT  115400.0 31400.000000000004 116200.0 32200.000000000004 ;
      RECT  120200.0 31400.000000000004 121000.0 32200.000000000004 ;
      RECT  125000.00000000001 31400.000000000004 125800.00000000001 32200.000000000004 ;
      RECT  129799.99999999999 31400.000000000004 130600.0 32200.000000000004 ;
      RECT  134600.0 31400.000000000004 135400.0 32200.000000000004 ;
      RECT  139399.99999999997 31400.000000000004 140200.0 32200.000000000004 ;
      RECT  144200.0 31400.000000000004 145000.0 32200.000000000004 ;
      RECT  149000.0 31400.000000000004 149800.0 32200.000000000004 ;
      RECT  153800.0 31400.000000000004 154600.00000000003 32200.000000000004 ;
      RECT  158600.0 31400.000000000004 159400.0 32200.000000000004 ;
      RECT  163399.99999999997 31400.000000000004 164200.0 32200.000000000004 ;
      RECT  168200.0 31400.000000000004 169000.0 32200.000000000004 ;
      RECT  173000.0 31400.000000000004 173800.0 32200.000000000004 ;
      RECT  177800.0 31400.000000000004 178600.00000000003 32200.000000000004 ;
      RECT  182600.0 31400.000000000004 183400.0 32200.000000000004 ;
      RECT  187399.99999999997 31400.000000000004 188200.0 32200.000000000004 ;
      RECT  192200.0 31400.000000000004 193000.0 32200.000000000004 ;
      RECT  197000.0 31400.000000000004 197800.0 32200.000000000004 ;
      RECT  201800.0 31400.000000000004 202600.00000000003 32200.000000000004 ;
      RECT  206600.0 31400.000000000004 207400.0 32200.000000000004 ;
      RECT  4999.999999999997 36200.0 5799.999999999997 37000.0 ;
      RECT  9799.999999999993 36200.0 10599.999999999995 37000.0 ;
      RECT  14599.999999999998 36200.0 15399.999999999998 37000.0 ;
      RECT  19399.999999999996 36200.0 20199.999999999996 37000.0 ;
      RECT  24200.0 36200.0 25000.0 37000.0 ;
      RECT  28999.999999999996 36200.0 29799.999999999996 37000.0 ;
      RECT  33800.0 36200.0 34599.99999999999 37000.0 ;
      RECT  62600.0 36200.0 63400.0 37000.0 ;
      RECT  67400.0 36200.0 68200.0 37000.0 ;
      RECT  72200.0 36200.0 73000.0 37000.0 ;
      RECT  77000.0 36200.0 77800.0 37000.0 ;
      RECT  81800.0 36200.0 82600.0 37000.0 ;
      RECT  86600.00000000001 36200.0 87400.0 37000.0 ;
      RECT  91400.0 36200.0 92200.0 37000.0 ;
      RECT  96200.0 36200.0 97000.0 37000.0 ;
      RECT  101000.0 36200.0 101800.0 37000.0 ;
      RECT  105800.0 36200.0 106600.0 37000.0 ;
      RECT  110600.00000000001 36200.0 111400.0 37000.0 ;
      RECT  115400.0 36200.0 116200.0 37000.0 ;
      RECT  120200.0 36200.0 121000.0 37000.0 ;
      RECT  125000.00000000001 36200.0 125800.00000000001 37000.0 ;
      RECT  129799.99999999999 36200.0 130600.0 37000.0 ;
      RECT  134600.0 36200.0 135400.0 37000.0 ;
      RECT  139399.99999999997 36200.0 140200.0 37000.0 ;
      RECT  144200.0 36200.0 145000.0 37000.0 ;
      RECT  149000.0 36200.0 149800.0 37000.0 ;
      RECT  153800.0 36200.0 154600.00000000003 37000.0 ;
      RECT  158600.0 36200.0 159400.0 37000.0 ;
      RECT  163399.99999999997 36200.0 164200.0 37000.0 ;
      RECT  168200.0 36200.0 169000.0 37000.0 ;
      RECT  173000.0 36200.0 173800.0 37000.0 ;
      RECT  177800.0 36200.0 178600.00000000003 37000.0 ;
      RECT  182600.0 36200.0 183400.0 37000.0 ;
      RECT  187399.99999999997 36200.0 188200.0 37000.0 ;
      RECT  192200.0 36200.0 193000.0 37000.0 ;
      RECT  197000.0 36200.0 197800.0 37000.0 ;
      RECT  201800.0 36200.0 202600.00000000003 37000.0 ;
      RECT  206600.0 36200.0 207400.0 37000.0 ;
      RECT  9799.999999999993 41000.0 10599.999999999995 41800.0 ;
      RECT  14599.999999999998 41000.0 15399.999999999998 41800.0 ;
      RECT  19399.999999999996 41000.0 20199.999999999996 41800.0 ;
      RECT  24200.0 41000.0 25000.0 41800.0 ;
      RECT  28999.999999999996 41000.0 29799.999999999996 41800.0 ;
      RECT  33800.0 41000.0 34599.99999999999 41800.0 ;
      RECT  38600.0 41000.0 39400.0 41800.0 ;
      RECT  43400.00000000001 41000.0 44200.0 41800.0 ;
      RECT  48200.0 41000.0 49000.0 41800.0 ;
      RECT  53000.0 41000.0 53800.0 41800.0 ;
      RECT  57800.0 41000.0 58599.99999999999 41800.0 ;
      RECT  62600.0 41000.0 63400.0 41800.0 ;
      RECT  77000.0 41000.0 77800.0 41800.0 ;
      RECT  81800.0 41000.0 82600.0 41800.0 ;
      RECT  86600.00000000001 41000.0 87400.0 41800.0 ;
      RECT  91400.0 41000.0 92200.0 41800.0 ;
      RECT  96200.0 41000.0 97000.0 41800.0 ;
      RECT  101000.0 41000.0 101800.0 41800.0 ;
      RECT  105800.0 41000.0 106600.0 41800.0 ;
      RECT  110600.00000000001 41000.0 111400.0 41800.0 ;
      RECT  115400.0 41000.0 116200.0 41800.0 ;
      RECT  120200.0 41000.0 121000.0 41800.0 ;
      RECT  125000.00000000001 41000.0 125800.00000000001 41800.0 ;
      RECT  129799.99999999999 41000.0 130600.0 41800.0 ;
      RECT  134600.0 41000.0 135400.0 41800.0 ;
      RECT  139399.99999999997 41000.0 140200.0 41800.0 ;
      RECT  144200.0 41000.0 145000.0 41800.0 ;
      RECT  149000.0 41000.0 149800.0 41800.0 ;
      RECT  153800.0 41000.0 154600.00000000003 41800.0 ;
      RECT  158600.0 41000.0 159400.0 41800.0 ;
      RECT  163399.99999999997 41000.0 164200.0 41800.0 ;
      RECT  168200.0 41000.0 169000.0 41800.0 ;
      RECT  173000.0 41000.0 173800.0 41800.0 ;
      RECT  4999.999999999997 45800.00000000001 5799.999999999997 46600.0 ;
      RECT  9799.999999999993 45800.00000000001 10599.999999999995 46600.0 ;
      RECT  14599.999999999998 45800.00000000001 15399.999999999998 46600.0 ;
      RECT  19399.999999999996 45800.00000000001 20199.999999999996 46600.0 ;
      RECT  24200.0 45800.00000000001 25000.0 46600.0 ;
      RECT  28999.999999999996 45800.00000000001 29799.999999999996 46600.0 ;
      RECT  33800.0 45800.00000000001 34599.99999999999 46600.0 ;
      RECT  38600.0 45800.00000000001 39400.0 46600.0 ;
      RECT  43400.00000000001 45800.00000000001 44200.0 46600.0 ;
      RECT  48200.0 45800.00000000001 49000.0 46600.0 ;
      RECT  53000.0 45800.00000000001 53800.0 46600.0 ;
      RECT  57800.0 45800.00000000001 58599.99999999999 46600.0 ;
      RECT  62600.0 45800.00000000001 63400.0 46600.0 ;
      RECT  67400.0 45800.00000000001 68200.0 46600.0 ;
      RECT  72200.0 45800.00000000001 73000.0 46600.0 ;
      RECT  77000.0 45800.00000000001 77800.0 46600.0 ;
      RECT  81800.0 45800.00000000001 82600.0 46600.0 ;
      RECT  86600.00000000001 45800.00000000001 87400.0 46600.0 ;
      RECT  91400.0 45800.00000000001 92200.0 46600.0 ;
      RECT  96200.0 45800.00000000001 97000.0 46600.0 ;
      RECT  101000.0 45800.00000000001 101800.0 46600.0 ;
      RECT  105800.0 45800.00000000001 106600.0 46600.0 ;
      RECT  110600.00000000001 45800.00000000001 111400.0 46600.0 ;
      RECT  115400.0 45800.00000000001 116200.0 46600.0 ;
      RECT  120200.0 45800.00000000001 121000.0 46600.0 ;
      RECT  125000.00000000001 45800.00000000001 125800.00000000001 46600.0 ;
      RECT  129799.99999999999 45800.00000000001 130600.0 46600.0 ;
      RECT  134600.0 45800.00000000001 135400.0 46600.0 ;
      RECT  139399.99999999997 45800.00000000001 140200.0 46600.0 ;
      RECT  144200.0 45800.00000000001 145000.0 46600.0 ;
      RECT  149000.0 45800.00000000001 149800.0 46600.0 ;
      RECT  153800.0 45800.00000000001 154600.00000000003 46600.0 ;
      RECT  158600.0 45800.00000000001 159400.0 46600.0 ;
      RECT  163399.99999999997 45800.00000000001 164200.0 46600.0 ;
      RECT  168200.0 45800.00000000001 169000.0 46600.0 ;
      RECT  173000.0 45800.00000000001 173800.0 46600.0 ;
      RECT  177800.0 45800.00000000001 178600.00000000003 46600.0 ;
      RECT  182600.0 45800.00000000001 183400.0 46600.0 ;
      RECT  187399.99999999997 45800.00000000001 188200.0 46600.0 ;
      RECT  192200.0 45800.00000000001 193000.0 46600.0 ;
      RECT  197000.0 45800.00000000001 197800.0 46600.0 ;
      RECT  201800.0 45800.00000000001 202600.00000000003 46600.0 ;
      RECT  206600.0 45800.00000000001 207400.0 46600.0 ;
      RECT  4999.999999999997 50600.00000000001 5799.999999999997 51400.00000000001 ;
      RECT  9799.999999999993 50600.00000000001 10599.999999999995 51400.00000000001 ;
      RECT  14599.999999999998 50600.00000000001 15399.999999999998 51400.00000000001 ;
      RECT  19399.999999999996 50600.00000000001 20199.999999999996 51400.00000000001 ;
      RECT  24200.0 50600.00000000001 25000.0 51400.00000000001 ;
      RECT  28999.999999999996 50600.00000000001 29799.999999999996 51400.00000000001 ;
      RECT  67400.0 50600.00000000001 68200.0 51400.00000000001 ;
      RECT  72200.0 50600.00000000001 73000.0 51400.00000000001 ;
      RECT  77000.0 50600.00000000001 77800.0 51400.00000000001 ;
      RECT  81800.0 50600.00000000001 82600.0 51400.00000000001 ;
      RECT  86600.00000000001 50600.00000000001 87400.0 51400.00000000001 ;
      RECT  91400.0 50600.00000000001 92200.0 51400.00000000001 ;
      RECT  96200.0 50600.00000000001 97000.0 51400.00000000001 ;
      RECT  101000.0 50600.00000000001 101800.0 51400.00000000001 ;
      RECT  105800.0 50600.00000000001 106600.0 51400.00000000001 ;
      RECT  110600.00000000001 50600.00000000001 111400.0 51400.00000000001 ;
      RECT  115400.0 50600.00000000001 116200.0 51400.00000000001 ;
      RECT  120200.0 50600.00000000001 121000.0 51400.00000000001 ;
      RECT  125000.00000000001 50600.00000000001 125800.00000000001 51400.00000000001 ;
      RECT  129799.99999999999 50600.00000000001 130600.0 51400.00000000001 ;
      RECT  134600.0 50600.00000000001 135400.0 51400.00000000001 ;
      RECT  139399.99999999997 50600.00000000001 140200.0 51400.00000000001 ;
      RECT  144200.0 50600.00000000001 145000.0 51400.00000000001 ;
      RECT  149000.0 50600.00000000001 149800.0 51400.00000000001 ;
      RECT  153800.0 50600.00000000001 154600.00000000003 51400.00000000001 ;
      RECT  158600.0 50600.00000000001 159400.0 51400.00000000001 ;
      RECT  163399.99999999997 50600.00000000001 164200.0 51400.00000000001 ;
      RECT  168200.0 50600.00000000001 169000.0 51400.00000000001 ;
      RECT  173000.0 50600.00000000001 173800.0 51400.00000000001 ;
      RECT  177800.0 50600.00000000001 178600.00000000003 51400.00000000001 ;
      RECT  182600.0 50600.00000000001 183400.0 51400.00000000001 ;
      RECT  187399.99999999997 50600.00000000001 188200.0 51400.00000000001 ;
      RECT  192200.0 50600.00000000001 193000.0 51400.00000000001 ;
      RECT  197000.0 50600.00000000001 197800.0 51400.00000000001 ;
      RECT  201800.0 50600.00000000001 202600.00000000003 51400.00000000001 ;
      RECT  206600.0 50600.00000000001 207400.0 51400.00000000001 ;
      RECT  4999.999999999997 55400.00000000001 5799.999999999997 56200.0 ;
      RECT  9799.999999999993 55400.00000000001 10599.999999999995 56200.0 ;
      RECT  14599.999999999998 55400.00000000001 15399.999999999998 56200.0 ;
      RECT  19399.999999999996 55400.00000000001 20199.999999999996 56200.0 ;
      RECT  24200.0 55400.00000000001 25000.0 56200.0 ;
      RECT  28999.999999999996 55400.00000000001 29799.999999999996 56200.0 ;
      RECT  33800.0 55400.00000000001 34599.99999999999 56200.0 ;
      RECT  38600.0 55400.00000000001 39400.0 56200.0 ;
      RECT  43400.00000000001 55400.00000000001 44200.0 56200.0 ;
      RECT  48200.0 55400.00000000001 49000.0 56200.0 ;
      RECT  53000.0 55400.00000000001 53800.0 56200.0 ;
      RECT  57800.0 55400.00000000001 58599.99999999999 56200.0 ;
      RECT  62600.0 55400.00000000001 63400.0 56200.0 ;
      RECT  67400.0 55400.00000000001 68200.0 56200.0 ;
      RECT  72200.0 55400.00000000001 73000.0 56200.0 ;
      RECT  77000.0 55400.00000000001 77800.0 56200.0 ;
      RECT  81800.0 55400.00000000001 82600.0 56200.0 ;
      RECT  86600.00000000001 55400.00000000001 87400.0 56200.0 ;
      RECT  91400.0 55400.00000000001 92200.0 56200.0 ;
      RECT  96200.0 55400.00000000001 97000.0 56200.0 ;
      RECT  101000.0 55400.00000000001 101800.0 56200.0 ;
      RECT  105800.0 55400.00000000001 106600.0 56200.0 ;
      RECT  110600.00000000001 55400.00000000001 111400.0 56200.0 ;
      RECT  115400.0 55400.00000000001 116200.0 56200.0 ;
      RECT  120200.0 55400.00000000001 121000.0 56200.0 ;
      RECT  125000.00000000001 55400.00000000001 125800.00000000001 56200.0 ;
      RECT  129799.99999999999 55400.00000000001 130600.0 56200.0 ;
      RECT  134600.0 55400.00000000001 135400.0 56200.0 ;
      RECT  139399.99999999997 55400.00000000001 140200.0 56200.0 ;
      RECT  144200.0 55400.00000000001 145000.0 56200.0 ;
      RECT  149000.0 55400.00000000001 149800.0 56200.0 ;
      RECT  153800.0 55400.00000000001 154600.00000000003 56200.0 ;
      RECT  158600.0 55400.00000000001 159400.0 56200.0 ;
      RECT  163399.99999999997 55400.00000000001 164200.0 56200.0 ;
      RECT  168200.0 55400.00000000001 169000.0 56200.0 ;
      RECT  173000.0 55400.00000000001 173800.0 56200.0 ;
      RECT  177800.0 55400.00000000001 178600.00000000003 56200.0 ;
      RECT  182600.0 55400.00000000001 183400.0 56200.0 ;
      RECT  187399.99999999997 55400.00000000001 188200.0 56200.0 ;
      RECT  192200.0 55400.00000000001 193000.0 56200.0 ;
      RECT  197000.0 55400.00000000001 197800.0 56200.0 ;
      RECT  201800.0 55400.00000000001 202600.00000000003 56200.0 ;
      RECT  206600.0 55400.00000000001 207400.0 56200.0 ;
      RECT  4999.999999999997 60200.0 5799.999999999997 61000.0 ;
      RECT  9799.999999999993 60200.0 10599.999999999995 61000.0 ;
      RECT  14599.999999999998 60200.0 15399.999999999998 61000.0 ;
      RECT  19399.999999999996 60200.0 20199.999999999996 61000.0 ;
      RECT  24200.0 60200.0 25000.0 61000.0 ;
      RECT  28999.999999999996 60200.0 29799.999999999996 61000.0 ;
      RECT  33800.0 60200.0 34599.99999999999 61000.0 ;
      RECT  38600.0 60200.0 39400.0 61000.0 ;
      RECT  43400.00000000001 60200.0 44200.0 61000.0 ;
      RECT  48200.0 60200.0 49000.0 61000.0 ;
      RECT  53000.0 60200.0 53800.0 61000.0 ;
      RECT  57800.0 60200.0 58599.99999999999 61000.0 ;
      RECT  62600.0 60200.0 63400.0 61000.0 ;
      RECT  67400.0 60200.0 68200.0 61000.0 ;
      RECT  72200.0 60200.0 73000.0 61000.0 ;
      RECT  77000.0 60200.0 77800.0 61000.0 ;
      RECT  81800.0 60200.0 82600.0 61000.0 ;
      RECT  86600.00000000001 60200.0 87400.0 61000.0 ;
      RECT  91400.0 60200.0 92200.0 61000.0 ;
      RECT  96200.0 60200.0 97000.0 61000.0 ;
      RECT  101000.0 60200.0 101800.0 61000.0 ;
      RECT  105800.0 60200.0 106600.0 61000.0 ;
      RECT  110600.00000000001 60200.0 111400.0 61000.0 ;
      RECT  115400.0 60200.0 116200.0 61000.0 ;
      RECT  120200.0 60200.0 121000.0 61000.0 ;
      RECT  125000.00000000001 60200.0 125800.00000000001 61000.0 ;
      RECT  129799.99999999999 60200.0 130600.0 61000.0 ;
      RECT  134600.0 60200.0 135400.0 61000.0 ;
      RECT  139399.99999999997 60200.0 140200.0 61000.0 ;
      RECT  144200.0 60200.0 145000.0 61000.0 ;
      RECT  149000.0 60200.0 149800.0 61000.0 ;
      RECT  153800.0 60200.0 154600.00000000003 61000.0 ;
      RECT  158600.0 60200.0 159400.0 61000.0 ;
      RECT  163399.99999999997 60200.0 164200.0 61000.0 ;
      RECT  168200.0 60200.0 169000.0 61000.0 ;
      RECT  173000.0 60200.0 173800.0 61000.0 ;
      RECT  177800.0 60200.0 178600.00000000003 61000.0 ;
      RECT  182600.0 60200.0 183400.0 61000.0 ;
      RECT  187399.99999999997 60200.0 188200.0 61000.0 ;
      RECT  192200.0 60200.0 193000.0 61000.0 ;
      RECT  197000.0 60200.0 197800.0 61000.0 ;
      RECT  201800.0 60200.0 202600.00000000003 61000.0 ;
      RECT  206600.0 60200.0 207400.0 61000.0 ;
      RECT  4999.999999999997 65000.0 5799.999999999997 65800.0 ;
      RECT  9799.999999999993 65000.0 10599.999999999995 65800.0 ;
      RECT  14599.999999999998 65000.0 15399.999999999998 65800.0 ;
      RECT  19399.999999999996 65000.0 20199.999999999996 65800.0 ;
      RECT  24200.0 65000.0 25000.0 65800.0 ;
      RECT  28999.999999999996 65000.0 29799.999999999996 65800.0 ;
      RECT  33800.0 65000.0 34599.99999999999 65800.0 ;
      RECT  38600.0 65000.0 39400.0 65800.0 ;
      RECT  43400.00000000001 65000.0 44200.0 65800.0 ;
      RECT  48200.0 65000.0 49000.0 65800.0 ;
      RECT  53000.0 65000.0 53800.0 65800.0 ;
      RECT  57800.0 65000.0 58599.99999999999 65800.0 ;
      RECT  62600.0 65000.0 63400.0 65800.0 ;
      RECT  67400.0 65000.0 68200.0 65800.0 ;
      RECT  72200.0 65000.0 73000.0 65800.0 ;
      RECT  77000.0 65000.0 77800.0 65800.0 ;
      RECT  81800.0 65000.0 82600.0 65800.0 ;
      RECT  86600.00000000001 65000.0 87400.0 65800.0 ;
      RECT  91400.0 65000.0 92200.0 65800.0 ;
      RECT  96200.0 65000.0 97000.0 65800.0 ;
      RECT  101000.0 65000.0 101800.0 65800.0 ;
      RECT  105800.0 65000.0 106600.0 65800.0 ;
      RECT  110600.00000000001 65000.0 111400.0 65800.0 ;
      RECT  115400.0 65000.0 116200.0 65800.0 ;
      RECT  120200.0 65000.0 121000.0 65800.0 ;
      RECT  125000.00000000001 65000.0 125800.00000000001 65800.0 ;
      RECT  129799.99999999999 65000.0 130600.0 65800.0 ;
      RECT  134600.0 65000.0 135400.0 65800.0 ;
      RECT  139399.99999999997 65000.0 140200.0 65800.0 ;
      RECT  144200.0 65000.0 145000.0 65800.0 ;
      RECT  149000.0 65000.0 149800.0 65800.0 ;
      RECT  153800.0 65000.0 154600.00000000003 65800.0 ;
      RECT  158600.0 65000.0 159400.0 65800.0 ;
      RECT  163399.99999999997 65000.0 164200.0 65800.0 ;
      RECT  168200.0 65000.0 169000.0 65800.0 ;
      RECT  173000.0 65000.0 173800.0 65800.0 ;
      RECT  177800.0 65000.0 178600.00000000003 65800.0 ;
      RECT  182600.0 65000.0 183400.0 65800.0 ;
      RECT  187399.99999999997 65000.0 188200.0 65800.0 ;
      RECT  192200.0 65000.0 193000.0 65800.0 ;
      RECT  197000.0 65000.0 197800.0 65800.0 ;
      RECT  201800.0 65000.0 202600.00000000003 65800.0 ;
      RECT  206600.0 65000.0 207400.0 65800.0 ;
      RECT  4999.999999999997 69800.00000000001 5799.999999999997 70600.00000000001 ;
      RECT  9799.999999999993 69800.00000000001 10599.999999999995 70600.00000000001 ;
      RECT  14599.999999999998 69800.00000000001 15399.999999999998 70600.00000000001 ;
      RECT  19399.999999999996 69800.00000000001 20199.999999999996 70600.00000000001 ;
      RECT  24200.0 69800.00000000001 25000.0 70600.00000000001 ;
      RECT  28999.999999999996 69800.00000000001 29799.999999999996 70600.00000000001 ;
      RECT  33800.0 69800.00000000001 34599.99999999999 70600.00000000001 ;
      RECT  38600.0 69800.00000000001 39400.0 70600.00000000001 ;
      RECT  43400.00000000001 69800.00000000001 44200.0 70600.00000000001 ;
      RECT  48200.0 69800.00000000001 49000.0 70600.00000000001 ;
      RECT  53000.0 69800.00000000001 53800.0 70600.00000000001 ;
      RECT  57800.0 69800.00000000001 58599.99999999999 70600.00000000001 ;
      RECT  62600.0 69800.00000000001 63400.0 70600.00000000001 ;
      RECT  67400.0 69800.00000000001 68200.0 70600.00000000001 ;
      RECT  72200.0 69800.00000000001 73000.0 70600.00000000001 ;
      RECT  77000.0 69800.00000000001 77800.0 70600.00000000001 ;
      RECT  81800.0 69800.00000000001 82600.0 70600.00000000001 ;
      RECT  86600.00000000001 69800.00000000001 87400.0 70600.00000000001 ;
      RECT  91400.0 69800.00000000001 92200.0 70600.00000000001 ;
      RECT  96200.0 69800.00000000001 97000.0 70600.00000000001 ;
      RECT  101000.0 69800.00000000001 101800.0 70600.00000000001 ;
      RECT  105800.0 69800.00000000001 106600.0 70600.00000000001 ;
      RECT  110600.00000000001 69800.00000000001 111400.0 70600.00000000001 ;
      RECT  115400.0 69800.00000000001 116200.0 70600.00000000001 ;
      RECT  120200.0 69800.00000000001 121000.0 70600.00000000001 ;
      RECT  125000.00000000001 69800.00000000001 125800.00000000001 70600.00000000001 ;
      RECT  129799.99999999999 69800.00000000001 130600.0 70600.00000000001 ;
      RECT  134600.0 69800.00000000001 135400.0 70600.00000000001 ;
      RECT  139399.99999999997 69800.00000000001 140200.0 70600.00000000001 ;
      RECT  144200.0 69800.00000000001 145000.0 70600.00000000001 ;
      RECT  149000.0 69800.00000000001 149800.0 70600.00000000001 ;
      RECT  153800.0 69800.00000000001 154600.00000000003 70600.00000000001 ;
      RECT  158600.0 69800.00000000001 159400.0 70600.00000000001 ;
      RECT  163399.99999999997 69800.00000000001 164200.0 70600.00000000001 ;
      RECT  168200.0 69800.00000000001 169000.0 70600.00000000001 ;
      RECT  173000.0 69800.00000000001 173800.0 70600.00000000001 ;
      RECT  177800.0 69800.00000000001 178600.00000000003 70600.00000000001 ;
      RECT  182600.0 69800.00000000001 183400.0 70600.00000000001 ;
      RECT  187399.99999999997 69800.00000000001 188200.0 70600.00000000001 ;
      RECT  192200.0 69800.00000000001 193000.0 70600.00000000001 ;
      RECT  197000.0 69800.00000000001 197800.0 70600.00000000001 ;
      RECT  201800.0 69800.00000000001 202600.00000000003 70600.00000000001 ;
      RECT  206600.0 69800.00000000001 207400.0 70600.00000000001 ;
      RECT  4999.999999999997 74600.00000000001 5799.999999999997 75400.0 ;
      RECT  9799.999999999993 74600.00000000001 10599.999999999995 75400.0 ;
      RECT  14599.999999999998 74600.00000000001 15399.999999999998 75400.0 ;
      RECT  19399.999999999996 74600.00000000001 20199.999999999996 75400.0 ;
      RECT  24200.0 74600.00000000001 25000.0 75400.0 ;
      RECT  28999.999999999996 74600.00000000001 29799.999999999996 75400.0 ;
      RECT  33800.0 74600.00000000001 34599.99999999999 75400.0 ;
      RECT  38600.0 74600.00000000001 39400.0 75400.0 ;
      RECT  43400.00000000001 74600.00000000001 44200.0 75400.0 ;
      RECT  48200.0 74600.00000000001 49000.0 75400.0 ;
      RECT  53000.0 74600.00000000001 53800.0 75400.0 ;
      RECT  57800.0 74600.00000000001 58599.99999999999 75400.0 ;
      RECT  62600.0 74600.00000000001 63400.0 75400.0 ;
      RECT  67400.0 74600.00000000001 68200.0 75400.0 ;
      RECT  72200.0 74600.00000000001 73000.0 75400.0 ;
      RECT  77000.0 74600.00000000001 77800.0 75400.0 ;
      RECT  81800.0 74600.00000000001 82600.0 75400.0 ;
      RECT  86600.00000000001 74600.00000000001 87400.0 75400.0 ;
      RECT  91400.0 74600.00000000001 92200.0 75400.0 ;
      RECT  96200.0 74600.00000000001 97000.0 75400.0 ;
      RECT  101000.0 74600.00000000001 101800.0 75400.0 ;
      RECT  105800.0 74600.00000000001 106600.0 75400.0 ;
      RECT  110600.00000000001 74600.00000000001 111400.0 75400.0 ;
      RECT  115400.0 74600.00000000001 116200.0 75400.0 ;
      RECT  120200.0 74600.00000000001 121000.0 75400.0 ;
      RECT  125000.00000000001 74600.00000000001 125800.00000000001 75400.0 ;
      RECT  129799.99999999999 74600.00000000001 130600.0 75400.0 ;
      RECT  134600.0 74600.00000000001 135400.0 75400.0 ;
      RECT  139399.99999999997 74600.00000000001 140200.0 75400.0 ;
      RECT  144200.0 74600.00000000001 145000.0 75400.0 ;
      RECT  149000.0 74600.00000000001 149800.0 75400.0 ;
      RECT  153800.0 74600.00000000001 154600.00000000003 75400.0 ;
      RECT  158600.0 74600.00000000001 159400.0 75400.0 ;
      RECT  163399.99999999997 74600.00000000001 164200.0 75400.0 ;
      RECT  168200.0 74600.00000000001 169000.0 75400.0 ;
      RECT  173000.0 74600.00000000001 173800.0 75400.0 ;
      RECT  177800.0 74600.00000000001 178600.00000000003 75400.0 ;
      RECT  182600.0 74600.00000000001 183400.0 75400.0 ;
      RECT  187399.99999999997 74600.00000000001 188200.0 75400.0 ;
      RECT  192200.0 74600.00000000001 193000.0 75400.0 ;
      RECT  197000.0 74600.00000000001 197800.0 75400.0 ;
      RECT  201800.0 74600.00000000001 202600.00000000003 75400.0 ;
      RECT  206600.0 74600.00000000001 207400.0 75400.0 ;
      RECT  4999.999999999997 79400.0 5799.999999999997 80200.0 ;
      RECT  9799.999999999993 79400.0 10599.999999999995 80200.0 ;
      RECT  14599.999999999998 79400.0 15399.999999999998 80200.0 ;
      RECT  19399.999999999996 79400.0 20199.999999999996 80200.0 ;
      RECT  24200.0 79400.0 25000.0 80200.0 ;
      RECT  28999.999999999996 79400.0 29799.999999999996 80200.0 ;
      RECT  33800.0 79400.0 34599.99999999999 80200.0 ;
      RECT  38600.0 79400.0 39400.0 80200.0 ;
      RECT  43400.00000000001 79400.0 44200.0 80200.0 ;
      RECT  48200.0 79400.0 49000.0 80200.0 ;
      RECT  53000.0 79400.0 53800.0 80200.0 ;
      RECT  57800.0 79400.0 58599.99999999999 80200.0 ;
      RECT  62600.0 79400.0 63400.0 80200.0 ;
      RECT  77000.0 79400.0 77800.0 80200.0 ;
      RECT  81800.0 79400.0 82600.0 80200.0 ;
      RECT  86600.00000000001 79400.0 87400.0 80200.0 ;
      RECT  91400.0 79400.0 92200.0 80200.0 ;
      RECT  96200.0 79400.0 97000.0 80200.0 ;
      RECT  101000.0 79400.0 101800.0 80200.0 ;
      RECT  105800.0 79400.0 106600.0 80200.0 ;
      RECT  110600.00000000001 79400.0 111400.0 80200.0 ;
      RECT  115400.0 79400.0 116200.0 80200.0 ;
      RECT  120200.0 79400.0 121000.0 80200.0 ;
      RECT  125000.00000000001 79400.0 125800.00000000001 80200.0 ;
      RECT  129799.99999999999 79400.0 130600.0 80200.0 ;
      RECT  134600.0 79400.0 135400.0 80200.0 ;
      RECT  139399.99999999997 79400.0 140200.0 80200.0 ;
      RECT  144200.0 79400.0 145000.0 80200.0 ;
      RECT  149000.0 79400.0 149800.0 80200.0 ;
      RECT  153800.0 79400.0 154600.00000000003 80200.0 ;
      RECT  158600.0 79400.0 159400.0 80200.0 ;
      RECT  163399.99999999997 79400.0 164200.0 80200.0 ;
      RECT  168200.0 79400.0 169000.0 80200.0 ;
      RECT  173000.0 79400.0 173800.0 80200.0 ;
      RECT  177800.0 79400.0 178600.00000000003 80200.0 ;
      RECT  182600.0 79400.0 183400.0 80200.0 ;
      RECT  187399.99999999997 79400.0 188200.0 80200.0 ;
      RECT  192200.0 79400.0 193000.0 80200.0 ;
      RECT  197000.0 79400.0 197800.0 80200.0 ;
      RECT  201800.0 79400.0 202600.00000000003 80200.0 ;
      RECT  206600.0 79400.0 207400.0 80200.0 ;
      RECT  4999.999999999997 84200.0 5799.999999999997 85000.0 ;
      RECT  9799.999999999993 84200.0 10599.999999999995 85000.0 ;
      RECT  14599.999999999998 84200.0 15399.999999999998 85000.0 ;
      RECT  19399.999999999996 84200.0 20199.999999999996 85000.0 ;
      RECT  24200.0 84200.0 25000.0 85000.0 ;
      RECT  28999.999999999996 84200.0 29799.999999999996 85000.0 ;
      RECT  33800.0 84200.0 34599.99999999999 85000.0 ;
      RECT  38600.0 84200.0 39400.0 85000.0 ;
      RECT  43400.00000000001 84200.0 44200.0 85000.0 ;
      RECT  48200.0 84200.0 49000.0 85000.0 ;
      RECT  53000.0 84200.0 53800.0 85000.0 ;
      RECT  57800.0 84200.0 58599.99999999999 85000.0 ;
      RECT  62600.0 84200.0 63400.0 85000.0 ;
      RECT  67400.0 84200.0 68200.0 85000.0 ;
      RECT  72200.0 84200.0 73000.0 85000.0 ;
      RECT  77000.0 84200.0 77800.0 85000.0 ;
      RECT  81800.0 84200.0 82600.0 85000.0 ;
      RECT  86600.00000000001 84200.0 87400.0 85000.0 ;
      RECT  91400.0 84200.0 92200.0 85000.0 ;
      RECT  96200.0 84200.0 97000.0 85000.0 ;
      RECT  101000.0 84200.0 101800.0 85000.0 ;
      RECT  105800.0 84200.0 106600.0 85000.0 ;
      RECT  110600.00000000001 84200.0 111400.0 85000.0 ;
      RECT  115400.0 84200.0 116200.0 85000.0 ;
      RECT  120200.0 84200.0 121000.0 85000.0 ;
      RECT  125000.00000000001 84200.0 125800.00000000001 85000.0 ;
      RECT  129799.99999999999 84200.0 130600.0 85000.0 ;
      RECT  134600.0 84200.0 135400.0 85000.0 ;
      RECT  139399.99999999997 84200.0 140200.0 85000.0 ;
      RECT  144200.0 84200.0 145000.0 85000.0 ;
      RECT  149000.0 84200.0 149800.0 85000.0 ;
      RECT  153800.0 84200.0 154600.00000000003 85000.0 ;
      RECT  158600.0 84200.0 159400.0 85000.0 ;
      RECT  163399.99999999997 84200.0 164200.0 85000.0 ;
      RECT  4999.999999999997 89000.00000000001 5799.999999999997 89800.00000000001 ;
      RECT  9799.999999999993 89000.00000000001 10599.999999999995 89800.00000000001 ;
      RECT  14599.999999999998 89000.00000000001 15399.999999999998 89800.00000000001 ;
      RECT  19399.999999999996 89000.00000000001 20199.999999999996 89800.00000000001 ;
      RECT  24200.0 89000.00000000001 25000.0 89800.00000000001 ;
      RECT  28999.999999999996 89000.00000000001 29799.999999999996 89800.00000000001 ;
      RECT  33800.0 89000.00000000001 34599.99999999999 89800.00000000001 ;
      RECT  38600.0 89000.00000000001 39400.0 89800.00000000001 ;
      RECT  43400.00000000001 89000.00000000001 44200.0 89800.00000000001 ;
      RECT  48200.0 89000.00000000001 49000.0 89800.00000000001 ;
      RECT  53000.0 89000.00000000001 53800.0 89800.00000000001 ;
      RECT  57800.0 89000.00000000001 58599.99999999999 89800.00000000001 ;
      RECT  62600.0 89000.00000000001 63400.0 89800.00000000001 ;
      RECT  4999.999999999997 93800.00000000001 5799.999999999997 94600.00000000001 ;
      RECT  9799.999999999993 93800.00000000001 10599.999999999995 94600.00000000001 ;
      RECT  14599.999999999998 93800.00000000001 15399.999999999998 94600.00000000001 ;
      RECT  19399.999999999996 93800.00000000001 20199.999999999996 94600.00000000001 ;
      RECT  24200.0 93800.00000000001 25000.0 94600.00000000001 ;
      RECT  28999.999999999996 93800.00000000001 29799.999999999996 94600.00000000001 ;
      RECT  33800.0 93800.00000000001 34599.99999999999 94600.00000000001 ;
      RECT  38600.0 93800.00000000001 39400.0 94600.00000000001 ;
      RECT  43400.00000000001 93800.00000000001 44200.0 94600.00000000001 ;
      RECT  48200.0 93800.00000000001 49000.0 94600.00000000001 ;
      RECT  53000.0 93800.00000000001 53800.0 94600.00000000001 ;
      RECT  57800.0 93800.00000000001 58599.99999999999 94600.00000000001 ;
      RECT  62600.0 93800.00000000001 63400.0 94600.00000000001 ;
      RECT  67400.0 93800.00000000001 68200.0 94600.00000000001 ;
      RECT  72200.0 93800.00000000001 73000.0 94600.00000000001 ;
      RECT  77000.0 93800.00000000001 77800.0 94600.00000000001 ;
      RECT  81800.0 93800.00000000001 82600.0 94600.00000000001 ;
      RECT  86600.00000000001 93800.00000000001 87400.0 94600.00000000001 ;
      RECT  91400.0 93800.00000000001 92200.0 94600.00000000001 ;
      RECT  96200.0 93800.00000000001 97000.0 94600.00000000001 ;
      RECT  101000.0 93800.00000000001 101800.0 94600.00000000001 ;
      RECT  105800.0 93800.00000000001 106600.0 94600.00000000001 ;
      RECT  110600.00000000001 93800.00000000001 111400.0 94600.00000000001 ;
      RECT  115400.0 93800.00000000001 116200.0 94600.00000000001 ;
      RECT  120200.0 93800.00000000001 121000.0 94600.00000000001 ;
      RECT  125000.00000000001 93800.00000000001 125800.00000000001 94600.00000000001 ;
      RECT  129799.99999999999 93800.00000000001 130600.0 94600.00000000001 ;
      RECT  134600.0 93800.00000000001 135400.0 94600.00000000001 ;
      RECT  139399.99999999997 93800.00000000001 140200.0 94600.00000000001 ;
      RECT  144200.0 93800.00000000001 145000.0 94600.00000000001 ;
      RECT  149000.0 93800.00000000001 149800.0 94600.00000000001 ;
      RECT  153800.0 93800.00000000001 154600.00000000003 94600.00000000001 ;
      RECT  158600.0 93800.00000000001 159400.0 94600.00000000001 ;
      RECT  163399.99999999997 93800.00000000001 164200.0 94600.00000000001 ;
      RECT  168200.0 93800.00000000001 169000.0 94600.00000000001 ;
      RECT  173000.0 93800.00000000001 173800.0 94600.00000000001 ;
      RECT  177800.0 93800.00000000001 178600.00000000003 94600.00000000001 ;
      RECT  182600.0 93800.00000000001 183400.0 94600.00000000001 ;
      RECT  187399.99999999997 93800.00000000001 188200.0 94600.00000000001 ;
      RECT  192200.0 93800.00000000001 193000.0 94600.00000000001 ;
      RECT  197000.0 93800.00000000001 197800.0 94600.00000000001 ;
      RECT  201800.0 93800.00000000001 202600.00000000003 94600.00000000001 ;
      RECT  206600.0 93800.00000000001 207400.0 94600.00000000001 ;
      RECT  4999.999999999997 98600.00000000001 5799.999999999997 99400.0 ;
      RECT  9799.999999999993 98600.00000000001 10599.999999999995 99400.0 ;
      RECT  14599.999999999998 98600.00000000001 15399.999999999998 99400.0 ;
      RECT  19399.999999999996 98600.00000000001 20199.999999999996 99400.0 ;
      RECT  24200.0 98600.00000000001 25000.0 99400.0 ;
      RECT  28999.999999999996 98600.00000000001 29799.999999999996 99400.0 ;
      RECT  33800.0 98600.00000000001 34599.99999999999 99400.0 ;
      RECT  38600.0 98600.00000000001 39400.0 99400.0 ;
      RECT  43400.00000000001 98600.00000000001 44200.0 99400.0 ;
      RECT  48200.0 98600.00000000001 49000.0 99400.0 ;
      RECT  53000.0 98600.00000000001 53800.0 99400.0 ;
      RECT  57800.0 98600.00000000001 58599.99999999999 99400.0 ;
      RECT  62600.0 98600.00000000001 63400.0 99400.0 ;
      RECT  67400.0 98600.00000000001 68200.0 99400.0 ;
      RECT  72200.0 98600.00000000001 73000.0 99400.0 ;
      RECT  77000.0 98600.00000000001 77800.0 99400.0 ;
      RECT  81800.0 98600.00000000001 82600.0 99400.0 ;
      RECT  86600.00000000001 98600.00000000001 87400.0 99400.0 ;
      RECT  91400.0 98600.00000000001 92200.0 99400.0 ;
      RECT  96200.0 98600.00000000001 97000.0 99400.0 ;
      RECT  101000.0 98600.00000000001 101800.0 99400.0 ;
      RECT  105800.0 98600.00000000001 106600.0 99400.0 ;
      RECT  110600.00000000001 98600.00000000001 111400.0 99400.0 ;
      RECT  115400.0 98600.00000000001 116200.0 99400.0 ;
      RECT  120200.0 98600.00000000001 121000.0 99400.0 ;
      RECT  125000.00000000001 98600.00000000001 125800.00000000001 99400.0 ;
      RECT  129799.99999999999 98600.00000000001 130600.0 99400.0 ;
      RECT  134600.0 98600.00000000001 135400.0 99400.0 ;
      RECT  139399.99999999997 98600.00000000001 140200.0 99400.0 ;
      RECT  144200.0 98600.00000000001 145000.0 99400.0 ;
      RECT  149000.0 98600.00000000001 149800.0 99400.0 ;
      RECT  153800.0 98600.00000000001 154600.00000000003 99400.0 ;
      RECT  158600.0 98600.00000000001 159400.0 99400.0 ;
      RECT  163399.99999999997 98600.00000000001 164200.0 99400.0 ;
      RECT  168200.0 98600.00000000001 169000.0 99400.0 ;
      RECT  187399.99999999997 98600.00000000001 188200.0 99400.0 ;
      RECT  192200.0 98600.00000000001 193000.0 99400.0 ;
      RECT  197000.0 98600.00000000001 197800.0 99400.0 ;
      RECT  201800.0 98600.00000000001 202600.00000000003 99400.0 ;
      RECT  206600.0 98600.00000000001 207400.0 99400.0 ;
      RECT  4999.999999999997 103400.0 5799.999999999997 104200.0 ;
      RECT  9799.999999999993 103400.0 10599.999999999995 104200.0 ;
      RECT  14599.999999999998 103400.0 15399.999999999998 104200.0 ;
      RECT  19399.999999999996 103400.0 20199.999999999996 104200.0 ;
      RECT  24200.0 103400.0 25000.0 104200.0 ;
      RECT  28999.999999999996 103400.0 29799.999999999996 104200.0 ;
      RECT  33800.0 103400.0 34599.99999999999 104200.0 ;
      RECT  38600.0 103400.0 39400.0 104200.0 ;
      RECT  43400.00000000001 103400.0 44200.0 104200.0 ;
      RECT  48200.0 103400.0 49000.0 104200.0 ;
      RECT  53000.0 103400.0 53800.0 104200.0 ;
      RECT  57800.0 103400.0 58599.99999999999 104200.0 ;
      RECT  62600.0 103400.0 63400.0 104200.0 ;
      RECT  67400.0 103400.0 68200.0 104200.0 ;
      RECT  72200.0 103400.0 73000.0 104200.0 ;
      RECT  77000.0 103400.0 77800.0 104200.0 ;
      RECT  81800.0 103400.0 82600.0 104200.0 ;
      RECT  86600.00000000001 103400.0 87400.0 104200.0 ;
      RECT  91400.0 103400.0 92200.0 104200.0 ;
      RECT  96200.0 103400.0 97000.0 104200.0 ;
      RECT  101000.0 103400.0 101800.0 104200.0 ;
      RECT  105800.0 103400.0 106600.0 104200.0 ;
      RECT  110600.00000000001 103400.0 111400.0 104200.0 ;
      RECT  115400.0 103400.0 116200.0 104200.0 ;
      RECT  120200.0 103400.0 121000.0 104200.0 ;
      RECT  125000.00000000001 103400.0 125800.00000000001 104200.0 ;
      RECT  129799.99999999999 103400.0 130600.0 104200.0 ;
      RECT  134600.0 103400.0 135400.0 104200.0 ;
      RECT  139399.99999999997 103400.0 140200.0 104200.0 ;
      RECT  144200.0 103400.0 145000.0 104200.0 ;
      RECT  149000.0 103400.0 149800.0 104200.0 ;
      RECT  153800.0 103400.0 154600.00000000003 104200.0 ;
      RECT  158600.0 103400.0 159400.0 104200.0 ;
      RECT  163399.99999999997 103400.0 164200.0 104200.0 ;
      RECT  168200.0 103400.0 169000.0 104200.0 ;
      RECT  173000.0 103400.0 173800.0 104200.0 ;
      RECT  177800.0 103400.0 178600.00000000003 104200.0 ;
      RECT  182600.0 103400.0 183400.0 104200.0 ;
      RECT  187399.99999999997 103400.0 188200.0 104200.0 ;
      RECT  192200.0 103400.0 193000.0 104200.0 ;
      RECT  197000.0 103400.0 197800.0 104200.0 ;
      RECT  201800.0 103400.0 202600.00000000003 104200.0 ;
      RECT  206600.0 103400.0 207400.0 104200.0 ;
      RECT  4999.999999999997 108200.0 5799.999999999997 109000.0 ;
      RECT  9799.999999999993 108200.0 10599.999999999995 109000.0 ;
      RECT  14599.999999999998 108200.0 15399.999999999998 109000.0 ;
      RECT  19399.999999999996 108200.0 20199.999999999996 109000.0 ;
      RECT  24200.0 108200.0 25000.0 109000.0 ;
      RECT  28999.999999999996 108200.0 29799.999999999996 109000.0 ;
      RECT  33800.0 108200.0 34599.99999999999 109000.0 ;
      RECT  38600.0 108200.0 39400.0 109000.0 ;
      RECT  43400.00000000001 108200.0 44200.0 109000.0 ;
      RECT  48200.0 108200.0 49000.0 109000.0 ;
      RECT  53000.0 108200.0 53800.0 109000.0 ;
      RECT  57800.0 108200.0 58599.99999999999 109000.0 ;
      RECT  62600.0 108200.0 63400.0 109000.0 ;
      RECT  67400.0 108200.0 68200.0 109000.0 ;
      RECT  72200.0 108200.0 73000.0 109000.0 ;
      RECT  77000.0 108200.0 77800.0 109000.0 ;
      RECT  81800.0 108200.0 82600.0 109000.0 ;
      RECT  86600.00000000001 108200.0 87400.0 109000.0 ;
      RECT  91400.0 108200.0 92200.0 109000.0 ;
      RECT  96200.0 108200.0 97000.0 109000.0 ;
      RECT  101000.0 108200.0 101800.0 109000.0 ;
      RECT  105800.0 108200.0 106600.0 109000.0 ;
      RECT  110600.00000000001 108200.0 111400.0 109000.0 ;
      RECT  115400.0 108200.0 116200.0 109000.0 ;
      RECT  120200.0 108200.0 121000.0 109000.0 ;
      RECT  125000.00000000001 108200.0 125800.00000000001 109000.0 ;
      RECT  129799.99999999999 108200.0 130600.0 109000.0 ;
      RECT  134600.0 108200.0 135400.0 109000.0 ;
      RECT  139399.99999999997 108200.0 140200.0 109000.0 ;
      RECT  144200.0 108200.0 145000.0 109000.0 ;
      RECT  149000.0 108200.0 149800.0 109000.0 ;
      RECT  153800.0 108200.0 154600.00000000003 109000.0 ;
      RECT  158600.0 108200.0 159400.0 109000.0 ;
      RECT  163399.99999999997 108200.0 164200.0 109000.0 ;
      RECT  168200.0 108200.0 169000.0 109000.0 ;
      RECT  173000.0 108200.0 173800.0 109000.0 ;
      RECT  177800.0 108200.0 178600.00000000003 109000.0 ;
      RECT  182600.0 108200.0 183400.0 109000.0 ;
      RECT  187399.99999999997 108200.0 188200.0 109000.0 ;
      RECT  192200.0 108200.0 193000.0 109000.0 ;
      RECT  197000.0 108200.0 197800.0 109000.0 ;
      RECT  201800.0 108200.0 202600.00000000003 109000.0 ;
      RECT  206600.0 108200.0 207400.0 109000.0 ;
      RECT  67400.0 113000.00000000001 68200.0 113800.00000000001 ;
      RECT  72200.0 113000.00000000001 73000.0 113800.00000000001 ;
      RECT  77000.0 113000.00000000001 77800.0 113800.00000000001 ;
      RECT  81800.0 113000.00000000001 82600.0 113800.00000000001 ;
      RECT  86600.00000000001 113000.00000000001 87400.0 113800.00000000001 ;
      RECT  91400.0 113000.00000000001 92200.0 113800.00000000001 ;
      RECT  96200.0 113000.00000000001 97000.0 113800.00000000001 ;
      RECT  101000.0 113000.00000000001 101800.0 113800.00000000001 ;
      RECT  105800.0 113000.00000000001 106600.0 113800.00000000001 ;
      RECT  110600.00000000001 113000.00000000001 111400.0 113800.00000000001 ;
      RECT  115400.0 113000.00000000001 116200.0 113800.00000000001 ;
      RECT  120200.0 113000.00000000001 121000.0 113800.00000000001 ;
      RECT  125000.00000000001 113000.00000000001 125800.00000000001 113800.00000000001 ;
      RECT  129799.99999999999 113000.00000000001 130600.0 113800.00000000001 ;
      RECT  134600.0 113000.00000000001 135400.0 113800.00000000001 ;
      RECT  139399.99999999997 113000.00000000001 140200.0 113800.00000000001 ;
      RECT  144200.0 113000.00000000001 145000.0 113800.00000000001 ;
      RECT  149000.0 113000.00000000001 149800.0 113800.00000000001 ;
      RECT  153800.0 113000.00000000001 154600.00000000003 113800.00000000001 ;
      RECT  158600.0 113000.00000000001 159400.0 113800.00000000001 ;
      RECT  163399.99999999997 113000.00000000001 164200.0 113800.00000000001 ;
      RECT  168200.0 113000.00000000001 169000.0 113800.00000000001 ;
      RECT  173000.0 113000.00000000001 173800.0 113800.00000000001 ;
      RECT  177800.0 113000.00000000001 178600.00000000003 113800.00000000001 ;
      RECT  182600.0 113000.00000000001 183400.0 113800.00000000001 ;
      RECT  187399.99999999997 113000.00000000001 188200.0 113800.00000000001 ;
      RECT  192200.0 113000.00000000001 193000.0 113800.00000000001 ;
      RECT  197000.0 113000.00000000001 197800.0 113800.00000000001 ;
      RECT  201800.0 113000.00000000001 202600.00000000003 113800.00000000001 ;
      RECT  206600.0 113000.00000000001 207400.0 113800.00000000001 ;
      RECT  4999.999999999997 117800.00000000001 5799.999999999997 118600.00000000001 ;
      RECT  9799.999999999993 117800.00000000001 10599.999999999995 118600.00000000001 ;
      RECT  14599.999999999998 117800.00000000001 15399.999999999998 118600.00000000001 ;
      RECT  19399.999999999996 117800.00000000001 20199.999999999996 118600.00000000001 ;
      RECT  24200.0 117800.00000000001 25000.0 118600.00000000001 ;
      RECT  28999.999999999996 117800.00000000001 29799.999999999996 118600.00000000001 ;
      RECT  33800.0 117800.00000000001 34599.99999999999 118600.00000000001 ;
      RECT  38600.0 117800.00000000001 39400.0 118600.00000000001 ;
      RECT  43400.00000000001 117800.00000000001 44200.0 118600.00000000001 ;
      RECT  48200.0 117800.00000000001 49000.0 118600.00000000001 ;
      RECT  53000.0 117800.00000000001 53800.0 118600.00000000001 ;
      RECT  57800.0 117800.00000000001 58599.99999999999 118600.00000000001 ;
      RECT  62600.0 117800.00000000001 63400.0 118600.00000000001 ;
      RECT  67400.0 117800.00000000001 68200.0 118600.00000000001 ;
      RECT  72200.0 117800.00000000001 73000.0 118600.00000000001 ;
      RECT  77000.0 117800.00000000001 77800.0 118600.00000000001 ;
      RECT  81800.0 117800.00000000001 82600.0 118600.00000000001 ;
      RECT  86600.00000000001 117800.00000000001 87400.0 118600.00000000001 ;
      RECT  91400.0 117800.00000000001 92200.0 118600.00000000001 ;
      RECT  96200.0 117800.00000000001 97000.0 118600.00000000001 ;
      RECT  101000.0 117800.00000000001 101800.0 118600.00000000001 ;
      RECT  105800.0 117800.00000000001 106600.0 118600.00000000001 ;
      RECT  110600.00000000001 117800.00000000001 111400.0 118600.00000000001 ;
      RECT  115400.0 117800.00000000001 116200.0 118600.00000000001 ;
      RECT  120200.0 117800.00000000001 121000.0 118600.00000000001 ;
      RECT  125000.00000000001 117800.00000000001 125800.00000000001 118600.00000000001 ;
      RECT  129799.99999999999 117800.00000000001 130600.0 118600.00000000001 ;
      RECT  134600.0 117800.00000000001 135400.0 118600.00000000001 ;
      RECT  139399.99999999997 117800.00000000001 140200.0 118600.00000000001 ;
      RECT  144200.0 117800.00000000001 145000.0 118600.00000000001 ;
      RECT  149000.0 117800.00000000001 149800.0 118600.00000000001 ;
      RECT  153800.0 117800.00000000001 154600.00000000003 118600.00000000001 ;
      RECT  158600.0 117800.00000000001 159400.0 118600.00000000001 ;
      RECT  163399.99999999997 117800.00000000001 164200.0 118600.00000000001 ;
      RECT  168200.0 117800.00000000001 169000.0 118600.00000000001 ;
      RECT  173000.0 117800.00000000001 173800.0 118600.00000000001 ;
      RECT  177800.0 117800.00000000001 178600.00000000003 118600.00000000001 ;
      RECT  182600.0 117800.00000000001 183400.0 118600.00000000001 ;
      RECT  187399.99999999997 117800.00000000001 188200.0 118600.00000000001 ;
      RECT  192200.0 117800.00000000001 193000.0 118600.00000000001 ;
      RECT  197000.0 117800.00000000001 197800.0 118600.00000000001 ;
      RECT  201800.0 117800.00000000001 202600.00000000003 118600.00000000001 ;
      RECT  206600.0 117800.00000000001 207400.0 118600.00000000001 ;
      RECT  4999.999999999997 122600.00000000001 5799.999999999997 123400.0 ;
      RECT  9799.999999999993 122600.00000000001 10599.999999999995 123400.0 ;
      RECT  14599.999999999998 122600.00000000001 15399.999999999998 123400.0 ;
      RECT  19399.999999999996 122600.00000000001 20199.999999999996 123400.0 ;
      RECT  24200.0 122600.00000000001 25000.0 123400.0 ;
      RECT  28999.999999999996 122600.00000000001 29799.999999999996 123400.0 ;
      RECT  33800.0 122600.00000000001 34599.99999999999 123400.0 ;
      RECT  38600.0 122600.00000000001 39400.0 123400.0 ;
      RECT  43400.00000000001 122600.00000000001 44200.0 123400.0 ;
      RECT  48200.0 122600.00000000001 49000.0 123400.0 ;
      RECT  53000.0 122600.00000000001 53800.0 123400.0 ;
      RECT  57800.0 122600.00000000001 58599.99999999999 123400.0 ;
      RECT  62600.0 122600.00000000001 63400.0 123400.0 ;
      RECT  77000.0 122600.00000000001 77800.0 123400.0 ;
      RECT  81800.0 122600.00000000001 82600.0 123400.0 ;
      RECT  86600.00000000001 122600.00000000001 87400.0 123400.0 ;
      RECT  91400.0 122600.00000000001 92200.0 123400.0 ;
      RECT  96200.0 122600.00000000001 97000.0 123400.0 ;
      RECT  101000.0 122600.00000000001 101800.0 123400.0 ;
      RECT  105800.0 122600.00000000001 106600.0 123400.0 ;
      RECT  110600.00000000001 122600.00000000001 111400.0 123400.0 ;
      RECT  115400.0 122600.00000000001 116200.0 123400.0 ;
      RECT  120200.0 122600.00000000001 121000.0 123400.0 ;
      RECT  125000.00000000001 122600.00000000001 125800.00000000001 123400.0 ;
      RECT  129799.99999999999 122600.00000000001 130600.0 123400.0 ;
      RECT  134600.0 122600.00000000001 135400.0 123400.0 ;
      RECT  139399.99999999997 122600.00000000001 140200.0 123400.0 ;
      RECT  144200.0 122600.00000000001 145000.0 123400.0 ;
      RECT  149000.0 122600.00000000001 149800.0 123400.0 ;
      RECT  153800.0 122600.00000000001 154600.00000000003 123400.0 ;
      RECT  158600.0 122600.00000000001 159400.0 123400.0 ;
      RECT  163399.99999999997 122600.00000000001 164200.0 123400.0 ;
      RECT  168200.0 122600.00000000001 169000.0 123400.0 ;
      RECT  173000.0 122600.00000000001 173800.0 123400.0 ;
      RECT  177800.0 122600.00000000001 178600.00000000003 123400.0 ;
      RECT  182600.0 122600.00000000001 183400.0 123400.0 ;
      RECT  187399.99999999997 122600.00000000001 188200.0 123400.0 ;
      RECT  192200.0 122600.00000000001 193000.0 123400.0 ;
      RECT  197000.0 122600.00000000001 197800.0 123400.0 ;
      RECT  201800.0 122600.00000000001 202600.00000000003 123400.0 ;
      RECT  206600.0 122600.00000000001 207400.0 123400.0 ;
      RECT  4999.999999999997 127400.0 5799.999999999997 128199.99999999999 ;
      RECT  9799.999999999993 127400.0 10599.999999999995 128199.99999999999 ;
      RECT  14599.999999999998 127400.0 15399.999999999998 128199.99999999999 ;
      RECT  19399.999999999996 127400.0 20199.999999999996 128199.99999999999 ;
      RECT  24200.0 127400.0 25000.0 128199.99999999999 ;
      RECT  28999.999999999996 127400.0 29799.999999999996 128199.99999999999 ;
      RECT  33800.0 127400.0 34599.99999999999 128199.99999999999 ;
      RECT  38600.0 127400.0 39400.0 128199.99999999999 ;
      RECT  43400.00000000001 127400.0 44200.0 128199.99999999999 ;
      RECT  48200.0 127400.0 49000.0 128199.99999999999 ;
      RECT  53000.0 127400.0 53800.0 128199.99999999999 ;
      RECT  57800.0 127400.0 58599.99999999999 128199.99999999999 ;
      RECT  62600.0 127400.0 63400.0 128199.99999999999 ;
      RECT  67400.0 127400.0 68200.0 128199.99999999999 ;
      RECT  72200.0 127400.0 73000.0 128199.99999999999 ;
      RECT  77000.0 127400.0 77800.0 128199.99999999999 ;
      RECT  81800.0 127400.0 82600.0 128199.99999999999 ;
      RECT  86600.00000000001 127400.0 87400.0 128199.99999999999 ;
      RECT  91400.0 127400.0 92200.0 128199.99999999999 ;
      RECT  96200.0 127400.0 97000.0 128199.99999999999 ;
      RECT  101000.0 127400.0 101800.0 128199.99999999999 ;
      RECT  105800.0 127400.0 106600.0 128199.99999999999 ;
      RECT  110600.00000000001 127400.0 111400.0 128199.99999999999 ;
      RECT  115400.0 127400.0 116200.0 128199.99999999999 ;
      RECT  120200.0 127400.0 121000.0 128199.99999999999 ;
      RECT  125000.00000000001 127400.0 125800.00000000001 128199.99999999999 ;
      RECT  129799.99999999999 127400.0 130600.0 128199.99999999999 ;
      RECT  134600.0 127400.0 135400.0 128199.99999999999 ;
      RECT  139399.99999999997 127400.0 140200.0 128199.99999999999 ;
      RECT  144200.0 127400.0 145000.0 128199.99999999999 ;
      RECT  149000.0 127400.0 149800.0 128199.99999999999 ;
      RECT  153800.0 127400.0 154600.00000000003 128199.99999999999 ;
      RECT  158600.0 127400.0 159400.0 128199.99999999999 ;
      RECT  163399.99999999997 127400.0 164200.0 128199.99999999999 ;
      RECT  168200.0 127400.0 169000.0 128199.99999999999 ;
      RECT  173000.0 127400.0 173800.0 128199.99999999999 ;
      RECT  177800.0 127400.0 178600.00000000003 128199.99999999999 ;
      RECT  182600.0 127400.0 183400.0 128199.99999999999 ;
      RECT  187399.99999999997 127400.0 188200.0 128199.99999999999 ;
      RECT  192200.0 127400.0 193000.0 128199.99999999999 ;
      RECT  197000.0 127400.0 197800.0 128199.99999999999 ;
      RECT  201800.0 127400.0 202600.00000000003 128199.99999999999 ;
      RECT  206600.0 127400.0 207400.0 128199.99999999999 ;
      RECT  4999.999999999997 132200.0 5799.999999999997 133000.0 ;
      RECT  9799.999999999993 132200.0 10599.999999999995 133000.0 ;
      RECT  14599.999999999998 132200.0 15399.999999999998 133000.0 ;
      RECT  19399.999999999996 132200.0 20199.999999999996 133000.0 ;
      RECT  24200.0 132200.0 25000.0 133000.0 ;
      RECT  28999.999999999996 132200.0 29799.999999999996 133000.0 ;
      RECT  33800.0 132200.0 34599.99999999999 133000.0 ;
      RECT  38600.0 132200.0 39400.0 133000.0 ;
      RECT  43400.00000000001 132200.0 44200.0 133000.0 ;
      RECT  48200.0 132200.0 49000.0 133000.0 ;
      RECT  53000.0 132200.0 53800.0 133000.0 ;
      RECT  57800.0 132200.0 58599.99999999999 133000.0 ;
      RECT  62600.0 132200.0 63400.0 133000.0 ;
      RECT  67400.0 132200.0 68200.0 133000.0 ;
      RECT  72200.0 132200.0 73000.0 133000.0 ;
      RECT  77000.0 132200.0 77800.0 133000.0 ;
      RECT  81800.0 132200.0 82600.0 133000.0 ;
      RECT  86600.00000000001 132200.0 87400.0 133000.0 ;
      RECT  91400.0 132200.0 92200.0 133000.0 ;
      RECT  96200.0 132200.0 97000.0 133000.0 ;
      RECT  101000.0 132200.0 101800.0 133000.0 ;
      RECT  105800.0 132200.0 106600.0 133000.0 ;
      RECT  110600.00000000001 132200.0 111400.0 133000.0 ;
      RECT  115400.0 132200.0 116200.0 133000.0 ;
      RECT  120200.0 132200.0 121000.0 133000.0 ;
      RECT  125000.00000000001 132200.0 125800.00000000001 133000.0 ;
      RECT  129799.99999999999 132200.0 130600.0 133000.0 ;
      RECT  134600.0 132200.0 135400.0 133000.0 ;
      RECT  139399.99999999997 132200.0 140200.0 133000.0 ;
      RECT  144200.0 132200.0 145000.0 133000.0 ;
      RECT  149000.0 132200.0 149800.0 133000.0 ;
      RECT  153800.0 132200.0 154600.00000000003 133000.0 ;
      RECT  158600.0 132200.0 159400.0 133000.0 ;
      RECT  163399.99999999997 132200.0 164200.0 133000.0 ;
      RECT  168200.0 132200.0 169000.0 133000.0 ;
      RECT  173000.0 132200.0 173800.0 133000.0 ;
      RECT  177800.0 132200.0 178600.00000000003 133000.0 ;
      RECT  182600.0 132200.0 183400.0 133000.0 ;
      RECT  187399.99999999997 132200.0 188200.0 133000.0 ;
      RECT  192200.0 132200.0 193000.0 133000.0 ;
      RECT  197000.0 132200.0 197800.0 133000.0 ;
      RECT  201800.0 132200.0 202600.00000000003 133000.0 ;
      RECT  206600.0 132200.0 207400.0 133000.0 ;
      RECT  4999.999999999997 137000.0 5799.999999999997 137800.0 ;
      RECT  9799.999999999993 137000.0 10599.999999999995 137800.0 ;
      RECT  14599.999999999998 137000.0 15399.999999999998 137800.0 ;
      RECT  19399.999999999996 137000.0 20199.999999999996 137800.0 ;
      RECT  24200.0 137000.0 25000.0 137800.0 ;
      RECT  28999.999999999996 137000.0 29799.999999999996 137800.0 ;
      RECT  33800.0 137000.0 34599.99999999999 137800.0 ;
      RECT  38600.0 137000.0 39400.0 137800.0 ;
      RECT  43400.00000000001 137000.0 44200.0 137800.0 ;
      RECT  48200.0 137000.0 49000.0 137800.0 ;
      RECT  53000.0 137000.0 53800.0 137800.0 ;
      RECT  57800.0 137000.0 58599.99999999999 137800.0 ;
      RECT  62600.0 137000.0 63400.0 137800.0 ;
      RECT  67400.0 137000.0 68200.0 137800.0 ;
      RECT  72200.0 137000.0 73000.0 137800.0 ;
      RECT  77000.0 137000.0 77800.0 137800.0 ;
      RECT  81800.0 137000.0 82600.0 137800.0 ;
      RECT  86600.00000000001 137000.0 87400.0 137800.0 ;
      RECT  91400.0 137000.0 92200.0 137800.0 ;
      RECT  96200.0 137000.0 97000.0 137800.0 ;
      RECT  101000.0 137000.0 101800.0 137800.0 ;
      RECT  105800.0 137000.0 106600.0 137800.0 ;
      RECT  110600.00000000001 137000.0 111400.0 137800.0 ;
      RECT  115400.0 137000.0 116200.0 137800.0 ;
      RECT  120200.0 137000.0 121000.0 137800.0 ;
      RECT  125000.00000000001 137000.0 125800.00000000001 137800.0 ;
      RECT  129799.99999999999 137000.0 130600.0 137800.0 ;
      RECT  134600.0 137000.0 135400.0 137800.0 ;
      RECT  139399.99999999997 137000.0 140200.0 137800.0 ;
      RECT  144200.0 137000.0 145000.0 137800.0 ;
      RECT  149000.0 137000.0 149800.0 137800.0 ;
      RECT  153800.0 137000.0 154600.00000000003 137800.0 ;
      RECT  158600.0 137000.0 159400.0 137800.0 ;
      RECT  163399.99999999997 137000.0 164200.0 137800.0 ;
      RECT  168200.0 137000.0 169000.0 137800.0 ;
      RECT  173000.0 137000.0 173800.0 137800.0 ;
      RECT  177800.0 137000.0 178600.00000000003 137800.0 ;
      RECT  182600.0 137000.0 183400.0 137800.0 ;
      RECT  187399.99999999997 137000.0 188200.0 137800.0 ;
      RECT  192200.0 137000.0 193000.0 137800.0 ;
      RECT  197000.0 137000.0 197800.0 137800.0 ;
      RECT  201800.0 137000.0 202600.00000000003 137800.0 ;
      RECT  206600.0 137000.0 207400.0 137800.0 ;
      RECT  4999.999999999997 141800.0 5799.999999999997 142600.00000000003 ;
      RECT  9799.999999999993 141800.0 10599.999999999995 142600.00000000003 ;
      RECT  14599.999999999998 141800.0 15399.999999999998 142600.00000000003 ;
      RECT  19399.999999999996 141800.0 20199.999999999996 142600.00000000003 ;
      RECT  24200.0 141800.0 25000.0 142600.00000000003 ;
      RECT  28999.999999999996 141800.0 29799.999999999996 142600.00000000003 ;
      RECT  33800.0 141800.0 34599.99999999999 142600.00000000003 ;
      RECT  38600.0 141800.0 39400.0 142600.00000000003 ;
      RECT  43400.00000000001 141800.0 44200.0 142600.00000000003 ;
      RECT  48200.0 141800.0 49000.0 142600.00000000003 ;
      RECT  53000.0 141800.0 53800.0 142600.00000000003 ;
      RECT  57800.0 141800.0 58599.99999999999 142600.00000000003 ;
      RECT  62600.0 141800.0 63400.0 142600.00000000003 ;
      RECT  67400.0 141800.0 68200.0 142600.00000000003 ;
      RECT  72200.0 141800.0 73000.0 142600.00000000003 ;
      RECT  77000.0 141800.0 77800.0 142600.00000000003 ;
      RECT  81800.0 141800.0 82600.0 142600.00000000003 ;
      RECT  86600.00000000001 141800.0 87400.0 142600.00000000003 ;
      RECT  91400.0 141800.0 92200.0 142600.00000000003 ;
      RECT  96200.0 141800.0 97000.0 142600.00000000003 ;
      RECT  101000.0 141800.0 101800.0 142600.00000000003 ;
      RECT  105800.0 141800.0 106600.0 142600.00000000003 ;
      RECT  110600.00000000001 141800.0 111400.0 142600.00000000003 ;
      RECT  115400.0 141800.0 116200.0 142600.00000000003 ;
      RECT  120200.0 141800.0 121000.0 142600.00000000003 ;
      RECT  125000.00000000001 141800.0 125800.00000000001 142600.00000000003 ;
      RECT  129799.99999999999 141800.0 130600.0 142600.00000000003 ;
      RECT  134600.0 141800.0 135400.0 142600.00000000003 ;
      RECT  139399.99999999997 141800.0 140200.0 142600.00000000003 ;
      RECT  144200.0 141800.0 145000.0 142600.00000000003 ;
      RECT  149000.0 141800.0 149800.0 142600.00000000003 ;
      RECT  153800.0 141800.0 154600.00000000003 142600.00000000003 ;
      RECT  158600.0 141800.0 159400.0 142600.00000000003 ;
      RECT  163399.99999999997 141800.0 164200.0 142600.00000000003 ;
      RECT  168200.0 141800.0 169000.0 142600.00000000003 ;
      RECT  4999.999999999997 146600.0 5799.999999999997 147400.0 ;
      RECT  9799.999999999993 146600.0 10599.999999999995 147400.0 ;
      RECT  14599.999999999998 146600.0 15399.999999999998 147400.0 ;
      RECT  19399.999999999996 146600.0 20199.999999999996 147400.0 ;
      RECT  24200.0 146600.0 25000.0 147400.0 ;
      RECT  28999.999999999996 146600.0 29799.999999999996 147400.0 ;
      RECT  33800.0 146600.0 34599.99999999999 147400.0 ;
      RECT  38600.0 146600.0 39400.0 147400.0 ;
      RECT  43400.00000000001 146600.0 44200.0 147400.0 ;
      RECT  48200.0 146600.0 49000.0 147400.0 ;
      RECT  53000.0 146600.0 53800.0 147400.0 ;
      RECT  57800.0 146600.0 58599.99999999999 147400.0 ;
      RECT  62600.0 146600.0 63400.0 147400.0 ;
      RECT  67400.0 146600.0 68200.0 147400.0 ;
      RECT  72200.0 146600.0 73000.0 147400.0 ;
      RECT  77000.0 146600.0 77800.0 147400.0 ;
      RECT  81800.0 146600.0 82600.0 147400.0 ;
      RECT  86600.00000000001 146600.0 87400.0 147400.0 ;
      RECT  91400.0 146600.0 92200.0 147400.0 ;
      RECT  96200.0 146600.0 97000.0 147400.0 ;
      RECT  101000.0 146600.0 101800.0 147400.0 ;
      RECT  105800.0 146600.0 106600.0 147400.0 ;
      RECT  110600.00000000001 146600.0 111400.0 147400.0 ;
      RECT  115400.0 146600.0 116200.0 147400.0 ;
      RECT  120200.0 146600.0 121000.0 147400.0 ;
      RECT  125000.00000000001 146600.0 125800.00000000001 147400.0 ;
      RECT  129799.99999999999 146600.0 130600.0 147400.0 ;
      RECT  134600.0 146600.0 135400.0 147400.0 ;
      RECT  139399.99999999997 146600.0 140200.0 147400.0 ;
      RECT  144200.0 146600.0 145000.0 147400.0 ;
      RECT  149000.0 146600.0 149800.0 147400.0 ;
      RECT  153800.0 146600.0 154600.00000000003 147400.0 ;
      RECT  158600.0 146600.0 159400.0 147400.0 ;
      RECT  163399.99999999997 146600.0 164200.0 147400.0 ;
      RECT  168200.0 146600.0 169000.0 147400.0 ;
      RECT  173000.0 146600.0 173800.0 147400.0 ;
      RECT  177800.0 146600.0 178600.00000000003 147400.0 ;
      RECT  182600.0 146600.0 183400.0 147400.0 ;
      RECT  187399.99999999997 146600.0 188200.0 147400.0 ;
      RECT  192200.0 146600.0 193000.0 147400.0 ;
      RECT  197000.0 146600.0 197800.0 147400.0 ;
      RECT  201800.0 146600.0 202600.00000000003 147400.0 ;
      RECT  206600.0 146600.0 207400.0 147400.0 ;
      RECT  4999.999999999997 151399.99999999997 5799.999999999997 152200.0 ;
      RECT  9799.999999999993 151399.99999999997 10599.999999999995 152200.0 ;
      RECT  14599.999999999998 151399.99999999997 15399.999999999998 152200.0 ;
      RECT  19399.999999999996 151399.99999999997 20199.999999999996 152200.0 ;
      RECT  24200.0 151399.99999999997 25000.0 152200.0 ;
      RECT  28999.999999999996 151399.99999999997 29799.999999999996 152200.0 ;
      RECT  33800.0 151399.99999999997 34599.99999999999 152200.0 ;
      RECT  38600.0 151399.99999999997 39400.0 152200.0 ;
      RECT  43400.00000000001 151399.99999999997 44200.0 152200.0 ;
      RECT  48200.0 151399.99999999997 49000.0 152200.0 ;
      RECT  53000.0 151399.99999999997 53800.0 152200.0 ;
      RECT  57800.0 151399.99999999997 58599.99999999999 152200.0 ;
      RECT  62600.0 151399.99999999997 63400.0 152200.0 ;
      RECT  177800.0 151399.99999999997 178600.00000000003 152200.0 ;
      RECT  182600.0 151399.99999999997 183400.0 152200.0 ;
      RECT  187399.99999999997 151399.99999999997 188200.0 152200.0 ;
      RECT  192200.0 151399.99999999997 193000.0 152200.0 ;
      RECT  197000.0 151399.99999999997 197800.0 152200.0 ;
      RECT  201800.0 151399.99999999997 202600.00000000003 152200.0 ;
      RECT  206600.0 151399.99999999997 207400.0 152200.0 ;
      RECT  4999.999999999997 156200.0 5799.999999999997 157000.0 ;
      RECT  9799.999999999993 156200.0 10599.999999999995 157000.0 ;
      RECT  14599.999999999998 156200.0 15399.999999999998 157000.0 ;
      RECT  19399.999999999996 156200.0 20199.999999999996 157000.0 ;
      RECT  24200.0 156200.0 25000.0 157000.0 ;
      RECT  28999.999999999996 156200.0 29799.999999999996 157000.0 ;
      RECT  33800.0 156200.0 34599.99999999999 157000.0 ;
      RECT  38600.0 156200.0 39400.0 157000.0 ;
      RECT  43400.00000000001 156200.0 44200.0 157000.0 ;
      RECT  48200.0 156200.0 49000.0 157000.0 ;
      RECT  53000.0 156200.0 53800.0 157000.0 ;
      RECT  57800.0 156200.0 58599.99999999999 157000.0 ;
      RECT  62600.0 156200.0 63400.0 157000.0 ;
      RECT  67400.0 156200.0 68200.0 157000.0 ;
      RECT  72200.0 156200.0 73000.0 157000.0 ;
      RECT  77000.0 156200.0 77800.0 157000.0 ;
      RECT  81800.0 156200.0 82600.0 157000.0 ;
      RECT  86600.00000000001 156200.0 87400.0 157000.0 ;
      RECT  91400.0 156200.0 92200.0 157000.0 ;
      RECT  96200.0 156200.0 97000.0 157000.0 ;
      RECT  101000.0 156200.0 101800.0 157000.0 ;
      RECT  105800.0 156200.0 106600.0 157000.0 ;
      RECT  110600.00000000001 156200.0 111400.0 157000.0 ;
      RECT  115400.0 156200.0 116200.0 157000.0 ;
      RECT  120200.0 156200.0 121000.0 157000.0 ;
      RECT  125000.00000000001 156200.0 125800.00000000001 157000.0 ;
      RECT  129799.99999999999 156200.0 130600.0 157000.0 ;
      RECT  134600.0 156200.0 135400.0 157000.0 ;
      RECT  139399.99999999997 156200.0 140200.0 157000.0 ;
      RECT  144200.0 156200.0 145000.0 157000.0 ;
      RECT  149000.0 156200.0 149800.0 157000.0 ;
      RECT  153800.0 156200.0 154600.00000000003 157000.0 ;
      RECT  158600.0 156200.0 159400.0 157000.0 ;
      RECT  163399.99999999997 156200.0 164200.0 157000.0 ;
      RECT  168200.0 156200.0 169000.0 157000.0 ;
      RECT  173000.0 156200.0 173800.0 157000.0 ;
      RECT  177800.0 156200.0 178600.00000000003 157000.0 ;
      RECT  182600.0 156200.0 183400.0 157000.0 ;
      RECT  187399.99999999997 156200.0 188200.0 157000.0 ;
      RECT  192200.0 156200.0 193000.0 157000.0 ;
      RECT  197000.0 156200.0 197800.0 157000.0 ;
      RECT  201800.0 156200.0 202600.00000000003 157000.0 ;
      RECT  206600.0 156200.0 207400.0 157000.0 ;
      RECT  4999.999999999997 161000.0 5799.999999999997 161800.0 ;
      RECT  9799.999999999993 161000.0 10599.999999999995 161800.0 ;
      RECT  14599.999999999998 161000.0 15399.999999999998 161800.0 ;
      RECT  19399.999999999996 161000.0 20199.999999999996 161800.0 ;
      RECT  24200.0 161000.0 25000.0 161800.0 ;
      RECT  28999.999999999996 161000.0 29799.999999999996 161800.0 ;
      RECT  33800.0 161000.0 34599.99999999999 161800.0 ;
      RECT  38600.0 161000.0 39400.0 161800.0 ;
      RECT  43400.00000000001 161000.0 44200.0 161800.0 ;
      RECT  48200.0 161000.0 49000.0 161800.0 ;
      RECT  53000.0 161000.0 53800.0 161800.0 ;
      RECT  57800.0 161000.0 58599.99999999999 161800.0 ;
      RECT  62600.0 161000.0 63400.0 161800.0 ;
      RECT  77000.0 161000.0 77800.0 161800.0 ;
      RECT  81800.0 161000.0 82600.0 161800.0 ;
      RECT  86600.00000000001 161000.0 87400.0 161800.0 ;
      RECT  91400.0 161000.0 92200.0 161800.0 ;
      RECT  96200.0 161000.0 97000.0 161800.0 ;
      RECT  101000.0 161000.0 101800.0 161800.0 ;
      RECT  105800.0 161000.0 106600.0 161800.0 ;
      RECT  110600.00000000001 161000.0 111400.0 161800.0 ;
      RECT  115400.0 161000.0 116200.0 161800.0 ;
      RECT  120200.0 161000.0 121000.0 161800.0 ;
      RECT  125000.00000000001 161000.0 125800.00000000001 161800.0 ;
      RECT  129799.99999999999 161000.0 130600.0 161800.0 ;
      RECT  134600.0 161000.0 135400.0 161800.0 ;
      RECT  139399.99999999997 161000.0 140200.0 161800.0 ;
      RECT  144200.0 161000.0 145000.0 161800.0 ;
      RECT  149000.0 161000.0 149800.0 161800.0 ;
      RECT  153800.0 161000.0 154600.00000000003 161800.0 ;
      RECT  158600.0 161000.0 159400.0 161800.0 ;
      RECT  163399.99999999997 161000.0 164200.0 161800.0 ;
      RECT  168200.0 161000.0 169000.0 161800.0 ;
      RECT  173000.0 161000.0 173800.0 161800.0 ;
      RECT  177800.0 161000.0 178600.00000000003 161800.0 ;
      RECT  182600.0 161000.0 183400.0 161800.0 ;
      RECT  187399.99999999997 161000.0 188200.0 161800.0 ;
      RECT  192200.0 161000.0 193000.0 161800.0 ;
      RECT  197000.0 161000.0 197800.0 161800.0 ;
      RECT  201800.0 161000.0 202600.00000000003 161800.0 ;
      RECT  206600.0 161000.0 207400.0 161800.0 ;
      RECT  4999.999999999997 165800.0 5799.999999999997 166600.00000000003 ;
      RECT  9799.999999999993 165800.0 10599.999999999995 166600.00000000003 ;
      RECT  14599.999999999998 165800.0 15399.999999999998 166600.00000000003 ;
      RECT  19399.999999999996 165800.0 20199.999999999996 166600.00000000003 ;
      RECT  24200.0 165800.0 25000.0 166600.00000000003 ;
      RECT  28999.999999999996 165800.0 29799.999999999996 166600.00000000003 ;
      RECT  33800.0 165800.0 34599.99999999999 166600.00000000003 ;
      RECT  38600.0 165800.0 39400.0 166600.00000000003 ;
      RECT  43400.00000000001 165800.0 44200.0 166600.00000000003 ;
      RECT  48200.0 165800.0 49000.0 166600.00000000003 ;
      RECT  53000.0 165800.0 53800.0 166600.00000000003 ;
      RECT  57800.0 165800.0 58599.99999999999 166600.00000000003 ;
      RECT  62600.0 165800.0 63400.0 166600.00000000003 ;
      RECT  67400.0 165800.0 68200.0 166600.00000000003 ;
      RECT  72200.0 165800.0 73000.0 166600.00000000003 ;
      RECT  77000.0 165800.0 77800.0 166600.00000000003 ;
      RECT  81800.0 165800.0 82600.0 166600.00000000003 ;
      RECT  86600.00000000001 165800.0 87400.0 166600.00000000003 ;
      RECT  91400.0 165800.0 92200.0 166600.00000000003 ;
      RECT  96200.0 165800.0 97000.0 166600.00000000003 ;
      RECT  101000.0 165800.0 101800.0 166600.00000000003 ;
      RECT  105800.0 165800.0 106600.0 166600.00000000003 ;
      RECT  110600.00000000001 165800.0 111400.0 166600.00000000003 ;
      RECT  115400.0 165800.0 116200.0 166600.00000000003 ;
      RECT  120200.0 165800.0 121000.0 166600.00000000003 ;
      RECT  125000.00000000001 165800.0 125800.00000000001 166600.00000000003 ;
      RECT  129799.99999999999 165800.0 130600.0 166600.00000000003 ;
      RECT  134600.0 165800.0 135400.0 166600.00000000003 ;
      RECT  139399.99999999997 165800.0 140200.0 166600.00000000003 ;
      RECT  144200.0 165800.0 145000.0 166600.00000000003 ;
      RECT  149000.0 165800.0 149800.0 166600.00000000003 ;
      RECT  153800.0 165800.0 154600.00000000003 166600.00000000003 ;
      RECT  158600.0 165800.0 159400.0 166600.00000000003 ;
      RECT  163399.99999999997 165800.0 164200.0 166600.00000000003 ;
      RECT  168200.0 165800.0 169000.0 166600.00000000003 ;
      RECT  173000.0 165800.0 173800.0 166600.00000000003 ;
      RECT  177800.0 165800.0 178600.00000000003 166600.00000000003 ;
      RECT  182600.0 165800.0 183400.0 166600.00000000003 ;
      RECT  187399.99999999997 165800.0 188200.0 166600.00000000003 ;
      RECT  192200.0 165800.0 193000.0 166600.00000000003 ;
      RECT  197000.0 165800.0 197800.0 166600.00000000003 ;
      RECT  201800.0 165800.0 202600.00000000003 166600.00000000003 ;
      RECT  206600.0 165800.0 207400.0 166600.00000000003 ;
      RECT  43400.00000000001 170600.0 44200.0 171400.0 ;
      RECT  48200.0 170600.0 49000.0 171400.0 ;
      RECT  53000.0 170600.0 53800.0 171400.0 ;
      RECT  57800.0 170600.0 58599.99999999999 171400.0 ;
      RECT  62600.0 170600.0 63400.0 171400.0 ;
      RECT  67400.0 170600.0 68200.0 171400.0 ;
      RECT  72200.0 170600.0 73000.0 171400.0 ;
      RECT  77000.0 170600.0 77800.0 171400.0 ;
      RECT  81800.0 170600.0 82600.0 171400.0 ;
      RECT  48200.0 175399.99999999997 49000.0 176200.0 ;
      RECT  53000.0 175399.99999999997 53800.0 176200.0 ;
      RECT  57800.0 175399.99999999997 58599.99999999999 176200.0 ;
      RECT  62600.0 175399.99999999997 63400.0 176200.0 ;
      RECT  67400.0 175399.99999999997 68200.0 176200.0 ;
      RECT  72200.0 175399.99999999997 73000.0 176200.0 ;
      RECT  77000.0 175399.99999999997 77800.0 176200.0 ;
      RECT  81800.0 175399.99999999997 82600.0 176200.0 ;
      RECT  86600.00000000001 175399.99999999997 87400.0 176200.0 ;
      RECT  91400.0 175399.99999999997 92200.0 176200.0 ;
      RECT  96200.0 175399.99999999997 97000.0 176200.0 ;
      RECT  101000.0 175399.99999999997 101800.0 176200.0 ;
      RECT  105800.0 175399.99999999997 106600.0 176200.0 ;
      RECT  110600.00000000001 175399.99999999997 111400.0 176200.0 ;
      RECT  115400.0 175399.99999999997 116200.0 176200.0 ;
      RECT  120200.0 175399.99999999997 121000.0 176200.0 ;
      RECT  125000.00000000001 175399.99999999997 125800.00000000001 176200.0 ;
      RECT  129799.99999999999 175399.99999999997 130600.0 176200.0 ;
      RECT  134600.0 175399.99999999997 135400.0 176200.0 ;
      RECT  139399.99999999997 175399.99999999997 140200.0 176200.0 ;
      RECT  144200.0 175399.99999999997 145000.0 176200.0 ;
      RECT  149000.0 175399.99999999997 149800.0 176200.0 ;
      RECT  153800.0 175399.99999999997 154600.00000000003 176200.0 ;
      RECT  158600.0 175399.99999999997 159400.0 176200.0 ;
      RECT  163399.99999999997 175399.99999999997 164200.0 176200.0 ;
      RECT  168200.0 175399.99999999997 169000.0 176200.0 ;
      RECT  173000.0 175399.99999999997 173800.0 176200.0 ;
      RECT  177800.0 175399.99999999997 178600.00000000003 176200.0 ;
      RECT  182600.0 175399.99999999997 183400.0 176200.0 ;
      RECT  187399.99999999997 175399.99999999997 188200.0 176200.0 ;
      RECT  192200.0 175399.99999999997 193000.0 176200.0 ;
      RECT  197000.0 175399.99999999997 197800.0 176200.0 ;
      RECT  201800.0 175399.99999999997 202600.00000000003 176200.0 ;
      RECT  206600.0 175399.99999999997 207400.0 176200.0 ;
      RECT  43400.00000000001 180200.0 44200.0 181000.0 ;
      RECT  48200.0 180200.0 49000.0 181000.0 ;
      RECT  53000.0 180200.0 53800.0 181000.0 ;
      RECT  57800.0 180200.0 58599.99999999999 181000.0 ;
      RECT  62600.0 180200.0 63400.0 181000.0 ;
      RECT  67400.0 180200.0 68200.0 181000.0 ;
      RECT  91400.0 180200.0 92200.0 181000.0 ;
      RECT  96200.0 180200.0 97000.0 181000.0 ;
      RECT  101000.0 180200.0 101800.0 181000.0 ;
      RECT  105800.0 180200.0 106600.0 181000.0 ;
      RECT  110600.00000000001 180200.0 111400.0 181000.0 ;
      RECT  115400.0 180200.0 116200.0 181000.0 ;
      RECT  120200.0 180200.0 121000.0 181000.0 ;
      RECT  125000.00000000001 180200.0 125800.00000000001 181000.0 ;
      RECT  129799.99999999999 180200.0 130600.0 181000.0 ;
      RECT  134600.0 180200.0 135400.0 181000.0 ;
      RECT  139399.99999999997 180200.0 140200.0 181000.0 ;
      RECT  144200.0 180200.0 145000.0 181000.0 ;
      RECT  149000.0 180200.0 149800.0 181000.0 ;
      RECT  153800.0 180200.0 154600.00000000003 181000.0 ;
      RECT  158600.0 180200.0 159400.0 181000.0 ;
      RECT  163399.99999999997 180200.0 164200.0 181000.0 ;
      RECT  4999.999999999997 185000.0 5799.999999999997 185800.0 ;
      RECT  9799.999999999993 185000.0 10599.999999999995 185800.0 ;
      RECT  14599.999999999998 185000.0 15399.999999999998 185800.0 ;
      RECT  19399.999999999996 185000.0 20199.999999999996 185800.0 ;
      RECT  24200.0 185000.0 25000.0 185800.0 ;
      RECT  28999.999999999996 185000.0 29799.999999999996 185800.0 ;
      RECT  33800.0 185000.0 34599.99999999999 185800.0 ;
      RECT  38600.0 185000.0 39400.0 185800.0 ;
      RECT  43400.00000000001 185000.0 44200.0 185800.0 ;
      RECT  48200.0 185000.0 49000.0 185800.0 ;
      RECT  53000.0 185000.0 53800.0 185800.0 ;
      RECT  57800.0 185000.0 58599.99999999999 185800.0 ;
      RECT  62600.0 185000.0 63400.0 185800.0 ;
      RECT  67400.0 185000.0 68200.0 185800.0 ;
      RECT  72200.0 185000.0 73000.0 185800.0 ;
      RECT  77000.0 185000.0 77800.0 185800.0 ;
      RECT  81800.0 185000.0 82600.0 185800.0 ;
      RECT  168200.0 185000.0 169000.0 185800.0 ;
      RECT  173000.0 185000.0 173800.0 185800.0 ;
      RECT  177800.0 185000.0 178600.00000000003 185800.0 ;
      RECT  182600.0 185000.0 183400.0 185800.0 ;
      RECT  187399.99999999997 185000.0 188200.0 185800.0 ;
      RECT  192200.0 185000.0 193000.0 185800.0 ;
      RECT  197000.0 185000.0 197800.0 185800.0 ;
      RECT  201800.0 185000.0 202600.00000000003 185800.0 ;
      RECT  206600.0 185000.0 207400.0 185800.0 ;
      RECT  43400.00000000001 189800.0 44200.0 190600.00000000003 ;
      RECT  48200.0 189800.0 49000.0 190600.00000000003 ;
      RECT  53000.0 189800.0 53800.0 190600.00000000003 ;
      RECT  57800.0 189800.0 58599.99999999999 190600.00000000003 ;
      RECT  62600.0 189800.0 63400.0 190600.00000000003 ;
      RECT  67400.0 189800.0 68200.0 190600.00000000003 ;
      RECT  91400.0 189800.0 92200.0 190600.00000000003 ;
      RECT  96200.0 189800.0 97000.0 190600.00000000003 ;
      RECT  101000.0 189800.0 101800.0 190600.00000000003 ;
      RECT  105800.0 189800.0 106600.0 190600.00000000003 ;
      RECT  110600.00000000001 189800.0 111400.0 190600.00000000003 ;
      RECT  115400.0 189800.0 116200.0 190600.00000000003 ;
      RECT  120200.0 189800.0 121000.0 190600.00000000003 ;
      RECT  125000.00000000001 189800.0 125800.00000000001 190600.00000000003 ;
      RECT  129799.99999999999 189800.0 130600.0 190600.00000000003 ;
      RECT  134600.0 189800.0 135400.0 190600.00000000003 ;
      RECT  139399.99999999997 189800.0 140200.0 190600.00000000003 ;
      RECT  144200.0 189800.0 145000.0 190600.00000000003 ;
      RECT  149000.0 189800.0 149800.0 190600.00000000003 ;
      RECT  153800.0 189800.0 154600.00000000003 190600.00000000003 ;
      RECT  158600.0 189800.0 159400.0 190600.00000000003 ;
      RECT  163399.99999999997 189800.0 164200.0 190600.00000000003 ;
      RECT  48200.0 194600.0 49000.0 195400.0 ;
      RECT  53000.0 194600.0 53800.0 195400.0 ;
      RECT  57800.0 194600.0 58599.99999999999 195400.0 ;
      RECT  62600.0 194600.0 63400.0 195400.0 ;
      RECT  67400.0 194600.0 68200.0 195400.0 ;
      RECT  72200.0 194600.0 73000.0 195400.0 ;
      RECT  77000.0 194600.0 77800.0 195400.0 ;
      RECT  81800.0 194600.0 82600.0 195400.0 ;
      RECT  86600.00000000001 194600.0 87400.0 195400.0 ;
      RECT  91400.0 194600.0 92200.0 195400.0 ;
      RECT  96200.0 194600.0 97000.0 195400.0 ;
      RECT  101000.0 194600.0 101800.0 195400.0 ;
      RECT  105800.0 194600.0 106600.0 195400.0 ;
      RECT  129799.99999999999 194600.0 130600.0 195400.0 ;
      RECT  134600.0 194600.0 135400.0 195400.0 ;
      RECT  139399.99999999997 194600.0 140200.0 195400.0 ;
      RECT  144200.0 194600.0 145000.0 195400.0 ;
      RECT  149000.0 194600.0 149800.0 195400.0 ;
      RECT  153800.0 194600.0 154600.00000000003 195400.0 ;
      RECT  158600.0 194600.0 159400.0 195400.0 ;
      RECT  163399.99999999997 194600.0 164200.0 195400.0 ;
      RECT  168200.0 194600.0 169000.0 195400.0 ;
      RECT  173000.0 194600.0 173800.0 195400.0 ;
      RECT  177800.0 194600.0 178600.00000000003 195400.0 ;
      RECT  182600.0 194600.0 183400.0 195400.0 ;
      RECT  187399.99999999997 194600.0 188200.0 195400.0 ;
      RECT  192200.0 194600.0 193000.0 195400.0 ;
      RECT  197000.0 194600.0 197800.0 195400.0 ;
      RECT  201800.0 194600.0 202600.00000000003 195400.0 ;
      RECT  206600.0 194600.0 207400.0 195400.0 ;
      RECT  43400.00000000001 199399.99999999997 44200.0 200200.0 ;
      RECT  48200.0 199399.99999999997 49000.0 200200.0 ;
      RECT  53000.0 199399.99999999997 53800.0 200200.0 ;
      RECT  57800.0 199399.99999999997 58599.99999999999 200200.0 ;
      RECT  62600.0 199399.99999999997 63400.0 200200.0 ;
      RECT  67400.0 199399.99999999997 68200.0 200200.0 ;
      RECT  72200.0 199399.99999999997 73000.0 200200.0 ;
      RECT  77000.0 199399.99999999997 77800.0 200200.0 ;
      RECT  81800.0 199399.99999999997 82600.0 200200.0 ;
      RECT  86600.00000000001 199399.99999999997 87400.0 200200.0 ;
      RECT  91400.0 199399.99999999997 92200.0 200200.0 ;
      RECT  96200.0 199399.99999999997 97000.0 200200.0 ;
      RECT  101000.0 199399.99999999997 101800.0 200200.0 ;
      RECT  105800.0 199399.99999999997 106600.0 200200.0 ;
      RECT  110600.00000000001 199399.99999999997 111400.0 200200.0 ;
      RECT  115400.0 199399.99999999997 116200.0 200200.0 ;
      RECT  120200.0 199399.99999999997 121000.0 200200.0 ;
      RECT  125000.00000000001 199399.99999999997 125800.00000000001 200200.0 ;
      RECT  129799.99999999999 199399.99999999997 130600.0 200200.0 ;
      RECT  134600.0 199399.99999999997 135400.0 200200.0 ;
      RECT  139399.99999999997 199399.99999999997 140200.0 200200.0 ;
      RECT  144200.0 199399.99999999997 145000.0 200200.0 ;
      RECT  149000.0 199399.99999999997 149800.0 200200.0 ;
      RECT  153800.0 199399.99999999997 154600.00000000003 200200.0 ;
      RECT  158600.0 199399.99999999997 159400.0 200200.0 ;
      RECT  163399.99999999997 199399.99999999997 164200.0 200200.0 ;
      RECT  4999.999999999997 204200.0 5799.999999999997 205000.0 ;
      RECT  9799.999999999993 204200.0 10599.999999999995 205000.0 ;
      RECT  14599.999999999998 204200.0 15399.999999999998 205000.0 ;
      RECT  19399.999999999996 204200.0 20199.999999999996 205000.0 ;
      RECT  24200.0 204200.0 25000.0 205000.0 ;
      RECT  28999.999999999996 204200.0 29799.999999999996 205000.0 ;
      RECT  33800.0 204200.0 34599.99999999999 205000.0 ;
      RECT  38600.0 204200.0 39400.0 205000.0 ;
      RECT  43400.00000000001 204200.0 44200.0 205000.0 ;
      RECT  48200.0 204200.0 49000.0 205000.0 ;
      RECT  53000.0 204200.0 53800.0 205000.0 ;
      RECT  57800.0 204200.0 58599.99999999999 205000.0 ;
      RECT  62600.0 204200.0 63400.0 205000.0 ;
      RECT  67400.0 204200.0 68200.0 205000.0 ;
      RECT  72200.0 204200.0 73000.0 205000.0 ;
      RECT  77000.0 204200.0 77800.0 205000.0 ;
      RECT  81800.0 204200.0 82600.0 205000.0 ;
      RECT  168200.0 204200.0 169000.0 205000.0 ;
      RECT  173000.0 204200.0 173800.0 205000.0 ;
      RECT  177800.0 204200.0 178600.00000000003 205000.0 ;
      RECT  182600.0 204200.0 183400.0 205000.0 ;
      RECT  187399.99999999997 204200.0 188200.0 205000.0 ;
      RECT  192200.0 204200.0 193000.0 205000.0 ;
      RECT  197000.0 204200.0 197800.0 205000.0 ;
      RECT  201800.0 204200.0 202600.00000000003 205000.0 ;
      RECT  206600.0 204200.0 207400.0 205000.0 ;
      RECT  48200.0 209000.0 49000.0 209800.0 ;
      RECT  53000.0 209000.0 53800.0 209800.0 ;
      RECT  57800.0 209000.0 58599.99999999999 209800.0 ;
      RECT  62600.0 209000.0 63400.0 209800.0 ;
      RECT  67400.0 209000.0 68200.0 209800.0 ;
      RECT  72200.0 209000.0 73000.0 209800.0 ;
      RECT  77000.0 209000.0 77800.0 209800.0 ;
      RECT  81800.0 209000.0 82600.0 209800.0 ;
      RECT  86600.00000000001 209000.0 87400.0 209800.0 ;
      RECT  91400.0 209000.0 92200.0 209800.0 ;
      RECT  96200.0 209000.0 97000.0 209800.0 ;
      RECT  101000.0 209000.0 101800.0 209800.0 ;
      RECT  105800.0 209000.0 106600.0 209800.0 ;
      RECT  110600.00000000001 209000.0 111400.0 209800.0 ;
      RECT  115400.0 209000.0 116200.0 209800.0 ;
      RECT  120200.0 209000.0 121000.0 209800.0 ;
      RECT  125000.00000000001 209000.0 125800.00000000001 209800.0 ;
      RECT  129799.99999999999 209000.0 130600.0 209800.0 ;
      RECT  134600.0 209000.0 135400.0 209800.0 ;
      RECT  139399.99999999997 209000.0 140200.0 209800.0 ;
      RECT  144200.0 209000.0 145000.0 209800.0 ;
      RECT  149000.0 209000.0 149800.0 209800.0 ;
      RECT  153800.0 209000.0 154600.00000000003 209800.0 ;
      RECT  158600.0 209000.0 159400.0 209800.0 ;
      RECT  163399.99999999997 209000.0 164200.0 209800.0 ;
      RECT  48200.0 213800.0 49000.0 214600.00000000003 ;
      RECT  53000.0 213800.0 53800.0 214600.00000000003 ;
      RECT  57800.0 213800.0 58599.99999999999 214600.00000000003 ;
      RECT  62600.0 213800.0 63400.0 214600.00000000003 ;
      RECT  67400.0 213800.0 68200.0 214600.00000000003 ;
      RECT  129799.99999999999 213800.0 130600.0 214600.00000000003 ;
      RECT  134600.0 213800.0 135400.0 214600.00000000003 ;
      RECT  139399.99999999997 213800.0 140200.0 214600.00000000003 ;
      RECT  144200.0 213800.0 145000.0 214600.00000000003 ;
      RECT  149000.0 213800.0 149800.0 214600.00000000003 ;
      RECT  153800.0 213800.0 154600.00000000003 214600.00000000003 ;
      RECT  158600.0 213800.0 159400.0 214600.00000000003 ;
      RECT  163399.99999999997 213800.0 164200.0 214600.00000000003 ;
      RECT  168200.0 213800.0 169000.0 214600.00000000003 ;
      RECT  173000.0 213800.0 173800.0 214600.00000000003 ;
      RECT  177800.0 213800.0 178600.00000000003 214600.00000000003 ;
      RECT  182600.0 213800.0 183400.0 214600.00000000003 ;
      RECT  187399.99999999997 213800.0 188200.0 214600.00000000003 ;
      RECT  192200.0 213800.0 193000.0 214600.00000000003 ;
      RECT  197000.0 213800.0 197800.0 214600.00000000003 ;
      RECT  201800.0 213800.0 202600.00000000003 214600.00000000003 ;
      RECT  206600.0 213800.0 207400.0 214600.00000000003 ;
      RECT  43400.00000000001 218600.00000000003 44200.0 219400.00000000003 ;
      RECT  48200.0 218600.00000000003 49000.0 219400.00000000003 ;
      RECT  53000.0 218600.00000000003 53800.0 219400.00000000003 ;
      RECT  57800.0 218600.00000000003 58599.99999999999 219400.00000000003 ;
      RECT  62600.0 218600.00000000003 63400.0 219400.00000000003 ;
      RECT  67400.0 218600.00000000003 68200.0 219400.00000000003 ;
      RECT  72200.0 218600.00000000003 73000.0 219400.00000000003 ;
      RECT  77000.0 218600.00000000003 77800.0 219400.00000000003 ;
      RECT  81800.0 218600.00000000003 82600.0 219400.00000000003 ;
      RECT  86600.00000000001 218600.00000000003 87400.0 219400.00000000003 ;
      RECT  91400.0 218600.00000000003 92200.0 219400.00000000003 ;
      RECT  96200.0 218600.00000000003 97000.0 219400.00000000003 ;
      RECT  101000.0 218600.00000000003 101800.0 219400.00000000003 ;
      RECT  105800.0 218600.00000000003 106600.0 219400.00000000003 ;
      RECT  110600.00000000001 218600.00000000003 111400.0 219400.00000000003 ;
      RECT  115400.0 218600.00000000003 116200.0 219400.00000000003 ;
      RECT  120200.0 218600.00000000003 121000.0 219400.00000000003 ;
      RECT  125000.00000000001 218600.00000000003 125800.00000000001 219400.00000000003 ;
      RECT  129799.99999999999 218600.00000000003 130600.0 219400.00000000003 ;
      RECT  134600.0 218600.00000000003 135400.0 219400.00000000003 ;
      RECT  139399.99999999997 218600.00000000003 140200.0 219400.00000000003 ;
      RECT  144200.0 218600.00000000003 145000.0 219400.00000000003 ;
      RECT  149000.0 218600.00000000003 149800.0 219400.00000000003 ;
      RECT  153800.0 218600.00000000003 154600.00000000003 219400.00000000003 ;
      RECT  158600.0 218600.00000000003 159400.0 219400.00000000003 ;
      RECT  163399.99999999997 218600.00000000003 164200.0 219400.00000000003 ;
      RECT  4999.999999999997 223399.99999999997 5799.999999999997 224200.0 ;
      RECT  9799.999999999993 223399.99999999997 10599.999999999995 224200.0 ;
      RECT  14599.999999999998 223399.99999999997 15399.999999999998 224200.0 ;
      RECT  19399.999999999996 223399.99999999997 20199.999999999996 224200.0 ;
      RECT  24200.0 223399.99999999997 25000.0 224200.0 ;
      RECT  28999.999999999996 223399.99999999997 29799.999999999996 224200.0 ;
      RECT  33800.0 223399.99999999997 34599.99999999999 224200.0 ;
      RECT  38600.0 223399.99999999997 39400.0 224200.0 ;
      RECT  43400.00000000001 223399.99999999997 44200.0 224200.0 ;
      RECT  48200.0 223399.99999999997 49000.0 224200.0 ;
      RECT  53000.0 223399.99999999997 53800.0 224200.0 ;
      RECT  57800.0 223399.99999999997 58599.99999999999 224200.0 ;
      RECT  62600.0 223399.99999999997 63400.0 224200.0 ;
      RECT  67400.0 223399.99999999997 68200.0 224200.0 ;
      RECT  72200.0 223399.99999999997 73000.0 224200.0 ;
      RECT  168200.0 223399.99999999997 169000.0 224200.0 ;
      RECT  173000.0 223399.99999999997 173800.0 224200.0 ;
      RECT  177800.0 223399.99999999997 178600.00000000003 224200.0 ;
      RECT  182600.0 223399.99999999997 183400.0 224200.0 ;
      RECT  187399.99999999997 223399.99999999997 188200.0 224200.0 ;
      RECT  192200.0 223399.99999999997 193000.0 224200.0 ;
      RECT  197000.0 223399.99999999997 197800.0 224200.0 ;
      RECT  201800.0 223399.99999999997 202600.00000000003 224200.0 ;
      RECT  206600.0 223399.99999999997 207400.0 224200.0 ;
      RECT  4999.999999999997 228200.0 5799.999999999997 229000.0 ;
      RECT  9799.999999999993 228200.0 10599.999999999995 229000.0 ;
      RECT  14599.999999999998 228200.0 15399.999999999998 229000.0 ;
      RECT  19399.999999999996 228200.0 20199.999999999996 229000.0 ;
      RECT  24200.0 228200.0 25000.0 229000.0 ;
      RECT  28999.999999999996 228200.0 29799.999999999996 229000.0 ;
      RECT  48200.0 228200.0 49000.0 229000.0 ;
      RECT  53000.0 228200.0 53800.0 229000.0 ;
      RECT  57800.0 228200.0 58599.99999999999 229000.0 ;
      RECT  62600.0 228200.0 63400.0 229000.0 ;
      RECT  67400.0 228200.0 68200.0 229000.0 ;
      RECT  72200.0 228200.0 73000.0 229000.0 ;
      RECT  77000.0 228200.0 77800.0 229000.0 ;
      RECT  81800.0 228200.0 82600.0 229000.0 ;
      RECT  86600.00000000001 228200.0 87400.0 229000.0 ;
      RECT  91400.0 228200.0 92200.0 229000.0 ;
      RECT  96200.0 228200.0 97000.0 229000.0 ;
      RECT  101000.0 228200.0 101800.0 229000.0 ;
      RECT  105800.0 228200.0 106600.0 229000.0 ;
      RECT  110600.00000000001 228200.0 111400.0 229000.0 ;
      RECT  115400.0 228200.0 116200.0 229000.0 ;
      RECT  120200.0 228200.0 121000.0 229000.0 ;
      RECT  125000.00000000001 228200.0 125800.00000000001 229000.0 ;
      RECT  129799.99999999999 228200.0 130600.0 229000.0 ;
      RECT  134600.0 228200.0 135400.0 229000.0 ;
      RECT  139399.99999999997 228200.0 140200.0 229000.0 ;
      RECT  144200.0 228200.0 145000.0 229000.0 ;
      RECT  149000.0 228200.0 149800.0 229000.0 ;
      RECT  153800.0 228200.0 154600.00000000003 229000.0 ;
      RECT  158600.0 228200.0 159400.0 229000.0 ;
      RECT  163399.99999999997 228200.0 164200.0 229000.0 ;
      RECT  48200.0 233000.0 49000.0 233800.0 ;
      RECT  53000.0 233000.0 53800.0 233800.0 ;
      RECT  57800.0 233000.0 58599.99999999999 233800.0 ;
      RECT  62600.0 233000.0 63400.0 233800.0 ;
      RECT  67400.0 233000.0 68200.0 233800.0 ;
      RECT  72200.0 233000.0 73000.0 233800.0 ;
      RECT  77000.0 233000.0 77800.0 233800.0 ;
      RECT  81800.0 233000.0 82600.0 233800.0 ;
      RECT  86600.00000000001 233000.0 87400.0 233800.0 ;
      RECT  91400.0 233000.0 92200.0 233800.0 ;
      RECT  96200.0 233000.0 97000.0 233800.0 ;
      RECT  101000.0 233000.0 101800.0 233800.0 ;
      RECT  105800.0 233000.0 106600.0 233800.0 ;
      RECT  134600.0 233000.0 135400.0 233800.0 ;
      RECT  139399.99999999997 233000.0 140200.0 233800.0 ;
      RECT  144200.0 233000.0 145000.0 233800.0 ;
      RECT  149000.0 233000.0 149800.0 233800.0 ;
      RECT  153800.0 233000.0 154600.00000000003 233800.0 ;
      RECT  158600.0 233000.0 159400.0 233800.0 ;
      RECT  163399.99999999997 233000.0 164200.0 233800.0 ;
      RECT  168200.0 233000.0 169000.0 233800.0 ;
      RECT  173000.0 233000.0 173800.0 233800.0 ;
      RECT  177800.0 233000.0 178600.00000000003 233800.0 ;
      RECT  182600.0 233000.0 183400.0 233800.0 ;
      RECT  187399.99999999997 233000.0 188200.0 233800.0 ;
      RECT  192200.0 233000.0 193000.0 233800.0 ;
      RECT  197000.0 233000.0 197800.0 233800.0 ;
      RECT  201800.0 233000.0 202600.00000000003 233800.0 ;
      RECT  206600.0 233000.0 207400.0 233800.0 ;
      RECT  4999.999999999997 237800.0 5799.999999999997 238600.00000000003 ;
      RECT  9799.999999999993 237800.0 10599.999999999995 238600.00000000003 ;
      RECT  14599.999999999998 237800.0 15399.999999999998 238600.00000000003 ;
      RECT  19399.999999999996 237800.0 20199.999999999996 238600.00000000003 ;
      RECT  24200.0 237800.0 25000.0 238600.00000000003 ;
      RECT  28999.999999999996 237800.0 29799.999999999996 238600.00000000003 ;
      RECT  33800.0 237800.0 34599.99999999999 238600.00000000003 ;
      RECT  38600.0 237800.0 39400.0 238600.00000000003 ;
      RECT  43400.00000000001 237800.0 44200.0 238600.00000000003 ;
      RECT  48200.0 237800.0 49000.0 238600.00000000003 ;
      RECT  53000.0 237800.0 53800.0 238600.00000000003 ;
      RECT  57800.0 237800.0 58599.99999999999 238600.00000000003 ;
      RECT  62600.0 237800.0 63400.0 238600.00000000003 ;
      RECT  67400.0 237800.0 68200.0 238600.00000000003 ;
      RECT  72200.0 237800.0 73000.0 238600.00000000003 ;
      RECT  77000.0 237800.0 77800.0 238600.00000000003 ;
      RECT  81800.0 237800.0 82600.0 238600.00000000003 ;
      RECT  86600.00000000001 237800.0 87400.0 238600.00000000003 ;
      RECT  91400.0 237800.0 92200.0 238600.00000000003 ;
      RECT  96200.0 237800.0 97000.0 238600.00000000003 ;
      RECT  101000.0 237800.0 101800.0 238600.00000000003 ;
      RECT  105800.0 237800.0 106600.0 238600.00000000003 ;
      RECT  110600.00000000001 237800.0 111400.0 238600.00000000003 ;
      RECT  115400.0 237800.0 116200.0 238600.00000000003 ;
      RECT  120200.0 237800.0 121000.0 238600.00000000003 ;
      RECT  125000.00000000001 237800.0 125800.00000000001 238600.00000000003 ;
      RECT  129799.99999999999 237800.0 130600.0 238600.00000000003 ;
      RECT  134600.0 237800.0 135400.0 238600.00000000003 ;
      RECT  139399.99999999997 237800.0 140200.0 238600.00000000003 ;
      RECT  144200.0 237800.0 145000.0 238600.00000000003 ;
      RECT  149000.0 237800.0 149800.0 238600.00000000003 ;
      RECT  153800.0 237800.0 154600.00000000003 238600.00000000003 ;
      RECT  158600.0 237800.0 159400.0 238600.00000000003 ;
      RECT  163399.99999999997 237800.0 164200.0 238600.00000000003 ;
      RECT  43400.00000000001 242600.00000000003 44200.0 243400.00000000003 ;
      RECT  48200.0 242600.00000000003 49000.0 243400.00000000003 ;
      RECT  53000.0 242600.00000000003 53800.0 243400.00000000003 ;
      RECT  57800.0 242600.00000000003 58599.99999999999 243400.00000000003 ;
      RECT  62600.0 242600.00000000003 63400.0 243400.00000000003 ;
      RECT  67400.0 242600.00000000003 68200.0 243400.00000000003 ;
      RECT  72200.0 242600.00000000003 73000.0 243400.00000000003 ;
      RECT  77000.0 242600.00000000003 77800.0 243400.00000000003 ;
      RECT  81800.0 242600.00000000003 82600.0 243400.00000000003 ;
      RECT  168200.0 242600.00000000003 169000.0 243400.00000000003 ;
      RECT  173000.0 242600.00000000003 173800.0 243400.00000000003 ;
      RECT  177800.0 242600.00000000003 178600.00000000003 243400.00000000003 ;
      RECT  182600.0 242600.00000000003 183400.0 243400.00000000003 ;
      RECT  187399.99999999997 242600.00000000003 188200.0 243400.00000000003 ;
      RECT  192200.0 242600.00000000003 193000.0 243400.00000000003 ;
      RECT  197000.0 242600.00000000003 197800.0 243400.00000000003 ;
      RECT  201800.0 242600.00000000003 202600.00000000003 243400.00000000003 ;
      RECT  206600.0 242600.00000000003 207400.0 243400.00000000003 ;
      RECT  4999.999999999997 247399.99999999997 5799.999999999997 248200.0 ;
      RECT  9799.999999999993 247399.99999999997 10599.999999999995 248200.0 ;
      RECT  14599.999999999998 247399.99999999997 15399.999999999998 248200.0 ;
      RECT  19399.999999999996 247399.99999999997 20199.999999999996 248200.0 ;
      RECT  24200.0 247399.99999999997 25000.0 248200.0 ;
      RECT  28999.999999999996 247399.99999999997 29799.999999999996 248200.0 ;
      RECT  48200.0 247399.99999999997 49000.0 248200.0 ;
      RECT  53000.0 247399.99999999997 53800.0 248200.0 ;
      RECT  57800.0 247399.99999999997 58599.99999999999 248200.0 ;
      RECT  62600.0 247399.99999999997 63400.0 248200.0 ;
      RECT  67400.0 247399.99999999997 68200.0 248200.0 ;
      RECT  72200.0 247399.99999999997 73000.0 248200.0 ;
      RECT  77000.0 247399.99999999997 77800.0 248200.0 ;
      RECT  81800.0 247399.99999999997 82600.0 248200.0 ;
      RECT  86600.00000000001 247399.99999999997 87400.0 248200.0 ;
      RECT  91400.0 247399.99999999997 92200.0 248200.0 ;
      RECT  96200.0 247399.99999999997 97000.0 248200.0 ;
      RECT  101000.0 247399.99999999997 101800.0 248200.0 ;
      RECT  105800.0 247399.99999999997 106600.0 248200.0 ;
      RECT  110600.00000000001 247399.99999999997 111400.0 248200.0 ;
      RECT  115400.0 247399.99999999997 116200.0 248200.0 ;
      RECT  120200.0 247399.99999999997 121000.0 248200.0 ;
      RECT  125000.00000000001 247399.99999999997 125800.00000000001 248200.0 ;
      RECT  129799.99999999999 247399.99999999997 130600.0 248200.0 ;
      RECT  134600.0 247399.99999999997 135400.0 248200.0 ;
      RECT  139399.99999999997 247399.99999999997 140200.0 248200.0 ;
      RECT  144200.0 247399.99999999997 145000.0 248200.0 ;
      RECT  149000.0 247399.99999999997 149800.0 248200.0 ;
      RECT  153800.0 247399.99999999997 154600.00000000003 248200.0 ;
      RECT  158600.0 247399.99999999997 159400.0 248200.0 ;
      RECT  163399.99999999997 247399.99999999997 164200.0 248200.0 ;
      RECT  4999.999999999997 252200.0 5799.999999999997 253000.0 ;
      RECT  9799.999999999993 252200.0 10599.999999999995 253000.0 ;
      RECT  14599.999999999998 252200.0 15399.999999999998 253000.0 ;
      RECT  19399.999999999996 252200.0 20199.999999999996 253000.0 ;
      RECT  24200.0 252200.0 25000.0 253000.0 ;
      RECT  28999.999999999996 252200.0 29799.999999999996 253000.0 ;
      RECT  33800.0 252200.0 34599.99999999999 253000.0 ;
      RECT  38600.0 252200.0 39400.0 253000.0 ;
      RECT  43400.00000000001 252200.0 44200.0 253000.0 ;
      RECT  48200.0 252200.0 49000.0 253000.0 ;
      RECT  53000.0 252200.0 53800.0 253000.0 ;
      RECT  57800.0 252200.0 58599.99999999999 253000.0 ;
      RECT  62600.0 252200.0 63400.0 253000.0 ;
      RECT  67400.0 252200.0 68200.0 253000.0 ;
      RECT  72200.0 252200.0 73000.0 253000.0 ;
      RECT  77000.0 252200.0 77800.0 253000.0 ;
      RECT  81800.0 252200.0 82600.0 253000.0 ;
      RECT  86600.00000000001 252200.0 87400.0 253000.0 ;
      RECT  91400.0 252200.0 92200.0 253000.0 ;
      RECT  96200.0 252200.0 97000.0 253000.0 ;
      RECT  101000.0 252200.0 101800.0 253000.0 ;
      RECT  105800.0 252200.0 106600.0 253000.0 ;
      RECT  110600.00000000001 252200.0 111400.0 253000.0 ;
      RECT  115400.0 252200.0 116200.0 253000.0 ;
      RECT  120200.0 252200.0 121000.0 253000.0 ;
      RECT  125000.00000000001 252200.0 125800.00000000001 253000.0 ;
      RECT  129799.99999999999 252200.0 130600.0 253000.0 ;
      RECT  134600.0 252200.0 135400.0 253000.0 ;
      RECT  139399.99999999997 252200.0 140200.0 253000.0 ;
      RECT  144200.0 252200.0 145000.0 253000.0 ;
      RECT  149000.0 252200.0 149800.0 253000.0 ;
      RECT  153800.0 252200.0 154600.00000000003 253000.0 ;
      RECT  158600.0 252200.0 159400.0 253000.0 ;
      RECT  163399.99999999997 252200.0 164200.0 253000.0 ;
      RECT  168200.0 252200.0 169000.0 253000.0 ;
      RECT  173000.0 252200.0 173800.0 253000.0 ;
      RECT  177800.0 252200.0 178600.00000000003 253000.0 ;
      RECT  182600.0 252200.0 183400.0 253000.0 ;
      RECT  187399.99999999997 252200.0 188200.0 253000.0 ;
      RECT  192200.0 252200.0 193000.0 253000.0 ;
      RECT  197000.0 252200.0 197800.0 253000.0 ;
      RECT  201800.0 252200.0 202600.00000000003 253000.0 ;
      RECT  206600.0 252200.0 207400.0 253000.0 ;
      RECT  4999.999999999997 257000.0 5799.999999999997 257800.0 ;
      RECT  9799.999999999993 257000.0 10599.999999999995 257800.0 ;
      RECT  14599.999999999998 257000.0 15399.999999999998 257800.0 ;
      RECT  19399.999999999996 257000.0 20199.999999999996 257800.0 ;
      RECT  24200.0 257000.0 25000.0 257800.0 ;
      RECT  28999.999999999996 257000.0 29799.999999999996 257800.0 ;
      RECT  33800.0 257000.0 34599.99999999999 257800.0 ;
      RECT  38600.0 257000.0 39400.0 257800.0 ;
      RECT  43400.00000000001 257000.0 44200.0 257800.0 ;
      RECT  48200.0 257000.0 49000.0 257800.0 ;
      RECT  53000.0 257000.0 53800.0 257800.0 ;
      RECT  67400.0 257000.0 68200.0 257800.0 ;
      RECT  72200.0 257000.0 73000.0 257800.0 ;
      RECT  77000.0 257000.0 77800.0 257800.0 ;
      RECT  81800.0 257000.0 82600.0 257800.0 ;
      RECT  86600.00000000001 257000.0 87400.0 257800.0 ;
      RECT  91400.0 257000.0 92200.0 257800.0 ;
      RECT  96200.0 257000.0 97000.0 257800.0 ;
      RECT  101000.0 257000.0 101800.0 257800.0 ;
      RECT  105800.0 257000.0 106600.0 257800.0 ;
      RECT  110600.00000000001 257000.0 111400.0 257800.0 ;
      RECT  115400.0 257000.0 116200.0 257800.0 ;
      RECT  120200.0 257000.0 121000.0 257800.0 ;
      RECT  125000.00000000001 257000.0 125800.00000000001 257800.0 ;
      RECT  129799.99999999999 257000.0 130600.0 257800.0 ;
      RECT  134600.0 257000.0 135400.0 257800.0 ;
      RECT  139399.99999999997 257000.0 140200.0 257800.0 ;
      RECT  144200.0 257000.0 145000.0 257800.0 ;
      RECT  149000.0 257000.0 149800.0 257800.0 ;
      RECT  153800.0 257000.0 154600.00000000003 257800.0 ;
      RECT  158600.0 257000.0 159400.0 257800.0 ;
      RECT  163399.99999999997 257000.0 164200.0 257800.0 ;
      RECT  4999.999999999997 261800.0 5799.999999999997 262600.0 ;
      RECT  9799.999999999993 261800.0 10599.999999999995 262600.0 ;
      RECT  14599.999999999998 261800.0 15399.999999999998 262600.0 ;
      RECT  19399.999999999996 261800.0 20199.999999999996 262600.0 ;
      RECT  24200.0 261800.0 25000.0 262600.0 ;
      RECT  28999.999999999996 261800.0 29799.999999999996 262600.0 ;
      RECT  33800.0 261800.0 34599.99999999999 262600.0 ;
      RECT  38600.0 261800.0 39400.0 262600.0 ;
      RECT  43400.00000000001 261800.0 44200.0 262600.0 ;
      RECT  81800.0 261800.0 82600.0 262600.0 ;
      RECT  86600.00000000001 261800.0 87400.0 262600.0 ;
      RECT  91400.0 261800.0 92200.0 262600.0 ;
      RECT  96200.0 261800.0 97000.0 262600.0 ;
      RECT  101000.0 261800.0 101800.0 262600.0 ;
      RECT  105800.0 261800.0 106600.0 262600.0 ;
      RECT  110600.00000000001 261800.0 111400.0 262600.0 ;
      RECT  115400.0 261800.0 116200.0 262600.0 ;
      RECT  120200.0 261800.0 121000.0 262600.0 ;
      RECT  168200.0 261800.0 169000.0 262600.0 ;
      RECT  173000.0 261800.0 173800.0 262600.0 ;
      RECT  177800.0 261800.0 178600.00000000003 262600.0 ;
      RECT  182600.0 261800.0 183400.0 262600.0 ;
      RECT  187399.99999999997 261800.0 188200.0 262600.0 ;
      RECT  192200.0 261800.0 193000.0 262600.0 ;
      RECT  197000.0 261800.0 197800.0 262600.0 ;
      RECT  201800.0 261800.0 202600.00000000003 262600.0 ;
      RECT  206600.0 261800.0 207400.0 262600.0 ;
      RECT  4999.999999999997 266600.0 5799.999999999997 267400.00000000006 ;
      RECT  9799.999999999993 266600.0 10599.999999999995 267400.00000000006 ;
      RECT  14599.999999999998 266600.0 15399.999999999998 267400.00000000006 ;
      RECT  19399.999999999996 266600.0 20199.999999999996 267400.00000000006 ;
      RECT  24200.0 266600.0 25000.0 267400.00000000006 ;
      RECT  28999.999999999996 266600.0 29799.999999999996 267400.00000000006 ;
      RECT  33800.0 266600.0 34599.99999999999 267400.00000000006 ;
      RECT  38600.0 266600.0 39400.0 267400.00000000006 ;
      RECT  43400.00000000001 266600.0 44200.0 267400.00000000006 ;
      RECT  48200.0 266600.0 49000.0 267400.00000000006 ;
      RECT  53000.0 266600.0 53800.0 267400.00000000006 ;
      RECT  57800.0 266600.0 58599.99999999999 267400.00000000006 ;
      RECT  81800.0 266600.0 82600.0 267400.00000000006 ;
      RECT  86600.00000000001 266600.0 87400.0 267400.00000000006 ;
      RECT  91400.0 266600.0 92200.0 267400.00000000006 ;
      RECT  96200.0 266600.0 97000.0 267400.00000000006 ;
      RECT  101000.0 266600.0 101800.0 267400.00000000006 ;
      RECT  105800.0 266600.0 106600.0 267400.00000000006 ;
      RECT  110600.00000000001 266600.0 111400.0 267400.00000000006 ;
      RECT  115400.0 266600.0 116200.0 267400.00000000006 ;
      RECT  120200.0 266600.0 121000.0 267400.00000000006 ;
      RECT  125000.00000000001 266600.0 125800.00000000001 267400.00000000006 ;
      RECT  129799.99999999999 266600.0 130600.0 267400.00000000006 ;
      RECT  134600.0 266600.0 135400.0 267400.00000000006 ;
      RECT  139399.99999999997 266600.0 140200.0 267400.00000000006 ;
      RECT  144200.0 266600.0 145000.0 267400.00000000006 ;
      RECT  149000.0 266600.0 149800.0 267400.00000000006 ;
      RECT  153800.0 266600.0 154600.00000000003 267400.00000000006 ;
      RECT  158600.0 266600.0 159400.0 267400.00000000006 ;
      RECT  163399.99999999997 266600.0 164200.0 267400.00000000006 ;
      RECT  4999.999999999997 271400.0 5799.999999999997 272200.0 ;
      RECT  9799.999999999993 271400.0 10599.999999999995 272200.0 ;
      RECT  14599.999999999998 271400.0 15399.999999999998 272200.0 ;
      RECT  19399.999999999996 271400.0 20199.999999999996 272200.0 ;
      RECT  24200.0 271400.0 25000.0 272200.0 ;
      RECT  28999.999999999996 271400.0 29799.999999999996 272200.0 ;
      RECT  33800.0 271400.0 34599.99999999999 272200.0 ;
      RECT  38600.0 271400.0 39400.0 272200.0 ;
      RECT  43400.00000000001 271400.0 44200.0 272200.0 ;
      RECT  48200.0 271400.0 49000.0 272200.0 ;
      RECT  53000.0 271400.0 53800.0 272200.0 ;
      RECT  57800.0 271400.0 58599.99999999999 272200.0 ;
      RECT  62600.0 271400.0 63400.0 272200.0 ;
      RECT  67400.0 271400.0 68200.0 272200.0 ;
      RECT  72200.0 271400.0 73000.0 272200.0 ;
      RECT  77000.0 271400.0 77800.0 272200.0 ;
      RECT  81800.0 271400.0 82600.0 272200.0 ;
      RECT  86600.00000000001 271400.0 87400.0 272200.0 ;
      RECT  91400.0 271400.0 92200.0 272200.0 ;
      RECT  96200.0 271400.0 97000.0 272200.0 ;
      RECT  101000.0 271400.0 101800.0 272200.0 ;
      RECT  105800.0 271400.0 106600.0 272200.0 ;
      RECT  110600.00000000001 271400.0 111400.0 272200.0 ;
      RECT  115400.0 271400.0 116200.0 272200.0 ;
      RECT  120200.0 271400.0 121000.0 272200.0 ;
      RECT  125000.00000000001 271400.0 125800.00000000001 272200.0 ;
      RECT  129799.99999999999 271400.0 130600.0 272200.0 ;
      RECT  134600.0 271400.0 135400.0 272200.0 ;
      RECT  139399.99999999997 271400.0 140200.0 272200.0 ;
      RECT  144200.0 271400.0 145000.0 272200.0 ;
      RECT  149000.0 271400.0 149800.0 272200.0 ;
      RECT  153800.0 271400.0 154600.00000000003 272200.0 ;
      RECT  158600.0 271400.0 159400.0 272200.0 ;
      RECT  163399.99999999997 271400.0 164200.0 272200.0 ;
      RECT  168200.0 271400.0 169000.0 272200.0 ;
      RECT  173000.0 271400.0 173800.0 272200.0 ;
      RECT  177800.0 271400.0 178600.00000000003 272200.0 ;
      RECT  182600.0 271400.0 183400.0 272200.0 ;
      RECT  187399.99999999997 271400.0 188200.0 272200.0 ;
      RECT  192200.0 271400.0 193000.0 272200.0 ;
      RECT  197000.0 271400.0 197800.0 272200.0 ;
      RECT  201800.0 271400.0 202600.00000000003 272200.0 ;
      RECT  206600.0 271400.0 207400.0 272200.0 ;
      RECT  4999.999999999997 276200.0 5799.999999999997 277000.0 ;
      RECT  9799.999999999993 276200.0 10599.999999999995 277000.0 ;
      RECT  14599.999999999998 276200.0 15399.999999999998 277000.0 ;
      RECT  19399.999999999996 276200.0 20199.999999999996 277000.0 ;
      RECT  24200.0 276200.0 25000.0 277000.0 ;
      RECT  28999.999999999996 276200.0 29799.999999999996 277000.0 ;
      RECT  33800.0 276200.0 34599.99999999999 277000.0 ;
      RECT  38600.0 276200.0 39400.0 277000.0 ;
      RECT  43400.00000000001 276200.0 44200.0 277000.0 ;
      RECT  48200.0 276200.0 49000.0 277000.0 ;
      RECT  53000.0 276200.0 53800.0 277000.0 ;
      RECT  57800.0 276200.0 58599.99999999999 277000.0 ;
      RECT  62600.0 276200.0 63400.0 277000.0 ;
      RECT  67400.0 276200.0 68200.0 277000.0 ;
      RECT  72200.0 276200.0 73000.0 277000.0 ;
      RECT  77000.0 276200.0 77800.0 277000.0 ;
      RECT  81800.0 276200.0 82600.0 277000.0 ;
      RECT  86600.00000000001 276200.0 87400.0 277000.0 ;
      RECT  91400.0 276200.0 92200.0 277000.0 ;
      RECT  96200.0 276200.0 97000.0 277000.0 ;
      RECT  101000.0 276200.0 101800.0 277000.0 ;
      RECT  105800.0 276200.0 106600.0 277000.0 ;
      RECT  110600.00000000001 276200.0 111400.0 277000.0 ;
      RECT  115400.0 276200.0 116200.0 277000.0 ;
      RECT  120200.0 276200.0 121000.0 277000.0 ;
      RECT  125000.00000000001 276200.0 125800.00000000001 277000.0 ;
      RECT  129799.99999999999 276200.0 130600.0 277000.0 ;
      RECT  134600.0 276200.0 135400.0 277000.0 ;
      RECT  139399.99999999997 276200.0 140200.0 277000.0 ;
      RECT  144200.0 276200.0 145000.0 277000.0 ;
      RECT  149000.0 276200.0 149800.0 277000.0 ;
      RECT  153800.0 276200.0 154600.00000000003 277000.0 ;
      RECT  158600.0 276200.0 159400.0 277000.0 ;
      RECT  163399.99999999997 276200.0 164200.0 277000.0 ;
      RECT  168200.0 276200.0 169000.0 277000.0 ;
      RECT  173000.0 276200.0 173800.0 277000.0 ;
      RECT  177800.0 276200.0 178600.00000000003 277000.0 ;
      RECT  182600.0 276200.0 183400.0 277000.0 ;
      RECT  187399.99999999997 276200.0 188200.0 277000.0 ;
      RECT  192200.0 276200.0 193000.0 277000.0 ;
      RECT  197000.0 276200.0 197800.0 277000.0 ;
      RECT  201800.0 276200.0 202600.00000000003 277000.0 ;
      RECT  206600.0 276200.0 207400.0 277000.0 ;
      RECT  4999.999999999997 281000.0 5799.999999999997 281800.0 ;
      RECT  9799.999999999993 281000.0 10599.999999999995 281800.0 ;
      RECT  14599.999999999998 281000.0 15399.999999999998 281800.0 ;
      RECT  19399.999999999996 281000.0 20199.999999999996 281800.0 ;
      RECT  24200.0 281000.0 25000.0 281800.0 ;
      RECT  28999.999999999996 281000.0 29799.999999999996 281800.0 ;
      RECT  33800.0 281000.0 34599.99999999999 281800.0 ;
      RECT  38600.0 281000.0 39400.0 281800.0 ;
      RECT  43400.00000000001 281000.0 44200.0 281800.0 ;
      RECT  48200.0 281000.0 49000.0 281800.0 ;
      RECT  53000.0 281000.0 53800.0 281800.0 ;
      RECT  57800.0 281000.0 58599.99999999999 281800.0 ;
      RECT  62600.0 281000.0 63400.0 281800.0 ;
      RECT  67400.0 281000.0 68200.0 281800.0 ;
      RECT  72200.0 281000.0 73000.0 281800.0 ;
      RECT  77000.0 281000.0 77800.0 281800.0 ;
      RECT  81800.0 281000.0 82600.0 281800.0 ;
      RECT  86600.00000000001 281000.0 87400.0 281800.0 ;
      RECT  91400.0 281000.0 92200.0 281800.0 ;
      RECT  96200.0 281000.0 97000.0 281800.0 ;
      RECT  101000.0 281000.0 101800.0 281800.0 ;
      RECT  105800.0 281000.0 106600.0 281800.0 ;
      RECT  110600.00000000001 281000.0 111400.0 281800.0 ;
      RECT  115400.0 281000.0 116200.0 281800.0 ;
      RECT  120200.0 281000.0 121000.0 281800.0 ;
      RECT  4999.999999999997 285800.0 5799.999999999997 286600.0 ;
      RECT  9799.999999999993 285800.0 10599.999999999995 286600.0 ;
      RECT  14599.999999999998 285800.0 15399.999999999998 286600.0 ;
      RECT  19399.999999999996 285800.0 20199.999999999996 286600.0 ;
      RECT  24200.0 285800.0 25000.0 286600.0 ;
      RECT  28999.999999999996 285800.0 29799.999999999996 286600.0 ;
      RECT  33800.0 285800.0 34599.99999999999 286600.0 ;
      RECT  38600.0 285800.0 39400.0 286600.0 ;
      RECT  43400.00000000001 285800.0 44200.0 286600.0 ;
      RECT  48200.0 285800.0 49000.0 286600.0 ;
      RECT  53000.0 285800.0 53800.0 286600.0 ;
      RECT  57800.0 285800.0 58599.99999999999 286600.0 ;
      RECT  86600.00000000001 285800.0 87400.0 286600.0 ;
      RECT  91400.0 285800.0 92200.0 286600.0 ;
      RECT  96200.0 285800.0 97000.0 286600.0 ;
      RECT  101000.0 285800.0 101800.0 286600.0 ;
      RECT  105800.0 285800.0 106600.0 286600.0 ;
      RECT  110600.00000000001 285800.0 111400.0 286600.0 ;
      RECT  115400.0 285800.0 116200.0 286600.0 ;
      RECT  120200.0 285800.0 121000.0 286600.0 ;
      RECT  125000.00000000001 285800.0 125800.00000000001 286600.0 ;
      RECT  129799.99999999999 285800.0 130600.0 286600.0 ;
      RECT  134600.0 285800.0 135400.0 286600.0 ;
      RECT  139399.99999999997 285800.0 140200.0 286600.0 ;
      RECT  144200.0 285800.0 145000.0 286600.0 ;
      RECT  149000.0 285800.0 149800.0 286600.0 ;
      RECT  153800.0 285800.0 154600.00000000003 286600.0 ;
      RECT  158600.0 285800.0 159400.0 286600.0 ;
      RECT  163399.99999999997 285800.0 164200.0 286600.0 ;
      RECT  168200.0 285800.0 169000.0 286600.0 ;
      RECT  173000.0 285800.0 173800.0 286600.0 ;
      RECT  177800.0 285800.0 178600.00000000003 286600.0 ;
      RECT  182600.0 285800.0 183400.0 286600.0 ;
      RECT  187399.99999999997 285800.0 188200.0 286600.0 ;
      RECT  192200.0 285800.0 193000.0 286600.0 ;
      RECT  197000.0 285800.0 197800.0 286600.0 ;
      RECT  201800.0 285800.0 202600.00000000003 286600.0 ;
      RECT  206600.0 285800.0 207400.0 286600.0 ;
      RECT  4999.999999999997 290600.0 5799.999999999997 291400.00000000006 ;
      RECT  9799.999999999993 290600.0 10599.999999999995 291400.00000000006 ;
      RECT  14599.999999999998 290600.0 15399.999999999998 291400.00000000006 ;
      RECT  19399.999999999996 290600.0 20199.999999999996 291400.00000000006 ;
      RECT  24200.0 290600.0 25000.0 291400.00000000006 ;
      RECT  28999.999999999996 290600.0 29799.999999999996 291400.00000000006 ;
      RECT  33800.0 290600.0 34599.99999999999 291400.00000000006 ;
      RECT  38600.0 290600.0 39400.0 291400.00000000006 ;
      RECT  43400.00000000001 290600.0 44200.0 291400.00000000006 ;
      RECT  48200.0 290600.0 49000.0 291400.00000000006 ;
      RECT  53000.0 290600.0 53800.0 291400.00000000006 ;
      RECT  57800.0 290600.0 58599.99999999999 291400.00000000006 ;
      RECT  62600.0 290600.0 63400.0 291400.00000000006 ;
      RECT  67400.0 290600.0 68200.0 291400.00000000006 ;
      RECT  72200.0 290600.0 73000.0 291400.00000000006 ;
      RECT  77000.0 290600.0 77800.0 291400.00000000006 ;
      RECT  81800.0 290600.0 82600.0 291400.00000000006 ;
      RECT  86600.00000000001 290600.0 87400.0 291400.00000000006 ;
      RECT  91400.0 290600.0 92200.0 291400.00000000006 ;
      RECT  96200.0 290600.0 97000.0 291400.00000000006 ;
      RECT  101000.0 290600.0 101800.0 291400.00000000006 ;
      RECT  105800.0 290600.0 106600.0 291400.00000000006 ;
      RECT  110600.00000000001 290600.0 111400.0 291400.00000000006 ;
      RECT  115400.0 290600.0 116200.0 291400.00000000006 ;
      RECT  120200.0 290600.0 121000.0 291400.00000000006 ;
      RECT  125000.00000000001 290600.0 125800.00000000001 291400.00000000006 ;
      RECT  129799.99999999999 290600.0 130600.0 291400.00000000006 ;
      RECT  134600.0 290600.0 135400.0 291400.00000000006 ;
      RECT  139399.99999999997 290600.0 140200.0 291400.00000000006 ;
      RECT  144200.0 290600.0 145000.0 291400.00000000006 ;
      RECT  149000.0 290600.0 149800.0 291400.00000000006 ;
      RECT  153800.0 290600.0 154600.00000000003 291400.00000000006 ;
      RECT  158600.0 290600.0 159400.0 291400.00000000006 ;
      RECT  163399.99999999997 290600.0 164200.0 291400.00000000006 ;
      RECT  4999.999999999997 295400.0 5799.999999999997 296200.0 ;
      RECT  9799.999999999993 295400.0 10599.999999999995 296200.0 ;
      RECT  14599.999999999998 295400.0 15399.999999999998 296200.0 ;
      RECT  19399.999999999996 295400.0 20199.999999999996 296200.0 ;
      RECT  24200.0 295400.0 25000.0 296200.0 ;
      RECT  28999.999999999996 295400.0 29799.999999999996 296200.0 ;
      RECT  33800.0 295400.0 34599.99999999999 296200.0 ;
      RECT  38600.0 295400.0 39400.0 296200.0 ;
      RECT  43400.00000000001 295400.0 44200.0 296200.0 ;
      RECT  48200.0 295400.0 49000.0 296200.0 ;
      RECT  53000.0 295400.0 53800.0 296200.0 ;
      RECT  67400.0 295400.0 68200.0 296200.0 ;
      RECT  72200.0 295400.0 73000.0 296200.0 ;
      RECT  77000.0 295400.0 77800.0 296200.0 ;
      RECT  81800.0 295400.0 82600.0 296200.0 ;
      RECT  86600.00000000001 295400.0 87400.0 296200.0 ;
      RECT  91400.0 295400.0 92200.0 296200.0 ;
      RECT  96200.0 295400.0 97000.0 296200.0 ;
      RECT  101000.0 295400.0 101800.0 296200.0 ;
      RECT  105800.0 295400.0 106600.0 296200.0 ;
      RECT  110600.00000000001 295400.0 111400.0 296200.0 ;
      RECT  115400.0 295400.0 116200.0 296200.0 ;
      RECT  120200.0 295400.0 121000.0 296200.0 ;
      RECT  168200.0 295400.0 169000.0 296200.0 ;
      RECT  173000.0 295400.0 173800.0 296200.0 ;
      RECT  177800.0 295400.0 178600.00000000003 296200.0 ;
      RECT  182600.0 295400.0 183400.0 296200.0 ;
      RECT  187399.99999999997 295400.0 188200.0 296200.0 ;
      RECT  192200.0 295400.0 193000.0 296200.0 ;
      RECT  197000.0 295400.0 197800.0 296200.0 ;
      RECT  201800.0 295400.0 202600.00000000003 296200.0 ;
      RECT  206600.0 295400.0 207400.0 296200.0 ;
      RECT  4999.999999999997 300200.0 5799.999999999997 301000.0 ;
      RECT  9799.999999999993 300200.0 10599.999999999995 301000.0 ;
      RECT  14599.999999999998 300200.0 15399.999999999998 301000.0 ;
      RECT  19399.999999999996 300200.0 20199.999999999996 301000.0 ;
      RECT  24200.0 300200.0 25000.0 301000.0 ;
      RECT  28999.999999999996 300200.0 29799.999999999996 301000.0 ;
      RECT  33800.0 300200.0 34599.99999999999 301000.0 ;
      RECT  38600.0 300200.0 39400.0 301000.0 ;
      RECT  43400.00000000001 300200.0 44200.0 301000.0 ;
      RECT  48200.0 300200.0 49000.0 301000.0 ;
      RECT  53000.0 300200.0 53800.0 301000.0 ;
      RECT  57800.0 300200.0 58599.99999999999 301000.0 ;
      RECT  62600.0 300200.0 63400.0 301000.0 ;
      RECT  67400.0 300200.0 68200.0 301000.0 ;
      RECT  72200.0 300200.0 73000.0 301000.0 ;
      RECT  77000.0 300200.0 77800.0 301000.0 ;
      RECT  81800.0 300200.0 82600.0 301000.0 ;
      RECT  86600.00000000001 300200.0 87400.0 301000.0 ;
      RECT  91400.0 300200.0 92200.0 301000.0 ;
      RECT  96200.0 300200.0 97000.0 301000.0 ;
      RECT  101000.0 300200.0 101800.0 301000.0 ;
      RECT  105800.0 300200.0 106600.0 301000.0 ;
      RECT  110600.00000000001 300200.0 111400.0 301000.0 ;
      RECT  115400.0 300200.0 116200.0 301000.0 ;
      RECT  120200.0 300200.0 121000.0 301000.0 ;
      RECT  125000.00000000001 300200.0 125800.00000000001 301000.0 ;
      RECT  129799.99999999999 300200.0 130600.0 301000.0 ;
      RECT  134600.0 300200.0 135400.0 301000.0 ;
      RECT  139399.99999999997 300200.0 140200.0 301000.0 ;
      RECT  144200.0 300200.0 145000.0 301000.0 ;
      RECT  149000.0 300200.0 149800.0 301000.0 ;
      RECT  153800.0 300200.0 154600.00000000003 301000.0 ;
      RECT  158600.0 300200.0 159400.0 301000.0 ;
      RECT  163399.99999999997 300200.0 164200.0 301000.0 ;
      RECT  4999.999999999997 305000.0 5799.999999999997 305800.0 ;
      RECT  9799.999999999993 305000.0 10599.999999999995 305800.0 ;
      RECT  14599.999999999998 305000.0 15399.999999999998 305800.0 ;
      RECT  19399.999999999996 305000.0 20199.999999999996 305800.0 ;
      RECT  24200.0 305000.0 25000.0 305800.0 ;
      RECT  28999.999999999996 305000.0 29799.999999999996 305800.0 ;
      RECT  33800.0 305000.0 34599.99999999999 305800.0 ;
      RECT  38600.0 305000.0 39400.0 305800.0 ;
      RECT  43400.00000000001 305000.0 44200.0 305800.0 ;
      RECT  48200.0 305000.0 49000.0 305800.0 ;
      RECT  53000.0 305000.0 53800.0 305800.0 ;
      RECT  57800.0 305000.0 58599.99999999999 305800.0 ;
      RECT  86600.00000000001 305000.0 87400.0 305800.0 ;
      RECT  91400.0 305000.0 92200.0 305800.0 ;
      RECT  96200.0 305000.0 97000.0 305800.0 ;
      RECT  101000.0 305000.0 101800.0 305800.0 ;
      RECT  105800.0 305000.0 106600.0 305800.0 ;
      RECT  110600.00000000001 305000.0 111400.0 305800.0 ;
      RECT  115400.0 305000.0 116200.0 305800.0 ;
      RECT  120200.0 305000.0 121000.0 305800.0 ;
      RECT  125000.00000000001 305000.0 125800.00000000001 305800.0 ;
      RECT  129799.99999999999 305000.0 130600.0 305800.0 ;
      RECT  134600.0 305000.0 135400.0 305800.0 ;
      RECT  139399.99999999997 305000.0 140200.0 305800.0 ;
      RECT  144200.0 305000.0 145000.0 305800.0 ;
      RECT  149000.0 305000.0 149800.0 305800.0 ;
      RECT  153800.0 305000.0 154600.00000000003 305800.0 ;
      RECT  158600.0 305000.0 159400.0 305800.0 ;
      RECT  163399.99999999997 305000.0 164200.0 305800.0 ;
      RECT  168200.0 305000.0 169000.0 305800.0 ;
      RECT  173000.0 305000.0 173800.0 305800.0 ;
      RECT  177800.0 305000.0 178600.00000000003 305800.0 ;
      RECT  182600.0 305000.0 183400.0 305800.0 ;
      RECT  187399.99999999997 305000.0 188200.0 305800.0 ;
      RECT  192200.0 305000.0 193000.0 305800.0 ;
      RECT  197000.0 305000.0 197800.0 305800.0 ;
      RECT  201800.0 305000.0 202600.00000000003 305800.0 ;
      RECT  206600.0 305000.0 207400.0 305800.0 ;
      RECT  4999.999999999997 309800.0 5799.999999999997 310600.0 ;
      RECT  9799.999999999993 309800.0 10599.999999999995 310600.0 ;
      RECT  14599.999999999998 309800.0 15399.999999999998 310600.0 ;
      RECT  19399.999999999996 309800.0 20199.999999999996 310600.0 ;
      RECT  24200.0 309800.0 25000.0 310600.0 ;
      RECT  28999.999999999996 309800.0 29799.999999999996 310600.0 ;
      RECT  33800.0 309800.0 34599.99999999999 310600.0 ;
      RECT  38600.0 309800.0 39400.0 310600.0 ;
      RECT  43400.00000000001 309800.0 44200.0 310600.0 ;
      RECT  48200.0 309800.0 49000.0 310600.0 ;
      RECT  53000.0 309800.0 53800.0 310600.0 ;
      RECT  57800.0 309800.0 58599.99999999999 310600.0 ;
      RECT  62600.0 309800.0 63400.0 310600.0 ;
      RECT  67400.0 309800.0 68200.0 310600.0 ;
      RECT  72200.0 309800.0 73000.0 310600.0 ;
      RECT  77000.0 309800.0 77800.0 310600.0 ;
      RECT  81800.0 309800.0 82600.0 310600.0 ;
      RECT  86600.00000000001 309800.0 87400.0 310600.0 ;
      RECT  91400.0 309800.0 92200.0 310600.0 ;
      RECT  96200.0 309800.0 97000.0 310600.0 ;
      RECT  101000.0 309800.0 101800.0 310600.0 ;
      RECT  105800.0 309800.0 106600.0 310600.0 ;
      RECT  110600.00000000001 309800.0 111400.0 310600.0 ;
      RECT  115400.0 309800.0 116200.0 310600.0 ;
      RECT  120200.0 309800.0 121000.0 310600.0 ;
      RECT  125000.00000000001 309800.0 125800.00000000001 310600.0 ;
      RECT  129799.99999999999 309800.0 130600.0 310600.0 ;
      RECT  134600.0 309800.0 135400.0 310600.0 ;
      RECT  139399.99999999997 309800.0 140200.0 310600.0 ;
      RECT  144200.0 309800.0 145000.0 310600.0 ;
      RECT  149000.0 309800.0 149800.0 310600.0 ;
      RECT  153800.0 309800.0 154600.00000000003 310600.0 ;
      RECT  158600.0 309800.0 159400.0 310600.0 ;
      RECT  163399.99999999997 309800.0 164200.0 310600.0 ;
      RECT  4999.999999999997 314600.0 5799.999999999997 315400.00000000006 ;
      RECT  9799.999999999993 314600.0 10599.999999999995 315400.00000000006 ;
      RECT  14599.999999999998 314600.0 15399.999999999998 315400.00000000006 ;
      RECT  19399.999999999996 314600.0 20199.999999999996 315400.00000000006 ;
      RECT  24200.0 314600.0 25000.0 315400.00000000006 ;
      RECT  28999.999999999996 314600.0 29799.999999999996 315400.00000000006 ;
      RECT  33800.0 314600.0 34599.99999999999 315400.00000000006 ;
      RECT  38600.0 314600.0 39400.0 315400.00000000006 ;
      RECT  43400.00000000001 314600.0 44200.0 315400.00000000006 ;
      RECT  48200.0 314600.0 49000.0 315400.00000000006 ;
      RECT  53000.0 314600.0 53800.0 315400.00000000006 ;
      RECT  57800.0 314600.0 58599.99999999999 315400.00000000006 ;
      RECT  62600.0 314600.0 63400.0 315400.00000000006 ;
      RECT  67400.0 314600.0 68200.0 315400.00000000006 ;
      RECT  72200.0 314600.0 73000.0 315400.00000000006 ;
      RECT  77000.0 314600.0 77800.0 315400.00000000006 ;
      RECT  81800.0 314600.0 82600.0 315400.00000000006 ;
      RECT  86600.00000000001 314600.0 87400.0 315400.00000000006 ;
      RECT  91400.0 314600.0 92200.0 315400.00000000006 ;
      RECT  96200.0 314600.0 97000.0 315400.00000000006 ;
      RECT  101000.0 314600.0 101800.0 315400.00000000006 ;
      RECT  105800.0 314600.0 106600.0 315400.00000000006 ;
      RECT  110600.00000000001 314600.0 111400.0 315400.00000000006 ;
      RECT  115400.0 314600.0 116200.0 315400.00000000006 ;
      RECT  120200.0 314600.0 121000.0 315400.00000000006 ;
      RECT  168200.0 314600.0 169000.0 315400.00000000006 ;
      RECT  173000.0 314600.0 173800.0 315400.00000000006 ;
      RECT  177800.0 314600.0 178600.00000000003 315400.00000000006 ;
      RECT  182600.0 314600.0 183400.0 315400.00000000006 ;
      RECT  187399.99999999997 314600.0 188200.0 315400.00000000006 ;
      RECT  192200.0 314600.0 193000.0 315400.00000000006 ;
      RECT  197000.0 314600.0 197800.0 315400.00000000006 ;
      RECT  201800.0 314600.0 202600.00000000003 315400.00000000006 ;
      RECT  206600.0 314600.0 207400.0 315400.00000000006 ;
      RECT  4999.999999999997 319400.0 5799.999999999997 320200.0 ;
      RECT  9799.999999999993 319400.0 10599.999999999995 320200.0 ;
      RECT  14599.999999999998 319400.0 15399.999999999998 320200.0 ;
      RECT  19399.999999999996 319400.0 20199.999999999996 320200.0 ;
      RECT  24200.0 319400.0 25000.0 320200.0 ;
      RECT  28999.999999999996 319400.0 29799.999999999996 320200.0 ;
      RECT  33800.0 319400.0 34599.99999999999 320200.0 ;
      RECT  38600.0 319400.0 39400.0 320200.0 ;
      RECT  43400.00000000001 319400.0 44200.0 320200.0 ;
      RECT  48200.0 319400.0 49000.0 320200.0 ;
      RECT  53000.0 319400.0 53800.0 320200.0 ;
      RECT  57800.0 319400.0 58599.99999999999 320200.0 ;
      RECT  62600.0 319400.0 63400.0 320200.0 ;
      RECT  67400.0 319400.0 68200.0 320200.0 ;
      RECT  72200.0 319400.0 73000.0 320200.0 ;
      RECT  77000.0 319400.0 77800.0 320200.0 ;
      RECT  81800.0 319400.0 82600.0 320200.0 ;
      RECT  86600.00000000001 319400.0 87400.0 320200.0 ;
      RECT  91400.0 319400.0 92200.0 320200.0 ;
      RECT  96200.0 319400.0 97000.0 320200.0 ;
      RECT  101000.0 319400.0 101800.0 320200.0 ;
      RECT  105800.0 319400.0 106600.0 320200.0 ;
      RECT  110600.00000000001 319400.0 111400.0 320200.0 ;
      RECT  115400.0 319400.0 116200.0 320200.0 ;
      RECT  120200.0 319400.0 121000.0 320200.0 ;
      RECT  125000.00000000001 319400.0 125800.00000000001 320200.0 ;
      RECT  129799.99999999999 319400.0 130600.0 320200.0 ;
      RECT  134600.0 319400.0 135400.0 320200.0 ;
      RECT  139399.99999999997 319400.0 140200.0 320200.0 ;
      RECT  144200.0 319400.0 145000.0 320200.0 ;
      RECT  149000.0 319400.0 149800.0 320200.0 ;
      RECT  153800.0 319400.0 154600.00000000003 320200.0 ;
      RECT  158600.0 319400.0 159400.0 320200.0 ;
      RECT  163399.99999999997 319400.0 164200.0 320200.0 ;
      RECT  168200.0 319400.0 169000.0 320200.0 ;
      RECT  173000.0 319400.0 173800.0 320200.0 ;
      RECT  177800.0 319400.0 178600.00000000003 320200.0 ;
      RECT  182600.0 319400.0 183400.0 320200.0 ;
      RECT  187399.99999999997 319400.0 188200.0 320200.0 ;
      RECT  192200.0 319400.0 193000.0 320200.0 ;
      RECT  197000.0 319400.0 197800.0 320200.0 ;
      RECT  201800.0 319400.0 202600.00000000003 320200.0 ;
      RECT  206600.0 319400.0 207400.0 320200.0 ;
      RECT  4999.999999999997 324200.0 5799.999999999997 325000.0 ;
      RECT  9799.999999999993 324200.0 10599.999999999995 325000.0 ;
      RECT  14599.999999999998 324200.0 15399.999999999998 325000.0 ;
      RECT  19399.999999999996 324200.0 20199.999999999996 325000.0 ;
      RECT  24200.0 324200.0 25000.0 325000.0 ;
      RECT  28999.999999999996 324200.0 29799.999999999996 325000.0 ;
      RECT  33800.0 324200.0 34599.99999999999 325000.0 ;
      RECT  38600.0 324200.0 39400.0 325000.0 ;
      RECT  43400.00000000001 324200.0 44200.0 325000.0 ;
      RECT  48200.0 324200.0 49000.0 325000.0 ;
      RECT  53000.0 324200.0 53800.0 325000.0 ;
      RECT  57800.0 324200.0 58599.99999999999 325000.0 ;
      RECT  86600.00000000001 324200.0 87400.0 325000.0 ;
      RECT  91400.0 324200.0 92200.0 325000.0 ;
      RECT  96200.0 324200.0 97000.0 325000.0 ;
      RECT  101000.0 324200.0 101800.0 325000.0 ;
      RECT  105800.0 324200.0 106600.0 325000.0 ;
      RECT  110600.00000000001 324200.0 111400.0 325000.0 ;
      RECT  115400.0 324200.0 116200.0 325000.0 ;
      RECT  120200.0 324200.0 121000.0 325000.0 ;
      RECT  125000.00000000001 324200.0 125800.00000000001 325000.0 ;
      RECT  129799.99999999999 324200.0 130600.0 325000.0 ;
      RECT  134600.0 324200.0 135400.0 325000.0 ;
      RECT  139399.99999999997 324200.0 140200.0 325000.0 ;
      RECT  144200.0 324200.0 145000.0 325000.0 ;
      RECT  149000.0 324200.0 149800.0 325000.0 ;
      RECT  153800.0 324200.0 154600.00000000003 325000.0 ;
      RECT  158600.0 324200.0 159400.0 325000.0 ;
      RECT  163399.99999999997 324200.0 164200.0 325000.0 ;
      RECT  168200.0 324200.0 169000.0 325000.0 ;
      RECT  173000.0 324200.0 173800.0 325000.0 ;
      RECT  177800.0 324200.0 178600.00000000003 325000.0 ;
      RECT  182600.0 324200.0 183400.0 325000.0 ;
      RECT  187399.99999999997 324200.0 188200.0 325000.0 ;
      RECT  192200.0 324200.0 193000.0 325000.0 ;
      RECT  197000.0 324200.0 197800.0 325000.0 ;
      RECT  201800.0 324200.0 202600.00000000003 325000.0 ;
      RECT  206600.0 324200.0 207400.0 325000.0 ;
      RECT  4999.999999999997 329000.0 5799.999999999997 329800.0 ;
      RECT  9799.999999999993 329000.0 10599.999999999995 329800.0 ;
      RECT  14599.999999999998 329000.0 15399.999999999998 329800.0 ;
      RECT  19399.999999999996 329000.0 20199.999999999996 329800.0 ;
      RECT  24200.0 329000.0 25000.0 329800.0 ;
      RECT  28999.999999999996 329000.0 29799.999999999996 329800.0 ;
      RECT  33800.0 329000.0 34599.99999999999 329800.0 ;
      RECT  38600.0 329000.0 39400.0 329800.0 ;
      RECT  43400.00000000001 329000.0 44200.0 329800.0 ;
      RECT  48200.0 329000.0 49000.0 329800.0 ;
      RECT  53000.0 329000.0 53800.0 329800.0 ;
      RECT  57800.0 329000.0 58599.99999999999 329800.0 ;
      RECT  62600.0 329000.0 63400.0 329800.0 ;
      RECT  67400.0 329000.0 68200.0 329800.0 ;
      RECT  72200.0 329000.0 73000.0 329800.0 ;
      RECT  77000.0 329000.0 77800.0 329800.0 ;
      RECT  81800.0 329000.0 82600.0 329800.0 ;
      RECT  86600.00000000001 329000.0 87400.0 329800.0 ;
      RECT  91400.0 329000.0 92200.0 329800.0 ;
      RECT  96200.0 329000.0 97000.0 329800.0 ;
      RECT  101000.0 329000.0 101800.0 329800.0 ;
      RECT  105800.0 329000.0 106600.0 329800.0 ;
      RECT  110600.00000000001 329000.0 111400.0 329800.0 ;
      RECT  115400.0 329000.0 116200.0 329800.0 ;
      RECT  120200.0 329000.0 121000.0 329800.0 ;
      RECT  125000.00000000001 329000.0 125800.00000000001 329800.0 ;
      RECT  129799.99999999999 329000.0 130600.0 329800.0 ;
      RECT  134600.0 329000.0 135400.0 329800.0 ;
      RECT  139399.99999999997 329000.0 140200.0 329800.0 ;
      RECT  144200.0 329000.0 145000.0 329800.0 ;
      RECT  149000.0 329000.0 149800.0 329800.0 ;
      RECT  153800.0 329000.0 154600.00000000003 329800.0 ;
      RECT  158600.0 329000.0 159400.0 329800.0 ;
      RECT  163399.99999999997 329000.0 164200.0 329800.0 ;
      RECT  168200.0 329000.0 169000.0 329800.0 ;
      RECT  173000.0 329000.0 173800.0 329800.0 ;
      RECT  177800.0 329000.0 178600.00000000003 329800.0 ;
      RECT  182600.0 329000.0 183400.0 329800.0 ;
      RECT  187399.99999999997 329000.0 188200.0 329800.0 ;
      RECT  192200.0 329000.0 193000.0 329800.0 ;
      RECT  197000.0 329000.0 197800.0 329800.0 ;
      RECT  201800.0 329000.0 202600.00000000003 329800.0 ;
      RECT  206600.0 329000.0 207400.0 329800.0 ;
      RECT  20200.0 170600.0 19400.0 171400.0 ;
      RECT  92200.0 213800.0 91400.0 214600.00000000003 ;
      RECT  17800.0 173000.0 17000.0 173800.0 ;
      RECT  22599.999999999996 175399.99999999997 21799.999999999996 176200.0 ;
      RECT  70600.0 200.0 69800.0 1000.0 ;
      RECT  89800.0 187399.99999999997 89000.0 188200.0 ;
      RECT  109000.0 187399.99999999997 108200.0 188200.0 ;
   END
   END    sram_2_16_scn4m_subm
END    LIBRARY
