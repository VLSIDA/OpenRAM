
.SUBCKT cell 
.ENDS cell
