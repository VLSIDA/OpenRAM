VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 148050.0 by 461850.0 ;
END  MacroSite
MACRO sram_2_16_1_scn3me_subm
   CLASS BLOCK ;
   SIZE 148050.0 BY 461850.0 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN DATA[0]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  120900.0 0.0 121800.0 1800.0 ;
      END
   END DATA[0]
   PIN DATA[1]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  131100.0 0.0 132000.0 1800.0 ;
      END
   END DATA[1]
   PIN ADDR[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 87600.0 10800.0 89100.0 ;
      END
   END ADDR[0]
   PIN ADDR[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 77400.0 10800.0 78900.0 ;
      END
   END ADDR[1]
   PIN ADDR[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 67200.0 10800.0 68700.0 ;
      END
   END ADDR[2]
   PIN ADDR[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 57000.0 10800.0 58500.0 ;
      END
   END ADDR[3]
   PIN CSb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  -38400.0 182700.0 -36600.0 184500.0 ;
      END
   END CSb
   PIN WEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  -28200.0 182700.0 -26400.0 184500.0 ;
      END
   END WEb
   PIN OEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  -48600.0 182700.0 -46800.0 184500.0 ;
      END
   END OEb
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER metal1 ;
         RECT  -10200.0 181800.0 -9000.0 185400.0 ;
      END
   END clk
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal2 ;
         RECT  4950.0 0.0 8550.0 461850.0 ;
         LAYER metal2 ;
         RECT  144450.0 0.0 148050.0 461850.0 ;
         LAYER metal1 ;
         RECT  0.0 4950.0 148050.0 8550.0 ;
         LAYER metal1 ;
         RECT  0.0 458250.0 148050.0 461850.0 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal2 ;
         RECT  0.0 0.0 3600.0 461850.0 ;
         LAYER metal2 ;
         RECT  139500.0 0.0 143100.0 461850.0 ;
         LAYER metal1 ;
         RECT  0.0 0.0 148050.0 3600.0 ;
         LAYER metal1 ;
         RECT  0.0 453300.0 148050.0 456900.0 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  48300.0 215550.0 49200.0 216450.0 ;
      RECT  48300.0 213150.0 49200.0 214050.0 ;
      RECT  46950.0 215550.0 48750.0 216450.0 ;
      RECT  48300.0 213600.0 49200.0 216000.0 ;
      RECT  48750.0 213150.0 50700.0 214050.0 ;
      RECT  100800.0 215550.0 101700.0 216450.0 ;
      RECT  100800.0 211050.0 101700.0 211950.0 ;
      RECT  86850.0 215550.0 101250.0 216450.0 ;
      RECT  100800.0 211500.0 101700.0 216000.0 ;
      RECT  101250.0 211050.0 115800.0 211950.0 ;
      RECT  48300.0 229950.0 49200.0 230850.0 ;
      RECT  48300.0 232350.0 49200.0 233250.0 ;
      RECT  46950.0 229950.0 48750.0 230850.0 ;
      RECT  48300.0 230400.0 49200.0 232800.0 ;
      RECT  48750.0 232350.0 50700.0 233250.0 ;
      RECT  100800.0 229950.0 101700.0 230850.0 ;
      RECT  100800.0 234450.0 101700.0 235350.0 ;
      RECT  86850.0 229950.0 101250.0 230850.0 ;
      RECT  100800.0 230400.0 101700.0 234900.0 ;
      RECT  101250.0 234450.0 115800.0 235350.0 ;
      RECT  48300.0 243150.0 49200.0 244050.0 ;
      RECT  48300.0 240750.0 49200.0 241650.0 ;
      RECT  46950.0 243150.0 48750.0 244050.0 ;
      RECT  48300.0 241200.0 49200.0 243600.0 ;
      RECT  48750.0 240750.0 50700.0 241650.0 ;
      RECT  100800.0 243150.0 101700.0 244050.0 ;
      RECT  100800.0 238650.0 101700.0 239550.0 ;
      RECT  86850.0 243150.0 101250.0 244050.0 ;
      RECT  100800.0 239100.0 101700.0 243600.0 ;
      RECT  101250.0 238650.0 115800.0 239550.0 ;
      RECT  48300.0 257550.0 49200.0 258450.0 ;
      RECT  48300.0 259950.0 49200.0 260850.0 ;
      RECT  46950.0 257550.0 48750.0 258450.0 ;
      RECT  48300.0 258000.0 49200.0 260400.0 ;
      RECT  48750.0 259950.0 50700.0 260850.0 ;
      RECT  100800.0 257550.0 101700.0 258450.0 ;
      RECT  100800.0 262050.0 101700.0 262950.0 ;
      RECT  86850.0 257550.0 101250.0 258450.0 ;
      RECT  100800.0 258000.0 101700.0 262500.0 ;
      RECT  101250.0 262050.0 115800.0 262950.0 ;
      RECT  48300.0 270750.0 49200.0 271650.0 ;
      RECT  48300.0 268350.0 49200.0 269250.0 ;
      RECT  46950.0 270750.0 48750.0 271650.0 ;
      RECT  48300.0 268800.0 49200.0 271200.0 ;
      RECT  48750.0 268350.0 50700.0 269250.0 ;
      RECT  100800.0 270750.0 101700.0 271650.0 ;
      RECT  100800.0 266250.0 101700.0 267150.0 ;
      RECT  86850.0 270750.0 101250.0 271650.0 ;
      RECT  100800.0 266700.0 101700.0 271200.0 ;
      RECT  101250.0 266250.0 115800.0 267150.0 ;
      RECT  48300.0 285150.0 49200.0 286050.0 ;
      RECT  48300.0 287550.0 49200.0 288450.0 ;
      RECT  46950.0 285150.0 48750.0 286050.0 ;
      RECT  48300.0 285600.0 49200.0 288000.0 ;
      RECT  48750.0 287550.0 50700.0 288450.0 ;
      RECT  100800.0 285150.0 101700.0 286050.0 ;
      RECT  100800.0 289650.0 101700.0 290550.0 ;
      RECT  86850.0 285150.0 101250.0 286050.0 ;
      RECT  100800.0 285600.0 101700.0 290100.0 ;
      RECT  101250.0 289650.0 115800.0 290550.0 ;
      RECT  48300.0 298350.0 49200.0 299250.0 ;
      RECT  48300.0 295950.0 49200.0 296850.0 ;
      RECT  46950.0 298350.0 48750.0 299250.0 ;
      RECT  48300.0 296400.0 49200.0 298800.0 ;
      RECT  48750.0 295950.0 50700.0 296850.0 ;
      RECT  100800.0 298350.0 101700.0 299250.0 ;
      RECT  100800.0 293850.0 101700.0 294750.0 ;
      RECT  86850.0 298350.0 101250.0 299250.0 ;
      RECT  100800.0 294300.0 101700.0 298800.0 ;
      RECT  101250.0 293850.0 115800.0 294750.0 ;
      RECT  48300.0 312750.0 49200.0 313650.0 ;
      RECT  48300.0 315150.0 49200.0 316050.0 ;
      RECT  46950.0 312750.0 48750.0 313650.0 ;
      RECT  48300.0 313200.0 49200.0 315600.0 ;
      RECT  48750.0 315150.0 50700.0 316050.0 ;
      RECT  100800.0 312750.0 101700.0 313650.0 ;
      RECT  100800.0 317250.0 101700.0 318150.0 ;
      RECT  86850.0 312750.0 101250.0 313650.0 ;
      RECT  100800.0 313200.0 101700.0 317700.0 ;
      RECT  101250.0 317250.0 115800.0 318150.0 ;
      RECT  48300.0 325950.0 49200.0 326850.0 ;
      RECT  48300.0 323550.0 49200.0 324450.0 ;
      RECT  46950.0 325950.0 48750.0 326850.0 ;
      RECT  48300.0 324000.0 49200.0 326400.0 ;
      RECT  48750.0 323550.0 50700.0 324450.0 ;
      RECT  100800.0 325950.0 101700.0 326850.0 ;
      RECT  100800.0 321450.0 101700.0 322350.0 ;
      RECT  86850.0 325950.0 101250.0 326850.0 ;
      RECT  100800.0 321900.0 101700.0 326400.0 ;
      RECT  101250.0 321450.0 115800.0 322350.0 ;
      RECT  48300.0 340350.0 49200.0 341250.0 ;
      RECT  48300.0 342750.0 49200.0 343650.0 ;
      RECT  46950.0 340350.0 48750.0 341250.0 ;
      RECT  48300.0 340800.0 49200.0 343200.0 ;
      RECT  48750.0 342750.0 50700.0 343650.0 ;
      RECT  100800.0 340350.0 101700.0 341250.0 ;
      RECT  100800.0 344850.0 101700.0 345750.0 ;
      RECT  86850.0 340350.0 101250.0 341250.0 ;
      RECT  100800.0 340800.0 101700.0 345300.0 ;
      RECT  101250.0 344850.0 115800.0 345750.0 ;
      RECT  48300.0 353550.0 49200.0 354450.0 ;
      RECT  48300.0 351150.0 49200.0 352050.0 ;
      RECT  46950.0 353550.0 48750.0 354450.0 ;
      RECT  48300.0 351600.0 49200.0 354000.0 ;
      RECT  48750.0 351150.0 50700.0 352050.0 ;
      RECT  100800.0 353550.0 101700.0 354450.0 ;
      RECT  100800.0 349050.0 101700.0 349950.0 ;
      RECT  86850.0 353550.0 101250.0 354450.0 ;
      RECT  100800.0 349500.0 101700.0 354000.0 ;
      RECT  101250.0 349050.0 115800.0 349950.0 ;
      RECT  48300.0 367950.0 49200.0 368850.0 ;
      RECT  48300.0 370350.0 49200.0 371250.0 ;
      RECT  46950.0 367950.0 48750.0 368850.0 ;
      RECT  48300.0 368400.0 49200.0 370800.0 ;
      RECT  48750.0 370350.0 50700.0 371250.0 ;
      RECT  100800.0 367950.0 101700.0 368850.0 ;
      RECT  100800.0 372450.0 101700.0 373350.0 ;
      RECT  86850.0 367950.0 101250.0 368850.0 ;
      RECT  100800.0 368400.0 101700.0 372900.0 ;
      RECT  101250.0 372450.0 115800.0 373350.0 ;
      RECT  48300.0 381150.0 49200.0 382050.0 ;
      RECT  48300.0 378750.0 49200.0 379650.0 ;
      RECT  46950.0 381150.0 48750.0 382050.0 ;
      RECT  48300.0 379200.0 49200.0 381600.0 ;
      RECT  48750.0 378750.0 50700.0 379650.0 ;
      RECT  100800.0 381150.0 101700.0 382050.0 ;
      RECT  100800.0 376650.0 101700.0 377550.0 ;
      RECT  86850.0 381150.0 101250.0 382050.0 ;
      RECT  100800.0 377100.0 101700.0 381600.0 ;
      RECT  101250.0 376650.0 115800.0 377550.0 ;
      RECT  48300.0 395550.0 49200.0 396450.0 ;
      RECT  48300.0 397950.0 49200.0 398850.0 ;
      RECT  46950.0 395550.0 48750.0 396450.0 ;
      RECT  48300.0 396000.0 49200.0 398400.0 ;
      RECT  48750.0 397950.0 50700.0 398850.0 ;
      RECT  100800.0 395550.0 101700.0 396450.0 ;
      RECT  100800.0 400050.0 101700.0 400950.0 ;
      RECT  86850.0 395550.0 101250.0 396450.0 ;
      RECT  100800.0 396000.0 101700.0 400500.0 ;
      RECT  101250.0 400050.0 115800.0 400950.0 ;
      RECT  48300.0 408750.0 49200.0 409650.0 ;
      RECT  48300.0 406350.0 49200.0 407250.0 ;
      RECT  46950.0 408750.0 48750.0 409650.0 ;
      RECT  48300.0 406800.0 49200.0 409200.0 ;
      RECT  48750.0 406350.0 50700.0 407250.0 ;
      RECT  100800.0 408750.0 101700.0 409650.0 ;
      RECT  100800.0 404250.0 101700.0 405150.0 ;
      RECT  86850.0 408750.0 101250.0 409650.0 ;
      RECT  100800.0 404700.0 101700.0 409200.0 ;
      RECT  101250.0 404250.0 115800.0 405150.0 ;
      RECT  48300.0 423150.0 49200.0 424050.0 ;
      RECT  48300.0 425550.0 49200.0 426450.0 ;
      RECT  46950.0 423150.0 48750.0 424050.0 ;
      RECT  48300.0 423600.0 49200.0 426000.0 ;
      RECT  48750.0 425550.0 50700.0 426450.0 ;
      RECT  100800.0 423150.0 101700.0 424050.0 ;
      RECT  100800.0 427650.0 101700.0 428550.0 ;
      RECT  86850.0 423150.0 101250.0 424050.0 ;
      RECT  100800.0 423600.0 101700.0 428100.0 ;
      RECT  101250.0 427650.0 115800.0 428550.0 ;
      RECT  81300.0 101250.0 85800.0 102150.0 ;
      RECT  78300.0 115050.0 88500.0 115950.0 ;
      RECT  81300.0 156450.0 91200.0 157350.0 ;
      RECT  78300.0 170250.0 93900.0 171150.0 ;
      RECT  1800.0 98550.0 81300.0 99450.0 ;
      RECT  1800.0 126150.0 81300.0 127050.0 ;
      RECT  1800.0 153750.0 81300.0 154650.0 ;
      RECT  1800.0 181350.0 81300.0 182250.0 ;
      RECT  6750.0 112350.0 81300.0 113250.0 ;
      RECT  6750.0 139950.0 81300.0 140850.0 ;
      RECT  6750.0 167550.0 81300.0 168450.0 ;
      RECT  6750.0 195150.0 81300.0 196050.0 ;
      RECT  68700.0 87300.0 85800.0 88200.0 ;
      RECT  68700.0 78600.0 88500.0 79500.0 ;
      RECT  68700.0 66900.0 91200.0 67800.0 ;
      RECT  68700.0 58200.0 93900.0 59100.0 ;
      RECT  1800.0 82950.0 9900.0 83850.0 ;
      RECT  1800.0 62550.0 9900.0 63450.0 ;
      RECT  66300.0 50250.0 67200.0 51150.0 ;
      RECT  66300.0 50700.0 67200.0 52800.0 ;
      RECT  6750.0 50250.0 66750.0 51150.0 ;
      RECT  104700.0 42300.0 116400.0 43200.0 ;
      RECT  99300.0 37800.0 116400.0 38700.0 ;
      RECT  102000.0 35400.0 116400.0 36300.0 ;
      RECT  104700.0 438600.0 116400.0 439500.0 ;
      RECT  107400.0 107100.0 116400.0 108000.0 ;
      RECT  110100.0 205200.0 116400.0 206100.0 ;
      RECT  12300.0 95250.0 13200.0 96150.0 ;
      RECT  12300.0 93600.0 13200.0 95700.0 ;
      RECT  12750.0 95250.0 96600.0 96150.0 ;
      RECT  53850.0 431850.0 97500.0 432750.0 ;
      RECT  116400.0 449700.0 146250.0 450600.0 ;
      RECT  116400.0 177900.0 146250.0 178800.0 ;
      RECT  116400.0 109200.0 146250.0 110100.0 ;
      RECT  116400.0 96300.0 146250.0 97200.0 ;
      RECT  116400.0 19500.0 146250.0 20400.0 ;
      RECT  6750.0 222750.0 146250.0 223650.0 ;
      RECT  6750.0 250350.0 146250.0 251250.0 ;
      RECT  6750.0 277950.0 146250.0 278850.0 ;
      RECT  6750.0 305550.0 146250.0 306450.0 ;
      RECT  6750.0 333150.0 146250.0 334050.0 ;
      RECT  6750.0 360750.0 146250.0 361650.0 ;
      RECT  6750.0 388350.0 146250.0 389250.0 ;
      RECT  6750.0 415950.0 146250.0 416850.0 ;
      RECT  116400.0 33300.0 143100.0 34200.0 ;
      RECT  116400.0 203100.0 143100.0 204000.0 ;
      RECT  116400.0 105000.0 143100.0 105900.0 ;
      RECT  1800.0 208950.0 57000.0 209850.0 ;
      RECT  1800.0 236550.0 57000.0 237450.0 ;
      RECT  1800.0 264150.0 57000.0 265050.0 ;
      RECT  1800.0 291750.0 57000.0 292650.0 ;
      RECT  1800.0 319350.0 57000.0 320250.0 ;
      RECT  1800.0 346950.0 57000.0 347850.0 ;
      RECT  1800.0 374550.0 57000.0 375450.0 ;
      RECT  1800.0 402150.0 57000.0 403050.0 ;
      RECT  1800.0 429750.0 57000.0 430650.0 ;
      RECT  116400.0 209400.0 126600.0 223200.0 ;
      RECT  116400.0 237000.0 126600.0 223200.0 ;
      RECT  116400.0 237000.0 126600.0 250800.0 ;
      RECT  116400.0 264600.0 126600.0 250800.0 ;
      RECT  116400.0 264600.0 126600.0 278400.0 ;
      RECT  116400.0 292200.0 126600.0 278400.0 ;
      RECT  116400.0 292200.0 126600.0 306000.0 ;
      RECT  116400.0 319800.0 126600.0 306000.0 ;
      RECT  116400.0 319800.0 126600.0 333600.0 ;
      RECT  116400.0 347400.0 126600.0 333600.0 ;
      RECT  116400.0 347400.0 126600.0 361200.0 ;
      RECT  116400.0 375000.0 126600.0 361200.0 ;
      RECT  116400.0 375000.0 126600.0 388800.0 ;
      RECT  116400.0 402600.0 126600.0 388800.0 ;
      RECT  116400.0 402600.0 126600.0 416400.0 ;
      RECT  116400.0 430200.0 126600.0 416400.0 ;
      RECT  126600.0 209400.0 136800.0 223200.0 ;
      RECT  126600.0 237000.0 136800.0 223200.0 ;
      RECT  126600.0 237000.0 136800.0 250800.0 ;
      RECT  126600.0 264600.0 136800.0 250800.0 ;
      RECT  126600.0 264600.0 136800.0 278400.0 ;
      RECT  126600.0 292200.0 136800.0 278400.0 ;
      RECT  126600.0 292200.0 136800.0 306000.0 ;
      RECT  126600.0 319800.0 136800.0 306000.0 ;
      RECT  126600.0 319800.0 136800.0 333600.0 ;
      RECT  126600.0 347400.0 136800.0 333600.0 ;
      RECT  126600.0 347400.0 136800.0 361200.0 ;
      RECT  126600.0 375000.0 136800.0 361200.0 ;
      RECT  126600.0 375000.0 136800.0 388800.0 ;
      RECT  126600.0 402600.0 136800.0 388800.0 ;
      RECT  126600.0 402600.0 136800.0 416400.0 ;
      RECT  126600.0 430200.0 136800.0 416400.0 ;
      RECT  115800.0 210900.0 137400.0 212100.0 ;
      RECT  115800.0 234300.0 137400.0 235500.0 ;
      RECT  115800.0 238500.0 137400.0 239700.0 ;
      RECT  115800.0 261900.0 137400.0 263100.0 ;
      RECT  115800.0 266100.0 137400.0 267300.0 ;
      RECT  115800.0 289500.0 137400.0 290700.0 ;
      RECT  115800.0 293700.0 137400.0 294900.0 ;
      RECT  115800.0 317100.0 137400.0 318300.0 ;
      RECT  115800.0 321300.0 137400.0 322500.0 ;
      RECT  115800.0 344700.0 137400.0 345900.0 ;
      RECT  115800.0 348900.0 137400.0 350100.0 ;
      RECT  115800.0 372300.0 137400.0 373500.0 ;
      RECT  115800.0 376500.0 137400.0 377700.0 ;
      RECT  115800.0 399900.0 137400.0 401100.0 ;
      RECT  115800.0 404100.0 137400.0 405300.0 ;
      RECT  115800.0 427500.0 137400.0 428700.0 ;
      RECT  115800.0 222600.0 137400.0 223500.0 ;
      RECT  115800.0 250200.0 137400.0 251100.0 ;
      RECT  115800.0 277800.0 137400.0 278700.0 ;
      RECT  115800.0 305400.0 137400.0 306300.0 ;
      RECT  115800.0 333000.0 137400.0 333900.0 ;
      RECT  115800.0 360600.0 137400.0 361500.0 ;
      RECT  115800.0 388200.0 137400.0 389100.0 ;
      RECT  115800.0 415800.0 137400.0 416700.0 ;
      RECT  121800.0 443400.0 123000.0 450600.0 ;
      RECT  119400.0 436200.0 120600.0 437400.0 ;
      RECT  121800.0 436200.0 123000.0 437400.0 ;
      RECT  121800.0 436200.0 123000.0 437400.0 ;
      RECT  119400.0 436200.0 120600.0 437400.0 ;
      RECT  119400.0 443400.0 120600.0 444600.0 ;
      RECT  121800.0 443400.0 123000.0 444600.0 ;
      RECT  121800.0 443400.0 123000.0 444600.0 ;
      RECT  119400.0 443400.0 120600.0 444600.0 ;
      RECT  121800.0 443400.0 123000.0 444600.0 ;
      RECT  124200.0 443400.0 125400.0 444600.0 ;
      RECT  124200.0 443400.0 125400.0 444600.0 ;
      RECT  121800.0 443400.0 123000.0 444600.0 ;
      RECT  121500.0 438450.0 120300.0 439650.0 ;
      RECT  121800.0 448800.0 123000.0 450000.0 ;
      RECT  119400.0 436200.0 120600.0 437400.0 ;
      RECT  121800.0 436200.0 123000.0 437400.0 ;
      RECT  119400.0 443400.0 120600.0 444600.0 ;
      RECT  124200.0 443400.0 125400.0 444600.0 ;
      RECT  116400.0 438600.0 126600.0 439500.0 ;
      RECT  116400.0 449700.0 126600.0 450600.0 ;
      RECT  132000.0 443400.0 133200.0 450600.0 ;
      RECT  129600.0 436200.0 130800.0 437400.0 ;
      RECT  132000.0 436200.0 133200.0 437400.0 ;
      RECT  132000.0 436200.0 133200.0 437400.0 ;
      RECT  129600.0 436200.0 130800.0 437400.0 ;
      RECT  129600.0 443400.0 130800.0 444600.0 ;
      RECT  132000.0 443400.0 133200.0 444600.0 ;
      RECT  132000.0 443400.0 133200.0 444600.0 ;
      RECT  129600.0 443400.0 130800.0 444600.0 ;
      RECT  132000.0 443400.0 133200.0 444600.0 ;
      RECT  134400.0 443400.0 135600.0 444600.0 ;
      RECT  134400.0 443400.0 135600.0 444600.0 ;
      RECT  132000.0 443400.0 133200.0 444600.0 ;
      RECT  131700.0 438450.0 130500.0 439650.0 ;
      RECT  132000.0 448800.0 133200.0 450000.0 ;
      RECT  129600.0 436200.0 130800.0 437400.0 ;
      RECT  132000.0 436200.0 133200.0 437400.0 ;
      RECT  129600.0 443400.0 130800.0 444600.0 ;
      RECT  134400.0 443400.0 135600.0 444600.0 ;
      RECT  126600.0 438600.0 136800.0 439500.0 ;
      RECT  126600.0 449700.0 136800.0 450600.0 ;
      RECT  116400.0 438600.0 136800.0 439500.0 ;
      RECT  116400.0 449700.0 136800.0 450600.0 ;
      RECT  116400.0 160500.0 126600.0 209400.0 ;
      RECT  126600.0 160500.0 136800.0 209400.0 ;
      RECT  116400.0 205200.0 136800.0 206100.0 ;
      RECT  116400.0 177900.0 136800.0 178800.0 ;
      RECT  116400.0 203100.0 136800.0 204000.0 ;
      RECT  116400.0 99900.0 126600.0 160500.0 ;
      RECT  126600.0 99900.0 136800.0 160500.0 ;
      RECT  116400.0 107100.0 136800.0 108000.0 ;
      RECT  116400.0 109200.0 136800.0 110100.0 ;
      RECT  116400.0 105000.0 136800.0 105900.0 ;
      RECT  116400.0 39900.0 126600.0 99900.0 ;
      RECT  136800.0 39900.0 126600.0 99900.0 ;
      RECT  116400.0 42300.0 136800.0 43200.0 ;
      RECT  116400.0 96300.0 136800.0 97200.0 ;
      RECT  116400.0 39900.0 126600.0 18000.0 ;
      RECT  126600.0 39900.0 136800.0 18000.0 ;
      RECT  116400.0 36300.0 136800.0 35400.0 ;
      RECT  116400.0 38700.0 136800.0 37800.0 ;
      RECT  116400.0 20400.0 136800.0 19500.0 ;
      RECT  116400.0 34200.0 136800.0 33300.0 ;
      RECT  38550.0 216750.0 39450.0 217650.0 ;
      RECT  38550.0 215550.0 39450.0 216450.0 ;
      RECT  34500.0 216750.0 39000.0 217650.0 ;
      RECT  38550.0 216000.0 39450.0 217200.0 ;
      RECT  39000.0 215550.0 43500.0 216450.0 ;
      RECT  38550.0 228750.0 39450.0 229650.0 ;
      RECT  38550.0 229950.0 39450.0 230850.0 ;
      RECT  34500.0 228750.0 39000.0 229650.0 ;
      RECT  38550.0 229200.0 39450.0 230400.0 ;
      RECT  39000.0 229950.0 43500.0 230850.0 ;
      RECT  38550.0 244350.0 39450.0 245250.0 ;
      RECT  38550.0 243150.0 39450.0 244050.0 ;
      RECT  34500.0 244350.0 39000.0 245250.0 ;
      RECT  38550.0 243600.0 39450.0 244800.0 ;
      RECT  39000.0 243150.0 43500.0 244050.0 ;
      RECT  38550.0 256350.0 39450.0 257250.0 ;
      RECT  38550.0 257550.0 39450.0 258450.0 ;
      RECT  34500.0 256350.0 39000.0 257250.0 ;
      RECT  38550.0 256800.0 39450.0 258000.0 ;
      RECT  39000.0 257550.0 43500.0 258450.0 ;
      RECT  38550.0 271950.0 39450.0 272850.0 ;
      RECT  38550.0 270750.0 39450.0 271650.0 ;
      RECT  34500.0 271950.0 39000.0 272850.0 ;
      RECT  38550.0 271200.0 39450.0 272400.0 ;
      RECT  39000.0 270750.0 43500.0 271650.0 ;
      RECT  38550.0 283950.0 39450.0 284850.0 ;
      RECT  38550.0 285150.0 39450.0 286050.0 ;
      RECT  34500.0 283950.0 39000.0 284850.0 ;
      RECT  38550.0 284400.0 39450.0 285600.0 ;
      RECT  39000.0 285150.0 43500.0 286050.0 ;
      RECT  38550.0 299550.0 39450.0 300450.0 ;
      RECT  38550.0 298350.0 39450.0 299250.0 ;
      RECT  34500.0 299550.0 39000.0 300450.0 ;
      RECT  38550.0 298800.0 39450.0 300000.0 ;
      RECT  39000.0 298350.0 43500.0 299250.0 ;
      RECT  38550.0 311550.0 39450.0 312450.0 ;
      RECT  38550.0 312750.0 39450.0 313650.0 ;
      RECT  34500.0 311550.0 39000.0 312450.0 ;
      RECT  38550.0 312000.0 39450.0 313200.0 ;
      RECT  39000.0 312750.0 43500.0 313650.0 ;
      RECT  38550.0 327150.0 39450.0 328050.0 ;
      RECT  38550.0 325950.0 39450.0 326850.0 ;
      RECT  34500.0 327150.0 39000.0 328050.0 ;
      RECT  38550.0 326400.0 39450.0 327600.0 ;
      RECT  39000.0 325950.0 43500.0 326850.0 ;
      RECT  38550.0 339150.0 39450.0 340050.0 ;
      RECT  38550.0 340350.0 39450.0 341250.0 ;
      RECT  34500.0 339150.0 39000.0 340050.0 ;
      RECT  38550.0 339600.0 39450.0 340800.0 ;
      RECT  39000.0 340350.0 43500.0 341250.0 ;
      RECT  38550.0 354750.0 39450.0 355650.0 ;
      RECT  38550.0 353550.0 39450.0 354450.0 ;
      RECT  34500.0 354750.0 39000.0 355650.0 ;
      RECT  38550.0 354000.0 39450.0 355200.0 ;
      RECT  39000.0 353550.0 43500.0 354450.0 ;
      RECT  38550.0 366750.0 39450.0 367650.0 ;
      RECT  38550.0 367950.0 39450.0 368850.0 ;
      RECT  34500.0 366750.0 39000.0 367650.0 ;
      RECT  38550.0 367200.0 39450.0 368400.0 ;
      RECT  39000.0 367950.0 43500.0 368850.0 ;
      RECT  38550.0 382350.0 39450.0 383250.0 ;
      RECT  38550.0 381150.0 39450.0 382050.0 ;
      RECT  34500.0 382350.0 39000.0 383250.0 ;
      RECT  38550.0 381600.0 39450.0 382800.0 ;
      RECT  39000.0 381150.0 43500.0 382050.0 ;
      RECT  38550.0 394350.0 39450.0 395250.0 ;
      RECT  38550.0 395550.0 39450.0 396450.0 ;
      RECT  34500.0 394350.0 39000.0 395250.0 ;
      RECT  38550.0 394800.0 39450.0 396000.0 ;
      RECT  39000.0 395550.0 43500.0 396450.0 ;
      RECT  38550.0 409950.0 39450.0 410850.0 ;
      RECT  38550.0 408750.0 39450.0 409650.0 ;
      RECT  34500.0 409950.0 39000.0 410850.0 ;
      RECT  38550.0 409200.0 39450.0 410400.0 ;
      RECT  39000.0 408750.0 43500.0 409650.0 ;
      RECT  38550.0 421950.0 39450.0 422850.0 ;
      RECT  38550.0 423150.0 39450.0 424050.0 ;
      RECT  34500.0 421950.0 39000.0 422850.0 ;
      RECT  38550.0 422400.0 39450.0 423600.0 ;
      RECT  39000.0 423150.0 43500.0 424050.0 ;
      RECT  10350.0 105150.0 26700.0 106050.0 ;
      RECT  12450.0 119550.0 26700.0 120450.0 ;
      RECT  14550.0 132750.0 26700.0 133650.0 ;
      RECT  16650.0 147150.0 26700.0 148050.0 ;
      RECT  18750.0 160350.0 26700.0 161250.0 ;
      RECT  20850.0 174750.0 26700.0 175650.0 ;
      RECT  22950.0 187950.0 26700.0 188850.0 ;
      RECT  25050.0 202350.0 26700.0 203250.0 ;
      RECT  10350.0 216750.0 29100.0 217650.0 ;
      RECT  18750.0 214050.0 32100.0 214950.0 ;
      RECT  10350.0 228750.0 29100.0 229650.0 ;
      RECT  20850.0 231450.0 32100.0 232350.0 ;
      RECT  10350.0 244350.0 29100.0 245250.0 ;
      RECT  22950.0 241650.0 32100.0 242550.0 ;
      RECT  10350.0 256350.0 29100.0 257250.0 ;
      RECT  25050.0 259050.0 32100.0 259950.0 ;
      RECT  12450.0 271950.0 29100.0 272850.0 ;
      RECT  18750.0 269250.0 32100.0 270150.0 ;
      RECT  12450.0 283950.0 29100.0 284850.0 ;
      RECT  20850.0 286650.0 32100.0 287550.0 ;
      RECT  12450.0 299550.0 29100.0 300450.0 ;
      RECT  22950.0 296850.0 32100.0 297750.0 ;
      RECT  12450.0 311550.0 29100.0 312450.0 ;
      RECT  25050.0 314250.0 32100.0 315150.0 ;
      RECT  14550.0 327150.0 29100.0 328050.0 ;
      RECT  18750.0 324450.0 32100.0 325350.0 ;
      RECT  14550.0 339150.0 29100.0 340050.0 ;
      RECT  20850.0 341850.0 32100.0 342750.0 ;
      RECT  14550.0 354750.0 29100.0 355650.0 ;
      RECT  22950.0 352050.0 32100.0 352950.0 ;
      RECT  14550.0 366750.0 29100.0 367650.0 ;
      RECT  25050.0 369450.0 32100.0 370350.0 ;
      RECT  16650.0 382350.0 29100.0 383250.0 ;
      RECT  18750.0 379650.0 32100.0 380550.0 ;
      RECT  16650.0 394350.0 29100.0 395250.0 ;
      RECT  20850.0 397050.0 32100.0 397950.0 ;
      RECT  16650.0 409950.0 29100.0 410850.0 ;
      RECT  22950.0 407250.0 32100.0 408150.0 ;
      RECT  16650.0 421950.0 29100.0 422850.0 ;
      RECT  25050.0 424650.0 32100.0 425550.0 ;
      RECT  65250.0 105150.0 64350.0 106050.0 ;
      RECT  65250.0 109650.0 64350.0 110550.0 ;
      RECT  69450.0 105150.0 64800.0 106050.0 ;
      RECT  65250.0 105600.0 64350.0 110100.0 ;
      RECT  64800.0 109650.0 62250.0 110550.0 ;
      RECT  80850.0 105150.0 72900.0 106050.0 ;
      RECT  65250.0 119550.0 64350.0 120450.0 ;
      RECT  65250.0 123450.0 64350.0 124350.0 ;
      RECT  69450.0 119550.0 64800.0 120450.0 ;
      RECT  65250.0 120000.0 64350.0 123900.0 ;
      RECT  64800.0 123450.0 59250.0 124350.0 ;
      RECT  77850.0 119550.0 72900.0 120450.0 ;
      RECT  80850.0 128250.0 56250.0 129150.0 ;
      RECT  77850.0 142050.0 53250.0 142950.0 ;
      RECT  62250.0 106350.0 48300.0 107250.0 ;
      RECT  59250.0 103650.0 45300.0 104550.0 ;
      RECT  56250.0 118350.0 48300.0 119250.0 ;
      RECT  59250.0 121050.0 45300.0 121950.0 ;
      RECT  62250.0 133950.0 48300.0 134850.0 ;
      RECT  53250.0 131250.0 45300.0 132150.0 ;
      RECT  56250.0 145950.0 48300.0 146850.0 ;
      RECT  53250.0 148650.0 45300.0 149550.0 ;
      RECT  38850.0 106350.0 37950.0 107250.0 ;
      RECT  38850.0 105150.0 37950.0 106050.0 ;
      RECT  42900.0 106350.0 38400.0 107250.0 ;
      RECT  38850.0 105600.0 37950.0 106800.0 ;
      RECT  38400.0 105150.0 33900.0 106050.0 ;
      RECT  38850.0 118350.0 37950.0 119250.0 ;
      RECT  38850.0 119550.0 37950.0 120450.0 ;
      RECT  42900.0 118350.0 38400.0 119250.0 ;
      RECT  38850.0 118800.0 37950.0 120000.0 ;
      RECT  38400.0 119550.0 33900.0 120450.0 ;
      RECT  38850.0 133950.0 37950.0 134850.0 ;
      RECT  38850.0 132750.0 37950.0 133650.0 ;
      RECT  42900.0 133950.0 38400.0 134850.0 ;
      RECT  38850.0 133200.0 37950.0 134400.0 ;
      RECT  38400.0 132750.0 33900.0 133650.0 ;
      RECT  38850.0 145950.0 37950.0 146850.0 ;
      RECT  38850.0 147150.0 37950.0 148050.0 ;
      RECT  42900.0 145950.0 38400.0 146850.0 ;
      RECT  38850.0 146400.0 37950.0 147600.0 ;
      RECT  38400.0 147150.0 33900.0 148050.0 ;
      RECT  68700.0 110850.0 67500.0 112800.0 ;
      RECT  68700.0 99000.0 67500.0 100950.0 ;
      RECT  73500.0 100350.0 72300.0 98550.0 ;
      RECT  73500.0 109650.0 72300.0 113250.0 ;
      RECT  70800.0 100350.0 69900.0 109650.0 ;
      RECT  73500.0 109650.0 72300.0 110850.0 ;
      RECT  71100.0 109650.0 69900.0 110850.0 ;
      RECT  71100.0 109650.0 69900.0 110850.0 ;
      RECT  73500.0 109650.0 72300.0 110850.0 ;
      RECT  73500.0 100350.0 72300.0 101550.0 ;
      RECT  71100.0 100350.0 69900.0 101550.0 ;
      RECT  71100.0 100350.0 69900.0 101550.0 ;
      RECT  73500.0 100350.0 72300.0 101550.0 ;
      RECT  68700.0 110250.0 67500.0 111450.0 ;
      RECT  68700.0 100350.0 67500.0 101550.0 ;
      RECT  72900.0 105000.0 71700.0 106200.0 ;
      RECT  72900.0 105000.0 71700.0 106200.0 ;
      RECT  70350.0 105150.0 69450.0 106050.0 ;
      RECT  75300.0 112350.0 65700.0 113250.0 ;
      RECT  75300.0 98550.0 65700.0 99450.0 ;
      RECT  68700.0 114750.0 67500.0 112800.0 ;
      RECT  68700.0 126600.0 67500.0 124650.0 ;
      RECT  73500.0 125250.0 72300.0 127050.0 ;
      RECT  73500.0 115950.0 72300.0 112350.0 ;
      RECT  70800.0 125250.0 69900.0 115950.0 ;
      RECT  73500.0 115950.0 72300.0 114750.0 ;
      RECT  71100.0 115950.0 69900.0 114750.0 ;
      RECT  71100.0 115950.0 69900.0 114750.0 ;
      RECT  73500.0 115950.0 72300.0 114750.0 ;
      RECT  73500.0 125250.0 72300.0 124050.0 ;
      RECT  71100.0 125250.0 69900.0 124050.0 ;
      RECT  71100.0 125250.0 69900.0 124050.0 ;
      RECT  73500.0 125250.0 72300.0 124050.0 ;
      RECT  68700.0 115350.0 67500.0 114150.0 ;
      RECT  68700.0 125250.0 67500.0 124050.0 ;
      RECT  72900.0 120600.0 71700.0 119400.0 ;
      RECT  72900.0 120600.0 71700.0 119400.0 ;
      RECT  70350.0 120450.0 69450.0 119550.0 ;
      RECT  75300.0 113250.0 65700.0 112350.0 ;
      RECT  75300.0 127050.0 65700.0 126150.0 ;
      RECT  29700.0 110850.0 28500.0 112800.0 ;
      RECT  29700.0 99000.0 28500.0 100950.0 ;
      RECT  34500.0 100350.0 33300.0 98550.0 ;
      RECT  34500.0 109650.0 33300.0 113250.0 ;
      RECT  31800.0 100350.0 30900.0 109650.0 ;
      RECT  34500.0 109650.0 33300.0 110850.0 ;
      RECT  32100.0 109650.0 30900.0 110850.0 ;
      RECT  32100.0 109650.0 30900.0 110850.0 ;
      RECT  34500.0 109650.0 33300.0 110850.0 ;
      RECT  34500.0 100350.0 33300.0 101550.0 ;
      RECT  32100.0 100350.0 30900.0 101550.0 ;
      RECT  32100.0 100350.0 30900.0 101550.0 ;
      RECT  34500.0 100350.0 33300.0 101550.0 ;
      RECT  29700.0 110250.0 28500.0 111450.0 ;
      RECT  29700.0 100350.0 28500.0 101550.0 ;
      RECT  33900.0 105000.0 32700.0 106200.0 ;
      RECT  33900.0 105000.0 32700.0 106200.0 ;
      RECT  31350.0 105150.0 30450.0 106050.0 ;
      RECT  36300.0 112350.0 26700.0 113250.0 ;
      RECT  36300.0 98550.0 26700.0 99450.0 ;
      RECT  29700.0 114750.0 28500.0 112800.0 ;
      RECT  29700.0 126600.0 28500.0 124650.0 ;
      RECT  34500.0 125250.0 33300.0 127050.0 ;
      RECT  34500.0 115950.0 33300.0 112350.0 ;
      RECT  31800.0 125250.0 30900.0 115950.0 ;
      RECT  34500.0 115950.0 33300.0 114750.0 ;
      RECT  32100.0 115950.0 30900.0 114750.0 ;
      RECT  32100.0 115950.0 30900.0 114750.0 ;
      RECT  34500.0 115950.0 33300.0 114750.0 ;
      RECT  34500.0 125250.0 33300.0 124050.0 ;
      RECT  32100.0 125250.0 30900.0 124050.0 ;
      RECT  32100.0 125250.0 30900.0 124050.0 ;
      RECT  34500.0 125250.0 33300.0 124050.0 ;
      RECT  29700.0 115350.0 28500.0 114150.0 ;
      RECT  29700.0 125250.0 28500.0 124050.0 ;
      RECT  33900.0 120600.0 32700.0 119400.0 ;
      RECT  33900.0 120600.0 32700.0 119400.0 ;
      RECT  31350.0 120450.0 30450.0 119550.0 ;
      RECT  36300.0 113250.0 26700.0 112350.0 ;
      RECT  36300.0 127050.0 26700.0 126150.0 ;
      RECT  29700.0 138450.0 28500.0 140400.0 ;
      RECT  29700.0 126600.0 28500.0 128550.0 ;
      RECT  34500.0 127950.0 33300.0 126150.0 ;
      RECT  34500.0 137250.0 33300.0 140850.0 ;
      RECT  31800.0 127950.0 30900.0 137250.0 ;
      RECT  34500.0 137250.0 33300.0 138450.0 ;
      RECT  32100.0 137250.0 30900.0 138450.0 ;
      RECT  32100.0 137250.0 30900.0 138450.0 ;
      RECT  34500.0 137250.0 33300.0 138450.0 ;
      RECT  34500.0 127950.0 33300.0 129150.0 ;
      RECT  32100.0 127950.0 30900.0 129150.0 ;
      RECT  32100.0 127950.0 30900.0 129150.0 ;
      RECT  34500.0 127950.0 33300.0 129150.0 ;
      RECT  29700.0 137850.0 28500.0 139050.0 ;
      RECT  29700.0 127950.0 28500.0 129150.0 ;
      RECT  33900.0 132600.0 32700.0 133800.0 ;
      RECT  33900.0 132600.0 32700.0 133800.0 ;
      RECT  31350.0 132750.0 30450.0 133650.0 ;
      RECT  36300.0 139950.0 26700.0 140850.0 ;
      RECT  36300.0 126150.0 26700.0 127050.0 ;
      RECT  29700.0 142350.0 28500.0 140400.0 ;
      RECT  29700.0 154200.0 28500.0 152250.0 ;
      RECT  34500.0 152850.0 33300.0 154650.0 ;
      RECT  34500.0 143550.0 33300.0 139950.0 ;
      RECT  31800.0 152850.0 30900.0 143550.0 ;
      RECT  34500.0 143550.0 33300.0 142350.0 ;
      RECT  32100.0 143550.0 30900.0 142350.0 ;
      RECT  32100.0 143550.0 30900.0 142350.0 ;
      RECT  34500.0 143550.0 33300.0 142350.0 ;
      RECT  34500.0 152850.0 33300.0 151650.0 ;
      RECT  32100.0 152850.0 30900.0 151650.0 ;
      RECT  32100.0 152850.0 30900.0 151650.0 ;
      RECT  34500.0 152850.0 33300.0 151650.0 ;
      RECT  29700.0 142950.0 28500.0 141750.0 ;
      RECT  29700.0 152850.0 28500.0 151650.0 ;
      RECT  33900.0 148200.0 32700.0 147000.0 ;
      RECT  33900.0 148200.0 32700.0 147000.0 ;
      RECT  31350.0 148050.0 30450.0 147150.0 ;
      RECT  36300.0 140850.0 26700.0 139950.0 ;
      RECT  36300.0 154650.0 26700.0 153750.0 ;
      RECT  48900.0 100950.0 47700.0 98550.0 ;
      RECT  48900.0 109650.0 47700.0 113250.0 ;
      RECT  44100.0 109650.0 42900.0 113250.0 ;
      RECT  41700.0 110850.0 40500.0 112800.0 ;
      RECT  41700.0 99000.0 40500.0 100950.0 ;
      RECT  48900.0 109650.0 47700.0 110850.0 ;
      RECT  46500.0 109650.0 45300.0 110850.0 ;
      RECT  46500.0 109650.0 45300.0 110850.0 ;
      RECT  48900.0 109650.0 47700.0 110850.0 ;
      RECT  46500.0 109650.0 45300.0 110850.0 ;
      RECT  44100.0 109650.0 42900.0 110850.0 ;
      RECT  44100.0 109650.0 42900.0 110850.0 ;
      RECT  46500.0 109650.0 45300.0 110850.0 ;
      RECT  48900.0 100950.0 47700.0 102150.0 ;
      RECT  46500.0 100950.0 45300.0 102150.0 ;
      RECT  46500.0 100950.0 45300.0 102150.0 ;
      RECT  48900.0 100950.0 47700.0 102150.0 ;
      RECT  46500.0 100950.0 45300.0 102150.0 ;
      RECT  44100.0 100950.0 42900.0 102150.0 ;
      RECT  44100.0 100950.0 42900.0 102150.0 ;
      RECT  46500.0 100950.0 45300.0 102150.0 ;
      RECT  41700.0 110250.0 40500.0 111450.0 ;
      RECT  41700.0 100350.0 40500.0 101550.0 ;
      RECT  44100.0 103500.0 45300.0 104700.0 ;
      RECT  47100.0 106200.0 48300.0 107400.0 ;
      RECT  46500.0 109650.0 45300.0 110850.0 ;
      RECT  44100.0 100950.0 42900.0 102150.0 ;
      RECT  42900.0 106200.0 44100.0 107400.0 ;
      RECT  48300.0 106200.0 47100.0 107400.0 ;
      RECT  45300.0 103500.0 44100.0 104700.0 ;
      RECT  44100.0 106200.0 42900.0 107400.0 ;
      RECT  50700.0 112350.0 36300.0 113250.0 ;
      RECT  50700.0 98550.0 36300.0 99450.0 ;
      RECT  48900.0 124650.0 47700.0 127050.0 ;
      RECT  48900.0 115950.0 47700.0 112350.0 ;
      RECT  44100.0 115950.0 42900.0 112350.0 ;
      RECT  41700.0 114750.0 40500.0 112800.0 ;
      RECT  41700.0 126600.0 40500.0 124650.0 ;
      RECT  48900.0 115950.0 47700.0 114750.0 ;
      RECT  46500.0 115950.0 45300.0 114750.0 ;
      RECT  46500.0 115950.0 45300.0 114750.0 ;
      RECT  48900.0 115950.0 47700.0 114750.0 ;
      RECT  46500.0 115950.0 45300.0 114750.0 ;
      RECT  44100.0 115950.0 42900.0 114750.0 ;
      RECT  44100.0 115950.0 42900.0 114750.0 ;
      RECT  46500.0 115950.0 45300.0 114750.0 ;
      RECT  48900.0 124650.0 47700.0 123450.0 ;
      RECT  46500.0 124650.0 45300.0 123450.0 ;
      RECT  46500.0 124650.0 45300.0 123450.0 ;
      RECT  48900.0 124650.0 47700.0 123450.0 ;
      RECT  46500.0 124650.0 45300.0 123450.0 ;
      RECT  44100.0 124650.0 42900.0 123450.0 ;
      RECT  44100.0 124650.0 42900.0 123450.0 ;
      RECT  46500.0 124650.0 45300.0 123450.0 ;
      RECT  41700.0 115350.0 40500.0 114150.0 ;
      RECT  41700.0 125250.0 40500.0 124050.0 ;
      RECT  44100.0 122100.0 45300.0 120900.0 ;
      RECT  47100.0 119400.0 48300.0 118200.0 ;
      RECT  46500.0 115950.0 45300.0 114750.0 ;
      RECT  44100.0 124650.0 42900.0 123450.0 ;
      RECT  42900.0 119400.0 44100.0 118200.0 ;
      RECT  48300.0 119400.0 47100.0 118200.0 ;
      RECT  45300.0 122100.0 44100.0 120900.0 ;
      RECT  44100.0 119400.0 42900.0 118200.0 ;
      RECT  50700.0 113250.0 36300.0 112350.0 ;
      RECT  50700.0 127050.0 36300.0 126150.0 ;
      RECT  48900.0 128550.0 47700.0 126150.0 ;
      RECT  48900.0 137250.0 47700.0 140850.0 ;
      RECT  44100.0 137250.0 42900.0 140850.0 ;
      RECT  41700.0 138450.0 40500.0 140400.0 ;
      RECT  41700.0 126600.0 40500.0 128550.0 ;
      RECT  48900.0 137250.0 47700.0 138450.0 ;
      RECT  46500.0 137250.0 45300.0 138450.0 ;
      RECT  46500.0 137250.0 45300.0 138450.0 ;
      RECT  48900.0 137250.0 47700.0 138450.0 ;
      RECT  46500.0 137250.0 45300.0 138450.0 ;
      RECT  44100.0 137250.0 42900.0 138450.0 ;
      RECT  44100.0 137250.0 42900.0 138450.0 ;
      RECT  46500.0 137250.0 45300.0 138450.0 ;
      RECT  48900.0 128550.0 47700.0 129750.0 ;
      RECT  46500.0 128550.0 45300.0 129750.0 ;
      RECT  46500.0 128550.0 45300.0 129750.0 ;
      RECT  48900.0 128550.0 47700.0 129750.0 ;
      RECT  46500.0 128550.0 45300.0 129750.0 ;
      RECT  44100.0 128550.0 42900.0 129750.0 ;
      RECT  44100.0 128550.0 42900.0 129750.0 ;
      RECT  46500.0 128550.0 45300.0 129750.0 ;
      RECT  41700.0 137850.0 40500.0 139050.0 ;
      RECT  41700.0 127950.0 40500.0 129150.0 ;
      RECT  44100.0 131100.0 45300.0 132300.0 ;
      RECT  47100.0 133800.0 48300.0 135000.0 ;
      RECT  46500.0 137250.0 45300.0 138450.0 ;
      RECT  44100.0 128550.0 42900.0 129750.0 ;
      RECT  42900.0 133800.0 44100.0 135000.0 ;
      RECT  48300.0 133800.0 47100.0 135000.0 ;
      RECT  45300.0 131100.0 44100.0 132300.0 ;
      RECT  44100.0 133800.0 42900.0 135000.0 ;
      RECT  50700.0 139950.0 36300.0 140850.0 ;
      RECT  50700.0 126150.0 36300.0 127050.0 ;
      RECT  48900.0 152250.0 47700.0 154650.0 ;
      RECT  48900.0 143550.0 47700.0 139950.0 ;
      RECT  44100.0 143550.0 42900.0 139950.0 ;
      RECT  41700.0 142350.0 40500.0 140400.0 ;
      RECT  41700.0 154200.0 40500.0 152250.0 ;
      RECT  48900.0 143550.0 47700.0 142350.0 ;
      RECT  46500.0 143550.0 45300.0 142350.0 ;
      RECT  46500.0 143550.0 45300.0 142350.0 ;
      RECT  48900.0 143550.0 47700.0 142350.0 ;
      RECT  46500.0 143550.0 45300.0 142350.0 ;
      RECT  44100.0 143550.0 42900.0 142350.0 ;
      RECT  44100.0 143550.0 42900.0 142350.0 ;
      RECT  46500.0 143550.0 45300.0 142350.0 ;
      RECT  48900.0 152250.0 47700.0 151050.0 ;
      RECT  46500.0 152250.0 45300.0 151050.0 ;
      RECT  46500.0 152250.0 45300.0 151050.0 ;
      RECT  48900.0 152250.0 47700.0 151050.0 ;
      RECT  46500.0 152250.0 45300.0 151050.0 ;
      RECT  44100.0 152250.0 42900.0 151050.0 ;
      RECT  44100.0 152250.0 42900.0 151050.0 ;
      RECT  46500.0 152250.0 45300.0 151050.0 ;
      RECT  41700.0 142950.0 40500.0 141750.0 ;
      RECT  41700.0 152850.0 40500.0 151650.0 ;
      RECT  44100.0 149700.0 45300.0 148500.0 ;
      RECT  47100.0 147000.0 48300.0 145800.0 ;
      RECT  46500.0 143550.0 45300.0 142350.0 ;
      RECT  44100.0 152250.0 42900.0 151050.0 ;
      RECT  42900.0 147000.0 44100.0 145800.0 ;
      RECT  48300.0 147000.0 47100.0 145800.0 ;
      RECT  45300.0 149700.0 44100.0 148500.0 ;
      RECT  44100.0 147000.0 42900.0 145800.0 ;
      RECT  50700.0 140850.0 36300.0 139950.0 ;
      RECT  50700.0 154650.0 36300.0 153750.0 ;
      RECT  61650.0 109500.0 62850.0 110700.0 ;
      RECT  80250.0 105000.0 81450.0 106200.0 ;
      RECT  58650.0 123300.0 59850.0 124500.0 ;
      RECT  77250.0 119400.0 78450.0 120600.0 ;
      RECT  80250.0 128100.0 81450.0 129300.0 ;
      RECT  55650.0 128100.0 56850.0 129300.0 ;
      RECT  77250.0 141900.0 78450.0 143100.0 ;
      RECT  52650.0 141900.0 53850.0 143100.0 ;
      RECT  61650.0 106200.0 62850.0 107400.0 ;
      RECT  58650.0 103500.0 59850.0 104700.0 ;
      RECT  55650.0 118200.0 56850.0 119400.0 ;
      RECT  58650.0 120900.0 59850.0 122100.0 ;
      RECT  61650.0 133800.0 62850.0 135000.0 ;
      RECT  52650.0 131100.0 53850.0 132300.0 ;
      RECT  55650.0 145800.0 56850.0 147000.0 ;
      RECT  52650.0 148500.0 53850.0 149700.0 ;
      RECT  30450.0 105150.0 26700.0 106050.0 ;
      RECT  30450.0 119550.0 26700.0 120450.0 ;
      RECT  30450.0 132750.0 26700.0 133650.0 ;
      RECT  30450.0 147150.0 26700.0 148050.0 ;
      RECT  81300.0 112350.0 26700.0 113250.0 ;
      RECT  81300.0 139950.0 26700.0 140850.0 ;
      RECT  81300.0 98550.0 26700.0 99450.0 ;
      RECT  81300.0 126150.0 26700.0 127050.0 ;
      RECT  81300.0 153750.0 26700.0 154650.0 ;
      RECT  65250.0 160350.0 64350.0 161250.0 ;
      RECT  65250.0 164850.0 64350.0 165750.0 ;
      RECT  69450.0 160350.0 64800.0 161250.0 ;
      RECT  65250.0 160800.0 64350.0 165300.0 ;
      RECT  64800.0 164850.0 62250.0 165750.0 ;
      RECT  80850.0 160350.0 72900.0 161250.0 ;
      RECT  65250.0 174750.0 64350.0 175650.0 ;
      RECT  65250.0 178650.0 64350.0 179550.0 ;
      RECT  69450.0 174750.0 64800.0 175650.0 ;
      RECT  65250.0 175200.0 64350.0 179100.0 ;
      RECT  64800.0 178650.0 59250.0 179550.0 ;
      RECT  77850.0 174750.0 72900.0 175650.0 ;
      RECT  80850.0 183450.0 56250.0 184350.0 ;
      RECT  77850.0 197250.0 53250.0 198150.0 ;
      RECT  62250.0 161550.0 48300.0 162450.0 ;
      RECT  59250.0 158850.0 45300.0 159750.0 ;
      RECT  56250.0 173550.0 48300.0 174450.0 ;
      RECT  59250.0 176250.0 45300.0 177150.0 ;
      RECT  62250.0 189150.0 48300.0 190050.0 ;
      RECT  53250.0 186450.0 45300.0 187350.0 ;
      RECT  56250.0 201150.0 48300.0 202050.0 ;
      RECT  53250.0 203850.0 45300.0 204750.0 ;
      RECT  38850.0 161550.0 37950.0 162450.0 ;
      RECT  38850.0 160350.0 37950.0 161250.0 ;
      RECT  42900.0 161550.0 38400.0 162450.0 ;
      RECT  38850.0 160800.0 37950.0 162000.0 ;
      RECT  38400.0 160350.0 33900.0 161250.0 ;
      RECT  38850.0 173550.0 37950.0 174450.0 ;
      RECT  38850.0 174750.0 37950.0 175650.0 ;
      RECT  42900.0 173550.0 38400.0 174450.0 ;
      RECT  38850.0 174000.0 37950.0 175200.0 ;
      RECT  38400.0 174750.0 33900.0 175650.0 ;
      RECT  38850.0 189150.0 37950.0 190050.0 ;
      RECT  38850.0 187950.0 37950.0 188850.0 ;
      RECT  42900.0 189150.0 38400.0 190050.0 ;
      RECT  38850.0 188400.0 37950.0 189600.0 ;
      RECT  38400.0 187950.0 33900.0 188850.0 ;
      RECT  38850.0 201150.0 37950.0 202050.0 ;
      RECT  38850.0 202350.0 37950.0 203250.0 ;
      RECT  42900.0 201150.0 38400.0 202050.0 ;
      RECT  38850.0 201600.0 37950.0 202800.0 ;
      RECT  38400.0 202350.0 33900.0 203250.0 ;
      RECT  68700.0 166050.0 67500.0 168000.0 ;
      RECT  68700.0 154200.0 67500.0 156150.0 ;
      RECT  73500.0 155550.0 72300.0 153750.0 ;
      RECT  73500.0 164850.0 72300.0 168450.0 ;
      RECT  70800.0 155550.0 69900.0 164850.0 ;
      RECT  73500.0 164850.0 72300.0 166050.0 ;
      RECT  71100.0 164850.0 69900.0 166050.0 ;
      RECT  71100.0 164850.0 69900.0 166050.0 ;
      RECT  73500.0 164850.0 72300.0 166050.0 ;
      RECT  73500.0 155550.0 72300.0 156750.0 ;
      RECT  71100.0 155550.0 69900.0 156750.0 ;
      RECT  71100.0 155550.0 69900.0 156750.0 ;
      RECT  73500.0 155550.0 72300.0 156750.0 ;
      RECT  68700.0 165450.0 67500.0 166650.0 ;
      RECT  68700.0 155550.0 67500.0 156750.0 ;
      RECT  72900.0 160200.0 71700.0 161400.0 ;
      RECT  72900.0 160200.0 71700.0 161400.0 ;
      RECT  70350.0 160350.0 69450.0 161250.0 ;
      RECT  75300.0 167550.0 65700.0 168450.0 ;
      RECT  75300.0 153750.0 65700.0 154650.0 ;
      RECT  68700.0 169950.0 67500.0 168000.0 ;
      RECT  68700.0 181800.0 67500.0 179850.0 ;
      RECT  73500.0 180450.0 72300.0 182250.0 ;
      RECT  73500.0 171150.0 72300.0 167550.0 ;
      RECT  70800.0 180450.0 69900.0 171150.0 ;
      RECT  73500.0 171150.0 72300.0 169950.0 ;
      RECT  71100.0 171150.0 69900.0 169950.0 ;
      RECT  71100.0 171150.0 69900.0 169950.0 ;
      RECT  73500.0 171150.0 72300.0 169950.0 ;
      RECT  73500.0 180450.0 72300.0 179250.0 ;
      RECT  71100.0 180450.0 69900.0 179250.0 ;
      RECT  71100.0 180450.0 69900.0 179250.0 ;
      RECT  73500.0 180450.0 72300.0 179250.0 ;
      RECT  68700.0 170550.0 67500.0 169350.0 ;
      RECT  68700.0 180450.0 67500.0 179250.0 ;
      RECT  72900.0 175800.0 71700.0 174600.0 ;
      RECT  72900.0 175800.0 71700.0 174600.0 ;
      RECT  70350.0 175650.0 69450.0 174750.0 ;
      RECT  75300.0 168450.0 65700.0 167550.0 ;
      RECT  75300.0 182250.0 65700.0 181350.0 ;
      RECT  29700.0 166050.0 28500.0 168000.0 ;
      RECT  29700.0 154200.0 28500.0 156150.0 ;
      RECT  34500.0 155550.0 33300.0 153750.0 ;
      RECT  34500.0 164850.0 33300.0 168450.0 ;
      RECT  31800.0 155550.0 30900.0 164850.0 ;
      RECT  34500.0 164850.0 33300.0 166050.0 ;
      RECT  32100.0 164850.0 30900.0 166050.0 ;
      RECT  32100.0 164850.0 30900.0 166050.0 ;
      RECT  34500.0 164850.0 33300.0 166050.0 ;
      RECT  34500.0 155550.0 33300.0 156750.0 ;
      RECT  32100.0 155550.0 30900.0 156750.0 ;
      RECT  32100.0 155550.0 30900.0 156750.0 ;
      RECT  34500.0 155550.0 33300.0 156750.0 ;
      RECT  29700.0 165450.0 28500.0 166650.0 ;
      RECT  29700.0 155550.0 28500.0 156750.0 ;
      RECT  33900.0 160200.0 32700.0 161400.0 ;
      RECT  33900.0 160200.0 32700.0 161400.0 ;
      RECT  31350.0 160350.0 30450.0 161250.0 ;
      RECT  36300.0 167550.0 26700.0 168450.0 ;
      RECT  36300.0 153750.0 26700.0 154650.0 ;
      RECT  29700.0 169950.0 28500.0 168000.0 ;
      RECT  29700.0 181800.0 28500.0 179850.0 ;
      RECT  34500.0 180450.0 33300.0 182250.0 ;
      RECT  34500.0 171150.0 33300.0 167550.0 ;
      RECT  31800.0 180450.0 30900.0 171150.0 ;
      RECT  34500.0 171150.0 33300.0 169950.0 ;
      RECT  32100.0 171150.0 30900.0 169950.0 ;
      RECT  32100.0 171150.0 30900.0 169950.0 ;
      RECT  34500.0 171150.0 33300.0 169950.0 ;
      RECT  34500.0 180450.0 33300.0 179250.0 ;
      RECT  32100.0 180450.0 30900.0 179250.0 ;
      RECT  32100.0 180450.0 30900.0 179250.0 ;
      RECT  34500.0 180450.0 33300.0 179250.0 ;
      RECT  29700.0 170550.0 28500.0 169350.0 ;
      RECT  29700.0 180450.0 28500.0 179250.0 ;
      RECT  33900.0 175800.0 32700.0 174600.0 ;
      RECT  33900.0 175800.0 32700.0 174600.0 ;
      RECT  31350.0 175650.0 30450.0 174750.0 ;
      RECT  36300.0 168450.0 26700.0 167550.0 ;
      RECT  36300.0 182250.0 26700.0 181350.0 ;
      RECT  29700.0 193650.0 28500.0 195600.0 ;
      RECT  29700.0 181800.0 28500.0 183750.0 ;
      RECT  34500.0 183150.0 33300.0 181350.0 ;
      RECT  34500.0 192450.0 33300.0 196050.0 ;
      RECT  31800.0 183150.0 30900.0 192450.0 ;
      RECT  34500.0 192450.0 33300.0 193650.0 ;
      RECT  32100.0 192450.0 30900.0 193650.0 ;
      RECT  32100.0 192450.0 30900.0 193650.0 ;
      RECT  34500.0 192450.0 33300.0 193650.0 ;
      RECT  34500.0 183150.0 33300.0 184350.0 ;
      RECT  32100.0 183150.0 30900.0 184350.0 ;
      RECT  32100.0 183150.0 30900.0 184350.0 ;
      RECT  34500.0 183150.0 33300.0 184350.0 ;
      RECT  29700.0 193050.0 28500.0 194250.0 ;
      RECT  29700.0 183150.0 28500.0 184350.0 ;
      RECT  33900.0 187800.0 32700.0 189000.0 ;
      RECT  33900.0 187800.0 32700.0 189000.0 ;
      RECT  31350.0 187950.0 30450.0 188850.0 ;
      RECT  36300.0 195150.0 26700.0 196050.0 ;
      RECT  36300.0 181350.0 26700.0 182250.0 ;
      RECT  29700.0 197550.0 28500.0 195600.0 ;
      RECT  29700.0 209400.0 28500.0 207450.0 ;
      RECT  34500.0 208050.0 33300.0 209850.0 ;
      RECT  34500.0 198750.0 33300.0 195150.0 ;
      RECT  31800.0 208050.0 30900.0 198750.0 ;
      RECT  34500.0 198750.0 33300.0 197550.0 ;
      RECT  32100.0 198750.0 30900.0 197550.0 ;
      RECT  32100.0 198750.0 30900.0 197550.0 ;
      RECT  34500.0 198750.0 33300.0 197550.0 ;
      RECT  34500.0 208050.0 33300.0 206850.0 ;
      RECT  32100.0 208050.0 30900.0 206850.0 ;
      RECT  32100.0 208050.0 30900.0 206850.0 ;
      RECT  34500.0 208050.0 33300.0 206850.0 ;
      RECT  29700.0 198150.0 28500.0 196950.0 ;
      RECT  29700.0 208050.0 28500.0 206850.0 ;
      RECT  33900.0 203400.0 32700.0 202200.0 ;
      RECT  33900.0 203400.0 32700.0 202200.0 ;
      RECT  31350.0 203250.0 30450.0 202350.0 ;
      RECT  36300.0 196050.0 26700.0 195150.0 ;
      RECT  36300.0 209850.0 26700.0 208950.0 ;
      RECT  48900.0 156150.0 47700.0 153750.0 ;
      RECT  48900.0 164850.0 47700.0 168450.0 ;
      RECT  44100.0 164850.0 42900.0 168450.0 ;
      RECT  41700.0 166050.0 40500.0 168000.0 ;
      RECT  41700.0 154200.0 40500.0 156150.0 ;
      RECT  48900.0 164850.0 47700.0 166050.0 ;
      RECT  46500.0 164850.0 45300.0 166050.0 ;
      RECT  46500.0 164850.0 45300.0 166050.0 ;
      RECT  48900.0 164850.0 47700.0 166050.0 ;
      RECT  46500.0 164850.0 45300.0 166050.0 ;
      RECT  44100.0 164850.0 42900.0 166050.0 ;
      RECT  44100.0 164850.0 42900.0 166050.0 ;
      RECT  46500.0 164850.0 45300.0 166050.0 ;
      RECT  48900.0 156150.0 47700.0 157350.0 ;
      RECT  46500.0 156150.0 45300.0 157350.0 ;
      RECT  46500.0 156150.0 45300.0 157350.0 ;
      RECT  48900.0 156150.0 47700.0 157350.0 ;
      RECT  46500.0 156150.0 45300.0 157350.0 ;
      RECT  44100.0 156150.0 42900.0 157350.0 ;
      RECT  44100.0 156150.0 42900.0 157350.0 ;
      RECT  46500.0 156150.0 45300.0 157350.0 ;
      RECT  41700.0 165450.0 40500.0 166650.0 ;
      RECT  41700.0 155550.0 40500.0 156750.0 ;
      RECT  44100.0 158700.0 45300.0 159900.0 ;
      RECT  47100.0 161400.0 48300.0 162600.0 ;
      RECT  46500.0 164850.0 45300.0 166050.0 ;
      RECT  44100.0 156150.0 42900.0 157350.0 ;
      RECT  42900.0 161400.0 44100.0 162600.0 ;
      RECT  48300.0 161400.0 47100.0 162600.0 ;
      RECT  45300.0 158700.0 44100.0 159900.0 ;
      RECT  44100.0 161400.0 42900.0 162600.0 ;
      RECT  50700.0 167550.0 36300.0 168450.0 ;
      RECT  50700.0 153750.0 36300.0 154650.0 ;
      RECT  48900.0 179850.0 47700.0 182250.0 ;
      RECT  48900.0 171150.0 47700.0 167550.0 ;
      RECT  44100.0 171150.0 42900.0 167550.0 ;
      RECT  41700.0 169950.0 40500.0 168000.0 ;
      RECT  41700.0 181800.0 40500.0 179850.0 ;
      RECT  48900.0 171150.0 47700.0 169950.0 ;
      RECT  46500.0 171150.0 45300.0 169950.0 ;
      RECT  46500.0 171150.0 45300.0 169950.0 ;
      RECT  48900.0 171150.0 47700.0 169950.0 ;
      RECT  46500.0 171150.0 45300.0 169950.0 ;
      RECT  44100.0 171150.0 42900.0 169950.0 ;
      RECT  44100.0 171150.0 42900.0 169950.0 ;
      RECT  46500.0 171150.0 45300.0 169950.0 ;
      RECT  48900.0 179850.0 47700.0 178650.0 ;
      RECT  46500.0 179850.0 45300.0 178650.0 ;
      RECT  46500.0 179850.0 45300.0 178650.0 ;
      RECT  48900.0 179850.0 47700.0 178650.0 ;
      RECT  46500.0 179850.0 45300.0 178650.0 ;
      RECT  44100.0 179850.0 42900.0 178650.0 ;
      RECT  44100.0 179850.0 42900.0 178650.0 ;
      RECT  46500.0 179850.0 45300.0 178650.0 ;
      RECT  41700.0 170550.0 40500.0 169350.0 ;
      RECT  41700.0 180450.0 40500.0 179250.0 ;
      RECT  44100.0 177300.0 45300.0 176100.0 ;
      RECT  47100.0 174600.0 48300.0 173400.0 ;
      RECT  46500.0 171150.0 45300.0 169950.0 ;
      RECT  44100.0 179850.0 42900.0 178650.0 ;
      RECT  42900.0 174600.0 44100.0 173400.0 ;
      RECT  48300.0 174600.0 47100.0 173400.0 ;
      RECT  45300.0 177300.0 44100.0 176100.0 ;
      RECT  44100.0 174600.0 42900.0 173400.0 ;
      RECT  50700.0 168450.0 36300.0 167550.0 ;
      RECT  50700.0 182250.0 36300.0 181350.0 ;
      RECT  48900.0 183750.0 47700.0 181350.0 ;
      RECT  48900.0 192450.0 47700.0 196050.0 ;
      RECT  44100.0 192450.0 42900.0 196050.0 ;
      RECT  41700.0 193650.0 40500.0 195600.0 ;
      RECT  41700.0 181800.0 40500.0 183750.0 ;
      RECT  48900.0 192450.0 47700.0 193650.0 ;
      RECT  46500.0 192450.0 45300.0 193650.0 ;
      RECT  46500.0 192450.0 45300.0 193650.0 ;
      RECT  48900.0 192450.0 47700.0 193650.0 ;
      RECT  46500.0 192450.0 45300.0 193650.0 ;
      RECT  44100.0 192450.0 42900.0 193650.0 ;
      RECT  44100.0 192450.0 42900.0 193650.0 ;
      RECT  46500.0 192450.0 45300.0 193650.0 ;
      RECT  48900.0 183750.0 47700.0 184950.0 ;
      RECT  46500.0 183750.0 45300.0 184950.0 ;
      RECT  46500.0 183750.0 45300.0 184950.0 ;
      RECT  48900.0 183750.0 47700.0 184950.0 ;
      RECT  46500.0 183750.0 45300.0 184950.0 ;
      RECT  44100.0 183750.0 42900.0 184950.0 ;
      RECT  44100.0 183750.0 42900.0 184950.0 ;
      RECT  46500.0 183750.0 45300.0 184950.0 ;
      RECT  41700.0 193050.0 40500.0 194250.0 ;
      RECT  41700.0 183150.0 40500.0 184350.0 ;
      RECT  44100.0 186300.0 45300.0 187500.0 ;
      RECT  47100.0 189000.0 48300.0 190200.0 ;
      RECT  46500.0 192450.0 45300.0 193650.0 ;
      RECT  44100.0 183750.0 42900.0 184950.0 ;
      RECT  42900.0 189000.0 44100.0 190200.0 ;
      RECT  48300.0 189000.0 47100.0 190200.0 ;
      RECT  45300.0 186300.0 44100.0 187500.0 ;
      RECT  44100.0 189000.0 42900.0 190200.0 ;
      RECT  50700.0 195150.0 36300.0 196050.0 ;
      RECT  50700.0 181350.0 36300.0 182250.0 ;
      RECT  48900.0 207450.0 47700.0 209850.0 ;
      RECT  48900.0 198750.0 47700.0 195150.0 ;
      RECT  44100.0 198750.0 42900.0 195150.0 ;
      RECT  41700.0 197550.0 40500.0 195600.0 ;
      RECT  41700.0 209400.0 40500.0 207450.0 ;
      RECT  48900.0 198750.0 47700.0 197550.0 ;
      RECT  46500.0 198750.0 45300.0 197550.0 ;
      RECT  46500.0 198750.0 45300.0 197550.0 ;
      RECT  48900.0 198750.0 47700.0 197550.0 ;
      RECT  46500.0 198750.0 45300.0 197550.0 ;
      RECT  44100.0 198750.0 42900.0 197550.0 ;
      RECT  44100.0 198750.0 42900.0 197550.0 ;
      RECT  46500.0 198750.0 45300.0 197550.0 ;
      RECT  48900.0 207450.0 47700.0 206250.0 ;
      RECT  46500.0 207450.0 45300.0 206250.0 ;
      RECT  46500.0 207450.0 45300.0 206250.0 ;
      RECT  48900.0 207450.0 47700.0 206250.0 ;
      RECT  46500.0 207450.0 45300.0 206250.0 ;
      RECT  44100.0 207450.0 42900.0 206250.0 ;
      RECT  44100.0 207450.0 42900.0 206250.0 ;
      RECT  46500.0 207450.0 45300.0 206250.0 ;
      RECT  41700.0 198150.0 40500.0 196950.0 ;
      RECT  41700.0 208050.0 40500.0 206850.0 ;
      RECT  44100.0 204900.0 45300.0 203700.0 ;
      RECT  47100.0 202200.0 48300.0 201000.0 ;
      RECT  46500.0 198750.0 45300.0 197550.0 ;
      RECT  44100.0 207450.0 42900.0 206250.0 ;
      RECT  42900.0 202200.0 44100.0 201000.0 ;
      RECT  48300.0 202200.0 47100.0 201000.0 ;
      RECT  45300.0 204900.0 44100.0 203700.0 ;
      RECT  44100.0 202200.0 42900.0 201000.0 ;
      RECT  50700.0 196050.0 36300.0 195150.0 ;
      RECT  50700.0 209850.0 36300.0 208950.0 ;
      RECT  61650.0 164700.0 62850.0 165900.0 ;
      RECT  80250.0 160200.0 81450.0 161400.0 ;
      RECT  58650.0 178500.0 59850.0 179700.0 ;
      RECT  77250.0 174600.0 78450.0 175800.0 ;
      RECT  80250.0 183300.0 81450.0 184500.0 ;
      RECT  55650.0 183300.0 56850.0 184500.0 ;
      RECT  77250.0 197100.0 78450.0 198300.0 ;
      RECT  52650.0 197100.0 53850.0 198300.0 ;
      RECT  61650.0 161400.0 62850.0 162600.0 ;
      RECT  58650.0 158700.0 59850.0 159900.0 ;
      RECT  55650.0 173400.0 56850.0 174600.0 ;
      RECT  58650.0 176100.0 59850.0 177300.0 ;
      RECT  61650.0 189000.0 62850.0 190200.0 ;
      RECT  52650.0 186300.0 53850.0 187500.0 ;
      RECT  55650.0 201000.0 56850.0 202200.0 ;
      RECT  52650.0 203700.0 53850.0 204900.0 ;
      RECT  30450.0 160350.0 26700.0 161250.0 ;
      RECT  30450.0 174750.0 26700.0 175650.0 ;
      RECT  30450.0 187950.0 26700.0 188850.0 ;
      RECT  30450.0 202350.0 26700.0 203250.0 ;
      RECT  81300.0 167550.0 26700.0 168450.0 ;
      RECT  81300.0 195150.0 26700.0 196050.0 ;
      RECT  81300.0 153750.0 26700.0 154650.0 ;
      RECT  81300.0 181350.0 26700.0 182250.0 ;
      RECT  81300.0 208950.0 26700.0 209850.0 ;
      RECT  28500.0 211350.0 29700.0 208950.0 ;
      RECT  28500.0 220050.0 29700.0 223650.0 ;
      RECT  33300.0 220050.0 34500.0 223650.0 ;
      RECT  35700.0 221250.0 36900.0 223200.0 ;
      RECT  35700.0 209400.0 36900.0 211350.0 ;
      RECT  28500.0 220050.0 29700.0 221250.0 ;
      RECT  30900.0 220050.0 32100.0 221250.0 ;
      RECT  30900.0 220050.0 32100.0 221250.0 ;
      RECT  28500.0 220050.0 29700.0 221250.0 ;
      RECT  30900.0 220050.0 32100.0 221250.0 ;
      RECT  33300.0 220050.0 34500.0 221250.0 ;
      RECT  33300.0 220050.0 34500.0 221250.0 ;
      RECT  30900.0 220050.0 32100.0 221250.0 ;
      RECT  28500.0 211350.0 29700.0 212550.0 ;
      RECT  30900.0 211350.0 32100.0 212550.0 ;
      RECT  30900.0 211350.0 32100.0 212550.0 ;
      RECT  28500.0 211350.0 29700.0 212550.0 ;
      RECT  30900.0 211350.0 32100.0 212550.0 ;
      RECT  33300.0 211350.0 34500.0 212550.0 ;
      RECT  33300.0 211350.0 34500.0 212550.0 ;
      RECT  30900.0 211350.0 32100.0 212550.0 ;
      RECT  35700.0 220650.0 36900.0 221850.0 ;
      RECT  35700.0 210750.0 36900.0 211950.0 ;
      RECT  33300.0 213900.0 32100.0 215100.0 ;
      RECT  30300.0 216600.0 29100.0 217800.0 ;
      RECT  30900.0 220050.0 32100.0 221250.0 ;
      RECT  33300.0 211350.0 34500.0 212550.0 ;
      RECT  34500.0 216600.0 33300.0 217800.0 ;
      RECT  29100.0 216600.0 30300.0 217800.0 ;
      RECT  32100.0 213900.0 33300.0 215100.0 ;
      RECT  33300.0 216600.0 34500.0 217800.0 ;
      RECT  26700.0 222750.0 41100.0 223650.0 ;
      RECT  26700.0 208950.0 41100.0 209850.0 ;
      RECT  28500.0 235050.0 29700.0 237450.0 ;
      RECT  28500.0 226350.0 29700.0 222750.0 ;
      RECT  33300.0 226350.0 34500.0 222750.0 ;
      RECT  35700.0 225150.0 36900.0 223200.0 ;
      RECT  35700.0 237000.0 36900.0 235050.0 ;
      RECT  28500.0 226350.0 29700.0 225150.0 ;
      RECT  30900.0 226350.0 32100.0 225150.0 ;
      RECT  30900.0 226350.0 32100.0 225150.0 ;
      RECT  28500.0 226350.0 29700.0 225150.0 ;
      RECT  30900.0 226350.0 32100.0 225150.0 ;
      RECT  33300.0 226350.0 34500.0 225150.0 ;
      RECT  33300.0 226350.0 34500.0 225150.0 ;
      RECT  30900.0 226350.0 32100.0 225150.0 ;
      RECT  28500.0 235050.0 29700.0 233850.0 ;
      RECT  30900.0 235050.0 32100.0 233850.0 ;
      RECT  30900.0 235050.0 32100.0 233850.0 ;
      RECT  28500.0 235050.0 29700.0 233850.0 ;
      RECT  30900.0 235050.0 32100.0 233850.0 ;
      RECT  33300.0 235050.0 34500.0 233850.0 ;
      RECT  33300.0 235050.0 34500.0 233850.0 ;
      RECT  30900.0 235050.0 32100.0 233850.0 ;
      RECT  35700.0 225750.0 36900.0 224550.0 ;
      RECT  35700.0 235650.0 36900.0 234450.0 ;
      RECT  33300.0 232500.0 32100.0 231300.0 ;
      RECT  30300.0 229800.0 29100.0 228600.0 ;
      RECT  30900.0 226350.0 32100.0 225150.0 ;
      RECT  33300.0 235050.0 34500.0 233850.0 ;
      RECT  34500.0 229800.0 33300.0 228600.0 ;
      RECT  29100.0 229800.0 30300.0 228600.0 ;
      RECT  32100.0 232500.0 33300.0 231300.0 ;
      RECT  33300.0 229800.0 34500.0 228600.0 ;
      RECT  26700.0 223650.0 41100.0 222750.0 ;
      RECT  26700.0 237450.0 41100.0 236550.0 ;
      RECT  28500.0 238950.0 29700.0 236550.0 ;
      RECT  28500.0 247650.0 29700.0 251250.0 ;
      RECT  33300.0 247650.0 34500.0 251250.0 ;
      RECT  35700.0 248850.0 36900.0 250800.0 ;
      RECT  35700.0 237000.0 36900.0 238950.0 ;
      RECT  28500.0 247650.0 29700.0 248850.0 ;
      RECT  30900.0 247650.0 32100.0 248850.0 ;
      RECT  30900.0 247650.0 32100.0 248850.0 ;
      RECT  28500.0 247650.0 29700.0 248850.0 ;
      RECT  30900.0 247650.0 32100.0 248850.0 ;
      RECT  33300.0 247650.0 34500.0 248850.0 ;
      RECT  33300.0 247650.0 34500.0 248850.0 ;
      RECT  30900.0 247650.0 32100.0 248850.0 ;
      RECT  28500.0 238950.0 29700.0 240150.0 ;
      RECT  30900.0 238950.0 32100.0 240150.0 ;
      RECT  30900.0 238950.0 32100.0 240150.0 ;
      RECT  28500.0 238950.0 29700.0 240150.0 ;
      RECT  30900.0 238950.0 32100.0 240150.0 ;
      RECT  33300.0 238950.0 34500.0 240150.0 ;
      RECT  33300.0 238950.0 34500.0 240150.0 ;
      RECT  30900.0 238950.0 32100.0 240150.0 ;
      RECT  35700.0 248250.0 36900.0 249450.0 ;
      RECT  35700.0 238350.0 36900.0 239550.0 ;
      RECT  33300.0 241500.0 32100.0 242700.0 ;
      RECT  30300.0 244200.0 29100.0 245400.0 ;
      RECT  30900.0 247650.0 32100.0 248850.0 ;
      RECT  33300.0 238950.0 34500.0 240150.0 ;
      RECT  34500.0 244200.0 33300.0 245400.0 ;
      RECT  29100.0 244200.0 30300.0 245400.0 ;
      RECT  32100.0 241500.0 33300.0 242700.0 ;
      RECT  33300.0 244200.0 34500.0 245400.0 ;
      RECT  26700.0 250350.0 41100.0 251250.0 ;
      RECT  26700.0 236550.0 41100.0 237450.0 ;
      RECT  28500.0 262650.0 29700.0 265050.0 ;
      RECT  28500.0 253950.0 29700.0 250350.0 ;
      RECT  33300.0 253950.0 34500.0 250350.0 ;
      RECT  35700.0 252750.0 36900.0 250800.0 ;
      RECT  35700.0 264600.0 36900.0 262650.0 ;
      RECT  28500.0 253950.0 29700.0 252750.0 ;
      RECT  30900.0 253950.0 32100.0 252750.0 ;
      RECT  30900.0 253950.0 32100.0 252750.0 ;
      RECT  28500.0 253950.0 29700.0 252750.0 ;
      RECT  30900.0 253950.0 32100.0 252750.0 ;
      RECT  33300.0 253950.0 34500.0 252750.0 ;
      RECT  33300.0 253950.0 34500.0 252750.0 ;
      RECT  30900.0 253950.0 32100.0 252750.0 ;
      RECT  28500.0 262650.0 29700.0 261450.0 ;
      RECT  30900.0 262650.0 32100.0 261450.0 ;
      RECT  30900.0 262650.0 32100.0 261450.0 ;
      RECT  28500.0 262650.0 29700.0 261450.0 ;
      RECT  30900.0 262650.0 32100.0 261450.0 ;
      RECT  33300.0 262650.0 34500.0 261450.0 ;
      RECT  33300.0 262650.0 34500.0 261450.0 ;
      RECT  30900.0 262650.0 32100.0 261450.0 ;
      RECT  35700.0 253350.0 36900.0 252150.0 ;
      RECT  35700.0 263250.0 36900.0 262050.0 ;
      RECT  33300.0 260100.0 32100.0 258900.0 ;
      RECT  30300.0 257400.0 29100.0 256200.0 ;
      RECT  30900.0 253950.0 32100.0 252750.0 ;
      RECT  33300.0 262650.0 34500.0 261450.0 ;
      RECT  34500.0 257400.0 33300.0 256200.0 ;
      RECT  29100.0 257400.0 30300.0 256200.0 ;
      RECT  32100.0 260100.0 33300.0 258900.0 ;
      RECT  33300.0 257400.0 34500.0 256200.0 ;
      RECT  26700.0 251250.0 41100.0 250350.0 ;
      RECT  26700.0 265050.0 41100.0 264150.0 ;
      RECT  28500.0 266550.0 29700.0 264150.0 ;
      RECT  28500.0 275250.0 29700.0 278850.0 ;
      RECT  33300.0 275250.0 34500.0 278850.0 ;
      RECT  35700.0 276450.0 36900.0 278400.0 ;
      RECT  35700.0 264600.0 36900.0 266550.0 ;
      RECT  28500.0 275250.0 29700.0 276450.0 ;
      RECT  30900.0 275250.0 32100.0 276450.0 ;
      RECT  30900.0 275250.0 32100.0 276450.0 ;
      RECT  28500.0 275250.0 29700.0 276450.0 ;
      RECT  30900.0 275250.0 32100.0 276450.0 ;
      RECT  33300.0 275250.0 34500.0 276450.0 ;
      RECT  33300.0 275250.0 34500.0 276450.0 ;
      RECT  30900.0 275250.0 32100.0 276450.0 ;
      RECT  28500.0 266550.0 29700.0 267750.0 ;
      RECT  30900.0 266550.0 32100.0 267750.0 ;
      RECT  30900.0 266550.0 32100.0 267750.0 ;
      RECT  28500.0 266550.0 29700.0 267750.0 ;
      RECT  30900.0 266550.0 32100.0 267750.0 ;
      RECT  33300.0 266550.0 34500.0 267750.0 ;
      RECT  33300.0 266550.0 34500.0 267750.0 ;
      RECT  30900.0 266550.0 32100.0 267750.0 ;
      RECT  35700.0 275850.0 36900.0 277050.0 ;
      RECT  35700.0 265950.0 36900.0 267150.0 ;
      RECT  33300.0 269100.0 32100.0 270300.0 ;
      RECT  30300.0 271800.0 29100.0 273000.0 ;
      RECT  30900.0 275250.0 32100.0 276450.0 ;
      RECT  33300.0 266550.0 34500.0 267750.0 ;
      RECT  34500.0 271800.0 33300.0 273000.0 ;
      RECT  29100.0 271800.0 30300.0 273000.0 ;
      RECT  32100.0 269100.0 33300.0 270300.0 ;
      RECT  33300.0 271800.0 34500.0 273000.0 ;
      RECT  26700.0 277950.0 41100.0 278850.0 ;
      RECT  26700.0 264150.0 41100.0 265050.0 ;
      RECT  28500.0 290250.0 29700.0 292650.0 ;
      RECT  28500.0 281550.0 29700.0 277950.0 ;
      RECT  33300.0 281550.0 34500.0 277950.0 ;
      RECT  35700.0 280350.0 36900.0 278400.0 ;
      RECT  35700.0 292200.0 36900.0 290250.0 ;
      RECT  28500.0 281550.0 29700.0 280350.0 ;
      RECT  30900.0 281550.0 32100.0 280350.0 ;
      RECT  30900.0 281550.0 32100.0 280350.0 ;
      RECT  28500.0 281550.0 29700.0 280350.0 ;
      RECT  30900.0 281550.0 32100.0 280350.0 ;
      RECT  33300.0 281550.0 34500.0 280350.0 ;
      RECT  33300.0 281550.0 34500.0 280350.0 ;
      RECT  30900.0 281550.0 32100.0 280350.0 ;
      RECT  28500.0 290250.0 29700.0 289050.0 ;
      RECT  30900.0 290250.0 32100.0 289050.0 ;
      RECT  30900.0 290250.0 32100.0 289050.0 ;
      RECT  28500.0 290250.0 29700.0 289050.0 ;
      RECT  30900.0 290250.0 32100.0 289050.0 ;
      RECT  33300.0 290250.0 34500.0 289050.0 ;
      RECT  33300.0 290250.0 34500.0 289050.0 ;
      RECT  30900.0 290250.0 32100.0 289050.0 ;
      RECT  35700.0 280950.0 36900.0 279750.0 ;
      RECT  35700.0 290850.0 36900.0 289650.0 ;
      RECT  33300.0 287700.0 32100.0 286500.0 ;
      RECT  30300.0 285000.0 29100.0 283800.0 ;
      RECT  30900.0 281550.0 32100.0 280350.0 ;
      RECT  33300.0 290250.0 34500.0 289050.0 ;
      RECT  34500.0 285000.0 33300.0 283800.0 ;
      RECT  29100.0 285000.0 30300.0 283800.0 ;
      RECT  32100.0 287700.0 33300.0 286500.0 ;
      RECT  33300.0 285000.0 34500.0 283800.0 ;
      RECT  26700.0 278850.0 41100.0 277950.0 ;
      RECT  26700.0 292650.0 41100.0 291750.0 ;
      RECT  28500.0 294150.0 29700.0 291750.0 ;
      RECT  28500.0 302850.0 29700.0 306450.0 ;
      RECT  33300.0 302850.0 34500.0 306450.0 ;
      RECT  35700.0 304050.0 36900.0 306000.0 ;
      RECT  35700.0 292200.0 36900.0 294150.0 ;
      RECT  28500.0 302850.0 29700.0 304050.0 ;
      RECT  30900.0 302850.0 32100.0 304050.0 ;
      RECT  30900.0 302850.0 32100.0 304050.0 ;
      RECT  28500.0 302850.0 29700.0 304050.0 ;
      RECT  30900.0 302850.0 32100.0 304050.0 ;
      RECT  33300.0 302850.0 34500.0 304050.0 ;
      RECT  33300.0 302850.0 34500.0 304050.0 ;
      RECT  30900.0 302850.0 32100.0 304050.0 ;
      RECT  28500.0 294150.0 29700.0 295350.0 ;
      RECT  30900.0 294150.0 32100.0 295350.0 ;
      RECT  30900.0 294150.0 32100.0 295350.0 ;
      RECT  28500.0 294150.0 29700.0 295350.0 ;
      RECT  30900.0 294150.0 32100.0 295350.0 ;
      RECT  33300.0 294150.0 34500.0 295350.0 ;
      RECT  33300.0 294150.0 34500.0 295350.0 ;
      RECT  30900.0 294150.0 32100.0 295350.0 ;
      RECT  35700.0 303450.0 36900.0 304650.0 ;
      RECT  35700.0 293550.0 36900.0 294750.0 ;
      RECT  33300.0 296700.0 32100.0 297900.0 ;
      RECT  30300.0 299400.0 29100.0 300600.0 ;
      RECT  30900.0 302850.0 32100.0 304050.0 ;
      RECT  33300.0 294150.0 34500.0 295350.0 ;
      RECT  34500.0 299400.0 33300.0 300600.0 ;
      RECT  29100.0 299400.0 30300.0 300600.0 ;
      RECT  32100.0 296700.0 33300.0 297900.0 ;
      RECT  33300.0 299400.0 34500.0 300600.0 ;
      RECT  26700.0 305550.0 41100.0 306450.0 ;
      RECT  26700.0 291750.0 41100.0 292650.0 ;
      RECT  28500.0 317850.0 29700.0 320250.0 ;
      RECT  28500.0 309150.0 29700.0 305550.0 ;
      RECT  33300.0 309150.0 34500.0 305550.0 ;
      RECT  35700.0 307950.0 36900.0 306000.0 ;
      RECT  35700.0 319800.0 36900.0 317850.0 ;
      RECT  28500.0 309150.0 29700.0 307950.0 ;
      RECT  30900.0 309150.0 32100.0 307950.0 ;
      RECT  30900.0 309150.0 32100.0 307950.0 ;
      RECT  28500.0 309150.0 29700.0 307950.0 ;
      RECT  30900.0 309150.0 32100.0 307950.0 ;
      RECT  33300.0 309150.0 34500.0 307950.0 ;
      RECT  33300.0 309150.0 34500.0 307950.0 ;
      RECT  30900.0 309150.0 32100.0 307950.0 ;
      RECT  28500.0 317850.0 29700.0 316650.0 ;
      RECT  30900.0 317850.0 32100.0 316650.0 ;
      RECT  30900.0 317850.0 32100.0 316650.0 ;
      RECT  28500.0 317850.0 29700.0 316650.0 ;
      RECT  30900.0 317850.0 32100.0 316650.0 ;
      RECT  33300.0 317850.0 34500.0 316650.0 ;
      RECT  33300.0 317850.0 34500.0 316650.0 ;
      RECT  30900.0 317850.0 32100.0 316650.0 ;
      RECT  35700.0 308550.0 36900.0 307350.0 ;
      RECT  35700.0 318450.0 36900.0 317250.0 ;
      RECT  33300.0 315300.0 32100.0 314100.0 ;
      RECT  30300.0 312600.0 29100.0 311400.0 ;
      RECT  30900.0 309150.0 32100.0 307950.0 ;
      RECT  33300.0 317850.0 34500.0 316650.0 ;
      RECT  34500.0 312600.0 33300.0 311400.0 ;
      RECT  29100.0 312600.0 30300.0 311400.0 ;
      RECT  32100.0 315300.0 33300.0 314100.0 ;
      RECT  33300.0 312600.0 34500.0 311400.0 ;
      RECT  26700.0 306450.0 41100.0 305550.0 ;
      RECT  26700.0 320250.0 41100.0 319350.0 ;
      RECT  28500.0 321750.0 29700.0 319350.0 ;
      RECT  28500.0 330450.0 29700.0 334050.0 ;
      RECT  33300.0 330450.0 34500.0 334050.0 ;
      RECT  35700.0 331650.0 36900.0 333600.0 ;
      RECT  35700.0 319800.0 36900.0 321750.0 ;
      RECT  28500.0 330450.0 29700.0 331650.0 ;
      RECT  30900.0 330450.0 32100.0 331650.0 ;
      RECT  30900.0 330450.0 32100.0 331650.0 ;
      RECT  28500.0 330450.0 29700.0 331650.0 ;
      RECT  30900.0 330450.0 32100.0 331650.0 ;
      RECT  33300.0 330450.0 34500.0 331650.0 ;
      RECT  33300.0 330450.0 34500.0 331650.0 ;
      RECT  30900.0 330450.0 32100.0 331650.0 ;
      RECT  28500.0 321750.0 29700.0 322950.0 ;
      RECT  30900.0 321750.0 32100.0 322950.0 ;
      RECT  30900.0 321750.0 32100.0 322950.0 ;
      RECT  28500.0 321750.0 29700.0 322950.0 ;
      RECT  30900.0 321750.0 32100.0 322950.0 ;
      RECT  33300.0 321750.0 34500.0 322950.0 ;
      RECT  33300.0 321750.0 34500.0 322950.0 ;
      RECT  30900.0 321750.0 32100.0 322950.0 ;
      RECT  35700.0 331050.0 36900.0 332250.0 ;
      RECT  35700.0 321150.0 36900.0 322350.0 ;
      RECT  33300.0 324300.0 32100.0 325500.0 ;
      RECT  30300.0 327000.0 29100.0 328200.0 ;
      RECT  30900.0 330450.0 32100.0 331650.0 ;
      RECT  33300.0 321750.0 34500.0 322950.0 ;
      RECT  34500.0 327000.0 33300.0 328200.0 ;
      RECT  29100.0 327000.0 30300.0 328200.0 ;
      RECT  32100.0 324300.0 33300.0 325500.0 ;
      RECT  33300.0 327000.0 34500.0 328200.0 ;
      RECT  26700.0 333150.0 41100.0 334050.0 ;
      RECT  26700.0 319350.0 41100.0 320250.0 ;
      RECT  28500.0 345450.0 29700.0 347850.0 ;
      RECT  28500.0 336750.0 29700.0 333150.0 ;
      RECT  33300.0 336750.0 34500.0 333150.0 ;
      RECT  35700.0 335550.0 36900.0 333600.0 ;
      RECT  35700.0 347400.0 36900.0 345450.0 ;
      RECT  28500.0 336750.0 29700.0 335550.0 ;
      RECT  30900.0 336750.0 32100.0 335550.0 ;
      RECT  30900.0 336750.0 32100.0 335550.0 ;
      RECT  28500.0 336750.0 29700.0 335550.0 ;
      RECT  30900.0 336750.0 32100.0 335550.0 ;
      RECT  33300.0 336750.0 34500.0 335550.0 ;
      RECT  33300.0 336750.0 34500.0 335550.0 ;
      RECT  30900.0 336750.0 32100.0 335550.0 ;
      RECT  28500.0 345450.0 29700.0 344250.0 ;
      RECT  30900.0 345450.0 32100.0 344250.0 ;
      RECT  30900.0 345450.0 32100.0 344250.0 ;
      RECT  28500.0 345450.0 29700.0 344250.0 ;
      RECT  30900.0 345450.0 32100.0 344250.0 ;
      RECT  33300.0 345450.0 34500.0 344250.0 ;
      RECT  33300.0 345450.0 34500.0 344250.0 ;
      RECT  30900.0 345450.0 32100.0 344250.0 ;
      RECT  35700.0 336150.0 36900.0 334950.0 ;
      RECT  35700.0 346050.0 36900.0 344850.0 ;
      RECT  33300.0 342900.0 32100.0 341700.0 ;
      RECT  30300.0 340200.0 29100.0 339000.0 ;
      RECT  30900.0 336750.0 32100.0 335550.0 ;
      RECT  33300.0 345450.0 34500.0 344250.0 ;
      RECT  34500.0 340200.0 33300.0 339000.0 ;
      RECT  29100.0 340200.0 30300.0 339000.0 ;
      RECT  32100.0 342900.0 33300.0 341700.0 ;
      RECT  33300.0 340200.0 34500.0 339000.0 ;
      RECT  26700.0 334050.0 41100.0 333150.0 ;
      RECT  26700.0 347850.0 41100.0 346950.0 ;
      RECT  28500.0 349350.0 29700.0 346950.0 ;
      RECT  28500.0 358050.0 29700.0 361650.0 ;
      RECT  33300.0 358050.0 34500.0 361650.0 ;
      RECT  35700.0 359250.0 36900.0 361200.0 ;
      RECT  35700.0 347400.0 36900.0 349350.0 ;
      RECT  28500.0 358050.0 29700.0 359250.0 ;
      RECT  30900.0 358050.0 32100.0 359250.0 ;
      RECT  30900.0 358050.0 32100.0 359250.0 ;
      RECT  28500.0 358050.0 29700.0 359250.0 ;
      RECT  30900.0 358050.0 32100.0 359250.0 ;
      RECT  33300.0 358050.0 34500.0 359250.0 ;
      RECT  33300.0 358050.0 34500.0 359250.0 ;
      RECT  30900.0 358050.0 32100.0 359250.0 ;
      RECT  28500.0 349350.0 29700.0 350550.0 ;
      RECT  30900.0 349350.0 32100.0 350550.0 ;
      RECT  30900.0 349350.0 32100.0 350550.0 ;
      RECT  28500.0 349350.0 29700.0 350550.0 ;
      RECT  30900.0 349350.0 32100.0 350550.0 ;
      RECT  33300.0 349350.0 34500.0 350550.0 ;
      RECT  33300.0 349350.0 34500.0 350550.0 ;
      RECT  30900.0 349350.0 32100.0 350550.0 ;
      RECT  35700.0 358650.0 36900.0 359850.0 ;
      RECT  35700.0 348750.0 36900.0 349950.0 ;
      RECT  33300.0 351900.0 32100.0 353100.0 ;
      RECT  30300.0 354600.0 29100.0 355800.0 ;
      RECT  30900.0 358050.0 32100.0 359250.0 ;
      RECT  33300.0 349350.0 34500.0 350550.0 ;
      RECT  34500.0 354600.0 33300.0 355800.0 ;
      RECT  29100.0 354600.0 30300.0 355800.0 ;
      RECT  32100.0 351900.0 33300.0 353100.0 ;
      RECT  33300.0 354600.0 34500.0 355800.0 ;
      RECT  26700.0 360750.0 41100.0 361650.0 ;
      RECT  26700.0 346950.0 41100.0 347850.0 ;
      RECT  28500.0 373050.0 29700.0 375450.0 ;
      RECT  28500.0 364350.0 29700.0 360750.0 ;
      RECT  33300.0 364350.0 34500.0 360750.0 ;
      RECT  35700.0 363150.0 36900.0 361200.0 ;
      RECT  35700.0 375000.0 36900.0 373050.0 ;
      RECT  28500.0 364350.0 29700.0 363150.0 ;
      RECT  30900.0 364350.0 32100.0 363150.0 ;
      RECT  30900.0 364350.0 32100.0 363150.0 ;
      RECT  28500.0 364350.0 29700.0 363150.0 ;
      RECT  30900.0 364350.0 32100.0 363150.0 ;
      RECT  33300.0 364350.0 34500.0 363150.0 ;
      RECT  33300.0 364350.0 34500.0 363150.0 ;
      RECT  30900.0 364350.0 32100.0 363150.0 ;
      RECT  28500.0 373050.0 29700.0 371850.0 ;
      RECT  30900.0 373050.0 32100.0 371850.0 ;
      RECT  30900.0 373050.0 32100.0 371850.0 ;
      RECT  28500.0 373050.0 29700.0 371850.0 ;
      RECT  30900.0 373050.0 32100.0 371850.0 ;
      RECT  33300.0 373050.0 34500.0 371850.0 ;
      RECT  33300.0 373050.0 34500.0 371850.0 ;
      RECT  30900.0 373050.0 32100.0 371850.0 ;
      RECT  35700.0 363750.0 36900.0 362550.0 ;
      RECT  35700.0 373650.0 36900.0 372450.0 ;
      RECT  33300.0 370500.0 32100.0 369300.0 ;
      RECT  30300.0 367800.0 29100.0 366600.0 ;
      RECT  30900.0 364350.0 32100.0 363150.0 ;
      RECT  33300.0 373050.0 34500.0 371850.0 ;
      RECT  34500.0 367800.0 33300.0 366600.0 ;
      RECT  29100.0 367800.0 30300.0 366600.0 ;
      RECT  32100.0 370500.0 33300.0 369300.0 ;
      RECT  33300.0 367800.0 34500.0 366600.0 ;
      RECT  26700.0 361650.0 41100.0 360750.0 ;
      RECT  26700.0 375450.0 41100.0 374550.0 ;
      RECT  28500.0 376950.0 29700.0 374550.0 ;
      RECT  28500.0 385650.0 29700.0 389250.0 ;
      RECT  33300.0 385650.0 34500.0 389250.0 ;
      RECT  35700.0 386850.0 36900.0 388800.0 ;
      RECT  35700.0 375000.0 36900.0 376950.0 ;
      RECT  28500.0 385650.0 29700.0 386850.0 ;
      RECT  30900.0 385650.0 32100.0 386850.0 ;
      RECT  30900.0 385650.0 32100.0 386850.0 ;
      RECT  28500.0 385650.0 29700.0 386850.0 ;
      RECT  30900.0 385650.0 32100.0 386850.0 ;
      RECT  33300.0 385650.0 34500.0 386850.0 ;
      RECT  33300.0 385650.0 34500.0 386850.0 ;
      RECT  30900.0 385650.0 32100.0 386850.0 ;
      RECT  28500.0 376950.0 29700.0 378150.0 ;
      RECT  30900.0 376950.0 32100.0 378150.0 ;
      RECT  30900.0 376950.0 32100.0 378150.0 ;
      RECT  28500.0 376950.0 29700.0 378150.0 ;
      RECT  30900.0 376950.0 32100.0 378150.0 ;
      RECT  33300.0 376950.0 34500.0 378150.0 ;
      RECT  33300.0 376950.0 34500.0 378150.0 ;
      RECT  30900.0 376950.0 32100.0 378150.0 ;
      RECT  35700.0 386250.0 36900.0 387450.0 ;
      RECT  35700.0 376350.0 36900.0 377550.0 ;
      RECT  33300.0 379500.0 32100.0 380700.0 ;
      RECT  30300.0 382200.0 29100.0 383400.0 ;
      RECT  30900.0 385650.0 32100.0 386850.0 ;
      RECT  33300.0 376950.0 34500.0 378150.0 ;
      RECT  34500.0 382200.0 33300.0 383400.0 ;
      RECT  29100.0 382200.0 30300.0 383400.0 ;
      RECT  32100.0 379500.0 33300.0 380700.0 ;
      RECT  33300.0 382200.0 34500.0 383400.0 ;
      RECT  26700.0 388350.0 41100.0 389250.0 ;
      RECT  26700.0 374550.0 41100.0 375450.0 ;
      RECT  28500.0 400650.0 29700.0 403050.0 ;
      RECT  28500.0 391950.0 29700.0 388350.0 ;
      RECT  33300.0 391950.0 34500.0 388350.0 ;
      RECT  35700.0 390750.0 36900.0 388800.0 ;
      RECT  35700.0 402600.0 36900.0 400650.0 ;
      RECT  28500.0 391950.0 29700.0 390750.0 ;
      RECT  30900.0 391950.0 32100.0 390750.0 ;
      RECT  30900.0 391950.0 32100.0 390750.0 ;
      RECT  28500.0 391950.0 29700.0 390750.0 ;
      RECT  30900.0 391950.0 32100.0 390750.0 ;
      RECT  33300.0 391950.0 34500.0 390750.0 ;
      RECT  33300.0 391950.0 34500.0 390750.0 ;
      RECT  30900.0 391950.0 32100.0 390750.0 ;
      RECT  28500.0 400650.0 29700.0 399450.0 ;
      RECT  30900.0 400650.0 32100.0 399450.0 ;
      RECT  30900.0 400650.0 32100.0 399450.0 ;
      RECT  28500.0 400650.0 29700.0 399450.0 ;
      RECT  30900.0 400650.0 32100.0 399450.0 ;
      RECT  33300.0 400650.0 34500.0 399450.0 ;
      RECT  33300.0 400650.0 34500.0 399450.0 ;
      RECT  30900.0 400650.0 32100.0 399450.0 ;
      RECT  35700.0 391350.0 36900.0 390150.0 ;
      RECT  35700.0 401250.0 36900.0 400050.0 ;
      RECT  33300.0 398100.0 32100.0 396900.0 ;
      RECT  30300.0 395400.0 29100.0 394200.0 ;
      RECT  30900.0 391950.0 32100.0 390750.0 ;
      RECT  33300.0 400650.0 34500.0 399450.0 ;
      RECT  34500.0 395400.0 33300.0 394200.0 ;
      RECT  29100.0 395400.0 30300.0 394200.0 ;
      RECT  32100.0 398100.0 33300.0 396900.0 ;
      RECT  33300.0 395400.0 34500.0 394200.0 ;
      RECT  26700.0 389250.0 41100.0 388350.0 ;
      RECT  26700.0 403050.0 41100.0 402150.0 ;
      RECT  28500.0 404550.0 29700.0 402150.0 ;
      RECT  28500.0 413250.0 29700.0 416850.0 ;
      RECT  33300.0 413250.0 34500.0 416850.0 ;
      RECT  35700.0 414450.0 36900.0 416400.0 ;
      RECT  35700.0 402600.0 36900.0 404550.0 ;
      RECT  28500.0 413250.0 29700.0 414450.0 ;
      RECT  30900.0 413250.0 32100.0 414450.0 ;
      RECT  30900.0 413250.0 32100.0 414450.0 ;
      RECT  28500.0 413250.0 29700.0 414450.0 ;
      RECT  30900.0 413250.0 32100.0 414450.0 ;
      RECT  33300.0 413250.0 34500.0 414450.0 ;
      RECT  33300.0 413250.0 34500.0 414450.0 ;
      RECT  30900.0 413250.0 32100.0 414450.0 ;
      RECT  28500.0 404550.0 29700.0 405750.0 ;
      RECT  30900.0 404550.0 32100.0 405750.0 ;
      RECT  30900.0 404550.0 32100.0 405750.0 ;
      RECT  28500.0 404550.0 29700.0 405750.0 ;
      RECT  30900.0 404550.0 32100.0 405750.0 ;
      RECT  33300.0 404550.0 34500.0 405750.0 ;
      RECT  33300.0 404550.0 34500.0 405750.0 ;
      RECT  30900.0 404550.0 32100.0 405750.0 ;
      RECT  35700.0 413850.0 36900.0 415050.0 ;
      RECT  35700.0 403950.0 36900.0 405150.0 ;
      RECT  33300.0 407100.0 32100.0 408300.0 ;
      RECT  30300.0 409800.0 29100.0 411000.0 ;
      RECT  30900.0 413250.0 32100.0 414450.0 ;
      RECT  33300.0 404550.0 34500.0 405750.0 ;
      RECT  34500.0 409800.0 33300.0 411000.0 ;
      RECT  29100.0 409800.0 30300.0 411000.0 ;
      RECT  32100.0 407100.0 33300.0 408300.0 ;
      RECT  33300.0 409800.0 34500.0 411000.0 ;
      RECT  26700.0 415950.0 41100.0 416850.0 ;
      RECT  26700.0 402150.0 41100.0 403050.0 ;
      RECT  28500.0 428250.0 29700.0 430650.0 ;
      RECT  28500.0 419550.0 29700.0 415950.0 ;
      RECT  33300.0 419550.0 34500.0 415950.0 ;
      RECT  35700.0 418350.0 36900.0 416400.0 ;
      RECT  35700.0 430200.0 36900.0 428250.0 ;
      RECT  28500.0 419550.0 29700.0 418350.0 ;
      RECT  30900.0 419550.0 32100.0 418350.0 ;
      RECT  30900.0 419550.0 32100.0 418350.0 ;
      RECT  28500.0 419550.0 29700.0 418350.0 ;
      RECT  30900.0 419550.0 32100.0 418350.0 ;
      RECT  33300.0 419550.0 34500.0 418350.0 ;
      RECT  33300.0 419550.0 34500.0 418350.0 ;
      RECT  30900.0 419550.0 32100.0 418350.0 ;
      RECT  28500.0 428250.0 29700.0 427050.0 ;
      RECT  30900.0 428250.0 32100.0 427050.0 ;
      RECT  30900.0 428250.0 32100.0 427050.0 ;
      RECT  28500.0 428250.0 29700.0 427050.0 ;
      RECT  30900.0 428250.0 32100.0 427050.0 ;
      RECT  33300.0 428250.0 34500.0 427050.0 ;
      RECT  33300.0 428250.0 34500.0 427050.0 ;
      RECT  30900.0 428250.0 32100.0 427050.0 ;
      RECT  35700.0 418950.0 36900.0 417750.0 ;
      RECT  35700.0 428850.0 36900.0 427650.0 ;
      RECT  33300.0 425700.0 32100.0 424500.0 ;
      RECT  30300.0 423000.0 29100.0 421800.0 ;
      RECT  30900.0 419550.0 32100.0 418350.0 ;
      RECT  33300.0 428250.0 34500.0 427050.0 ;
      RECT  34500.0 423000.0 33300.0 421800.0 ;
      RECT  29100.0 423000.0 30300.0 421800.0 ;
      RECT  32100.0 425700.0 33300.0 424500.0 ;
      RECT  33300.0 423000.0 34500.0 421800.0 ;
      RECT  26700.0 416850.0 41100.0 415950.0 ;
      RECT  26700.0 430650.0 41100.0 429750.0 ;
      RECT  47700.0 221250.0 48900.0 223200.0 ;
      RECT  47700.0 209400.0 48900.0 211350.0 ;
      RECT  42900.0 210750.0 44100.0 208950.0 ;
      RECT  42900.0 220050.0 44100.0 223650.0 ;
      RECT  45600.0 210750.0 46500.0 220050.0 ;
      RECT  42900.0 220050.0 44100.0 221250.0 ;
      RECT  45300.0 220050.0 46500.0 221250.0 ;
      RECT  45300.0 220050.0 46500.0 221250.0 ;
      RECT  42900.0 220050.0 44100.0 221250.0 ;
      RECT  42900.0 210750.0 44100.0 211950.0 ;
      RECT  45300.0 210750.0 46500.0 211950.0 ;
      RECT  45300.0 210750.0 46500.0 211950.0 ;
      RECT  42900.0 210750.0 44100.0 211950.0 ;
      RECT  47700.0 220650.0 48900.0 221850.0 ;
      RECT  47700.0 210750.0 48900.0 211950.0 ;
      RECT  43500.0 215400.0 44700.0 216600.0 ;
      RECT  43500.0 215400.0 44700.0 216600.0 ;
      RECT  46050.0 215550.0 46950.0 216450.0 ;
      RECT  41100.0 222750.0 50700.0 223650.0 ;
      RECT  41100.0 208950.0 50700.0 209850.0 ;
      RECT  47700.0 225150.0 48900.0 223200.0 ;
      RECT  47700.0 237000.0 48900.0 235050.0 ;
      RECT  42900.0 235650.0 44100.0 237450.0 ;
      RECT  42900.0 226350.0 44100.0 222750.0 ;
      RECT  45600.0 235650.0 46500.0 226350.0 ;
      RECT  42900.0 226350.0 44100.0 225150.0 ;
      RECT  45300.0 226350.0 46500.0 225150.0 ;
      RECT  45300.0 226350.0 46500.0 225150.0 ;
      RECT  42900.0 226350.0 44100.0 225150.0 ;
      RECT  42900.0 235650.0 44100.0 234450.0 ;
      RECT  45300.0 235650.0 46500.0 234450.0 ;
      RECT  45300.0 235650.0 46500.0 234450.0 ;
      RECT  42900.0 235650.0 44100.0 234450.0 ;
      RECT  47700.0 225750.0 48900.0 224550.0 ;
      RECT  47700.0 235650.0 48900.0 234450.0 ;
      RECT  43500.0 231000.0 44700.0 229800.0 ;
      RECT  43500.0 231000.0 44700.0 229800.0 ;
      RECT  46050.0 230850.0 46950.0 229950.0 ;
      RECT  41100.0 223650.0 50700.0 222750.0 ;
      RECT  41100.0 237450.0 50700.0 236550.0 ;
      RECT  47700.0 248850.0 48900.0 250800.0 ;
      RECT  47700.0 237000.0 48900.0 238950.0 ;
      RECT  42900.0 238350.0 44100.0 236550.0 ;
      RECT  42900.0 247650.0 44100.0 251250.0 ;
      RECT  45600.0 238350.0 46500.0 247650.0 ;
      RECT  42900.0 247650.0 44100.0 248850.0 ;
      RECT  45300.0 247650.0 46500.0 248850.0 ;
      RECT  45300.0 247650.0 46500.0 248850.0 ;
      RECT  42900.0 247650.0 44100.0 248850.0 ;
      RECT  42900.0 238350.0 44100.0 239550.0 ;
      RECT  45300.0 238350.0 46500.0 239550.0 ;
      RECT  45300.0 238350.0 46500.0 239550.0 ;
      RECT  42900.0 238350.0 44100.0 239550.0 ;
      RECT  47700.0 248250.0 48900.0 249450.0 ;
      RECT  47700.0 238350.0 48900.0 239550.0 ;
      RECT  43500.0 243000.0 44700.0 244200.0 ;
      RECT  43500.0 243000.0 44700.0 244200.0 ;
      RECT  46050.0 243150.0 46950.0 244050.0 ;
      RECT  41100.0 250350.0 50700.0 251250.0 ;
      RECT  41100.0 236550.0 50700.0 237450.0 ;
      RECT  47700.0 252750.0 48900.0 250800.0 ;
      RECT  47700.0 264600.0 48900.0 262650.0 ;
      RECT  42900.0 263250.0 44100.0 265050.0 ;
      RECT  42900.0 253950.0 44100.0 250350.0 ;
      RECT  45600.0 263250.0 46500.0 253950.0 ;
      RECT  42900.0 253950.0 44100.0 252750.0 ;
      RECT  45300.0 253950.0 46500.0 252750.0 ;
      RECT  45300.0 253950.0 46500.0 252750.0 ;
      RECT  42900.0 253950.0 44100.0 252750.0 ;
      RECT  42900.0 263250.0 44100.0 262050.0 ;
      RECT  45300.0 263250.0 46500.0 262050.0 ;
      RECT  45300.0 263250.0 46500.0 262050.0 ;
      RECT  42900.0 263250.0 44100.0 262050.0 ;
      RECT  47700.0 253350.0 48900.0 252150.0 ;
      RECT  47700.0 263250.0 48900.0 262050.0 ;
      RECT  43500.0 258600.0 44700.0 257400.0 ;
      RECT  43500.0 258600.0 44700.0 257400.0 ;
      RECT  46050.0 258450.0 46950.0 257550.0 ;
      RECT  41100.0 251250.0 50700.0 250350.0 ;
      RECT  41100.0 265050.0 50700.0 264150.0 ;
      RECT  47700.0 276450.0 48900.0 278400.0 ;
      RECT  47700.0 264600.0 48900.0 266550.0 ;
      RECT  42900.0 265950.0 44100.0 264150.0 ;
      RECT  42900.0 275250.0 44100.0 278850.0 ;
      RECT  45600.0 265950.0 46500.0 275250.0 ;
      RECT  42900.0 275250.0 44100.0 276450.0 ;
      RECT  45300.0 275250.0 46500.0 276450.0 ;
      RECT  45300.0 275250.0 46500.0 276450.0 ;
      RECT  42900.0 275250.0 44100.0 276450.0 ;
      RECT  42900.0 265950.0 44100.0 267150.0 ;
      RECT  45300.0 265950.0 46500.0 267150.0 ;
      RECT  45300.0 265950.0 46500.0 267150.0 ;
      RECT  42900.0 265950.0 44100.0 267150.0 ;
      RECT  47700.0 275850.0 48900.0 277050.0 ;
      RECT  47700.0 265950.0 48900.0 267150.0 ;
      RECT  43500.0 270600.0 44700.0 271800.0 ;
      RECT  43500.0 270600.0 44700.0 271800.0 ;
      RECT  46050.0 270750.0 46950.0 271650.0 ;
      RECT  41100.0 277950.0 50700.0 278850.0 ;
      RECT  41100.0 264150.0 50700.0 265050.0 ;
      RECT  47700.0 280350.0 48900.0 278400.0 ;
      RECT  47700.0 292200.0 48900.0 290250.0 ;
      RECT  42900.0 290850.0 44100.0 292650.0 ;
      RECT  42900.0 281550.0 44100.0 277950.0 ;
      RECT  45600.0 290850.0 46500.0 281550.0 ;
      RECT  42900.0 281550.0 44100.0 280350.0 ;
      RECT  45300.0 281550.0 46500.0 280350.0 ;
      RECT  45300.0 281550.0 46500.0 280350.0 ;
      RECT  42900.0 281550.0 44100.0 280350.0 ;
      RECT  42900.0 290850.0 44100.0 289650.0 ;
      RECT  45300.0 290850.0 46500.0 289650.0 ;
      RECT  45300.0 290850.0 46500.0 289650.0 ;
      RECT  42900.0 290850.0 44100.0 289650.0 ;
      RECT  47700.0 280950.0 48900.0 279750.0 ;
      RECT  47700.0 290850.0 48900.0 289650.0 ;
      RECT  43500.0 286200.0 44700.0 285000.0 ;
      RECT  43500.0 286200.0 44700.0 285000.0 ;
      RECT  46050.0 286050.0 46950.0 285150.0 ;
      RECT  41100.0 278850.0 50700.0 277950.0 ;
      RECT  41100.0 292650.0 50700.0 291750.0 ;
      RECT  47700.0 304050.0 48900.0 306000.0 ;
      RECT  47700.0 292200.0 48900.0 294150.0 ;
      RECT  42900.0 293550.0 44100.0 291750.0 ;
      RECT  42900.0 302850.0 44100.0 306450.0 ;
      RECT  45600.0 293550.0 46500.0 302850.0 ;
      RECT  42900.0 302850.0 44100.0 304050.0 ;
      RECT  45300.0 302850.0 46500.0 304050.0 ;
      RECT  45300.0 302850.0 46500.0 304050.0 ;
      RECT  42900.0 302850.0 44100.0 304050.0 ;
      RECT  42900.0 293550.0 44100.0 294750.0 ;
      RECT  45300.0 293550.0 46500.0 294750.0 ;
      RECT  45300.0 293550.0 46500.0 294750.0 ;
      RECT  42900.0 293550.0 44100.0 294750.0 ;
      RECT  47700.0 303450.0 48900.0 304650.0 ;
      RECT  47700.0 293550.0 48900.0 294750.0 ;
      RECT  43500.0 298200.0 44700.0 299400.0 ;
      RECT  43500.0 298200.0 44700.0 299400.0 ;
      RECT  46050.0 298350.0 46950.0 299250.0 ;
      RECT  41100.0 305550.0 50700.0 306450.0 ;
      RECT  41100.0 291750.0 50700.0 292650.0 ;
      RECT  47700.0 307950.0 48900.0 306000.0 ;
      RECT  47700.0 319800.0 48900.0 317850.0 ;
      RECT  42900.0 318450.0 44100.0 320250.0 ;
      RECT  42900.0 309150.0 44100.0 305550.0 ;
      RECT  45600.0 318450.0 46500.0 309150.0 ;
      RECT  42900.0 309150.0 44100.0 307950.0 ;
      RECT  45300.0 309150.0 46500.0 307950.0 ;
      RECT  45300.0 309150.0 46500.0 307950.0 ;
      RECT  42900.0 309150.0 44100.0 307950.0 ;
      RECT  42900.0 318450.0 44100.0 317250.0 ;
      RECT  45300.0 318450.0 46500.0 317250.0 ;
      RECT  45300.0 318450.0 46500.0 317250.0 ;
      RECT  42900.0 318450.0 44100.0 317250.0 ;
      RECT  47700.0 308550.0 48900.0 307350.0 ;
      RECT  47700.0 318450.0 48900.0 317250.0 ;
      RECT  43500.0 313800.0 44700.0 312600.0 ;
      RECT  43500.0 313800.0 44700.0 312600.0 ;
      RECT  46050.0 313650.0 46950.0 312750.0 ;
      RECT  41100.0 306450.0 50700.0 305550.0 ;
      RECT  41100.0 320250.0 50700.0 319350.0 ;
      RECT  47700.0 331650.0 48900.0 333600.0 ;
      RECT  47700.0 319800.0 48900.0 321750.0 ;
      RECT  42900.0 321150.0 44100.0 319350.0 ;
      RECT  42900.0 330450.0 44100.0 334050.0 ;
      RECT  45600.0 321150.0 46500.0 330450.0 ;
      RECT  42900.0 330450.0 44100.0 331650.0 ;
      RECT  45300.0 330450.0 46500.0 331650.0 ;
      RECT  45300.0 330450.0 46500.0 331650.0 ;
      RECT  42900.0 330450.0 44100.0 331650.0 ;
      RECT  42900.0 321150.0 44100.0 322350.0 ;
      RECT  45300.0 321150.0 46500.0 322350.0 ;
      RECT  45300.0 321150.0 46500.0 322350.0 ;
      RECT  42900.0 321150.0 44100.0 322350.0 ;
      RECT  47700.0 331050.0 48900.0 332250.0 ;
      RECT  47700.0 321150.0 48900.0 322350.0 ;
      RECT  43500.0 325800.0 44700.0 327000.0 ;
      RECT  43500.0 325800.0 44700.0 327000.0 ;
      RECT  46050.0 325950.0 46950.0 326850.0 ;
      RECT  41100.0 333150.0 50700.0 334050.0 ;
      RECT  41100.0 319350.0 50700.0 320250.0 ;
      RECT  47700.0 335550.0 48900.0 333600.0 ;
      RECT  47700.0 347400.0 48900.0 345450.0 ;
      RECT  42900.0 346050.0 44100.0 347850.0 ;
      RECT  42900.0 336750.0 44100.0 333150.0 ;
      RECT  45600.0 346050.0 46500.0 336750.0 ;
      RECT  42900.0 336750.0 44100.0 335550.0 ;
      RECT  45300.0 336750.0 46500.0 335550.0 ;
      RECT  45300.0 336750.0 46500.0 335550.0 ;
      RECT  42900.0 336750.0 44100.0 335550.0 ;
      RECT  42900.0 346050.0 44100.0 344850.0 ;
      RECT  45300.0 346050.0 46500.0 344850.0 ;
      RECT  45300.0 346050.0 46500.0 344850.0 ;
      RECT  42900.0 346050.0 44100.0 344850.0 ;
      RECT  47700.0 336150.0 48900.0 334950.0 ;
      RECT  47700.0 346050.0 48900.0 344850.0 ;
      RECT  43500.0 341400.0 44700.0 340200.0 ;
      RECT  43500.0 341400.0 44700.0 340200.0 ;
      RECT  46050.0 341250.0 46950.0 340350.0 ;
      RECT  41100.0 334050.0 50700.0 333150.0 ;
      RECT  41100.0 347850.0 50700.0 346950.0 ;
      RECT  47700.0 359250.0 48900.0 361200.0 ;
      RECT  47700.0 347400.0 48900.0 349350.0 ;
      RECT  42900.0 348750.0 44100.0 346950.0 ;
      RECT  42900.0 358050.0 44100.0 361650.0 ;
      RECT  45600.0 348750.0 46500.0 358050.0 ;
      RECT  42900.0 358050.0 44100.0 359250.0 ;
      RECT  45300.0 358050.0 46500.0 359250.0 ;
      RECT  45300.0 358050.0 46500.0 359250.0 ;
      RECT  42900.0 358050.0 44100.0 359250.0 ;
      RECT  42900.0 348750.0 44100.0 349950.0 ;
      RECT  45300.0 348750.0 46500.0 349950.0 ;
      RECT  45300.0 348750.0 46500.0 349950.0 ;
      RECT  42900.0 348750.0 44100.0 349950.0 ;
      RECT  47700.0 358650.0 48900.0 359850.0 ;
      RECT  47700.0 348750.0 48900.0 349950.0 ;
      RECT  43500.0 353400.0 44700.0 354600.0 ;
      RECT  43500.0 353400.0 44700.0 354600.0 ;
      RECT  46050.0 353550.0 46950.0 354450.0 ;
      RECT  41100.0 360750.0 50700.0 361650.0 ;
      RECT  41100.0 346950.0 50700.0 347850.0 ;
      RECT  47700.0 363150.0 48900.0 361200.0 ;
      RECT  47700.0 375000.0 48900.0 373050.0 ;
      RECT  42900.0 373650.0 44100.0 375450.0 ;
      RECT  42900.0 364350.0 44100.0 360750.0 ;
      RECT  45600.0 373650.0 46500.0 364350.0 ;
      RECT  42900.0 364350.0 44100.0 363150.0 ;
      RECT  45300.0 364350.0 46500.0 363150.0 ;
      RECT  45300.0 364350.0 46500.0 363150.0 ;
      RECT  42900.0 364350.0 44100.0 363150.0 ;
      RECT  42900.0 373650.0 44100.0 372450.0 ;
      RECT  45300.0 373650.0 46500.0 372450.0 ;
      RECT  45300.0 373650.0 46500.0 372450.0 ;
      RECT  42900.0 373650.0 44100.0 372450.0 ;
      RECT  47700.0 363750.0 48900.0 362550.0 ;
      RECT  47700.0 373650.0 48900.0 372450.0 ;
      RECT  43500.0 369000.0 44700.0 367800.0 ;
      RECT  43500.0 369000.0 44700.0 367800.0 ;
      RECT  46050.0 368850.0 46950.0 367950.0 ;
      RECT  41100.0 361650.0 50700.0 360750.0 ;
      RECT  41100.0 375450.0 50700.0 374550.0 ;
      RECT  47700.0 386850.0 48900.0 388800.0 ;
      RECT  47700.0 375000.0 48900.0 376950.0 ;
      RECT  42900.0 376350.0 44100.0 374550.0 ;
      RECT  42900.0 385650.0 44100.0 389250.0 ;
      RECT  45600.0 376350.0 46500.0 385650.0 ;
      RECT  42900.0 385650.0 44100.0 386850.0 ;
      RECT  45300.0 385650.0 46500.0 386850.0 ;
      RECT  45300.0 385650.0 46500.0 386850.0 ;
      RECT  42900.0 385650.0 44100.0 386850.0 ;
      RECT  42900.0 376350.0 44100.0 377550.0 ;
      RECT  45300.0 376350.0 46500.0 377550.0 ;
      RECT  45300.0 376350.0 46500.0 377550.0 ;
      RECT  42900.0 376350.0 44100.0 377550.0 ;
      RECT  47700.0 386250.0 48900.0 387450.0 ;
      RECT  47700.0 376350.0 48900.0 377550.0 ;
      RECT  43500.0 381000.0 44700.0 382200.0 ;
      RECT  43500.0 381000.0 44700.0 382200.0 ;
      RECT  46050.0 381150.0 46950.0 382050.0 ;
      RECT  41100.0 388350.0 50700.0 389250.0 ;
      RECT  41100.0 374550.0 50700.0 375450.0 ;
      RECT  47700.0 390750.0 48900.0 388800.0 ;
      RECT  47700.0 402600.0 48900.0 400650.0 ;
      RECT  42900.0 401250.0 44100.0 403050.0 ;
      RECT  42900.0 391950.0 44100.0 388350.0 ;
      RECT  45600.0 401250.0 46500.0 391950.0 ;
      RECT  42900.0 391950.0 44100.0 390750.0 ;
      RECT  45300.0 391950.0 46500.0 390750.0 ;
      RECT  45300.0 391950.0 46500.0 390750.0 ;
      RECT  42900.0 391950.0 44100.0 390750.0 ;
      RECT  42900.0 401250.0 44100.0 400050.0 ;
      RECT  45300.0 401250.0 46500.0 400050.0 ;
      RECT  45300.0 401250.0 46500.0 400050.0 ;
      RECT  42900.0 401250.0 44100.0 400050.0 ;
      RECT  47700.0 391350.0 48900.0 390150.0 ;
      RECT  47700.0 401250.0 48900.0 400050.0 ;
      RECT  43500.0 396600.0 44700.0 395400.0 ;
      RECT  43500.0 396600.0 44700.0 395400.0 ;
      RECT  46050.0 396450.0 46950.0 395550.0 ;
      RECT  41100.0 389250.0 50700.0 388350.0 ;
      RECT  41100.0 403050.0 50700.0 402150.0 ;
      RECT  47700.0 414450.0 48900.0 416400.0 ;
      RECT  47700.0 402600.0 48900.0 404550.0 ;
      RECT  42900.0 403950.0 44100.0 402150.0 ;
      RECT  42900.0 413250.0 44100.0 416850.0 ;
      RECT  45600.0 403950.0 46500.0 413250.0 ;
      RECT  42900.0 413250.0 44100.0 414450.0 ;
      RECT  45300.0 413250.0 46500.0 414450.0 ;
      RECT  45300.0 413250.0 46500.0 414450.0 ;
      RECT  42900.0 413250.0 44100.0 414450.0 ;
      RECT  42900.0 403950.0 44100.0 405150.0 ;
      RECT  45300.0 403950.0 46500.0 405150.0 ;
      RECT  45300.0 403950.0 46500.0 405150.0 ;
      RECT  42900.0 403950.0 44100.0 405150.0 ;
      RECT  47700.0 413850.0 48900.0 415050.0 ;
      RECT  47700.0 403950.0 48900.0 405150.0 ;
      RECT  43500.0 408600.0 44700.0 409800.0 ;
      RECT  43500.0 408600.0 44700.0 409800.0 ;
      RECT  46050.0 408750.0 46950.0 409650.0 ;
      RECT  41100.0 415950.0 50700.0 416850.0 ;
      RECT  41100.0 402150.0 50700.0 403050.0 ;
      RECT  47700.0 418350.0 48900.0 416400.0 ;
      RECT  47700.0 430200.0 48900.0 428250.0 ;
      RECT  42900.0 428850.0 44100.0 430650.0 ;
      RECT  42900.0 419550.0 44100.0 415950.0 ;
      RECT  45600.0 428850.0 46500.0 419550.0 ;
      RECT  42900.0 419550.0 44100.0 418350.0 ;
      RECT  45300.0 419550.0 46500.0 418350.0 ;
      RECT  45300.0 419550.0 46500.0 418350.0 ;
      RECT  42900.0 419550.0 44100.0 418350.0 ;
      RECT  42900.0 428850.0 44100.0 427650.0 ;
      RECT  45300.0 428850.0 46500.0 427650.0 ;
      RECT  45300.0 428850.0 46500.0 427650.0 ;
      RECT  42900.0 428850.0 44100.0 427650.0 ;
      RECT  47700.0 418950.0 48900.0 417750.0 ;
      RECT  47700.0 428850.0 48900.0 427650.0 ;
      RECT  43500.0 424200.0 44700.0 423000.0 ;
      RECT  43500.0 424200.0 44700.0 423000.0 ;
      RECT  46050.0 424050.0 46950.0 423150.0 ;
      RECT  41100.0 416850.0 50700.0 415950.0 ;
      RECT  41100.0 430650.0 50700.0 429750.0 ;
      RECT  10950.0 105000.0 9750.0 106200.0 ;
      RECT  13050.0 119400.0 11850.0 120600.0 ;
      RECT  15150.0 132600.0 13950.0 133800.0 ;
      RECT  17250.0 147000.0 16050.0 148200.0 ;
      RECT  19350.0 160200.0 18150.0 161400.0 ;
      RECT  21450.0 174600.0 20250.0 175800.0 ;
      RECT  23550.0 187800.0 22350.0 189000.0 ;
      RECT  25650.0 202200.0 24450.0 203400.0 ;
      RECT  10950.0 216600.0 9750.0 217800.0 ;
      RECT  19350.0 213900.0 18150.0 215100.0 ;
      RECT  10950.0 228600.0 9750.0 229800.0 ;
      RECT  21450.0 231300.0 20250.0 232500.0 ;
      RECT  10950.0 244200.0 9750.0 245400.0 ;
      RECT  23550.0 241500.0 22350.0 242700.0 ;
      RECT  10950.0 256200.0 9750.0 257400.0 ;
      RECT  25650.0 258900.0 24450.0 260100.0 ;
      RECT  13050.0 271800.0 11850.0 273000.0 ;
      RECT  19350.0 269100.0 18150.0 270300.0 ;
      RECT  13050.0 283800.0 11850.0 285000.0 ;
      RECT  21450.0 286500.0 20250.0 287700.0 ;
      RECT  13050.0 299400.0 11850.0 300600.0 ;
      RECT  23550.0 296700.0 22350.0 297900.0 ;
      RECT  13050.0 311400.0 11850.0 312600.0 ;
      RECT  25650.0 314100.0 24450.0 315300.0 ;
      RECT  15150.0 327000.0 13950.0 328200.0 ;
      RECT  19350.0 324300.0 18150.0 325500.0 ;
      RECT  15150.0 339000.0 13950.0 340200.0 ;
      RECT  21450.0 341700.0 20250.0 342900.0 ;
      RECT  15150.0 354600.0 13950.0 355800.0 ;
      RECT  23550.0 351900.0 22350.0 353100.0 ;
      RECT  15150.0 366600.0 13950.0 367800.0 ;
      RECT  25650.0 369300.0 24450.0 370500.0 ;
      RECT  17250.0 382200.0 16050.0 383400.0 ;
      RECT  19350.0 379500.0 18150.0 380700.0 ;
      RECT  17250.0 394200.0 16050.0 395400.0 ;
      RECT  21450.0 396900.0 20250.0 398100.0 ;
      RECT  17250.0 409800.0 16050.0 411000.0 ;
      RECT  23550.0 407100.0 22350.0 408300.0 ;
      RECT  17250.0 421800.0 16050.0 423000.0 ;
      RECT  25650.0 424500.0 24450.0 425700.0 ;
      RECT  46050.0 215550.0 46950.0 216450.0 ;
      RECT  46050.0 229950.0 46950.0 230850.0 ;
      RECT  46050.0 243150.0 46950.0 244050.0 ;
      RECT  46050.0 257550.0 46950.0 258450.0 ;
      RECT  46050.0 270750.0 46950.0 271650.0 ;
      RECT  46050.0 285150.0 46950.0 286050.0 ;
      RECT  46050.0 298350.0 46950.0 299250.0 ;
      RECT  46050.0 312750.0 46950.0 313650.0 ;
      RECT  46050.0 325950.0 46950.0 326850.0 ;
      RECT  46050.0 340350.0 46950.0 341250.0 ;
      RECT  46050.0 353550.0 46950.0 354450.0 ;
      RECT  46050.0 367950.0 46950.0 368850.0 ;
      RECT  46050.0 381150.0 46950.0 382050.0 ;
      RECT  46050.0 395550.0 46950.0 396450.0 ;
      RECT  46050.0 408750.0 46950.0 409650.0 ;
      RECT  46050.0 423150.0 46950.0 424050.0 ;
      RECT  9900.0 112350.0 81300.0 113250.0 ;
      RECT  9900.0 139950.0 81300.0 140850.0 ;
      RECT  9900.0 167550.0 81300.0 168450.0 ;
      RECT  9900.0 195150.0 81300.0 196050.0 ;
      RECT  9900.0 222750.0 81300.0 223650.0 ;
      RECT  9900.0 250350.0 81300.0 251250.0 ;
      RECT  9900.0 277950.0 81300.0 278850.0 ;
      RECT  9900.0 305550.0 81300.0 306450.0 ;
      RECT  9900.0 333150.0 81300.0 334050.0 ;
      RECT  9900.0 360750.0 81300.0 361650.0 ;
      RECT  9900.0 388350.0 81300.0 389250.0 ;
      RECT  9900.0 415950.0 81300.0 416850.0 ;
      RECT  9900.0 98550.0 81300.0 99450.0 ;
      RECT  9900.0 126150.0 81300.0 127050.0 ;
      RECT  9900.0 153750.0 81300.0 154650.0 ;
      RECT  9900.0 181350.0 81300.0 182250.0 ;
      RECT  9900.0 208950.0 81300.0 209850.0 ;
      RECT  9900.0 236550.0 81300.0 237450.0 ;
      RECT  9900.0 264150.0 81300.0 265050.0 ;
      RECT  9900.0 291750.0 81300.0 292650.0 ;
      RECT  9900.0 319350.0 81300.0 320250.0 ;
      RECT  9900.0 346950.0 81300.0 347850.0 ;
      RECT  9900.0 374550.0 81300.0 375450.0 ;
      RECT  9900.0 402150.0 81300.0 403050.0 ;
      RECT  9900.0 429750.0 81300.0 430650.0 ;
      RECT  53850.0 215550.0 59400.0 216450.0 ;
      RECT  61950.0 216750.0 62850.0 217650.0 ;
      RECT  61950.0 215550.0 62850.0 216450.0 ;
      RECT  61950.0 216450.0 62850.0 217200.0 ;
      RECT  62400.0 216750.0 69000.0 217650.0 ;
      RECT  69000.0 216750.0 70200.0 217650.0 ;
      RECT  78450.0 216750.0 79350.0 217650.0 ;
      RECT  78450.0 215550.0 79350.0 216450.0 ;
      RECT  74400.0 216750.0 78900.0 217650.0 ;
      RECT  78450.0 216000.0 79350.0 217200.0 ;
      RECT  78900.0 215550.0 83400.0 216450.0 ;
      RECT  53850.0 229950.0 59400.0 230850.0 ;
      RECT  61950.0 228750.0 62850.0 229650.0 ;
      RECT  61950.0 229950.0 62850.0 230850.0 ;
      RECT  61950.0 229200.0 62850.0 230850.0 ;
      RECT  62400.0 228750.0 69000.0 229650.0 ;
      RECT  69000.0 228750.0 70200.0 229650.0 ;
      RECT  78450.0 228750.0 79350.0 229650.0 ;
      RECT  78450.0 229950.0 79350.0 230850.0 ;
      RECT  74400.0 228750.0 78900.0 229650.0 ;
      RECT  78450.0 229200.0 79350.0 230400.0 ;
      RECT  78900.0 229950.0 83400.0 230850.0 ;
      RECT  53850.0 243150.0 59400.0 244050.0 ;
      RECT  61950.0 244350.0 62850.0 245250.0 ;
      RECT  61950.0 243150.0 62850.0 244050.0 ;
      RECT  61950.0 244050.0 62850.0 244800.0 ;
      RECT  62400.0 244350.0 69000.0 245250.0 ;
      RECT  69000.0 244350.0 70200.0 245250.0 ;
      RECT  78450.0 244350.0 79350.0 245250.0 ;
      RECT  78450.0 243150.0 79350.0 244050.0 ;
      RECT  74400.0 244350.0 78900.0 245250.0 ;
      RECT  78450.0 243600.0 79350.0 244800.0 ;
      RECT  78900.0 243150.0 83400.0 244050.0 ;
      RECT  53850.0 257550.0 59400.0 258450.0 ;
      RECT  61950.0 256350.0 62850.0 257250.0 ;
      RECT  61950.0 257550.0 62850.0 258450.0 ;
      RECT  61950.0 256800.0 62850.0 258450.0 ;
      RECT  62400.0 256350.0 69000.0 257250.0 ;
      RECT  69000.0 256350.0 70200.0 257250.0 ;
      RECT  78450.0 256350.0 79350.0 257250.0 ;
      RECT  78450.0 257550.0 79350.0 258450.0 ;
      RECT  74400.0 256350.0 78900.0 257250.0 ;
      RECT  78450.0 256800.0 79350.0 258000.0 ;
      RECT  78900.0 257550.0 83400.0 258450.0 ;
      RECT  53850.0 270750.0 59400.0 271650.0 ;
      RECT  61950.0 271950.0 62850.0 272850.0 ;
      RECT  61950.0 270750.0 62850.0 271650.0 ;
      RECT  61950.0 271650.0 62850.0 272400.0 ;
      RECT  62400.0 271950.0 69000.0 272850.0 ;
      RECT  69000.0 271950.0 70200.0 272850.0 ;
      RECT  78450.0 271950.0 79350.0 272850.0 ;
      RECT  78450.0 270750.0 79350.0 271650.0 ;
      RECT  74400.0 271950.0 78900.0 272850.0 ;
      RECT  78450.0 271200.0 79350.0 272400.0 ;
      RECT  78900.0 270750.0 83400.0 271650.0 ;
      RECT  53850.0 285150.0 59400.0 286050.0 ;
      RECT  61950.0 283950.0 62850.0 284850.0 ;
      RECT  61950.0 285150.0 62850.0 286050.0 ;
      RECT  61950.0 284400.0 62850.0 286050.0 ;
      RECT  62400.0 283950.0 69000.0 284850.0 ;
      RECT  69000.0 283950.0 70200.0 284850.0 ;
      RECT  78450.0 283950.0 79350.0 284850.0 ;
      RECT  78450.0 285150.0 79350.0 286050.0 ;
      RECT  74400.0 283950.0 78900.0 284850.0 ;
      RECT  78450.0 284400.0 79350.0 285600.0 ;
      RECT  78900.0 285150.0 83400.0 286050.0 ;
      RECT  53850.0 298350.0 59400.0 299250.0 ;
      RECT  61950.0 299550.0 62850.0 300450.0 ;
      RECT  61950.0 298350.0 62850.0 299250.0 ;
      RECT  61950.0 299250.0 62850.0 300000.0 ;
      RECT  62400.0 299550.0 69000.0 300450.0 ;
      RECT  69000.0 299550.0 70200.0 300450.0 ;
      RECT  78450.0 299550.0 79350.0 300450.0 ;
      RECT  78450.0 298350.0 79350.0 299250.0 ;
      RECT  74400.0 299550.0 78900.0 300450.0 ;
      RECT  78450.0 298800.0 79350.0 300000.0 ;
      RECT  78900.0 298350.0 83400.0 299250.0 ;
      RECT  53850.0 312750.0 59400.0 313650.0 ;
      RECT  61950.0 311550.0 62850.0 312450.0 ;
      RECT  61950.0 312750.0 62850.0 313650.0 ;
      RECT  61950.0 312000.0 62850.0 313650.0 ;
      RECT  62400.0 311550.0 69000.0 312450.0 ;
      RECT  69000.0 311550.0 70200.0 312450.0 ;
      RECT  78450.0 311550.0 79350.0 312450.0 ;
      RECT  78450.0 312750.0 79350.0 313650.0 ;
      RECT  74400.0 311550.0 78900.0 312450.0 ;
      RECT  78450.0 312000.0 79350.0 313200.0 ;
      RECT  78900.0 312750.0 83400.0 313650.0 ;
      RECT  53850.0 325950.0 59400.0 326850.0 ;
      RECT  61950.0 327150.0 62850.0 328050.0 ;
      RECT  61950.0 325950.0 62850.0 326850.0 ;
      RECT  61950.0 326850.0 62850.0 327600.0 ;
      RECT  62400.0 327150.0 69000.0 328050.0 ;
      RECT  69000.0 327150.0 70200.0 328050.0 ;
      RECT  78450.0 327150.0 79350.0 328050.0 ;
      RECT  78450.0 325950.0 79350.0 326850.0 ;
      RECT  74400.0 327150.0 78900.0 328050.0 ;
      RECT  78450.0 326400.0 79350.0 327600.0 ;
      RECT  78900.0 325950.0 83400.0 326850.0 ;
      RECT  53850.0 340350.0 59400.0 341250.0 ;
      RECT  61950.0 339150.0 62850.0 340050.0 ;
      RECT  61950.0 340350.0 62850.0 341250.0 ;
      RECT  61950.0 339600.0 62850.0 341250.0 ;
      RECT  62400.0 339150.0 69000.0 340050.0 ;
      RECT  69000.0 339150.0 70200.0 340050.0 ;
      RECT  78450.0 339150.0 79350.0 340050.0 ;
      RECT  78450.0 340350.0 79350.0 341250.0 ;
      RECT  74400.0 339150.0 78900.0 340050.0 ;
      RECT  78450.0 339600.0 79350.0 340800.0 ;
      RECT  78900.0 340350.0 83400.0 341250.0 ;
      RECT  53850.0 353550.0 59400.0 354450.0 ;
      RECT  61950.0 354750.0 62850.0 355650.0 ;
      RECT  61950.0 353550.0 62850.0 354450.0 ;
      RECT  61950.0 354450.0 62850.0 355200.0 ;
      RECT  62400.0 354750.0 69000.0 355650.0 ;
      RECT  69000.0 354750.0 70200.0 355650.0 ;
      RECT  78450.0 354750.0 79350.0 355650.0 ;
      RECT  78450.0 353550.0 79350.0 354450.0 ;
      RECT  74400.0 354750.0 78900.0 355650.0 ;
      RECT  78450.0 354000.0 79350.0 355200.0 ;
      RECT  78900.0 353550.0 83400.0 354450.0 ;
      RECT  53850.0 367950.0 59400.0 368850.0 ;
      RECT  61950.0 366750.0 62850.0 367650.0 ;
      RECT  61950.0 367950.0 62850.0 368850.0 ;
      RECT  61950.0 367200.0 62850.0 368850.0 ;
      RECT  62400.0 366750.0 69000.0 367650.0 ;
      RECT  69000.0 366750.0 70200.0 367650.0 ;
      RECT  78450.0 366750.0 79350.0 367650.0 ;
      RECT  78450.0 367950.0 79350.0 368850.0 ;
      RECT  74400.0 366750.0 78900.0 367650.0 ;
      RECT  78450.0 367200.0 79350.0 368400.0 ;
      RECT  78900.0 367950.0 83400.0 368850.0 ;
      RECT  53850.0 381150.0 59400.0 382050.0 ;
      RECT  61950.0 382350.0 62850.0 383250.0 ;
      RECT  61950.0 381150.0 62850.0 382050.0 ;
      RECT  61950.0 382050.0 62850.0 382800.0 ;
      RECT  62400.0 382350.0 69000.0 383250.0 ;
      RECT  69000.0 382350.0 70200.0 383250.0 ;
      RECT  78450.0 382350.0 79350.0 383250.0 ;
      RECT  78450.0 381150.0 79350.0 382050.0 ;
      RECT  74400.0 382350.0 78900.0 383250.0 ;
      RECT  78450.0 381600.0 79350.0 382800.0 ;
      RECT  78900.0 381150.0 83400.0 382050.0 ;
      RECT  53850.0 395550.0 59400.0 396450.0 ;
      RECT  61950.0 394350.0 62850.0 395250.0 ;
      RECT  61950.0 395550.0 62850.0 396450.0 ;
      RECT  61950.0 394800.0 62850.0 396450.0 ;
      RECT  62400.0 394350.0 69000.0 395250.0 ;
      RECT  69000.0 394350.0 70200.0 395250.0 ;
      RECT  78450.0 394350.0 79350.0 395250.0 ;
      RECT  78450.0 395550.0 79350.0 396450.0 ;
      RECT  74400.0 394350.0 78900.0 395250.0 ;
      RECT  78450.0 394800.0 79350.0 396000.0 ;
      RECT  78900.0 395550.0 83400.0 396450.0 ;
      RECT  53850.0 408750.0 59400.0 409650.0 ;
      RECT  61950.0 409950.0 62850.0 410850.0 ;
      RECT  61950.0 408750.0 62850.0 409650.0 ;
      RECT  61950.0 409650.0 62850.0 410400.0 ;
      RECT  62400.0 409950.0 69000.0 410850.0 ;
      RECT  69000.0 409950.0 70200.0 410850.0 ;
      RECT  78450.0 409950.0 79350.0 410850.0 ;
      RECT  78450.0 408750.0 79350.0 409650.0 ;
      RECT  74400.0 409950.0 78900.0 410850.0 ;
      RECT  78450.0 409200.0 79350.0 410400.0 ;
      RECT  78900.0 408750.0 83400.0 409650.0 ;
      RECT  53850.0 423150.0 59400.0 424050.0 ;
      RECT  61950.0 421950.0 62850.0 422850.0 ;
      RECT  61950.0 423150.0 62850.0 424050.0 ;
      RECT  61950.0 422400.0 62850.0 424050.0 ;
      RECT  62400.0 421950.0 69000.0 422850.0 ;
      RECT  69000.0 421950.0 70200.0 422850.0 ;
      RECT  78450.0 421950.0 79350.0 422850.0 ;
      RECT  78450.0 423150.0 79350.0 424050.0 ;
      RECT  74400.0 421950.0 78900.0 422850.0 ;
      RECT  78450.0 422400.0 79350.0 423600.0 ;
      RECT  78900.0 423150.0 83400.0 424050.0 ;
      RECT  63600.0 221250.0 64800.0 223200.0 ;
      RECT  63600.0 209400.0 64800.0 211350.0 ;
      RECT  58800.0 210750.0 60000.0 208950.0 ;
      RECT  58800.0 220050.0 60000.0 223650.0 ;
      RECT  61500.0 210750.0 62400.0 220050.0 ;
      RECT  58800.0 220050.0 60000.0 221250.0 ;
      RECT  61200.0 220050.0 62400.0 221250.0 ;
      RECT  61200.0 220050.0 62400.0 221250.0 ;
      RECT  58800.0 220050.0 60000.0 221250.0 ;
      RECT  58800.0 210750.0 60000.0 211950.0 ;
      RECT  61200.0 210750.0 62400.0 211950.0 ;
      RECT  61200.0 210750.0 62400.0 211950.0 ;
      RECT  58800.0 210750.0 60000.0 211950.0 ;
      RECT  63600.0 220650.0 64800.0 221850.0 ;
      RECT  63600.0 210750.0 64800.0 211950.0 ;
      RECT  59400.0 215400.0 60600.0 216600.0 ;
      RECT  59400.0 215400.0 60600.0 216600.0 ;
      RECT  61950.0 215550.0 62850.0 216450.0 ;
      RECT  57000.0 222750.0 66600.0 223650.0 ;
      RECT  57000.0 208950.0 66600.0 209850.0 ;
      RECT  68400.0 211350.0 69600.0 208950.0 ;
      RECT  68400.0 220050.0 69600.0 223650.0 ;
      RECT  73200.0 220050.0 74400.0 223650.0 ;
      RECT  75600.0 221250.0 76800.0 223200.0 ;
      RECT  75600.0 209400.0 76800.0 211350.0 ;
      RECT  68400.0 220050.0 69600.0 221250.0 ;
      RECT  70800.0 220050.0 72000.0 221250.0 ;
      RECT  70800.0 220050.0 72000.0 221250.0 ;
      RECT  68400.0 220050.0 69600.0 221250.0 ;
      RECT  70800.0 220050.0 72000.0 221250.0 ;
      RECT  73200.0 220050.0 74400.0 221250.0 ;
      RECT  73200.0 220050.0 74400.0 221250.0 ;
      RECT  70800.0 220050.0 72000.0 221250.0 ;
      RECT  68400.0 211350.0 69600.0 212550.0 ;
      RECT  70800.0 211350.0 72000.0 212550.0 ;
      RECT  70800.0 211350.0 72000.0 212550.0 ;
      RECT  68400.0 211350.0 69600.0 212550.0 ;
      RECT  70800.0 211350.0 72000.0 212550.0 ;
      RECT  73200.0 211350.0 74400.0 212550.0 ;
      RECT  73200.0 211350.0 74400.0 212550.0 ;
      RECT  70800.0 211350.0 72000.0 212550.0 ;
      RECT  75600.0 220650.0 76800.0 221850.0 ;
      RECT  75600.0 210750.0 76800.0 211950.0 ;
      RECT  73200.0 213900.0 72000.0 215100.0 ;
      RECT  70200.0 216600.0 69000.0 217800.0 ;
      RECT  70800.0 220050.0 72000.0 221250.0 ;
      RECT  73200.0 211350.0 74400.0 212550.0 ;
      RECT  74400.0 216600.0 73200.0 217800.0 ;
      RECT  69000.0 216600.0 70200.0 217800.0 ;
      RECT  72000.0 213900.0 73200.0 215100.0 ;
      RECT  73200.0 216600.0 74400.0 217800.0 ;
      RECT  66600.0 222750.0 81000.0 223650.0 ;
      RECT  66600.0 208950.0 81000.0 209850.0 ;
      RECT  87600.0 221250.0 88800.0 223200.0 ;
      RECT  87600.0 209400.0 88800.0 211350.0 ;
      RECT  82800.0 210750.0 84000.0 208950.0 ;
      RECT  82800.0 220050.0 84000.0 223650.0 ;
      RECT  85500.0 210750.0 86400.0 220050.0 ;
      RECT  82800.0 220050.0 84000.0 221250.0 ;
      RECT  85200.0 220050.0 86400.0 221250.0 ;
      RECT  85200.0 220050.0 86400.0 221250.0 ;
      RECT  82800.0 220050.0 84000.0 221250.0 ;
      RECT  82800.0 210750.0 84000.0 211950.0 ;
      RECT  85200.0 210750.0 86400.0 211950.0 ;
      RECT  85200.0 210750.0 86400.0 211950.0 ;
      RECT  82800.0 210750.0 84000.0 211950.0 ;
      RECT  87600.0 220650.0 88800.0 221850.0 ;
      RECT  87600.0 210750.0 88800.0 211950.0 ;
      RECT  83400.0 215400.0 84600.0 216600.0 ;
      RECT  83400.0 215400.0 84600.0 216600.0 ;
      RECT  85950.0 215550.0 86850.0 216450.0 ;
      RECT  81000.0 222750.0 90600.0 223650.0 ;
      RECT  81000.0 208950.0 90600.0 209850.0 ;
      RECT  53250.0 215400.0 54450.0 216600.0 ;
      RECT  55200.0 213000.0 56400.0 214200.0 ;
      RECT  72000.0 213900.0 70800.0 215100.0 ;
      RECT  63600.0 225150.0 64800.0 223200.0 ;
      RECT  63600.0 237000.0 64800.0 235050.0 ;
      RECT  58800.0 235650.0 60000.0 237450.0 ;
      RECT  58800.0 226350.0 60000.0 222750.0 ;
      RECT  61500.0 235650.0 62400.0 226350.0 ;
      RECT  58800.0 226350.0 60000.0 225150.0 ;
      RECT  61200.0 226350.0 62400.0 225150.0 ;
      RECT  61200.0 226350.0 62400.0 225150.0 ;
      RECT  58800.0 226350.0 60000.0 225150.0 ;
      RECT  58800.0 235650.0 60000.0 234450.0 ;
      RECT  61200.0 235650.0 62400.0 234450.0 ;
      RECT  61200.0 235650.0 62400.0 234450.0 ;
      RECT  58800.0 235650.0 60000.0 234450.0 ;
      RECT  63600.0 225750.0 64800.0 224550.0 ;
      RECT  63600.0 235650.0 64800.0 234450.0 ;
      RECT  59400.0 231000.0 60600.0 229800.0 ;
      RECT  59400.0 231000.0 60600.0 229800.0 ;
      RECT  61950.0 230850.0 62850.0 229950.0 ;
      RECT  57000.0 223650.0 66600.0 222750.0 ;
      RECT  57000.0 237450.0 66600.0 236550.0 ;
      RECT  68400.0 235050.0 69600.0 237450.0 ;
      RECT  68400.0 226350.0 69600.0 222750.0 ;
      RECT  73200.0 226350.0 74400.0 222750.0 ;
      RECT  75600.0 225150.0 76800.0 223200.0 ;
      RECT  75600.0 237000.0 76800.0 235050.0 ;
      RECT  68400.0 226350.0 69600.0 225150.0 ;
      RECT  70800.0 226350.0 72000.0 225150.0 ;
      RECT  70800.0 226350.0 72000.0 225150.0 ;
      RECT  68400.0 226350.0 69600.0 225150.0 ;
      RECT  70800.0 226350.0 72000.0 225150.0 ;
      RECT  73200.0 226350.0 74400.0 225150.0 ;
      RECT  73200.0 226350.0 74400.0 225150.0 ;
      RECT  70800.0 226350.0 72000.0 225150.0 ;
      RECT  68400.0 235050.0 69600.0 233850.0 ;
      RECT  70800.0 235050.0 72000.0 233850.0 ;
      RECT  70800.0 235050.0 72000.0 233850.0 ;
      RECT  68400.0 235050.0 69600.0 233850.0 ;
      RECT  70800.0 235050.0 72000.0 233850.0 ;
      RECT  73200.0 235050.0 74400.0 233850.0 ;
      RECT  73200.0 235050.0 74400.0 233850.0 ;
      RECT  70800.0 235050.0 72000.0 233850.0 ;
      RECT  75600.0 225750.0 76800.0 224550.0 ;
      RECT  75600.0 235650.0 76800.0 234450.0 ;
      RECT  73200.0 232500.0 72000.0 231300.0 ;
      RECT  70200.0 229800.0 69000.0 228600.0 ;
      RECT  70800.0 226350.0 72000.0 225150.0 ;
      RECT  73200.0 235050.0 74400.0 233850.0 ;
      RECT  74400.0 229800.0 73200.0 228600.0 ;
      RECT  69000.0 229800.0 70200.0 228600.0 ;
      RECT  72000.0 232500.0 73200.0 231300.0 ;
      RECT  73200.0 229800.0 74400.0 228600.0 ;
      RECT  66600.0 223650.0 81000.0 222750.0 ;
      RECT  66600.0 237450.0 81000.0 236550.0 ;
      RECT  87600.0 225150.0 88800.0 223200.0 ;
      RECT  87600.0 237000.0 88800.0 235050.0 ;
      RECT  82800.0 235650.0 84000.0 237450.0 ;
      RECT  82800.0 226350.0 84000.0 222750.0 ;
      RECT  85500.0 235650.0 86400.0 226350.0 ;
      RECT  82800.0 226350.0 84000.0 225150.0 ;
      RECT  85200.0 226350.0 86400.0 225150.0 ;
      RECT  85200.0 226350.0 86400.0 225150.0 ;
      RECT  82800.0 226350.0 84000.0 225150.0 ;
      RECT  82800.0 235650.0 84000.0 234450.0 ;
      RECT  85200.0 235650.0 86400.0 234450.0 ;
      RECT  85200.0 235650.0 86400.0 234450.0 ;
      RECT  82800.0 235650.0 84000.0 234450.0 ;
      RECT  87600.0 225750.0 88800.0 224550.0 ;
      RECT  87600.0 235650.0 88800.0 234450.0 ;
      RECT  83400.0 231000.0 84600.0 229800.0 ;
      RECT  83400.0 231000.0 84600.0 229800.0 ;
      RECT  85950.0 230850.0 86850.0 229950.0 ;
      RECT  81000.0 223650.0 90600.0 222750.0 ;
      RECT  81000.0 237450.0 90600.0 236550.0 ;
      RECT  53250.0 229800.0 54450.0 231000.0 ;
      RECT  55200.0 232200.0 56400.0 233400.0 ;
      RECT  72000.0 231300.0 70800.0 232500.0 ;
      RECT  63600.0 248850.0 64800.0 250800.0 ;
      RECT  63600.0 237000.0 64800.0 238950.0 ;
      RECT  58800.0 238350.0 60000.0 236550.0 ;
      RECT  58800.0 247650.0 60000.0 251250.0 ;
      RECT  61500.0 238350.0 62400.0 247650.0 ;
      RECT  58800.0 247650.0 60000.0 248850.0 ;
      RECT  61200.0 247650.0 62400.0 248850.0 ;
      RECT  61200.0 247650.0 62400.0 248850.0 ;
      RECT  58800.0 247650.0 60000.0 248850.0 ;
      RECT  58800.0 238350.0 60000.0 239550.0 ;
      RECT  61200.0 238350.0 62400.0 239550.0 ;
      RECT  61200.0 238350.0 62400.0 239550.0 ;
      RECT  58800.0 238350.0 60000.0 239550.0 ;
      RECT  63600.0 248250.0 64800.0 249450.0 ;
      RECT  63600.0 238350.0 64800.0 239550.0 ;
      RECT  59400.0 243000.0 60600.0 244200.0 ;
      RECT  59400.0 243000.0 60600.0 244200.0 ;
      RECT  61950.0 243150.0 62850.0 244050.0 ;
      RECT  57000.0 250350.0 66600.0 251250.0 ;
      RECT  57000.0 236550.0 66600.0 237450.0 ;
      RECT  68400.0 238950.0 69600.0 236550.0 ;
      RECT  68400.0 247650.0 69600.0 251250.0 ;
      RECT  73200.0 247650.0 74400.0 251250.0 ;
      RECT  75600.0 248850.0 76800.0 250800.0 ;
      RECT  75600.0 237000.0 76800.0 238950.0 ;
      RECT  68400.0 247650.0 69600.0 248850.0 ;
      RECT  70800.0 247650.0 72000.0 248850.0 ;
      RECT  70800.0 247650.0 72000.0 248850.0 ;
      RECT  68400.0 247650.0 69600.0 248850.0 ;
      RECT  70800.0 247650.0 72000.0 248850.0 ;
      RECT  73200.0 247650.0 74400.0 248850.0 ;
      RECT  73200.0 247650.0 74400.0 248850.0 ;
      RECT  70800.0 247650.0 72000.0 248850.0 ;
      RECT  68400.0 238950.0 69600.0 240150.0 ;
      RECT  70800.0 238950.0 72000.0 240150.0 ;
      RECT  70800.0 238950.0 72000.0 240150.0 ;
      RECT  68400.0 238950.0 69600.0 240150.0 ;
      RECT  70800.0 238950.0 72000.0 240150.0 ;
      RECT  73200.0 238950.0 74400.0 240150.0 ;
      RECT  73200.0 238950.0 74400.0 240150.0 ;
      RECT  70800.0 238950.0 72000.0 240150.0 ;
      RECT  75600.0 248250.0 76800.0 249450.0 ;
      RECT  75600.0 238350.0 76800.0 239550.0 ;
      RECT  73200.0 241500.0 72000.0 242700.0 ;
      RECT  70200.0 244200.0 69000.0 245400.0 ;
      RECT  70800.0 247650.0 72000.0 248850.0 ;
      RECT  73200.0 238950.0 74400.0 240150.0 ;
      RECT  74400.0 244200.0 73200.0 245400.0 ;
      RECT  69000.0 244200.0 70200.0 245400.0 ;
      RECT  72000.0 241500.0 73200.0 242700.0 ;
      RECT  73200.0 244200.0 74400.0 245400.0 ;
      RECT  66600.0 250350.0 81000.0 251250.0 ;
      RECT  66600.0 236550.0 81000.0 237450.0 ;
      RECT  87600.0 248850.0 88800.0 250800.0 ;
      RECT  87600.0 237000.0 88800.0 238950.0 ;
      RECT  82800.0 238350.0 84000.0 236550.0 ;
      RECT  82800.0 247650.0 84000.0 251250.0 ;
      RECT  85500.0 238350.0 86400.0 247650.0 ;
      RECT  82800.0 247650.0 84000.0 248850.0 ;
      RECT  85200.0 247650.0 86400.0 248850.0 ;
      RECT  85200.0 247650.0 86400.0 248850.0 ;
      RECT  82800.0 247650.0 84000.0 248850.0 ;
      RECT  82800.0 238350.0 84000.0 239550.0 ;
      RECT  85200.0 238350.0 86400.0 239550.0 ;
      RECT  85200.0 238350.0 86400.0 239550.0 ;
      RECT  82800.0 238350.0 84000.0 239550.0 ;
      RECT  87600.0 248250.0 88800.0 249450.0 ;
      RECT  87600.0 238350.0 88800.0 239550.0 ;
      RECT  83400.0 243000.0 84600.0 244200.0 ;
      RECT  83400.0 243000.0 84600.0 244200.0 ;
      RECT  85950.0 243150.0 86850.0 244050.0 ;
      RECT  81000.0 250350.0 90600.0 251250.0 ;
      RECT  81000.0 236550.0 90600.0 237450.0 ;
      RECT  53250.0 243000.0 54450.0 244200.0 ;
      RECT  55200.0 240600.0 56400.0 241800.0 ;
      RECT  72000.0 241500.0 70800.0 242700.0 ;
      RECT  63600.0 252750.0 64800.0 250800.0 ;
      RECT  63600.0 264600.0 64800.0 262650.0 ;
      RECT  58800.0 263250.0 60000.0 265050.0 ;
      RECT  58800.0 253950.0 60000.0 250350.0 ;
      RECT  61500.0 263250.0 62400.0 253950.0 ;
      RECT  58800.0 253950.0 60000.0 252750.0 ;
      RECT  61200.0 253950.0 62400.0 252750.0 ;
      RECT  61200.0 253950.0 62400.0 252750.0 ;
      RECT  58800.0 253950.0 60000.0 252750.0 ;
      RECT  58800.0 263250.0 60000.0 262050.0 ;
      RECT  61200.0 263250.0 62400.0 262050.0 ;
      RECT  61200.0 263250.0 62400.0 262050.0 ;
      RECT  58800.0 263250.0 60000.0 262050.0 ;
      RECT  63600.0 253350.0 64800.0 252150.0 ;
      RECT  63600.0 263250.0 64800.0 262050.0 ;
      RECT  59400.0 258600.0 60600.0 257400.0 ;
      RECT  59400.0 258600.0 60600.0 257400.0 ;
      RECT  61950.0 258450.0 62850.0 257550.0 ;
      RECT  57000.0 251250.0 66600.0 250350.0 ;
      RECT  57000.0 265050.0 66600.0 264150.0 ;
      RECT  68400.0 262650.0 69600.0 265050.0 ;
      RECT  68400.0 253950.0 69600.0 250350.0 ;
      RECT  73200.0 253950.0 74400.0 250350.0 ;
      RECT  75600.0 252750.0 76800.0 250800.0 ;
      RECT  75600.0 264600.0 76800.0 262650.0 ;
      RECT  68400.0 253950.0 69600.0 252750.0 ;
      RECT  70800.0 253950.0 72000.0 252750.0 ;
      RECT  70800.0 253950.0 72000.0 252750.0 ;
      RECT  68400.0 253950.0 69600.0 252750.0 ;
      RECT  70800.0 253950.0 72000.0 252750.0 ;
      RECT  73200.0 253950.0 74400.0 252750.0 ;
      RECT  73200.0 253950.0 74400.0 252750.0 ;
      RECT  70800.0 253950.0 72000.0 252750.0 ;
      RECT  68400.0 262650.0 69600.0 261450.0 ;
      RECT  70800.0 262650.0 72000.0 261450.0 ;
      RECT  70800.0 262650.0 72000.0 261450.0 ;
      RECT  68400.0 262650.0 69600.0 261450.0 ;
      RECT  70800.0 262650.0 72000.0 261450.0 ;
      RECT  73200.0 262650.0 74400.0 261450.0 ;
      RECT  73200.0 262650.0 74400.0 261450.0 ;
      RECT  70800.0 262650.0 72000.0 261450.0 ;
      RECT  75600.0 253350.0 76800.0 252150.0 ;
      RECT  75600.0 263250.0 76800.0 262050.0 ;
      RECT  73200.0 260100.0 72000.0 258900.0 ;
      RECT  70200.0 257400.0 69000.0 256200.0 ;
      RECT  70800.0 253950.0 72000.0 252750.0 ;
      RECT  73200.0 262650.0 74400.0 261450.0 ;
      RECT  74400.0 257400.0 73200.0 256200.0 ;
      RECT  69000.0 257400.0 70200.0 256200.0 ;
      RECT  72000.0 260100.0 73200.0 258900.0 ;
      RECT  73200.0 257400.0 74400.0 256200.0 ;
      RECT  66600.0 251250.0 81000.0 250350.0 ;
      RECT  66600.0 265050.0 81000.0 264150.0 ;
      RECT  87600.0 252750.0 88800.0 250800.0 ;
      RECT  87600.0 264600.0 88800.0 262650.0 ;
      RECT  82800.0 263250.0 84000.0 265050.0 ;
      RECT  82800.0 253950.0 84000.0 250350.0 ;
      RECT  85500.0 263250.0 86400.0 253950.0 ;
      RECT  82800.0 253950.0 84000.0 252750.0 ;
      RECT  85200.0 253950.0 86400.0 252750.0 ;
      RECT  85200.0 253950.0 86400.0 252750.0 ;
      RECT  82800.0 253950.0 84000.0 252750.0 ;
      RECT  82800.0 263250.0 84000.0 262050.0 ;
      RECT  85200.0 263250.0 86400.0 262050.0 ;
      RECT  85200.0 263250.0 86400.0 262050.0 ;
      RECT  82800.0 263250.0 84000.0 262050.0 ;
      RECT  87600.0 253350.0 88800.0 252150.0 ;
      RECT  87600.0 263250.0 88800.0 262050.0 ;
      RECT  83400.0 258600.0 84600.0 257400.0 ;
      RECT  83400.0 258600.0 84600.0 257400.0 ;
      RECT  85950.0 258450.0 86850.0 257550.0 ;
      RECT  81000.0 251250.0 90600.0 250350.0 ;
      RECT  81000.0 265050.0 90600.0 264150.0 ;
      RECT  53250.0 257400.0 54450.0 258600.0 ;
      RECT  55200.0 259800.0 56400.0 261000.0 ;
      RECT  72000.0 258900.0 70800.0 260100.0 ;
      RECT  63600.0 276450.0 64800.0 278400.0 ;
      RECT  63600.0 264600.0 64800.0 266550.0 ;
      RECT  58800.0 265950.0 60000.0 264150.0 ;
      RECT  58800.0 275250.0 60000.0 278850.0 ;
      RECT  61500.0 265950.0 62400.0 275250.0 ;
      RECT  58800.0 275250.0 60000.0 276450.0 ;
      RECT  61200.0 275250.0 62400.0 276450.0 ;
      RECT  61200.0 275250.0 62400.0 276450.0 ;
      RECT  58800.0 275250.0 60000.0 276450.0 ;
      RECT  58800.0 265950.0 60000.0 267150.0 ;
      RECT  61200.0 265950.0 62400.0 267150.0 ;
      RECT  61200.0 265950.0 62400.0 267150.0 ;
      RECT  58800.0 265950.0 60000.0 267150.0 ;
      RECT  63600.0 275850.0 64800.0 277050.0 ;
      RECT  63600.0 265950.0 64800.0 267150.0 ;
      RECT  59400.0 270600.0 60600.0 271800.0 ;
      RECT  59400.0 270600.0 60600.0 271800.0 ;
      RECT  61950.0 270750.0 62850.0 271650.0 ;
      RECT  57000.0 277950.0 66600.0 278850.0 ;
      RECT  57000.0 264150.0 66600.0 265050.0 ;
      RECT  68400.0 266550.0 69600.0 264150.0 ;
      RECT  68400.0 275250.0 69600.0 278850.0 ;
      RECT  73200.0 275250.0 74400.0 278850.0 ;
      RECT  75600.0 276450.0 76800.0 278400.0 ;
      RECT  75600.0 264600.0 76800.0 266550.0 ;
      RECT  68400.0 275250.0 69600.0 276450.0 ;
      RECT  70800.0 275250.0 72000.0 276450.0 ;
      RECT  70800.0 275250.0 72000.0 276450.0 ;
      RECT  68400.0 275250.0 69600.0 276450.0 ;
      RECT  70800.0 275250.0 72000.0 276450.0 ;
      RECT  73200.0 275250.0 74400.0 276450.0 ;
      RECT  73200.0 275250.0 74400.0 276450.0 ;
      RECT  70800.0 275250.0 72000.0 276450.0 ;
      RECT  68400.0 266550.0 69600.0 267750.0 ;
      RECT  70800.0 266550.0 72000.0 267750.0 ;
      RECT  70800.0 266550.0 72000.0 267750.0 ;
      RECT  68400.0 266550.0 69600.0 267750.0 ;
      RECT  70800.0 266550.0 72000.0 267750.0 ;
      RECT  73200.0 266550.0 74400.0 267750.0 ;
      RECT  73200.0 266550.0 74400.0 267750.0 ;
      RECT  70800.0 266550.0 72000.0 267750.0 ;
      RECT  75600.0 275850.0 76800.0 277050.0 ;
      RECT  75600.0 265950.0 76800.0 267150.0 ;
      RECT  73200.0 269100.0 72000.0 270300.0 ;
      RECT  70200.0 271800.0 69000.0 273000.0 ;
      RECT  70800.0 275250.0 72000.0 276450.0 ;
      RECT  73200.0 266550.0 74400.0 267750.0 ;
      RECT  74400.0 271800.0 73200.0 273000.0 ;
      RECT  69000.0 271800.0 70200.0 273000.0 ;
      RECT  72000.0 269100.0 73200.0 270300.0 ;
      RECT  73200.0 271800.0 74400.0 273000.0 ;
      RECT  66600.0 277950.0 81000.0 278850.0 ;
      RECT  66600.0 264150.0 81000.0 265050.0 ;
      RECT  87600.0 276450.0 88800.0 278400.0 ;
      RECT  87600.0 264600.0 88800.0 266550.0 ;
      RECT  82800.0 265950.0 84000.0 264150.0 ;
      RECT  82800.0 275250.0 84000.0 278850.0 ;
      RECT  85500.0 265950.0 86400.0 275250.0 ;
      RECT  82800.0 275250.0 84000.0 276450.0 ;
      RECT  85200.0 275250.0 86400.0 276450.0 ;
      RECT  85200.0 275250.0 86400.0 276450.0 ;
      RECT  82800.0 275250.0 84000.0 276450.0 ;
      RECT  82800.0 265950.0 84000.0 267150.0 ;
      RECT  85200.0 265950.0 86400.0 267150.0 ;
      RECT  85200.0 265950.0 86400.0 267150.0 ;
      RECT  82800.0 265950.0 84000.0 267150.0 ;
      RECT  87600.0 275850.0 88800.0 277050.0 ;
      RECT  87600.0 265950.0 88800.0 267150.0 ;
      RECT  83400.0 270600.0 84600.0 271800.0 ;
      RECT  83400.0 270600.0 84600.0 271800.0 ;
      RECT  85950.0 270750.0 86850.0 271650.0 ;
      RECT  81000.0 277950.0 90600.0 278850.0 ;
      RECT  81000.0 264150.0 90600.0 265050.0 ;
      RECT  53250.0 270600.0 54450.0 271800.0 ;
      RECT  55200.0 268200.0 56400.0 269400.0 ;
      RECT  72000.0 269100.0 70800.0 270300.0 ;
      RECT  63600.0 280350.0 64800.0 278400.0 ;
      RECT  63600.0 292200.0 64800.0 290250.0 ;
      RECT  58800.0 290850.0 60000.0 292650.0 ;
      RECT  58800.0 281550.0 60000.0 277950.0 ;
      RECT  61500.0 290850.0 62400.0 281550.0 ;
      RECT  58800.0 281550.0 60000.0 280350.0 ;
      RECT  61200.0 281550.0 62400.0 280350.0 ;
      RECT  61200.0 281550.0 62400.0 280350.0 ;
      RECT  58800.0 281550.0 60000.0 280350.0 ;
      RECT  58800.0 290850.0 60000.0 289650.0 ;
      RECT  61200.0 290850.0 62400.0 289650.0 ;
      RECT  61200.0 290850.0 62400.0 289650.0 ;
      RECT  58800.0 290850.0 60000.0 289650.0 ;
      RECT  63600.0 280950.0 64800.0 279750.0 ;
      RECT  63600.0 290850.0 64800.0 289650.0 ;
      RECT  59400.0 286200.0 60600.0 285000.0 ;
      RECT  59400.0 286200.0 60600.0 285000.0 ;
      RECT  61950.0 286050.0 62850.0 285150.0 ;
      RECT  57000.0 278850.0 66600.0 277950.0 ;
      RECT  57000.0 292650.0 66600.0 291750.0 ;
      RECT  68400.0 290250.0 69600.0 292650.0 ;
      RECT  68400.0 281550.0 69600.0 277950.0 ;
      RECT  73200.0 281550.0 74400.0 277950.0 ;
      RECT  75600.0 280350.0 76800.0 278400.0 ;
      RECT  75600.0 292200.0 76800.0 290250.0 ;
      RECT  68400.0 281550.0 69600.0 280350.0 ;
      RECT  70800.0 281550.0 72000.0 280350.0 ;
      RECT  70800.0 281550.0 72000.0 280350.0 ;
      RECT  68400.0 281550.0 69600.0 280350.0 ;
      RECT  70800.0 281550.0 72000.0 280350.0 ;
      RECT  73200.0 281550.0 74400.0 280350.0 ;
      RECT  73200.0 281550.0 74400.0 280350.0 ;
      RECT  70800.0 281550.0 72000.0 280350.0 ;
      RECT  68400.0 290250.0 69600.0 289050.0 ;
      RECT  70800.0 290250.0 72000.0 289050.0 ;
      RECT  70800.0 290250.0 72000.0 289050.0 ;
      RECT  68400.0 290250.0 69600.0 289050.0 ;
      RECT  70800.0 290250.0 72000.0 289050.0 ;
      RECT  73200.0 290250.0 74400.0 289050.0 ;
      RECT  73200.0 290250.0 74400.0 289050.0 ;
      RECT  70800.0 290250.0 72000.0 289050.0 ;
      RECT  75600.0 280950.0 76800.0 279750.0 ;
      RECT  75600.0 290850.0 76800.0 289650.0 ;
      RECT  73200.0 287700.0 72000.0 286500.0 ;
      RECT  70200.0 285000.0 69000.0 283800.0 ;
      RECT  70800.0 281550.0 72000.0 280350.0 ;
      RECT  73200.0 290250.0 74400.0 289050.0 ;
      RECT  74400.0 285000.0 73200.0 283800.0 ;
      RECT  69000.0 285000.0 70200.0 283800.0 ;
      RECT  72000.0 287700.0 73200.0 286500.0 ;
      RECT  73200.0 285000.0 74400.0 283800.0 ;
      RECT  66600.0 278850.0 81000.0 277950.0 ;
      RECT  66600.0 292650.0 81000.0 291750.0 ;
      RECT  87600.0 280350.0 88800.0 278400.0 ;
      RECT  87600.0 292200.0 88800.0 290250.0 ;
      RECT  82800.0 290850.0 84000.0 292650.0 ;
      RECT  82800.0 281550.0 84000.0 277950.0 ;
      RECT  85500.0 290850.0 86400.0 281550.0 ;
      RECT  82800.0 281550.0 84000.0 280350.0 ;
      RECT  85200.0 281550.0 86400.0 280350.0 ;
      RECT  85200.0 281550.0 86400.0 280350.0 ;
      RECT  82800.0 281550.0 84000.0 280350.0 ;
      RECT  82800.0 290850.0 84000.0 289650.0 ;
      RECT  85200.0 290850.0 86400.0 289650.0 ;
      RECT  85200.0 290850.0 86400.0 289650.0 ;
      RECT  82800.0 290850.0 84000.0 289650.0 ;
      RECT  87600.0 280950.0 88800.0 279750.0 ;
      RECT  87600.0 290850.0 88800.0 289650.0 ;
      RECT  83400.0 286200.0 84600.0 285000.0 ;
      RECT  83400.0 286200.0 84600.0 285000.0 ;
      RECT  85950.0 286050.0 86850.0 285150.0 ;
      RECT  81000.0 278850.0 90600.0 277950.0 ;
      RECT  81000.0 292650.0 90600.0 291750.0 ;
      RECT  53250.0 285000.0 54450.0 286200.0 ;
      RECT  55200.0 287400.0 56400.0 288600.0 ;
      RECT  72000.0 286500.0 70800.0 287700.0 ;
      RECT  63600.0 304050.0 64800.0 306000.0 ;
      RECT  63600.0 292200.0 64800.0 294150.0 ;
      RECT  58800.0 293550.0 60000.0 291750.0 ;
      RECT  58800.0 302850.0 60000.0 306450.0 ;
      RECT  61500.0 293550.0 62400.0 302850.0 ;
      RECT  58800.0 302850.0 60000.0 304050.0 ;
      RECT  61200.0 302850.0 62400.0 304050.0 ;
      RECT  61200.0 302850.0 62400.0 304050.0 ;
      RECT  58800.0 302850.0 60000.0 304050.0 ;
      RECT  58800.0 293550.0 60000.0 294750.0 ;
      RECT  61200.0 293550.0 62400.0 294750.0 ;
      RECT  61200.0 293550.0 62400.0 294750.0 ;
      RECT  58800.0 293550.0 60000.0 294750.0 ;
      RECT  63600.0 303450.0 64800.0 304650.0 ;
      RECT  63600.0 293550.0 64800.0 294750.0 ;
      RECT  59400.0 298200.0 60600.0 299400.0 ;
      RECT  59400.0 298200.0 60600.0 299400.0 ;
      RECT  61950.0 298350.0 62850.0 299250.0 ;
      RECT  57000.0 305550.0 66600.0 306450.0 ;
      RECT  57000.0 291750.0 66600.0 292650.0 ;
      RECT  68400.0 294150.0 69600.0 291750.0 ;
      RECT  68400.0 302850.0 69600.0 306450.0 ;
      RECT  73200.0 302850.0 74400.0 306450.0 ;
      RECT  75600.0 304050.0 76800.0 306000.0 ;
      RECT  75600.0 292200.0 76800.0 294150.0 ;
      RECT  68400.0 302850.0 69600.0 304050.0 ;
      RECT  70800.0 302850.0 72000.0 304050.0 ;
      RECT  70800.0 302850.0 72000.0 304050.0 ;
      RECT  68400.0 302850.0 69600.0 304050.0 ;
      RECT  70800.0 302850.0 72000.0 304050.0 ;
      RECT  73200.0 302850.0 74400.0 304050.0 ;
      RECT  73200.0 302850.0 74400.0 304050.0 ;
      RECT  70800.0 302850.0 72000.0 304050.0 ;
      RECT  68400.0 294150.0 69600.0 295350.0 ;
      RECT  70800.0 294150.0 72000.0 295350.0 ;
      RECT  70800.0 294150.0 72000.0 295350.0 ;
      RECT  68400.0 294150.0 69600.0 295350.0 ;
      RECT  70800.0 294150.0 72000.0 295350.0 ;
      RECT  73200.0 294150.0 74400.0 295350.0 ;
      RECT  73200.0 294150.0 74400.0 295350.0 ;
      RECT  70800.0 294150.0 72000.0 295350.0 ;
      RECT  75600.0 303450.0 76800.0 304650.0 ;
      RECT  75600.0 293550.0 76800.0 294750.0 ;
      RECT  73200.0 296700.0 72000.0 297900.0 ;
      RECT  70200.0 299400.0 69000.0 300600.0 ;
      RECT  70800.0 302850.0 72000.0 304050.0 ;
      RECT  73200.0 294150.0 74400.0 295350.0 ;
      RECT  74400.0 299400.0 73200.0 300600.0 ;
      RECT  69000.0 299400.0 70200.0 300600.0 ;
      RECT  72000.0 296700.0 73200.0 297900.0 ;
      RECT  73200.0 299400.0 74400.0 300600.0 ;
      RECT  66600.0 305550.0 81000.0 306450.0 ;
      RECT  66600.0 291750.0 81000.0 292650.0 ;
      RECT  87600.0 304050.0 88800.0 306000.0 ;
      RECT  87600.0 292200.0 88800.0 294150.0 ;
      RECT  82800.0 293550.0 84000.0 291750.0 ;
      RECT  82800.0 302850.0 84000.0 306450.0 ;
      RECT  85500.0 293550.0 86400.0 302850.0 ;
      RECT  82800.0 302850.0 84000.0 304050.0 ;
      RECT  85200.0 302850.0 86400.0 304050.0 ;
      RECT  85200.0 302850.0 86400.0 304050.0 ;
      RECT  82800.0 302850.0 84000.0 304050.0 ;
      RECT  82800.0 293550.0 84000.0 294750.0 ;
      RECT  85200.0 293550.0 86400.0 294750.0 ;
      RECT  85200.0 293550.0 86400.0 294750.0 ;
      RECT  82800.0 293550.0 84000.0 294750.0 ;
      RECT  87600.0 303450.0 88800.0 304650.0 ;
      RECT  87600.0 293550.0 88800.0 294750.0 ;
      RECT  83400.0 298200.0 84600.0 299400.0 ;
      RECT  83400.0 298200.0 84600.0 299400.0 ;
      RECT  85950.0 298350.0 86850.0 299250.0 ;
      RECT  81000.0 305550.0 90600.0 306450.0 ;
      RECT  81000.0 291750.0 90600.0 292650.0 ;
      RECT  53250.0 298200.0 54450.0 299400.0 ;
      RECT  55200.0 295800.0 56400.0 297000.0 ;
      RECT  72000.0 296700.0 70800.0 297900.0 ;
      RECT  63600.0 307950.0 64800.0 306000.0 ;
      RECT  63600.0 319800.0 64800.0 317850.0 ;
      RECT  58800.0 318450.0 60000.0 320250.0 ;
      RECT  58800.0 309150.0 60000.0 305550.0 ;
      RECT  61500.0 318450.0 62400.0 309150.0 ;
      RECT  58800.0 309150.0 60000.0 307950.0 ;
      RECT  61200.0 309150.0 62400.0 307950.0 ;
      RECT  61200.0 309150.0 62400.0 307950.0 ;
      RECT  58800.0 309150.0 60000.0 307950.0 ;
      RECT  58800.0 318450.0 60000.0 317250.0 ;
      RECT  61200.0 318450.0 62400.0 317250.0 ;
      RECT  61200.0 318450.0 62400.0 317250.0 ;
      RECT  58800.0 318450.0 60000.0 317250.0 ;
      RECT  63600.0 308550.0 64800.0 307350.0 ;
      RECT  63600.0 318450.0 64800.0 317250.0 ;
      RECT  59400.0 313800.0 60600.0 312600.0 ;
      RECT  59400.0 313800.0 60600.0 312600.0 ;
      RECT  61950.0 313650.0 62850.0 312750.0 ;
      RECT  57000.0 306450.0 66600.0 305550.0 ;
      RECT  57000.0 320250.0 66600.0 319350.0 ;
      RECT  68400.0 317850.0 69600.0 320250.0 ;
      RECT  68400.0 309150.0 69600.0 305550.0 ;
      RECT  73200.0 309150.0 74400.0 305550.0 ;
      RECT  75600.0 307950.0 76800.0 306000.0 ;
      RECT  75600.0 319800.0 76800.0 317850.0 ;
      RECT  68400.0 309150.0 69600.0 307950.0 ;
      RECT  70800.0 309150.0 72000.0 307950.0 ;
      RECT  70800.0 309150.0 72000.0 307950.0 ;
      RECT  68400.0 309150.0 69600.0 307950.0 ;
      RECT  70800.0 309150.0 72000.0 307950.0 ;
      RECT  73200.0 309150.0 74400.0 307950.0 ;
      RECT  73200.0 309150.0 74400.0 307950.0 ;
      RECT  70800.0 309150.0 72000.0 307950.0 ;
      RECT  68400.0 317850.0 69600.0 316650.0 ;
      RECT  70800.0 317850.0 72000.0 316650.0 ;
      RECT  70800.0 317850.0 72000.0 316650.0 ;
      RECT  68400.0 317850.0 69600.0 316650.0 ;
      RECT  70800.0 317850.0 72000.0 316650.0 ;
      RECT  73200.0 317850.0 74400.0 316650.0 ;
      RECT  73200.0 317850.0 74400.0 316650.0 ;
      RECT  70800.0 317850.0 72000.0 316650.0 ;
      RECT  75600.0 308550.0 76800.0 307350.0 ;
      RECT  75600.0 318450.0 76800.0 317250.0 ;
      RECT  73200.0 315300.0 72000.0 314100.0 ;
      RECT  70200.0 312600.0 69000.0 311400.0 ;
      RECT  70800.0 309150.0 72000.0 307950.0 ;
      RECT  73200.0 317850.0 74400.0 316650.0 ;
      RECT  74400.0 312600.0 73200.0 311400.0 ;
      RECT  69000.0 312600.0 70200.0 311400.0 ;
      RECT  72000.0 315300.0 73200.0 314100.0 ;
      RECT  73200.0 312600.0 74400.0 311400.0 ;
      RECT  66600.0 306450.0 81000.0 305550.0 ;
      RECT  66600.0 320250.0 81000.0 319350.0 ;
      RECT  87600.0 307950.0 88800.0 306000.0 ;
      RECT  87600.0 319800.0 88800.0 317850.0 ;
      RECT  82800.0 318450.0 84000.0 320250.0 ;
      RECT  82800.0 309150.0 84000.0 305550.0 ;
      RECT  85500.0 318450.0 86400.0 309150.0 ;
      RECT  82800.0 309150.0 84000.0 307950.0 ;
      RECT  85200.0 309150.0 86400.0 307950.0 ;
      RECT  85200.0 309150.0 86400.0 307950.0 ;
      RECT  82800.0 309150.0 84000.0 307950.0 ;
      RECT  82800.0 318450.0 84000.0 317250.0 ;
      RECT  85200.0 318450.0 86400.0 317250.0 ;
      RECT  85200.0 318450.0 86400.0 317250.0 ;
      RECT  82800.0 318450.0 84000.0 317250.0 ;
      RECT  87600.0 308550.0 88800.0 307350.0 ;
      RECT  87600.0 318450.0 88800.0 317250.0 ;
      RECT  83400.0 313800.0 84600.0 312600.0 ;
      RECT  83400.0 313800.0 84600.0 312600.0 ;
      RECT  85950.0 313650.0 86850.0 312750.0 ;
      RECT  81000.0 306450.0 90600.0 305550.0 ;
      RECT  81000.0 320250.0 90600.0 319350.0 ;
      RECT  53250.0 312600.0 54450.0 313800.0 ;
      RECT  55200.0 315000.0 56400.0 316200.0 ;
      RECT  72000.0 314100.0 70800.0 315300.0 ;
      RECT  63600.0 331650.0 64800.0 333600.0 ;
      RECT  63600.0 319800.0 64800.0 321750.0 ;
      RECT  58800.0 321150.0 60000.0 319350.0 ;
      RECT  58800.0 330450.0 60000.0 334050.0 ;
      RECT  61500.0 321150.0 62400.0 330450.0 ;
      RECT  58800.0 330450.0 60000.0 331650.0 ;
      RECT  61200.0 330450.0 62400.0 331650.0 ;
      RECT  61200.0 330450.0 62400.0 331650.0 ;
      RECT  58800.0 330450.0 60000.0 331650.0 ;
      RECT  58800.0 321150.0 60000.0 322350.0 ;
      RECT  61200.0 321150.0 62400.0 322350.0 ;
      RECT  61200.0 321150.0 62400.0 322350.0 ;
      RECT  58800.0 321150.0 60000.0 322350.0 ;
      RECT  63600.0 331050.0 64800.0 332250.0 ;
      RECT  63600.0 321150.0 64800.0 322350.0 ;
      RECT  59400.0 325800.0 60600.0 327000.0 ;
      RECT  59400.0 325800.0 60600.0 327000.0 ;
      RECT  61950.0 325950.0 62850.0 326850.0 ;
      RECT  57000.0 333150.0 66600.0 334050.0 ;
      RECT  57000.0 319350.0 66600.0 320250.0 ;
      RECT  68400.0 321750.0 69600.0 319350.0 ;
      RECT  68400.0 330450.0 69600.0 334050.0 ;
      RECT  73200.0 330450.0 74400.0 334050.0 ;
      RECT  75600.0 331650.0 76800.0 333600.0 ;
      RECT  75600.0 319800.0 76800.0 321750.0 ;
      RECT  68400.0 330450.0 69600.0 331650.0 ;
      RECT  70800.0 330450.0 72000.0 331650.0 ;
      RECT  70800.0 330450.0 72000.0 331650.0 ;
      RECT  68400.0 330450.0 69600.0 331650.0 ;
      RECT  70800.0 330450.0 72000.0 331650.0 ;
      RECT  73200.0 330450.0 74400.0 331650.0 ;
      RECT  73200.0 330450.0 74400.0 331650.0 ;
      RECT  70800.0 330450.0 72000.0 331650.0 ;
      RECT  68400.0 321750.0 69600.0 322950.0 ;
      RECT  70800.0 321750.0 72000.0 322950.0 ;
      RECT  70800.0 321750.0 72000.0 322950.0 ;
      RECT  68400.0 321750.0 69600.0 322950.0 ;
      RECT  70800.0 321750.0 72000.0 322950.0 ;
      RECT  73200.0 321750.0 74400.0 322950.0 ;
      RECT  73200.0 321750.0 74400.0 322950.0 ;
      RECT  70800.0 321750.0 72000.0 322950.0 ;
      RECT  75600.0 331050.0 76800.0 332250.0 ;
      RECT  75600.0 321150.0 76800.0 322350.0 ;
      RECT  73200.0 324300.0 72000.0 325500.0 ;
      RECT  70200.0 327000.0 69000.0 328200.0 ;
      RECT  70800.0 330450.0 72000.0 331650.0 ;
      RECT  73200.0 321750.0 74400.0 322950.0 ;
      RECT  74400.0 327000.0 73200.0 328200.0 ;
      RECT  69000.0 327000.0 70200.0 328200.0 ;
      RECT  72000.0 324300.0 73200.0 325500.0 ;
      RECT  73200.0 327000.0 74400.0 328200.0 ;
      RECT  66600.0 333150.0 81000.0 334050.0 ;
      RECT  66600.0 319350.0 81000.0 320250.0 ;
      RECT  87600.0 331650.0 88800.0 333600.0 ;
      RECT  87600.0 319800.0 88800.0 321750.0 ;
      RECT  82800.0 321150.0 84000.0 319350.0 ;
      RECT  82800.0 330450.0 84000.0 334050.0 ;
      RECT  85500.0 321150.0 86400.0 330450.0 ;
      RECT  82800.0 330450.0 84000.0 331650.0 ;
      RECT  85200.0 330450.0 86400.0 331650.0 ;
      RECT  85200.0 330450.0 86400.0 331650.0 ;
      RECT  82800.0 330450.0 84000.0 331650.0 ;
      RECT  82800.0 321150.0 84000.0 322350.0 ;
      RECT  85200.0 321150.0 86400.0 322350.0 ;
      RECT  85200.0 321150.0 86400.0 322350.0 ;
      RECT  82800.0 321150.0 84000.0 322350.0 ;
      RECT  87600.0 331050.0 88800.0 332250.0 ;
      RECT  87600.0 321150.0 88800.0 322350.0 ;
      RECT  83400.0 325800.0 84600.0 327000.0 ;
      RECT  83400.0 325800.0 84600.0 327000.0 ;
      RECT  85950.0 325950.0 86850.0 326850.0 ;
      RECT  81000.0 333150.0 90600.0 334050.0 ;
      RECT  81000.0 319350.0 90600.0 320250.0 ;
      RECT  53250.0 325800.0 54450.0 327000.0 ;
      RECT  55200.0 323400.0 56400.0 324600.0 ;
      RECT  72000.0 324300.0 70800.0 325500.0 ;
      RECT  63600.0 335550.0 64800.0 333600.0 ;
      RECT  63600.0 347400.0 64800.0 345450.0 ;
      RECT  58800.0 346050.0 60000.0 347850.0 ;
      RECT  58800.0 336750.0 60000.0 333150.0 ;
      RECT  61500.0 346050.0 62400.0 336750.0 ;
      RECT  58800.0 336750.0 60000.0 335550.0 ;
      RECT  61200.0 336750.0 62400.0 335550.0 ;
      RECT  61200.0 336750.0 62400.0 335550.0 ;
      RECT  58800.0 336750.0 60000.0 335550.0 ;
      RECT  58800.0 346050.0 60000.0 344850.0 ;
      RECT  61200.0 346050.0 62400.0 344850.0 ;
      RECT  61200.0 346050.0 62400.0 344850.0 ;
      RECT  58800.0 346050.0 60000.0 344850.0 ;
      RECT  63600.0 336150.0 64800.0 334950.0 ;
      RECT  63600.0 346050.0 64800.0 344850.0 ;
      RECT  59400.0 341400.0 60600.0 340200.0 ;
      RECT  59400.0 341400.0 60600.0 340200.0 ;
      RECT  61950.0 341250.0 62850.0 340350.0 ;
      RECT  57000.0 334050.0 66600.0 333150.0 ;
      RECT  57000.0 347850.0 66600.0 346950.0 ;
      RECT  68400.0 345450.0 69600.0 347850.0 ;
      RECT  68400.0 336750.0 69600.0 333150.0 ;
      RECT  73200.0 336750.0 74400.0 333150.0 ;
      RECT  75600.0 335550.0 76800.0 333600.0 ;
      RECT  75600.0 347400.0 76800.0 345450.0 ;
      RECT  68400.0 336750.0 69600.0 335550.0 ;
      RECT  70800.0 336750.0 72000.0 335550.0 ;
      RECT  70800.0 336750.0 72000.0 335550.0 ;
      RECT  68400.0 336750.0 69600.0 335550.0 ;
      RECT  70800.0 336750.0 72000.0 335550.0 ;
      RECT  73200.0 336750.0 74400.0 335550.0 ;
      RECT  73200.0 336750.0 74400.0 335550.0 ;
      RECT  70800.0 336750.0 72000.0 335550.0 ;
      RECT  68400.0 345450.0 69600.0 344250.0 ;
      RECT  70800.0 345450.0 72000.0 344250.0 ;
      RECT  70800.0 345450.0 72000.0 344250.0 ;
      RECT  68400.0 345450.0 69600.0 344250.0 ;
      RECT  70800.0 345450.0 72000.0 344250.0 ;
      RECT  73200.0 345450.0 74400.0 344250.0 ;
      RECT  73200.0 345450.0 74400.0 344250.0 ;
      RECT  70800.0 345450.0 72000.0 344250.0 ;
      RECT  75600.0 336150.0 76800.0 334950.0 ;
      RECT  75600.0 346050.0 76800.0 344850.0 ;
      RECT  73200.0 342900.0 72000.0 341700.0 ;
      RECT  70200.0 340200.0 69000.0 339000.0 ;
      RECT  70800.0 336750.0 72000.0 335550.0 ;
      RECT  73200.0 345450.0 74400.0 344250.0 ;
      RECT  74400.0 340200.0 73200.0 339000.0 ;
      RECT  69000.0 340200.0 70200.0 339000.0 ;
      RECT  72000.0 342900.0 73200.0 341700.0 ;
      RECT  73200.0 340200.0 74400.0 339000.0 ;
      RECT  66600.0 334050.0 81000.0 333150.0 ;
      RECT  66600.0 347850.0 81000.0 346950.0 ;
      RECT  87600.0 335550.0 88800.0 333600.0 ;
      RECT  87600.0 347400.0 88800.0 345450.0 ;
      RECT  82800.0 346050.0 84000.0 347850.0 ;
      RECT  82800.0 336750.0 84000.0 333150.0 ;
      RECT  85500.0 346050.0 86400.0 336750.0 ;
      RECT  82800.0 336750.0 84000.0 335550.0 ;
      RECT  85200.0 336750.0 86400.0 335550.0 ;
      RECT  85200.0 336750.0 86400.0 335550.0 ;
      RECT  82800.0 336750.0 84000.0 335550.0 ;
      RECT  82800.0 346050.0 84000.0 344850.0 ;
      RECT  85200.0 346050.0 86400.0 344850.0 ;
      RECT  85200.0 346050.0 86400.0 344850.0 ;
      RECT  82800.0 346050.0 84000.0 344850.0 ;
      RECT  87600.0 336150.0 88800.0 334950.0 ;
      RECT  87600.0 346050.0 88800.0 344850.0 ;
      RECT  83400.0 341400.0 84600.0 340200.0 ;
      RECT  83400.0 341400.0 84600.0 340200.0 ;
      RECT  85950.0 341250.0 86850.0 340350.0 ;
      RECT  81000.0 334050.0 90600.0 333150.0 ;
      RECT  81000.0 347850.0 90600.0 346950.0 ;
      RECT  53250.0 340200.0 54450.0 341400.0 ;
      RECT  55200.0 342600.0 56400.0 343800.0 ;
      RECT  72000.0 341700.0 70800.0 342900.0 ;
      RECT  63600.0 359250.0 64800.0 361200.0 ;
      RECT  63600.0 347400.0 64800.0 349350.0 ;
      RECT  58800.0 348750.0 60000.0 346950.0 ;
      RECT  58800.0 358050.0 60000.0 361650.0 ;
      RECT  61500.0 348750.0 62400.0 358050.0 ;
      RECT  58800.0 358050.0 60000.0 359250.0 ;
      RECT  61200.0 358050.0 62400.0 359250.0 ;
      RECT  61200.0 358050.0 62400.0 359250.0 ;
      RECT  58800.0 358050.0 60000.0 359250.0 ;
      RECT  58800.0 348750.0 60000.0 349950.0 ;
      RECT  61200.0 348750.0 62400.0 349950.0 ;
      RECT  61200.0 348750.0 62400.0 349950.0 ;
      RECT  58800.0 348750.0 60000.0 349950.0 ;
      RECT  63600.0 358650.0 64800.0 359850.0 ;
      RECT  63600.0 348750.0 64800.0 349950.0 ;
      RECT  59400.0 353400.0 60600.0 354600.0 ;
      RECT  59400.0 353400.0 60600.0 354600.0 ;
      RECT  61950.0 353550.0 62850.0 354450.0 ;
      RECT  57000.0 360750.0 66600.0 361650.0 ;
      RECT  57000.0 346950.0 66600.0 347850.0 ;
      RECT  68400.0 349350.0 69600.0 346950.0 ;
      RECT  68400.0 358050.0 69600.0 361650.0 ;
      RECT  73200.0 358050.0 74400.0 361650.0 ;
      RECT  75600.0 359250.0 76800.0 361200.0 ;
      RECT  75600.0 347400.0 76800.0 349350.0 ;
      RECT  68400.0 358050.0 69600.0 359250.0 ;
      RECT  70800.0 358050.0 72000.0 359250.0 ;
      RECT  70800.0 358050.0 72000.0 359250.0 ;
      RECT  68400.0 358050.0 69600.0 359250.0 ;
      RECT  70800.0 358050.0 72000.0 359250.0 ;
      RECT  73200.0 358050.0 74400.0 359250.0 ;
      RECT  73200.0 358050.0 74400.0 359250.0 ;
      RECT  70800.0 358050.0 72000.0 359250.0 ;
      RECT  68400.0 349350.0 69600.0 350550.0 ;
      RECT  70800.0 349350.0 72000.0 350550.0 ;
      RECT  70800.0 349350.0 72000.0 350550.0 ;
      RECT  68400.0 349350.0 69600.0 350550.0 ;
      RECT  70800.0 349350.0 72000.0 350550.0 ;
      RECT  73200.0 349350.0 74400.0 350550.0 ;
      RECT  73200.0 349350.0 74400.0 350550.0 ;
      RECT  70800.0 349350.0 72000.0 350550.0 ;
      RECT  75600.0 358650.0 76800.0 359850.0 ;
      RECT  75600.0 348750.0 76800.0 349950.0 ;
      RECT  73200.0 351900.0 72000.0 353100.0 ;
      RECT  70200.0 354600.0 69000.0 355800.0 ;
      RECT  70800.0 358050.0 72000.0 359250.0 ;
      RECT  73200.0 349350.0 74400.0 350550.0 ;
      RECT  74400.0 354600.0 73200.0 355800.0 ;
      RECT  69000.0 354600.0 70200.0 355800.0 ;
      RECT  72000.0 351900.0 73200.0 353100.0 ;
      RECT  73200.0 354600.0 74400.0 355800.0 ;
      RECT  66600.0 360750.0 81000.0 361650.0 ;
      RECT  66600.0 346950.0 81000.0 347850.0 ;
      RECT  87600.0 359250.0 88800.0 361200.0 ;
      RECT  87600.0 347400.0 88800.0 349350.0 ;
      RECT  82800.0 348750.0 84000.0 346950.0 ;
      RECT  82800.0 358050.0 84000.0 361650.0 ;
      RECT  85500.0 348750.0 86400.0 358050.0 ;
      RECT  82800.0 358050.0 84000.0 359250.0 ;
      RECT  85200.0 358050.0 86400.0 359250.0 ;
      RECT  85200.0 358050.0 86400.0 359250.0 ;
      RECT  82800.0 358050.0 84000.0 359250.0 ;
      RECT  82800.0 348750.0 84000.0 349950.0 ;
      RECT  85200.0 348750.0 86400.0 349950.0 ;
      RECT  85200.0 348750.0 86400.0 349950.0 ;
      RECT  82800.0 348750.0 84000.0 349950.0 ;
      RECT  87600.0 358650.0 88800.0 359850.0 ;
      RECT  87600.0 348750.0 88800.0 349950.0 ;
      RECT  83400.0 353400.0 84600.0 354600.0 ;
      RECT  83400.0 353400.0 84600.0 354600.0 ;
      RECT  85950.0 353550.0 86850.0 354450.0 ;
      RECT  81000.0 360750.0 90600.0 361650.0 ;
      RECT  81000.0 346950.0 90600.0 347850.0 ;
      RECT  53250.0 353400.0 54450.0 354600.0 ;
      RECT  55200.0 351000.0 56400.0 352200.0 ;
      RECT  72000.0 351900.0 70800.0 353100.0 ;
      RECT  63600.0 363150.0 64800.0 361200.0 ;
      RECT  63600.0 375000.0 64800.0 373050.0 ;
      RECT  58800.0 373650.0 60000.0 375450.0 ;
      RECT  58800.0 364350.0 60000.0 360750.0 ;
      RECT  61500.0 373650.0 62400.0 364350.0 ;
      RECT  58800.0 364350.0 60000.0 363150.0 ;
      RECT  61200.0 364350.0 62400.0 363150.0 ;
      RECT  61200.0 364350.0 62400.0 363150.0 ;
      RECT  58800.0 364350.0 60000.0 363150.0 ;
      RECT  58800.0 373650.0 60000.0 372450.0 ;
      RECT  61200.0 373650.0 62400.0 372450.0 ;
      RECT  61200.0 373650.0 62400.0 372450.0 ;
      RECT  58800.0 373650.0 60000.0 372450.0 ;
      RECT  63600.0 363750.0 64800.0 362550.0 ;
      RECT  63600.0 373650.0 64800.0 372450.0 ;
      RECT  59400.0 369000.0 60600.0 367800.0 ;
      RECT  59400.0 369000.0 60600.0 367800.0 ;
      RECT  61950.0 368850.0 62850.0 367950.0 ;
      RECT  57000.0 361650.0 66600.0 360750.0 ;
      RECT  57000.0 375450.0 66600.0 374550.0 ;
      RECT  68400.0 373050.0 69600.0 375450.0 ;
      RECT  68400.0 364350.0 69600.0 360750.0 ;
      RECT  73200.0 364350.0 74400.0 360750.0 ;
      RECT  75600.0 363150.0 76800.0 361200.0 ;
      RECT  75600.0 375000.0 76800.0 373050.0 ;
      RECT  68400.0 364350.0 69600.0 363150.0 ;
      RECT  70800.0 364350.0 72000.0 363150.0 ;
      RECT  70800.0 364350.0 72000.0 363150.0 ;
      RECT  68400.0 364350.0 69600.0 363150.0 ;
      RECT  70800.0 364350.0 72000.0 363150.0 ;
      RECT  73200.0 364350.0 74400.0 363150.0 ;
      RECT  73200.0 364350.0 74400.0 363150.0 ;
      RECT  70800.0 364350.0 72000.0 363150.0 ;
      RECT  68400.0 373050.0 69600.0 371850.0 ;
      RECT  70800.0 373050.0 72000.0 371850.0 ;
      RECT  70800.0 373050.0 72000.0 371850.0 ;
      RECT  68400.0 373050.0 69600.0 371850.0 ;
      RECT  70800.0 373050.0 72000.0 371850.0 ;
      RECT  73200.0 373050.0 74400.0 371850.0 ;
      RECT  73200.0 373050.0 74400.0 371850.0 ;
      RECT  70800.0 373050.0 72000.0 371850.0 ;
      RECT  75600.0 363750.0 76800.0 362550.0 ;
      RECT  75600.0 373650.0 76800.0 372450.0 ;
      RECT  73200.0 370500.0 72000.0 369300.0 ;
      RECT  70200.0 367800.0 69000.0 366600.0 ;
      RECT  70800.0 364350.0 72000.0 363150.0 ;
      RECT  73200.0 373050.0 74400.0 371850.0 ;
      RECT  74400.0 367800.0 73200.0 366600.0 ;
      RECT  69000.0 367800.0 70200.0 366600.0 ;
      RECT  72000.0 370500.0 73200.0 369300.0 ;
      RECT  73200.0 367800.0 74400.0 366600.0 ;
      RECT  66600.0 361650.0 81000.0 360750.0 ;
      RECT  66600.0 375450.0 81000.0 374550.0 ;
      RECT  87600.0 363150.0 88800.0 361200.0 ;
      RECT  87600.0 375000.0 88800.0 373050.0 ;
      RECT  82800.0 373650.0 84000.0 375450.0 ;
      RECT  82800.0 364350.0 84000.0 360750.0 ;
      RECT  85500.0 373650.0 86400.0 364350.0 ;
      RECT  82800.0 364350.0 84000.0 363150.0 ;
      RECT  85200.0 364350.0 86400.0 363150.0 ;
      RECT  85200.0 364350.0 86400.0 363150.0 ;
      RECT  82800.0 364350.0 84000.0 363150.0 ;
      RECT  82800.0 373650.0 84000.0 372450.0 ;
      RECT  85200.0 373650.0 86400.0 372450.0 ;
      RECT  85200.0 373650.0 86400.0 372450.0 ;
      RECT  82800.0 373650.0 84000.0 372450.0 ;
      RECT  87600.0 363750.0 88800.0 362550.0 ;
      RECT  87600.0 373650.0 88800.0 372450.0 ;
      RECT  83400.0 369000.0 84600.0 367800.0 ;
      RECT  83400.0 369000.0 84600.0 367800.0 ;
      RECT  85950.0 368850.0 86850.0 367950.0 ;
      RECT  81000.0 361650.0 90600.0 360750.0 ;
      RECT  81000.0 375450.0 90600.0 374550.0 ;
      RECT  53250.0 367800.0 54450.0 369000.0 ;
      RECT  55200.0 370200.0 56400.0 371400.0 ;
      RECT  72000.0 369300.0 70800.0 370500.0 ;
      RECT  63600.0 386850.0 64800.0 388800.0 ;
      RECT  63600.0 375000.0 64800.0 376950.0 ;
      RECT  58800.0 376350.0 60000.0 374550.0 ;
      RECT  58800.0 385650.0 60000.0 389250.0 ;
      RECT  61500.0 376350.0 62400.0 385650.0 ;
      RECT  58800.0 385650.0 60000.0 386850.0 ;
      RECT  61200.0 385650.0 62400.0 386850.0 ;
      RECT  61200.0 385650.0 62400.0 386850.0 ;
      RECT  58800.0 385650.0 60000.0 386850.0 ;
      RECT  58800.0 376350.0 60000.0 377550.0 ;
      RECT  61200.0 376350.0 62400.0 377550.0 ;
      RECT  61200.0 376350.0 62400.0 377550.0 ;
      RECT  58800.0 376350.0 60000.0 377550.0 ;
      RECT  63600.0 386250.0 64800.0 387450.0 ;
      RECT  63600.0 376350.0 64800.0 377550.0 ;
      RECT  59400.0 381000.0 60600.0 382200.0 ;
      RECT  59400.0 381000.0 60600.0 382200.0 ;
      RECT  61950.0 381150.0 62850.0 382050.0 ;
      RECT  57000.0 388350.0 66600.0 389250.0 ;
      RECT  57000.0 374550.0 66600.0 375450.0 ;
      RECT  68400.0 376950.0 69600.0 374550.0 ;
      RECT  68400.0 385650.0 69600.0 389250.0 ;
      RECT  73200.0 385650.0 74400.0 389250.0 ;
      RECT  75600.0 386850.0 76800.0 388800.0 ;
      RECT  75600.0 375000.0 76800.0 376950.0 ;
      RECT  68400.0 385650.0 69600.0 386850.0 ;
      RECT  70800.0 385650.0 72000.0 386850.0 ;
      RECT  70800.0 385650.0 72000.0 386850.0 ;
      RECT  68400.0 385650.0 69600.0 386850.0 ;
      RECT  70800.0 385650.0 72000.0 386850.0 ;
      RECT  73200.0 385650.0 74400.0 386850.0 ;
      RECT  73200.0 385650.0 74400.0 386850.0 ;
      RECT  70800.0 385650.0 72000.0 386850.0 ;
      RECT  68400.0 376950.0 69600.0 378150.0 ;
      RECT  70800.0 376950.0 72000.0 378150.0 ;
      RECT  70800.0 376950.0 72000.0 378150.0 ;
      RECT  68400.0 376950.0 69600.0 378150.0 ;
      RECT  70800.0 376950.0 72000.0 378150.0 ;
      RECT  73200.0 376950.0 74400.0 378150.0 ;
      RECT  73200.0 376950.0 74400.0 378150.0 ;
      RECT  70800.0 376950.0 72000.0 378150.0 ;
      RECT  75600.0 386250.0 76800.0 387450.0 ;
      RECT  75600.0 376350.0 76800.0 377550.0 ;
      RECT  73200.0 379500.0 72000.0 380700.0 ;
      RECT  70200.0 382200.0 69000.0 383400.0 ;
      RECT  70800.0 385650.0 72000.0 386850.0 ;
      RECT  73200.0 376950.0 74400.0 378150.0 ;
      RECT  74400.0 382200.0 73200.0 383400.0 ;
      RECT  69000.0 382200.0 70200.0 383400.0 ;
      RECT  72000.0 379500.0 73200.0 380700.0 ;
      RECT  73200.0 382200.0 74400.0 383400.0 ;
      RECT  66600.0 388350.0 81000.0 389250.0 ;
      RECT  66600.0 374550.0 81000.0 375450.0 ;
      RECT  87600.0 386850.0 88800.0 388800.0 ;
      RECT  87600.0 375000.0 88800.0 376950.0 ;
      RECT  82800.0 376350.0 84000.0 374550.0 ;
      RECT  82800.0 385650.0 84000.0 389250.0 ;
      RECT  85500.0 376350.0 86400.0 385650.0 ;
      RECT  82800.0 385650.0 84000.0 386850.0 ;
      RECT  85200.0 385650.0 86400.0 386850.0 ;
      RECT  85200.0 385650.0 86400.0 386850.0 ;
      RECT  82800.0 385650.0 84000.0 386850.0 ;
      RECT  82800.0 376350.0 84000.0 377550.0 ;
      RECT  85200.0 376350.0 86400.0 377550.0 ;
      RECT  85200.0 376350.0 86400.0 377550.0 ;
      RECT  82800.0 376350.0 84000.0 377550.0 ;
      RECT  87600.0 386250.0 88800.0 387450.0 ;
      RECT  87600.0 376350.0 88800.0 377550.0 ;
      RECT  83400.0 381000.0 84600.0 382200.0 ;
      RECT  83400.0 381000.0 84600.0 382200.0 ;
      RECT  85950.0 381150.0 86850.0 382050.0 ;
      RECT  81000.0 388350.0 90600.0 389250.0 ;
      RECT  81000.0 374550.0 90600.0 375450.0 ;
      RECT  53250.0 381000.0 54450.0 382200.0 ;
      RECT  55200.0 378600.0 56400.0 379800.0 ;
      RECT  72000.0 379500.0 70800.0 380700.0 ;
      RECT  63600.0 390750.0 64800.0 388800.0 ;
      RECT  63600.0 402600.0 64800.0 400650.0 ;
      RECT  58800.0 401250.0 60000.0 403050.0 ;
      RECT  58800.0 391950.0 60000.0 388350.0 ;
      RECT  61500.0 401250.0 62400.0 391950.0 ;
      RECT  58800.0 391950.0 60000.0 390750.0 ;
      RECT  61200.0 391950.0 62400.0 390750.0 ;
      RECT  61200.0 391950.0 62400.0 390750.0 ;
      RECT  58800.0 391950.0 60000.0 390750.0 ;
      RECT  58800.0 401250.0 60000.0 400050.0 ;
      RECT  61200.0 401250.0 62400.0 400050.0 ;
      RECT  61200.0 401250.0 62400.0 400050.0 ;
      RECT  58800.0 401250.0 60000.0 400050.0 ;
      RECT  63600.0 391350.0 64800.0 390150.0 ;
      RECT  63600.0 401250.0 64800.0 400050.0 ;
      RECT  59400.0 396600.0 60600.0 395400.0 ;
      RECT  59400.0 396600.0 60600.0 395400.0 ;
      RECT  61950.0 396450.0 62850.0 395550.0 ;
      RECT  57000.0 389250.0 66600.0 388350.0 ;
      RECT  57000.0 403050.0 66600.0 402150.0 ;
      RECT  68400.0 400650.0 69600.0 403050.0 ;
      RECT  68400.0 391950.0 69600.0 388350.0 ;
      RECT  73200.0 391950.0 74400.0 388350.0 ;
      RECT  75600.0 390750.0 76800.0 388800.0 ;
      RECT  75600.0 402600.0 76800.0 400650.0 ;
      RECT  68400.0 391950.0 69600.0 390750.0 ;
      RECT  70800.0 391950.0 72000.0 390750.0 ;
      RECT  70800.0 391950.0 72000.0 390750.0 ;
      RECT  68400.0 391950.0 69600.0 390750.0 ;
      RECT  70800.0 391950.0 72000.0 390750.0 ;
      RECT  73200.0 391950.0 74400.0 390750.0 ;
      RECT  73200.0 391950.0 74400.0 390750.0 ;
      RECT  70800.0 391950.0 72000.0 390750.0 ;
      RECT  68400.0 400650.0 69600.0 399450.0 ;
      RECT  70800.0 400650.0 72000.0 399450.0 ;
      RECT  70800.0 400650.0 72000.0 399450.0 ;
      RECT  68400.0 400650.0 69600.0 399450.0 ;
      RECT  70800.0 400650.0 72000.0 399450.0 ;
      RECT  73200.0 400650.0 74400.0 399450.0 ;
      RECT  73200.0 400650.0 74400.0 399450.0 ;
      RECT  70800.0 400650.0 72000.0 399450.0 ;
      RECT  75600.0 391350.0 76800.0 390150.0 ;
      RECT  75600.0 401250.0 76800.0 400050.0 ;
      RECT  73200.0 398100.0 72000.0 396900.0 ;
      RECT  70200.0 395400.0 69000.0 394200.0 ;
      RECT  70800.0 391950.0 72000.0 390750.0 ;
      RECT  73200.0 400650.0 74400.0 399450.0 ;
      RECT  74400.0 395400.0 73200.0 394200.0 ;
      RECT  69000.0 395400.0 70200.0 394200.0 ;
      RECT  72000.0 398100.0 73200.0 396900.0 ;
      RECT  73200.0 395400.0 74400.0 394200.0 ;
      RECT  66600.0 389250.0 81000.0 388350.0 ;
      RECT  66600.0 403050.0 81000.0 402150.0 ;
      RECT  87600.0 390750.0 88800.0 388800.0 ;
      RECT  87600.0 402600.0 88800.0 400650.0 ;
      RECT  82800.0 401250.0 84000.0 403050.0 ;
      RECT  82800.0 391950.0 84000.0 388350.0 ;
      RECT  85500.0 401250.0 86400.0 391950.0 ;
      RECT  82800.0 391950.0 84000.0 390750.0 ;
      RECT  85200.0 391950.0 86400.0 390750.0 ;
      RECT  85200.0 391950.0 86400.0 390750.0 ;
      RECT  82800.0 391950.0 84000.0 390750.0 ;
      RECT  82800.0 401250.0 84000.0 400050.0 ;
      RECT  85200.0 401250.0 86400.0 400050.0 ;
      RECT  85200.0 401250.0 86400.0 400050.0 ;
      RECT  82800.0 401250.0 84000.0 400050.0 ;
      RECT  87600.0 391350.0 88800.0 390150.0 ;
      RECT  87600.0 401250.0 88800.0 400050.0 ;
      RECT  83400.0 396600.0 84600.0 395400.0 ;
      RECT  83400.0 396600.0 84600.0 395400.0 ;
      RECT  85950.0 396450.0 86850.0 395550.0 ;
      RECT  81000.0 389250.0 90600.0 388350.0 ;
      RECT  81000.0 403050.0 90600.0 402150.0 ;
      RECT  53250.0 395400.0 54450.0 396600.0 ;
      RECT  55200.0 397800.0 56400.0 399000.0 ;
      RECT  72000.0 396900.0 70800.0 398100.0 ;
      RECT  63600.0 414450.0 64800.0 416400.0 ;
      RECT  63600.0 402600.0 64800.0 404550.0 ;
      RECT  58800.0 403950.0 60000.0 402150.0 ;
      RECT  58800.0 413250.0 60000.0 416850.0 ;
      RECT  61500.0 403950.0 62400.0 413250.0 ;
      RECT  58800.0 413250.0 60000.0 414450.0 ;
      RECT  61200.0 413250.0 62400.0 414450.0 ;
      RECT  61200.0 413250.0 62400.0 414450.0 ;
      RECT  58800.0 413250.0 60000.0 414450.0 ;
      RECT  58800.0 403950.0 60000.0 405150.0 ;
      RECT  61200.0 403950.0 62400.0 405150.0 ;
      RECT  61200.0 403950.0 62400.0 405150.0 ;
      RECT  58800.0 403950.0 60000.0 405150.0 ;
      RECT  63600.0 413850.0 64800.0 415050.0 ;
      RECT  63600.0 403950.0 64800.0 405150.0 ;
      RECT  59400.0 408600.0 60600.0 409800.0 ;
      RECT  59400.0 408600.0 60600.0 409800.0 ;
      RECT  61950.0 408750.0 62850.0 409650.0 ;
      RECT  57000.0 415950.0 66600.0 416850.0 ;
      RECT  57000.0 402150.0 66600.0 403050.0 ;
      RECT  68400.0 404550.0 69600.0 402150.0 ;
      RECT  68400.0 413250.0 69600.0 416850.0 ;
      RECT  73200.0 413250.0 74400.0 416850.0 ;
      RECT  75600.0 414450.0 76800.0 416400.0 ;
      RECT  75600.0 402600.0 76800.0 404550.0 ;
      RECT  68400.0 413250.0 69600.0 414450.0 ;
      RECT  70800.0 413250.0 72000.0 414450.0 ;
      RECT  70800.0 413250.0 72000.0 414450.0 ;
      RECT  68400.0 413250.0 69600.0 414450.0 ;
      RECT  70800.0 413250.0 72000.0 414450.0 ;
      RECT  73200.0 413250.0 74400.0 414450.0 ;
      RECT  73200.0 413250.0 74400.0 414450.0 ;
      RECT  70800.0 413250.0 72000.0 414450.0 ;
      RECT  68400.0 404550.0 69600.0 405750.0 ;
      RECT  70800.0 404550.0 72000.0 405750.0 ;
      RECT  70800.0 404550.0 72000.0 405750.0 ;
      RECT  68400.0 404550.0 69600.0 405750.0 ;
      RECT  70800.0 404550.0 72000.0 405750.0 ;
      RECT  73200.0 404550.0 74400.0 405750.0 ;
      RECT  73200.0 404550.0 74400.0 405750.0 ;
      RECT  70800.0 404550.0 72000.0 405750.0 ;
      RECT  75600.0 413850.0 76800.0 415050.0 ;
      RECT  75600.0 403950.0 76800.0 405150.0 ;
      RECT  73200.0 407100.0 72000.0 408300.0 ;
      RECT  70200.0 409800.0 69000.0 411000.0 ;
      RECT  70800.0 413250.0 72000.0 414450.0 ;
      RECT  73200.0 404550.0 74400.0 405750.0 ;
      RECT  74400.0 409800.0 73200.0 411000.0 ;
      RECT  69000.0 409800.0 70200.0 411000.0 ;
      RECT  72000.0 407100.0 73200.0 408300.0 ;
      RECT  73200.0 409800.0 74400.0 411000.0 ;
      RECT  66600.0 415950.0 81000.0 416850.0 ;
      RECT  66600.0 402150.0 81000.0 403050.0 ;
      RECT  87600.0 414450.0 88800.0 416400.0 ;
      RECT  87600.0 402600.0 88800.0 404550.0 ;
      RECT  82800.0 403950.0 84000.0 402150.0 ;
      RECT  82800.0 413250.0 84000.0 416850.0 ;
      RECT  85500.0 403950.0 86400.0 413250.0 ;
      RECT  82800.0 413250.0 84000.0 414450.0 ;
      RECT  85200.0 413250.0 86400.0 414450.0 ;
      RECT  85200.0 413250.0 86400.0 414450.0 ;
      RECT  82800.0 413250.0 84000.0 414450.0 ;
      RECT  82800.0 403950.0 84000.0 405150.0 ;
      RECT  85200.0 403950.0 86400.0 405150.0 ;
      RECT  85200.0 403950.0 86400.0 405150.0 ;
      RECT  82800.0 403950.0 84000.0 405150.0 ;
      RECT  87600.0 413850.0 88800.0 415050.0 ;
      RECT  87600.0 403950.0 88800.0 405150.0 ;
      RECT  83400.0 408600.0 84600.0 409800.0 ;
      RECT  83400.0 408600.0 84600.0 409800.0 ;
      RECT  85950.0 408750.0 86850.0 409650.0 ;
      RECT  81000.0 415950.0 90600.0 416850.0 ;
      RECT  81000.0 402150.0 90600.0 403050.0 ;
      RECT  53250.0 408600.0 54450.0 409800.0 ;
      RECT  55200.0 406200.0 56400.0 407400.0 ;
      RECT  72000.0 407100.0 70800.0 408300.0 ;
      RECT  63600.0 418350.0 64800.0 416400.0 ;
      RECT  63600.0 430200.0 64800.0 428250.0 ;
      RECT  58800.0 428850.0 60000.0 430650.0 ;
      RECT  58800.0 419550.0 60000.0 415950.0 ;
      RECT  61500.0 428850.0 62400.0 419550.0 ;
      RECT  58800.0 419550.0 60000.0 418350.0 ;
      RECT  61200.0 419550.0 62400.0 418350.0 ;
      RECT  61200.0 419550.0 62400.0 418350.0 ;
      RECT  58800.0 419550.0 60000.0 418350.0 ;
      RECT  58800.0 428850.0 60000.0 427650.0 ;
      RECT  61200.0 428850.0 62400.0 427650.0 ;
      RECT  61200.0 428850.0 62400.0 427650.0 ;
      RECT  58800.0 428850.0 60000.0 427650.0 ;
      RECT  63600.0 418950.0 64800.0 417750.0 ;
      RECT  63600.0 428850.0 64800.0 427650.0 ;
      RECT  59400.0 424200.0 60600.0 423000.0 ;
      RECT  59400.0 424200.0 60600.0 423000.0 ;
      RECT  61950.0 424050.0 62850.0 423150.0 ;
      RECT  57000.0 416850.0 66600.0 415950.0 ;
      RECT  57000.0 430650.0 66600.0 429750.0 ;
      RECT  68400.0 428250.0 69600.0 430650.0 ;
      RECT  68400.0 419550.0 69600.0 415950.0 ;
      RECT  73200.0 419550.0 74400.0 415950.0 ;
      RECT  75600.0 418350.0 76800.0 416400.0 ;
      RECT  75600.0 430200.0 76800.0 428250.0 ;
      RECT  68400.0 419550.0 69600.0 418350.0 ;
      RECT  70800.0 419550.0 72000.0 418350.0 ;
      RECT  70800.0 419550.0 72000.0 418350.0 ;
      RECT  68400.0 419550.0 69600.0 418350.0 ;
      RECT  70800.0 419550.0 72000.0 418350.0 ;
      RECT  73200.0 419550.0 74400.0 418350.0 ;
      RECT  73200.0 419550.0 74400.0 418350.0 ;
      RECT  70800.0 419550.0 72000.0 418350.0 ;
      RECT  68400.0 428250.0 69600.0 427050.0 ;
      RECT  70800.0 428250.0 72000.0 427050.0 ;
      RECT  70800.0 428250.0 72000.0 427050.0 ;
      RECT  68400.0 428250.0 69600.0 427050.0 ;
      RECT  70800.0 428250.0 72000.0 427050.0 ;
      RECT  73200.0 428250.0 74400.0 427050.0 ;
      RECT  73200.0 428250.0 74400.0 427050.0 ;
      RECT  70800.0 428250.0 72000.0 427050.0 ;
      RECT  75600.0 418950.0 76800.0 417750.0 ;
      RECT  75600.0 428850.0 76800.0 427650.0 ;
      RECT  73200.0 425700.0 72000.0 424500.0 ;
      RECT  70200.0 423000.0 69000.0 421800.0 ;
      RECT  70800.0 419550.0 72000.0 418350.0 ;
      RECT  73200.0 428250.0 74400.0 427050.0 ;
      RECT  74400.0 423000.0 73200.0 421800.0 ;
      RECT  69000.0 423000.0 70200.0 421800.0 ;
      RECT  72000.0 425700.0 73200.0 424500.0 ;
      RECT  73200.0 423000.0 74400.0 421800.0 ;
      RECT  66600.0 416850.0 81000.0 415950.0 ;
      RECT  66600.0 430650.0 81000.0 429750.0 ;
      RECT  87600.0 418350.0 88800.0 416400.0 ;
      RECT  87600.0 430200.0 88800.0 428250.0 ;
      RECT  82800.0 428850.0 84000.0 430650.0 ;
      RECT  82800.0 419550.0 84000.0 415950.0 ;
      RECT  85500.0 428850.0 86400.0 419550.0 ;
      RECT  82800.0 419550.0 84000.0 418350.0 ;
      RECT  85200.0 419550.0 86400.0 418350.0 ;
      RECT  85200.0 419550.0 86400.0 418350.0 ;
      RECT  82800.0 419550.0 84000.0 418350.0 ;
      RECT  82800.0 428850.0 84000.0 427650.0 ;
      RECT  85200.0 428850.0 86400.0 427650.0 ;
      RECT  85200.0 428850.0 86400.0 427650.0 ;
      RECT  82800.0 428850.0 84000.0 427650.0 ;
      RECT  87600.0 418950.0 88800.0 417750.0 ;
      RECT  87600.0 428850.0 88800.0 427650.0 ;
      RECT  83400.0 424200.0 84600.0 423000.0 ;
      RECT  83400.0 424200.0 84600.0 423000.0 ;
      RECT  85950.0 424050.0 86850.0 423150.0 ;
      RECT  81000.0 416850.0 90600.0 415950.0 ;
      RECT  81000.0 430650.0 90600.0 429750.0 ;
      RECT  53250.0 423000.0 54450.0 424200.0 ;
      RECT  55200.0 425400.0 56400.0 426600.0 ;
      RECT  72000.0 424500.0 70800.0 425700.0 ;
      RECT  50700.0 213150.0 55800.0 214050.0 ;
      RECT  50700.0 232350.0 55800.0 233250.0 ;
      RECT  50700.0 240750.0 55800.0 241650.0 ;
      RECT  50700.0 259950.0 55800.0 260850.0 ;
      RECT  50700.0 268350.0 55800.0 269250.0 ;
      RECT  50700.0 287550.0 55800.0 288450.0 ;
      RECT  50700.0 295950.0 55800.0 296850.0 ;
      RECT  50700.0 315150.0 55800.0 316050.0 ;
      RECT  50700.0 323550.0 55800.0 324450.0 ;
      RECT  50700.0 342750.0 55800.0 343650.0 ;
      RECT  50700.0 351150.0 55800.0 352050.0 ;
      RECT  50700.0 370350.0 55800.0 371250.0 ;
      RECT  50700.0 378750.0 55800.0 379650.0 ;
      RECT  50700.0 397950.0 55800.0 398850.0 ;
      RECT  50700.0 406350.0 55800.0 407250.0 ;
      RECT  50700.0 425550.0 55800.0 426450.0 ;
      RECT  85950.0 215550.0 86850.0 216450.0 ;
      RECT  85950.0 229950.0 86850.0 230850.0 ;
      RECT  85950.0 243150.0 86850.0 244050.0 ;
      RECT  85950.0 257550.0 86850.0 258450.0 ;
      RECT  85950.0 270750.0 86850.0 271650.0 ;
      RECT  85950.0 285150.0 86850.0 286050.0 ;
      RECT  85950.0 298350.0 86850.0 299250.0 ;
      RECT  85950.0 312750.0 86850.0 313650.0 ;
      RECT  85950.0 325950.0 86850.0 326850.0 ;
      RECT  85950.0 340350.0 86850.0 341250.0 ;
      RECT  85950.0 353550.0 86850.0 354450.0 ;
      RECT  85950.0 367950.0 86850.0 368850.0 ;
      RECT  85950.0 381150.0 86850.0 382050.0 ;
      RECT  85950.0 395550.0 86850.0 396450.0 ;
      RECT  85950.0 408750.0 86850.0 409650.0 ;
      RECT  85950.0 423150.0 86850.0 424050.0 ;
      RECT  50700.0 222750.0 57000.0 223650.0 ;
      RECT  50700.0 250350.0 57000.0 251250.0 ;
      RECT  50700.0 277950.0 57000.0 278850.0 ;
      RECT  50700.0 305550.0 57000.0 306450.0 ;
      RECT  50700.0 333150.0 57000.0 334050.0 ;
      RECT  50700.0 360750.0 57000.0 361650.0 ;
      RECT  50700.0 388350.0 57000.0 389250.0 ;
      RECT  50700.0 415950.0 57000.0 416850.0 ;
      RECT  50700.0 208950.0 57000.0 209850.0 ;
      RECT  50700.0 236550.0 57000.0 237450.0 ;
      RECT  50700.0 264150.0 57000.0 265050.0 ;
      RECT  50700.0 291750.0 57000.0 292650.0 ;
      RECT  50700.0 319350.0 57000.0 320250.0 ;
      RECT  50700.0 346950.0 57000.0 347850.0 ;
      RECT  50700.0 374550.0 57000.0 375450.0 ;
      RECT  50700.0 402150.0 57000.0 403050.0 ;
      RECT  50700.0 429750.0 57000.0 430650.0 ;
      RECT  9900.0 93600.0 69900.0 83400.0 ;
      RECT  9900.0 73200.0 69900.0 83400.0 ;
      RECT  9900.0 73200.0 69900.0 63000.0 ;
      RECT  9900.0 52800.0 69900.0 63000.0 ;
      RECT  12300.0 93600.0 13200.0 52800.0 ;
      RECT  66300.0 93600.0 67200.0 52800.0 ;
      RECT  0.0 0.0 3600.0 3600.0 ;
      RECT  0.0 453300.0 3600.0 456900.0 ;
      RECT  139500.0 0.0 143100.0 3600.0 ;
      RECT  139500.0 453300.0 143100.0 456900.0 ;
      RECT  4950.0 4950.0 8550.0 8550.0 ;
      RECT  4950.0 458250.0 8550.0 461850.0 ;
      RECT  144450.0 4950.0 148050.0 8550.0 ;
      RECT  144450.0 458250.0 148050.0 461850.0 ;
      RECT  81300.0 101250.0 80100.0 102450.0 ;
      RECT  86400.0 101100.0 85200.0 102300.0 ;
      RECT  78300.0 115050.0 77100.0 116250.0 ;
      RECT  89100.0 114900.0 87900.0 116100.0 ;
      RECT  81300.0 156450.0 80100.0 157650.0 ;
      RECT  91800.0 156300.0 90600.0 157500.0 ;
      RECT  78300.0 170250.0 77100.0 171450.0 ;
      RECT  94500.0 170100.0 93300.0 171300.0 ;
      RECT  3600.0 98400.0 -5.3290705182e-12 99600.0 ;
      RECT  3600.0 126000.0 -5.3290705182e-12 127200.0 ;
      RECT  3600.0 153600.0 -5.3290705182e-12 154800.0 ;
      RECT  3600.0 181200.0 -5.3290705182e-12 182400.0 ;
      RECT  8550.0 112200.0 4950.0 113400.0 ;
      RECT  8550.0 139800.0 4950.0 141000.0 ;
      RECT  8550.0 167400.0 4950.0 168600.0 ;
      RECT  8550.0 195000.0 4950.0 196200.0 ;
      RECT  69300.0 87150.0 68100.0 88350.0 ;
      RECT  86400.0 87150.0 85200.0 88350.0 ;
      RECT  69300.0 78450.0 68100.0 79650.0 ;
      RECT  89100.0 78450.0 87900.0 79650.0 ;
      RECT  69300.0 66750.0 68100.0 67950.0 ;
      RECT  91800.0 66750.0 90600.0 67950.0 ;
      RECT  69300.0 58050.0 68100.0 59250.0 ;
      RECT  94500.0 58050.0 93300.0 59250.0 ;
      RECT  11100.0 82800.0 9900.0 84000.0 ;
      RECT  3600.0 82800.0 -5.3290705182e-12 84000.0 ;
      RECT  11100.0 62400.0 9900.0 63600.0 ;
      RECT  3600.0 62400.0 -5.3290705182e-12 63600.0 ;
      RECT  8550.0 50100.0 4950.0 51300.0 ;
      RECT  105300.0 42150.0 104100.0 43350.0 ;
      RECT  99900.0 37650.0 98700.0 38850.0 ;
      RECT  102600.0 35250.0 101400.0 36450.0 ;
      RECT  105300.0 438450.0 104100.0 439650.0 ;
      RECT  108000.0 106950.0 106800.0 108150.0 ;
      RECT  110700.0 205050.0 109500.0 206250.0 ;
      RECT  97200.0 95100.0 96000.0 96300.0 ;
      RECT  54450.0 431700.0 53250.0 432900.0 ;
      RECT  97200.0 431700.0 96000.0 432900.0 ;
      RECT  148050.0 449550.0 144450.0 450750.0 ;
      RECT  148050.0 177750.0 144450.0 178950.0 ;
      RECT  148050.0 109050.0 144450.0 110250.0 ;
      RECT  148050.0 96150.0 144450.0 97350.0 ;
      RECT  148050.0 19350.0 144450.0 20550.0 ;
      RECT  8550.0 222600.0 4950.0 223800.0 ;
      RECT  148050.0 222600.0 144450.0 223800.0 ;
      RECT  8550.0 250200.0 4950.0 251400.0 ;
      RECT  148050.0 250200.0 144450.0 251400.0 ;
      RECT  8550.0 277800.0 4950.0 279000.0 ;
      RECT  148050.0 277800.0 144450.0 279000.0 ;
      RECT  8550.0 305400.0 4950.0 306600.0 ;
      RECT  148050.0 305400.0 144450.0 306600.0 ;
      RECT  8550.0 333000.0 4950.0 334200.0 ;
      RECT  148050.0 333000.0 144450.0 334200.0 ;
      RECT  8550.0 360600.0 4950.0 361800.0 ;
      RECT  148050.0 360600.0 144450.0 361800.0 ;
      RECT  8550.0 388200.0 4950.0 389400.0 ;
      RECT  148050.0 388200.0 144450.0 389400.0 ;
      RECT  8550.0 415800.0 4950.0 417000.0 ;
      RECT  148050.0 415800.0 144450.0 417000.0 ;
      RECT  143100.0 33150.0 139500.0 34350.0 ;
      RECT  143100.0 202950.0 139500.0 204150.0 ;
      RECT  143100.0 104850.0 139500.0 106050.0 ;
      RECT  3600.0 208800.0 -5.3290705182e-12 210000.0 ;
      RECT  3600.0 236400.0 -5.3290705182e-12 237600.0 ;
      RECT  3600.0 264000.0 -5.3290705182e-12 265200.0 ;
      RECT  3600.0 291600.0 -5.3290705182e-12 292800.0 ;
      RECT  3600.0 319200.0 -5.3290705182e-12 320400.0 ;
      RECT  3600.0 346800.0 -5.3290705182e-12 348000.0 ;
      RECT  3600.0 374400.0 -5.3290705182e-12 375600.0 ;
      RECT  3600.0 402000.0 -5.3290705182e-12 403200.0 ;
      RECT  3600.0 429600.0 -5.3290705182e-12 430800.0 ;
      RECT  0.0 4950.0 148050.0 8550.0 ;
      RECT  0.0 458250.0 148050.0 461850.0 ;
      RECT  0.0 0.0 148050.0 3600.0 ;
      RECT  0.0 453300.0 148050.0 456900.0 ;
      RECT  -9150.0 187200.0 -10050.0 196800.0 ;
      RECT  -9000.0 203400.0 -9900.0 204300.0 ;
      RECT  -9450.0 203400.0 -9600.0 204300.0 ;
      RECT  -9000.0 203850.0 -9900.0 211200.0 ;
      RECT  -9000.0 223050.0 -9900.0 230400.0 ;
      RECT  -17250.0 238200.0 -22200.0 239100.0 ;
      RECT  -9150.0 186750.0 -10050.0 187650.0 ;
      RECT  -9150.0 203400.0 -10050.0 204300.0 ;
      RECT  -23550.0 341700.0 -24450.0 355050.0 ;
      RECT  -9000.0 252300.0 -9900.0 264450.0 ;
      RECT  -19500.0 184200.0 -22200.0 185100.0 ;
      RECT  -23100.0 264450.0 -24000.0 291300.0 ;
      RECT  -25800.0 269850.0 -26700.0 294300.0 ;
      RECT  -11100.0 283350.0 -12000.0 291900.0 ;
      RECT  -9150.0 280650.0 -10050.0 294300.0 ;
      RECT  -7200.0 272550.0 -8100.0 296700.0 ;
      RECT  -11100.0 306450.0 -12000.0 307350.0 ;
      RECT  -11100.0 297900.0 -12000.0 306900.0 ;
      RECT  -9600.0 306450.0 -11550.0 307350.0 ;
      RECT  -9000.0 308850.0 -9900.0 309750.0 ;
      RECT  -9450.0 308850.0 -9600.0 309750.0 ;
      RECT  -9000.0 309300.0 -9900.0 366900.0 ;
      RECT  -38700.0 283350.0 -39600.0 301500.0 ;
      RECT  -36750.0 272550.0 -37650.0 303900.0 ;
      RECT  -34800.0 275250.0 -35700.0 306300.0 ;
      RECT  -38700.0 316050.0 -39600.0 316950.0 ;
      RECT  -38700.0 307500.0 -39600.0 316500.0 ;
      RECT  -37200.0 316050.0 -39150.0 316950.0 ;
      RECT  -36750.0 318900.0 -37650.0 326100.0 ;
      RECT  -36750.0 328500.0 -37650.0 335700.0 ;
      RECT  -23550.0 341250.0 -24450.0 342150.0 ;
      RECT  -24000.0 341250.0 -24450.0 342150.0 ;
      RECT  -23550.0 339300.0 -24450.0 341700.0 ;
      RECT  -23550.0 329100.0 -24450.0 336300.0 ;
      RECT  -23100.0 296400.0 -24000.0 302700.0 ;
      RECT  -22350.0 312600.0 -23250.0 319800.0 ;
      RECT  -36750.0 338100.0 -37650.0 342300.0 ;
      RECT  -23550.0 322500.0 -24450.0 326700.0 ;
      RECT  -2550.0 181800.0 -3450.0 341700.0 ;
      RECT  -2550.0 267150.0 -3450.0 288300.0 ;
      RECT  -16350.0 181800.0 -17250.0 341700.0 ;
      RECT  -16350.0 277950.0 -17250.0 288300.0 ;
      RECT  -30150.0 288300.0 -31050.0 341700.0 ;
      RECT  -30150.0 267150.0 -31050.0 288300.0 ;
      RECT  -43950.0 288300.0 -44850.0 341700.0 ;
      RECT  -43950.0 277950.0 -44850.0 288300.0 ;
      RECT  -43950.0 341250.0 -44850.0 342150.0 ;
      RECT  -43950.0 339600.0 -44850.0 341700.0 ;
      RECT  -44400.0 341250.0 -49200.0 342150.0 ;
      RECT  -52800.0 181800.0 -42600.0 241800.0 ;
      RECT  -32400.0 181800.0 -42600.0 241800.0 ;
      RECT  -32400.0 181800.0 -22200.0 241800.0 ;
      RECT  -52800.0 184200.0 -22200.0 185100.0 ;
      RECT  -52800.0 238200.0 -22200.0 239100.0 ;
      RECT  -14850.0 190800.0 -16800.0 192000.0 ;
      RECT  -3000.0 190800.0 -4950.0 192000.0 ;
      RECT  -4350.0 186300.0 -13650.0 187200.0 ;
      RECT  -14250.0 183750.0 -16200.0 184650.0 ;
      RECT  -14250.0 188550.0 -16200.0 189450.0 ;
      RECT  -13650.0 183600.0 -14850.0 184800.0 ;
      RECT  -13650.0 188400.0 -14850.0 189600.0 ;
      RECT  -13650.0 186000.0 -14850.0 187200.0 ;
      RECT  -13650.0 186000.0 -14850.0 187200.0 ;
      RECT  -15750.0 183750.0 -16650.0 189450.0 ;
      RECT  -3000.0 183750.0 -4950.0 184650.0 ;
      RECT  -3000.0 188550.0 -4950.0 189450.0 ;
      RECT  -4350.0 183600.0 -5550.0 184800.0 ;
      RECT  -4350.0 188400.0 -5550.0 189600.0 ;
      RECT  -4350.0 186000.0 -5550.0 187200.0 ;
      RECT  -4350.0 186000.0 -5550.0 187200.0 ;
      RECT  -2550.0 183750.0 -3450.0 189450.0 ;
      RECT  -14250.0 190800.0 -15450.0 192000.0 ;
      RECT  -4350.0 190800.0 -5550.0 192000.0 ;
      RECT  -9000.0 184200.0 -10200.0 185400.0 ;
      RECT  -9000.0 184200.0 -10200.0 185400.0 ;
      RECT  -9150.0 186750.0 -10050.0 187650.0 ;
      RECT  -16350.0 181800.0 -17250.0 193800.0 ;
      RECT  -2550.0 181800.0 -3450.0 193800.0 ;
      RECT  -14850.0 205200.0 -16800.0 206400.0 ;
      RECT  -3000.0 205200.0 -4950.0 206400.0 ;
      RECT  -15450.0 195750.0 -17250.0 201450.0 ;
      RECT  -6750.0 202950.0 -11550.0 203850.0 ;
      RECT  -13950.0 195750.0 -15900.0 196650.0 ;
      RECT  -13950.0 200550.0 -15900.0 201450.0 ;
      RECT  -12000.0 198150.0 -13950.0 199050.0 ;
      RECT  -12000.0 202950.0 -13950.0 203850.0 ;
      RECT  -13350.0 195600.0 -14550.0 196800.0 ;
      RECT  -13350.0 200400.0 -14550.0 201600.0 ;
      RECT  -13350.0 198000.0 -14550.0 199200.0 ;
      RECT  -13350.0 202800.0 -14550.0 204000.0 ;
      RECT  -11550.0 198150.0 -12450.0 203850.0 ;
      RECT  -15450.0 195750.0 -16350.0 201450.0 ;
      RECT  -3300.0 195750.0 -5250.0 196650.0 ;
      RECT  -3300.0 200550.0 -5250.0 201450.0 ;
      RECT  -5250.0 198150.0 -7200.0 199050.0 ;
      RECT  -5250.0 202950.0 -7200.0 203850.0 ;
      RECT  -4650.0 195600.0 -5850.0 196800.0 ;
      RECT  -4650.0 200400.0 -5850.0 201600.0 ;
      RECT  -4650.0 198000.0 -5850.0 199200.0 ;
      RECT  -4650.0 202800.0 -5850.0 204000.0 ;
      RECT  -6750.0 198150.0 -7650.0 203850.0 ;
      RECT  -2850.0 195750.0 -3750.0 201450.0 ;
      RECT  -14250.0 205200.0 -15450.0 206400.0 ;
      RECT  -4350.0 205200.0 -5550.0 206400.0 ;
      RECT  -9000.0 196200.0 -10200.0 197400.0 ;
      RECT  -9000.0 196200.0 -10200.0 197400.0 ;
      RECT  -9150.0 203400.0 -10050.0 204300.0 ;
      RECT  -16350.0 193800.0 -17250.0 208200.0 ;
      RECT  -2550.0 193800.0 -3450.0 208200.0 ;
      RECT  -14850.0 224400.0 -16800.0 225600.0 ;
      RECT  -3000.0 224400.0 -4950.0 225600.0 ;
      RECT  -15000.0 210150.0 -17250.0 220650.0 ;
      RECT  -6900.0 222150.0 -11100.0 223050.0 ;
      RECT  -13500.0 210150.0 -15450.0 211050.0 ;
      RECT  -13500.0 214950.0 -15450.0 215850.0 ;
      RECT  -13500.0 219750.0 -15450.0 220650.0 ;
      RECT  -11550.0 212550.0 -13500.0 213450.0 ;
      RECT  -11550.0 217350.0 -13500.0 218250.0 ;
      RECT  -11550.0 222150.0 -13500.0 223050.0 ;
      RECT  -12900.0 210000.0 -14100.0 211200.0 ;
      RECT  -12900.0 214800.0 -14100.0 216000.0 ;
      RECT  -12900.0 219600.0 -14100.0 220800.0 ;
      RECT  -12900.0 212400.0 -14100.0 213600.0 ;
      RECT  -12900.0 217200.0 -14100.0 218400.0 ;
      RECT  -12900.0 222000.0 -14100.0 223200.0 ;
      RECT  -11100.0 212550.0 -12000.0 223050.0 ;
      RECT  -15000.0 210150.0 -15900.0 220650.0 ;
      RECT  -3450.0 210150.0 -5400.0 211050.0 ;
      RECT  -3450.0 214950.0 -5400.0 215850.0 ;
      RECT  -3450.0 219750.0 -5400.0 220650.0 ;
      RECT  -5400.0 212550.0 -7350.0 213450.0 ;
      RECT  -5400.0 217350.0 -7350.0 218250.0 ;
      RECT  -5400.0 222150.0 -7350.0 223050.0 ;
      RECT  -4800.0 210000.0 -6000.0 211200.0 ;
      RECT  -4800.0 214800.0 -6000.0 216000.0 ;
      RECT  -4800.0 219600.0 -6000.0 220800.0 ;
      RECT  -4800.0 212400.0 -6000.0 213600.0 ;
      RECT  -4800.0 217200.0 -6000.0 218400.0 ;
      RECT  -4800.0 222000.0 -6000.0 223200.0 ;
      RECT  -6900.0 212550.0 -7800.0 223050.0 ;
      RECT  -3000.0 210150.0 -3900.0 220650.0 ;
      RECT  -14250.0 224400.0 -15450.0 225600.0 ;
      RECT  -4350.0 224400.0 -5550.0 225600.0 ;
      RECT  -8850.0 210600.0 -10050.0 211800.0 ;
      RECT  -8850.0 210600.0 -10050.0 211800.0 ;
      RECT  -9000.0 222600.0 -9900.0 223500.0 ;
      RECT  -16350.0 208200.0 -17250.0 227400.0 ;
      RECT  -2550.0 208200.0 -3450.0 227400.0 ;
      RECT  -14850.0 255600.0 -16800.0 256800.0 ;
      RECT  -3000.0 255600.0 -4950.0 256800.0 ;
      RECT  -15000.0 229350.0 -17250.0 254250.0 ;
      RECT  -6900.0 250950.0 -11100.0 251850.0 ;
      RECT  -13500.0 229350.0 -15450.0 230250.0 ;
      RECT  -13500.0 234150.0 -15450.0 235050.0 ;
      RECT  -13500.0 238950.0 -15450.0 239850.0 ;
      RECT  -13500.0 243750.0 -15450.0 244650.0 ;
      RECT  -13500.0 248550.0 -15450.0 249450.0 ;
      RECT  -13500.0 253350.0 -15450.0 254250.0 ;
      RECT  -11550.0 231750.0 -13500.0 232650.0 ;
      RECT  -11550.0 236550.0 -13500.0 237450.0 ;
      RECT  -11550.0 241350.0 -13500.0 242250.0 ;
      RECT  -11550.0 246150.0 -13500.0 247050.0 ;
      RECT  -11550.0 250950.0 -13500.0 251850.0 ;
      RECT  -12900.0 229200.0 -14100.0 230400.0 ;
      RECT  -12900.0 234000.0 -14100.0 235200.0 ;
      RECT  -12900.0 238800.0 -14100.0 240000.0 ;
      RECT  -12900.0 243600.0 -14100.0 244800.0 ;
      RECT  -12900.0 248400.0 -14100.0 249600.0 ;
      RECT  -12900.0 253200.0 -14100.0 254400.0 ;
      RECT  -12900.0 231600.0 -14100.0 232800.0 ;
      RECT  -12900.0 236400.0 -14100.0 237600.0 ;
      RECT  -12900.0 241200.0 -14100.0 242400.0 ;
      RECT  -12900.0 246000.0 -14100.0 247200.0 ;
      RECT  -12900.0 250800.0 -14100.0 252000.0 ;
      RECT  -11100.0 231750.0 -12000.0 251850.0 ;
      RECT  -15000.0 229350.0 -15900.0 254250.0 ;
      RECT  -3450.0 229350.0 -5400.0 230250.0 ;
      RECT  -3450.0 234150.0 -5400.0 235050.0 ;
      RECT  -3450.0 238950.0 -5400.0 239850.0 ;
      RECT  -3450.0 243750.0 -5400.0 244650.0 ;
      RECT  -3450.0 248550.0 -5400.0 249450.0 ;
      RECT  -3450.0 253350.0 -5400.0 254250.0 ;
      RECT  -5400.0 231750.0 -7350.0 232650.0 ;
      RECT  -5400.0 236550.0 -7350.0 237450.0 ;
      RECT  -5400.0 241350.0 -7350.0 242250.0 ;
      RECT  -5400.0 246150.0 -7350.0 247050.0 ;
      RECT  -5400.0 250950.0 -7350.0 251850.0 ;
      RECT  -4800.0 229200.0 -6000.0 230400.0 ;
      RECT  -4800.0 234000.0 -6000.0 235200.0 ;
      RECT  -4800.0 238800.0 -6000.0 240000.0 ;
      RECT  -4800.0 243600.0 -6000.0 244800.0 ;
      RECT  -4800.0 248400.0 -6000.0 249600.0 ;
      RECT  -4800.0 253200.0 -6000.0 254400.0 ;
      RECT  -4800.0 231600.0 -6000.0 232800.0 ;
      RECT  -4800.0 236400.0 -6000.0 237600.0 ;
      RECT  -4800.0 241200.0 -6000.0 242400.0 ;
      RECT  -4800.0 246000.0 -6000.0 247200.0 ;
      RECT  -4800.0 250800.0 -6000.0 252000.0 ;
      RECT  -6900.0 231750.0 -7800.0 251850.0 ;
      RECT  -3000.0 229350.0 -3900.0 254250.0 ;
      RECT  -14250.0 255600.0 -15450.0 256800.0 ;
      RECT  -4350.0 255600.0 -5550.0 256800.0 ;
      RECT  -8850.0 229800.0 -10050.0 231000.0 ;
      RECT  -8850.0 229800.0 -10050.0 231000.0 ;
      RECT  -9000.0 251400.0 -9900.0 252300.0 ;
      RECT  -16350.0 227400.0 -17250.0 258600.0 ;
      RECT  -2550.0 227400.0 -3450.0 258600.0 ;
      RECT  -4950.0 290100.0 -2550.0 291300.0 ;
      RECT  -13650.0 290100.0 -17250.0 291300.0 ;
      RECT  -13650.0 294900.0 -17250.0 296100.0 ;
      RECT  -14850.0 299700.0 -16800.0 300900.0 ;
      RECT  -3000.0 299700.0 -4950.0 300900.0 ;
      RECT  -13650.0 290100.0 -14850.0 291300.0 ;
      RECT  -13650.0 292500.0 -14850.0 293700.0 ;
      RECT  -13650.0 292500.0 -14850.0 293700.0 ;
      RECT  -13650.0 290100.0 -14850.0 291300.0 ;
      RECT  -13650.0 292500.0 -14850.0 293700.0 ;
      RECT  -13650.0 294900.0 -14850.0 296100.0 ;
      RECT  -13650.0 294900.0 -14850.0 296100.0 ;
      RECT  -13650.0 292500.0 -14850.0 293700.0 ;
      RECT  -13650.0 294900.0 -14850.0 296100.0 ;
      RECT  -13650.0 297300.0 -14850.0 298500.0 ;
      RECT  -13650.0 297300.0 -14850.0 298500.0 ;
      RECT  -13650.0 294900.0 -14850.0 296100.0 ;
      RECT  -4950.0 290100.0 -6150.0 291300.0 ;
      RECT  -4950.0 292500.0 -6150.0 293700.0 ;
      RECT  -4950.0 292500.0 -6150.0 293700.0 ;
      RECT  -4950.0 290100.0 -6150.0 291300.0 ;
      RECT  -4950.0 292500.0 -6150.0 293700.0 ;
      RECT  -4950.0 294900.0 -6150.0 296100.0 ;
      RECT  -4950.0 294900.0 -6150.0 296100.0 ;
      RECT  -4950.0 292500.0 -6150.0 293700.0 ;
      RECT  -4950.0 294900.0 -6150.0 296100.0 ;
      RECT  -4950.0 297300.0 -6150.0 298500.0 ;
      RECT  -4950.0 297300.0 -6150.0 298500.0 ;
      RECT  -4950.0 294900.0 -6150.0 296100.0 ;
      RECT  -14250.0 299700.0 -15450.0 300900.0 ;
      RECT  -4350.0 299700.0 -5550.0 300900.0 ;
      RECT  -7050.0 297300.0 -8250.0 296100.0 ;
      RECT  -9000.0 294900.0 -10200.0 293700.0 ;
      RECT  -10950.0 292500.0 -12150.0 291300.0 ;
      RECT  -13650.0 292500.0 -14850.0 293700.0 ;
      RECT  -13650.0 297300.0 -14850.0 298500.0 ;
      RECT  -4950.0 297300.0 -6150.0 298500.0 ;
      RECT  -10950.0 297300.0 -12150.0 298500.0 ;
      RECT  -10950.0 291300.0 -12150.0 292500.0 ;
      RECT  -9000.0 293700.0 -10200.0 294900.0 ;
      RECT  -7050.0 296100.0 -8250.0 297300.0 ;
      RECT  -10950.0 297300.0 -12150.0 298500.0 ;
      RECT  -16350.0 288300.0 -17250.0 303900.0 ;
      RECT  -2550.0 288300.0 -3450.0 303900.0 ;
      RECT  -14850.0 310500.0 -16800.0 311700.0 ;
      RECT  -3000.0 310500.0 -4950.0 311700.0 ;
      RECT  -4350.0 305700.0 -2550.0 306900.0 ;
      RECT  -13650.0 305700.0 -17250.0 306900.0 ;
      RECT  -4350.0 308400.0 -13650.0 309300.0 ;
      RECT  -13650.0 305700.0 -14850.0 306900.0 ;
      RECT  -13650.0 308100.0 -14850.0 309300.0 ;
      RECT  -13650.0 308100.0 -14850.0 309300.0 ;
      RECT  -13650.0 305700.0 -14850.0 306900.0 ;
      RECT  -4350.0 305700.0 -5550.0 306900.0 ;
      RECT  -4350.0 308100.0 -5550.0 309300.0 ;
      RECT  -4350.0 308100.0 -5550.0 309300.0 ;
      RECT  -4350.0 305700.0 -5550.0 306900.0 ;
      RECT  -14250.0 310500.0 -15450.0 311700.0 ;
      RECT  -4350.0 310500.0 -5550.0 311700.0 ;
      RECT  -9000.0 306300.0 -10200.0 307500.0 ;
      RECT  -9000.0 306300.0 -10200.0 307500.0 ;
      RECT  -9150.0 308850.0 -10050.0 309750.0 ;
      RECT  -16350.0 303900.0 -17250.0 313500.0 ;
      RECT  -2550.0 303900.0 -3450.0 313500.0 ;
      RECT  -29250.0 290100.0 -31050.0 291300.0 ;
      RECT  -29250.0 294900.0 -31050.0 296100.0 ;
      RECT  -20550.0 290100.0 -16350.0 291300.0 ;
      RECT  -18750.0 297300.0 -16800.0 298500.0 ;
      RECT  -30600.0 297300.0 -28650.0 298500.0 ;
      RECT  -20550.0 290100.0 -19350.0 291300.0 ;
      RECT  -20550.0 292500.0 -19350.0 293700.0 ;
      RECT  -20550.0 292500.0 -19350.0 293700.0 ;
      RECT  -20550.0 290100.0 -19350.0 291300.0 ;
      RECT  -20550.0 292500.0 -19350.0 293700.0 ;
      RECT  -20550.0 294900.0 -19350.0 296100.0 ;
      RECT  -20550.0 294900.0 -19350.0 296100.0 ;
      RECT  -20550.0 292500.0 -19350.0 293700.0 ;
      RECT  -29250.0 290100.0 -28050.0 291300.0 ;
      RECT  -29250.0 292500.0 -28050.0 293700.0 ;
      RECT  -29250.0 292500.0 -28050.0 293700.0 ;
      RECT  -29250.0 290100.0 -28050.0 291300.0 ;
      RECT  -29250.0 292500.0 -28050.0 293700.0 ;
      RECT  -29250.0 294900.0 -28050.0 296100.0 ;
      RECT  -29250.0 294900.0 -28050.0 296100.0 ;
      RECT  -29250.0 292500.0 -28050.0 293700.0 ;
      RECT  -19350.0 297300.0 -18150.0 298500.0 ;
      RECT  -29250.0 297300.0 -28050.0 298500.0 ;
      RECT  -26850.0 294900.0 -25650.0 293700.0 ;
      RECT  -24150.0 291900.0 -22950.0 290700.0 ;
      RECT  -20550.0 294900.0 -19350.0 296100.0 ;
      RECT  -29250.0 293700.0 -28050.0 292500.0 ;
      RECT  -24150.0 297000.0 -22950.0 295800.0 ;
      RECT  -24150.0 290700.0 -22950.0 291900.0 ;
      RECT  -26850.0 293700.0 -25650.0 294900.0 ;
      RECT  -24150.0 295800.0 -22950.0 297000.0 ;
      RECT  -17250.0 288300.0 -16350.0 302700.0 ;
      RECT  -31050.0 288300.0 -30150.0 302700.0 ;
      RECT  -28650.0 307200.0 -31050.0 308400.0 ;
      RECT  -19950.0 307200.0 -16350.0 308400.0 ;
      RECT  -19950.0 312000.0 -16350.0 313200.0 ;
      RECT  -18750.0 314400.0 -16800.0 315600.0 ;
      RECT  -30600.0 314400.0 -28650.0 315600.0 ;
      RECT  -19950.0 307200.0 -18750.0 308400.0 ;
      RECT  -19950.0 309600.0 -18750.0 310800.0 ;
      RECT  -19950.0 309600.0 -18750.0 310800.0 ;
      RECT  -19950.0 307200.0 -18750.0 308400.0 ;
      RECT  -19950.0 309600.0 -18750.0 310800.0 ;
      RECT  -19950.0 312000.0 -18750.0 313200.0 ;
      RECT  -19950.0 312000.0 -18750.0 313200.0 ;
      RECT  -19950.0 309600.0 -18750.0 310800.0 ;
      RECT  -28650.0 307200.0 -27450.0 308400.0 ;
      RECT  -28650.0 309600.0 -27450.0 310800.0 ;
      RECT  -28650.0 309600.0 -27450.0 310800.0 ;
      RECT  -28650.0 307200.0 -27450.0 308400.0 ;
      RECT  -28650.0 309600.0 -27450.0 310800.0 ;
      RECT  -28650.0 312000.0 -27450.0 313200.0 ;
      RECT  -28650.0 312000.0 -27450.0 313200.0 ;
      RECT  -28650.0 309600.0 -27450.0 310800.0 ;
      RECT  -19350.0 314400.0 -18150.0 315600.0 ;
      RECT  -29250.0 314400.0 -28050.0 315600.0 ;
      RECT  -26100.0 312000.0 -24900.0 310800.0 ;
      RECT  -23400.0 309000.0 -22200.0 307800.0 ;
      RECT  -19950.0 309600.0 -18750.0 310800.0 ;
      RECT  -28650.0 312000.0 -27450.0 313200.0 ;
      RECT  -23400.0 313200.0 -22200.0 312000.0 ;
      RECT  -23400.0 307800.0 -22200.0 309000.0 ;
      RECT  -26100.0 310800.0 -24900.0 312000.0 ;
      RECT  -23400.0 312000.0 -22200.0 313200.0 ;
      RECT  -17250.0 305400.0 -16350.0 319800.0 ;
      RECT  -31050.0 305400.0 -30150.0 319800.0 ;
      RECT  -18750.0 325500.0 -16800.0 324300.0 ;
      RECT  -30600.0 325500.0 -28650.0 324300.0 ;
      RECT  -29250.0 330300.0 -31050.0 329100.0 ;
      RECT  -19950.0 330300.0 -16350.0 329100.0 ;
      RECT  -29250.0 327600.0 -19950.0 326700.0 ;
      RECT  -19950.0 330300.0 -18750.0 329100.0 ;
      RECT  -19950.0 327900.0 -18750.0 326700.0 ;
      RECT  -19950.0 327900.0 -18750.0 326700.0 ;
      RECT  -19950.0 330300.0 -18750.0 329100.0 ;
      RECT  -29250.0 330300.0 -28050.0 329100.0 ;
      RECT  -29250.0 327900.0 -28050.0 326700.0 ;
      RECT  -29250.0 327900.0 -28050.0 326700.0 ;
      RECT  -29250.0 330300.0 -28050.0 329100.0 ;
      RECT  -19350.0 325500.0 -18150.0 324300.0 ;
      RECT  -29250.0 325500.0 -28050.0 324300.0 ;
      RECT  -24600.0 329700.0 -23400.0 328500.0 ;
      RECT  -24600.0 329700.0 -23400.0 328500.0 ;
      RECT  -24450.0 327150.0 -23550.0 326250.0 ;
      RECT  -17250.0 332100.0 -16350.0 322500.0 ;
      RECT  -31050.0 332100.0 -30150.0 322500.0 ;
      RECT  -18750.0 335100.0 -16800.0 333900.0 ;
      RECT  -30600.0 335100.0 -28650.0 333900.0 ;
      RECT  -29250.0 339900.0 -31050.0 338700.0 ;
      RECT  -19950.0 339900.0 -16350.0 338700.0 ;
      RECT  -29250.0 337200.0 -19950.0 336300.0 ;
      RECT  -19950.0 339900.0 -18750.0 338700.0 ;
      RECT  -19950.0 337500.0 -18750.0 336300.0 ;
      RECT  -19950.0 337500.0 -18750.0 336300.0 ;
      RECT  -19950.0 339900.0 -18750.0 338700.0 ;
      RECT  -29250.0 339900.0 -28050.0 338700.0 ;
      RECT  -29250.0 337500.0 -28050.0 336300.0 ;
      RECT  -29250.0 337500.0 -28050.0 336300.0 ;
      RECT  -29250.0 339900.0 -28050.0 338700.0 ;
      RECT  -19350.0 335100.0 -18150.0 333900.0 ;
      RECT  -29250.0 335100.0 -28050.0 333900.0 ;
      RECT  -24600.0 339300.0 -23400.0 338100.0 ;
      RECT  -24600.0 339300.0 -23400.0 338100.0 ;
      RECT  -24450.0 336750.0 -23550.0 335850.0 ;
      RECT  -17250.0 341700.0 -16350.0 332100.0 ;
      RECT  -31050.0 341700.0 -30150.0 332100.0 ;
      RECT  -32550.0 299700.0 -30150.0 300900.0 ;
      RECT  -41250.0 299700.0 -44850.0 300900.0 ;
      RECT  -41250.0 304500.0 -44850.0 305700.0 ;
      RECT  -42450.0 309300.0 -44400.0 310500.0 ;
      RECT  -30600.0 309300.0 -32550.0 310500.0 ;
      RECT  -41250.0 299700.0 -42450.0 300900.0 ;
      RECT  -41250.0 302100.0 -42450.0 303300.0 ;
      RECT  -41250.0 302100.0 -42450.0 303300.0 ;
      RECT  -41250.0 299700.0 -42450.0 300900.0 ;
      RECT  -41250.0 302100.0 -42450.0 303300.0 ;
      RECT  -41250.0 304500.0 -42450.0 305700.0 ;
      RECT  -41250.0 304500.0 -42450.0 305700.0 ;
      RECT  -41250.0 302100.0 -42450.0 303300.0 ;
      RECT  -41250.0 304500.0 -42450.0 305700.0 ;
      RECT  -41250.0 306900.0 -42450.0 308100.0 ;
      RECT  -41250.0 306900.0 -42450.0 308100.0 ;
      RECT  -41250.0 304500.0 -42450.0 305700.0 ;
      RECT  -32550.0 299700.0 -33750.0 300900.0 ;
      RECT  -32550.0 302100.0 -33750.0 303300.0 ;
      RECT  -32550.0 302100.0 -33750.0 303300.0 ;
      RECT  -32550.0 299700.0 -33750.0 300900.0 ;
      RECT  -32550.0 302100.0 -33750.0 303300.0 ;
      RECT  -32550.0 304500.0 -33750.0 305700.0 ;
      RECT  -32550.0 304500.0 -33750.0 305700.0 ;
      RECT  -32550.0 302100.0 -33750.0 303300.0 ;
      RECT  -32550.0 304500.0 -33750.0 305700.0 ;
      RECT  -32550.0 306900.0 -33750.0 308100.0 ;
      RECT  -32550.0 306900.0 -33750.0 308100.0 ;
      RECT  -32550.0 304500.0 -33750.0 305700.0 ;
      RECT  -41850.0 309300.0 -43050.0 310500.0 ;
      RECT  -31950.0 309300.0 -33150.0 310500.0 ;
      RECT  -34650.0 306900.0 -35850.0 305700.0 ;
      RECT  -36600.0 304500.0 -37800.0 303300.0 ;
      RECT  -38550.0 302100.0 -39750.0 300900.0 ;
      RECT  -41250.0 302100.0 -42450.0 303300.0 ;
      RECT  -41250.0 306900.0 -42450.0 308100.0 ;
      RECT  -32550.0 306900.0 -33750.0 308100.0 ;
      RECT  -38550.0 306900.0 -39750.0 308100.0 ;
      RECT  -38550.0 300900.0 -39750.0 302100.0 ;
      RECT  -36600.0 303300.0 -37800.0 304500.0 ;
      RECT  -34650.0 305700.0 -35850.0 306900.0 ;
      RECT  -38550.0 306900.0 -39750.0 308100.0 ;
      RECT  -43950.0 297900.0 -44850.0 313500.0 ;
      RECT  -30150.0 297900.0 -31050.0 313500.0 ;
      RECT  -42450.0 320100.0 -44400.0 321300.0 ;
      RECT  -30600.0 320100.0 -32550.0 321300.0 ;
      RECT  -31950.0 315300.0 -30150.0 316500.0 ;
      RECT  -41250.0 315300.0 -44850.0 316500.0 ;
      RECT  -31950.0 318000.0 -41250.0 318900.0 ;
      RECT  -41250.0 315300.0 -42450.0 316500.0 ;
      RECT  -41250.0 317700.0 -42450.0 318900.0 ;
      RECT  -41250.0 317700.0 -42450.0 318900.0 ;
      RECT  -41250.0 315300.0 -42450.0 316500.0 ;
      RECT  -31950.0 315300.0 -33150.0 316500.0 ;
      RECT  -31950.0 317700.0 -33150.0 318900.0 ;
      RECT  -31950.0 317700.0 -33150.0 318900.0 ;
      RECT  -31950.0 315300.0 -33150.0 316500.0 ;
      RECT  -41850.0 320100.0 -43050.0 321300.0 ;
      RECT  -31950.0 320100.0 -33150.0 321300.0 ;
      RECT  -36600.0 315900.0 -37800.0 317100.0 ;
      RECT  -36600.0 315900.0 -37800.0 317100.0 ;
      RECT  -36750.0 318450.0 -37650.0 319350.0 ;
      RECT  -43950.0 313500.0 -44850.0 323100.0 ;
      RECT  -30150.0 313500.0 -31050.0 323100.0 ;
      RECT  -42450.0 329700.0 -44400.0 330900.0 ;
      RECT  -30600.0 329700.0 -32550.0 330900.0 ;
      RECT  -31950.0 324900.0 -30150.0 326100.0 ;
      RECT  -41250.0 324900.0 -44850.0 326100.0 ;
      RECT  -31950.0 327600.0 -41250.0 328500.0 ;
      RECT  -41250.0 324900.0 -42450.0 326100.0 ;
      RECT  -41250.0 327300.0 -42450.0 328500.0 ;
      RECT  -41250.0 327300.0 -42450.0 328500.0 ;
      RECT  -41250.0 324900.0 -42450.0 326100.0 ;
      RECT  -31950.0 324900.0 -33150.0 326100.0 ;
      RECT  -31950.0 327300.0 -33150.0 328500.0 ;
      RECT  -31950.0 327300.0 -33150.0 328500.0 ;
      RECT  -31950.0 324900.0 -33150.0 326100.0 ;
      RECT  -41850.0 329700.0 -43050.0 330900.0 ;
      RECT  -31950.0 329700.0 -33150.0 330900.0 ;
      RECT  -36600.0 325500.0 -37800.0 326700.0 ;
      RECT  -36600.0 325500.0 -37800.0 326700.0 ;
      RECT  -36750.0 328050.0 -37650.0 328950.0 ;
      RECT  -43950.0 323100.0 -44850.0 332700.0 ;
      RECT  -30150.0 323100.0 -31050.0 332700.0 ;
      RECT  -42450.0 339300.0 -44400.0 340500.0 ;
      RECT  -30600.0 339300.0 -32550.0 340500.0 ;
      RECT  -31950.0 334500.0 -30150.0 335700.0 ;
      RECT  -41250.0 334500.0 -44850.0 335700.0 ;
      RECT  -31950.0 337200.0 -41250.0 338100.0 ;
      RECT  -41250.0 334500.0 -42450.0 335700.0 ;
      RECT  -41250.0 336900.0 -42450.0 338100.0 ;
      RECT  -41250.0 336900.0 -42450.0 338100.0 ;
      RECT  -41250.0 334500.0 -42450.0 335700.0 ;
      RECT  -31950.0 334500.0 -33150.0 335700.0 ;
      RECT  -31950.0 336900.0 -33150.0 338100.0 ;
      RECT  -31950.0 336900.0 -33150.0 338100.0 ;
      RECT  -31950.0 334500.0 -33150.0 335700.0 ;
      RECT  -41850.0 339300.0 -43050.0 340500.0 ;
      RECT  -31950.0 339300.0 -33150.0 340500.0 ;
      RECT  -36600.0 335100.0 -37800.0 336300.0 ;
      RECT  -36600.0 335100.0 -37800.0 336300.0 ;
      RECT  -36750.0 337650.0 -37650.0 338550.0 ;
      RECT  -43950.0 332700.0 -44850.0 342300.0 ;
      RECT  -30150.0 332700.0 -31050.0 342300.0 ;
      RECT  -30150.0 459150.0 -31050.0 437100.0 ;
      RECT  -31050.0 376350.0 -35400.0 377250.0 ;
      RECT  -31050.0 399750.0 -35400.0 400650.0 ;
      RECT  -31050.0 403950.0 -35400.0 404850.0 ;
      RECT  -31050.0 427350.0 -35400.0 428250.0 ;
      RECT  -30150.0 350850.0 -36000.0 351750.0 ;
      RECT  -36000.0 350850.0 -46200.0 351750.0 ;
      RECT  -48300.0 387900.0 -36000.0 388800.0 ;
      RECT  -48300.0 415500.0 -36000.0 416400.0 ;
      RECT  -48300.0 360300.0 -36000.0 361200.0 ;
      RECT  -23550.0 377100.0 -24450.0 389700.0 ;
      RECT  -23550.0 372150.0 -24450.0 373050.0 ;
      RECT  -23550.0 372600.0 -24450.0 377100.0 ;
      RECT  -24000.0 372150.0 -35400.0 373050.0 ;
      RECT  -16800.0 377850.0 -19050.0 378750.0 ;
      RECT  -19200.0 363150.0 -20100.0 364050.0 ;
      RECT  -23550.0 363150.0 -24450.0 364050.0 ;
      RECT  -19200.0 363600.0 -20100.0 375300.0 ;
      RECT  -19650.0 363150.0 -24000.0 364050.0 ;
      RECT  -23550.0 358500.0 -24450.0 363600.0 ;
      RECT  -24000.0 363150.0 -32850.0 364050.0 ;
      RECT  -32850.0 355050.0 -39600.0 355950.0 ;
      RECT  -23400.0 357300.0 -24600.0 358500.0 ;
      RECT  -23550.0 389700.0 -24450.0 393450.0 ;
      RECT  -18750.0 354300.0 -16800.0 353100.0 ;
      RECT  -30600.0 354300.0 -28650.0 353100.0 ;
      RECT  -29250.0 359100.0 -31050.0 357900.0 ;
      RECT  -19950.0 359100.0 -16350.0 357900.0 ;
      RECT  -29250.0 356400.0 -19950.0 355500.0 ;
      RECT  -19950.0 359100.0 -18750.0 357900.0 ;
      RECT  -19950.0 356700.0 -18750.0 355500.0 ;
      RECT  -19950.0 356700.0 -18750.0 355500.0 ;
      RECT  -19950.0 359100.0 -18750.0 357900.0 ;
      RECT  -29250.0 359100.0 -28050.0 357900.0 ;
      RECT  -29250.0 356700.0 -28050.0 355500.0 ;
      RECT  -29250.0 356700.0 -28050.0 355500.0 ;
      RECT  -29250.0 359100.0 -28050.0 357900.0 ;
      RECT  -19350.0 354300.0 -18150.0 353100.0 ;
      RECT  -29250.0 354300.0 -28050.0 353100.0 ;
      RECT  -24600.0 358500.0 -23400.0 357300.0 ;
      RECT  -24600.0 358500.0 -23400.0 357300.0 ;
      RECT  -24450.0 355950.0 -23550.0 355050.0 ;
      RECT  -17250.0 360900.0 -16350.0 351300.0 ;
      RECT  -31050.0 360900.0 -30150.0 351300.0 ;
      RECT  -20250.0 375300.0 -19050.0 376500.0 ;
      RECT  -20250.0 377700.0 -19050.0 378900.0 ;
      RECT  -20250.0 377700.0 -19050.0 378900.0 ;
      RECT  -20250.0 375300.0 -19050.0 376500.0 ;
      RECT  -31050.0 458250.0 -30150.0 459150.0 ;
      RECT  -3450.0 458250.0 -2550.0 459150.0 ;
      RECT  -31050.0 456900.0 -30150.0 458700.0 ;
      RECT  -30600.0 458250.0 -3000.0 459150.0 ;
      RECT  -3450.0 456900.0 -2550.0 458700.0 ;
      RECT  -14850.0 396300.0 -16800.0 397500.0 ;
      RECT  -3000.0 396300.0 -4950.0 397500.0 ;
      RECT  -4350.0 391500.0 -2550.0 392700.0 ;
      RECT  -13650.0 391500.0 -17250.0 392700.0 ;
      RECT  -4350.0 394200.0 -13650.0 395100.0 ;
      RECT  -13650.0 391500.0 -14850.0 392700.0 ;
      RECT  -13650.0 393900.0 -14850.0 395100.0 ;
      RECT  -13650.0 393900.0 -14850.0 395100.0 ;
      RECT  -13650.0 391500.0 -14850.0 392700.0 ;
      RECT  -4350.0 391500.0 -5550.0 392700.0 ;
      RECT  -4350.0 393900.0 -5550.0 395100.0 ;
      RECT  -4350.0 393900.0 -5550.0 395100.0 ;
      RECT  -4350.0 391500.0 -5550.0 392700.0 ;
      RECT  -14250.0 396300.0 -15450.0 397500.0 ;
      RECT  -4350.0 396300.0 -5550.0 397500.0 ;
      RECT  -9000.0 392100.0 -10200.0 393300.0 ;
      RECT  -9000.0 392100.0 -10200.0 393300.0 ;
      RECT  -9150.0 394650.0 -10050.0 395550.0 ;
      RECT  -16350.0 389700.0 -17250.0 399300.0 ;
      RECT  -2550.0 389700.0 -3450.0 399300.0 ;
      RECT  -14850.0 405900.0 -16800.0 407100.0 ;
      RECT  -3000.0 405900.0 -4950.0 407100.0 ;
      RECT  -4350.0 401100.0 -2550.0 402300.0 ;
      RECT  -13650.0 401100.0 -17250.0 402300.0 ;
      RECT  -4350.0 403800.0 -13650.0 404700.0 ;
      RECT  -13650.0 401100.0 -14850.0 402300.0 ;
      RECT  -13650.0 403500.0 -14850.0 404700.0 ;
      RECT  -13650.0 403500.0 -14850.0 404700.0 ;
      RECT  -13650.0 401100.0 -14850.0 402300.0 ;
      RECT  -4350.0 401100.0 -5550.0 402300.0 ;
      RECT  -4350.0 403500.0 -5550.0 404700.0 ;
      RECT  -4350.0 403500.0 -5550.0 404700.0 ;
      RECT  -4350.0 401100.0 -5550.0 402300.0 ;
      RECT  -14250.0 405900.0 -15450.0 407100.0 ;
      RECT  -4350.0 405900.0 -5550.0 407100.0 ;
      RECT  -9000.0 401700.0 -10200.0 402900.0 ;
      RECT  -9000.0 401700.0 -10200.0 402900.0 ;
      RECT  -9150.0 404250.0 -10050.0 405150.0 ;
      RECT  -16350.0 399300.0 -17250.0 408900.0 ;
      RECT  -2550.0 399300.0 -3450.0 408900.0 ;
      RECT  -10200.0 401700.0 -9000.0 402900.0 ;
      RECT  -14850.0 415500.0 -16800.0 416700.0 ;
      RECT  -3000.0 415500.0 -4950.0 416700.0 ;
      RECT  -4350.0 410700.0 -2550.0 411900.0 ;
      RECT  -13650.0 410700.0 -17250.0 411900.0 ;
      RECT  -4350.0 413400.0 -13650.0 414300.0 ;
      RECT  -13650.0 410700.0 -14850.0 411900.0 ;
      RECT  -13650.0 413100.0 -14850.0 414300.0 ;
      RECT  -13650.0 413100.0 -14850.0 414300.0 ;
      RECT  -13650.0 410700.0 -14850.0 411900.0 ;
      RECT  -4350.0 410700.0 -5550.0 411900.0 ;
      RECT  -4350.0 413100.0 -5550.0 414300.0 ;
      RECT  -4350.0 413100.0 -5550.0 414300.0 ;
      RECT  -4350.0 410700.0 -5550.0 411900.0 ;
      RECT  -14250.0 415500.0 -15450.0 416700.0 ;
      RECT  -4350.0 415500.0 -5550.0 416700.0 ;
      RECT  -9000.0 411300.0 -10200.0 412500.0 ;
      RECT  -9000.0 411300.0 -10200.0 412500.0 ;
      RECT  -9150.0 413850.0 -10050.0 414750.0 ;
      RECT  -16350.0 408900.0 -17250.0 418500.0 ;
      RECT  -2550.0 408900.0 -3450.0 418500.0 ;
      RECT  -10200.0 411300.0 -9000.0 412500.0 ;
      RECT  -14850.0 425100.0 -16800.0 426300.0 ;
      RECT  -3000.0 425100.0 -4950.0 426300.0 ;
      RECT  -4350.0 420300.0 -2550.0 421500.0 ;
      RECT  -13650.0 420300.0 -17250.0 421500.0 ;
      RECT  -4350.0 423000.0 -13650.0 423900.0 ;
      RECT  -13650.0 420300.0 -14850.0 421500.0 ;
      RECT  -13650.0 422700.0 -14850.0 423900.0 ;
      RECT  -13650.0 422700.0 -14850.0 423900.0 ;
      RECT  -13650.0 420300.0 -14850.0 421500.0 ;
      RECT  -4350.0 420300.0 -5550.0 421500.0 ;
      RECT  -4350.0 422700.0 -5550.0 423900.0 ;
      RECT  -4350.0 422700.0 -5550.0 423900.0 ;
      RECT  -4350.0 420300.0 -5550.0 421500.0 ;
      RECT  -14250.0 425100.0 -15450.0 426300.0 ;
      RECT  -4350.0 425100.0 -5550.0 426300.0 ;
      RECT  -9000.0 420900.0 -10200.0 422100.0 ;
      RECT  -9000.0 420900.0 -10200.0 422100.0 ;
      RECT  -9150.0 423450.0 -10050.0 424350.0 ;
      RECT  -16350.0 418500.0 -17250.0 428100.0 ;
      RECT  -2550.0 418500.0 -3450.0 428100.0 ;
      RECT  -10200.0 420900.0 -9000.0 422100.0 ;
      RECT  -14850.0 434700.0 -16800.0 435900.0 ;
      RECT  -3000.0 434700.0 -4950.0 435900.0 ;
      RECT  -4350.0 429900.0 -2550.0 431100.0 ;
      RECT  -13650.0 429900.0 -17250.0 431100.0 ;
      RECT  -4350.0 432600.0 -13650.0 433500.0 ;
      RECT  -13650.0 429900.0 -14850.0 431100.0 ;
      RECT  -13650.0 432300.0 -14850.0 433500.0 ;
      RECT  -13650.0 432300.0 -14850.0 433500.0 ;
      RECT  -13650.0 429900.0 -14850.0 431100.0 ;
      RECT  -4350.0 429900.0 -5550.0 431100.0 ;
      RECT  -4350.0 432300.0 -5550.0 433500.0 ;
      RECT  -4350.0 432300.0 -5550.0 433500.0 ;
      RECT  -4350.0 429900.0 -5550.0 431100.0 ;
      RECT  -14250.0 434700.0 -15450.0 435900.0 ;
      RECT  -4350.0 434700.0 -5550.0 435900.0 ;
      RECT  -9000.0 430500.0 -10200.0 431700.0 ;
      RECT  -9000.0 430500.0 -10200.0 431700.0 ;
      RECT  -9150.0 433050.0 -10050.0 433950.0 ;
      RECT  -16350.0 428100.0 -17250.0 437700.0 ;
      RECT  -2550.0 428100.0 -3450.0 437700.0 ;
      RECT  -10200.0 430500.0 -9000.0 431700.0 ;
      RECT  -14850.0 444300.0 -16800.0 445500.0 ;
      RECT  -3000.0 444300.0 -4950.0 445500.0 ;
      RECT  -4350.0 439500.0 -2550.0 440700.0 ;
      RECT  -13650.0 439500.0 -17250.0 440700.0 ;
      RECT  -4350.0 442200.0 -13650.0 443100.0 ;
      RECT  -13650.0 439500.0 -14850.0 440700.0 ;
      RECT  -13650.0 441900.0 -14850.0 443100.0 ;
      RECT  -13650.0 441900.0 -14850.0 443100.0 ;
      RECT  -13650.0 439500.0 -14850.0 440700.0 ;
      RECT  -4350.0 439500.0 -5550.0 440700.0 ;
      RECT  -4350.0 441900.0 -5550.0 443100.0 ;
      RECT  -4350.0 441900.0 -5550.0 443100.0 ;
      RECT  -4350.0 439500.0 -5550.0 440700.0 ;
      RECT  -14250.0 444300.0 -15450.0 445500.0 ;
      RECT  -4350.0 444300.0 -5550.0 445500.0 ;
      RECT  -9000.0 440100.0 -10200.0 441300.0 ;
      RECT  -9000.0 440100.0 -10200.0 441300.0 ;
      RECT  -9150.0 442650.0 -10050.0 443550.0 ;
      RECT  -16350.0 437700.0 -17250.0 447300.0 ;
      RECT  -2550.0 437700.0 -3450.0 447300.0 ;
      RECT  -10200.0 440100.0 -9000.0 441300.0 ;
      RECT  -14850.0 453900.0 -16800.0 455100.0 ;
      RECT  -3000.0 453900.0 -4950.0 455100.0 ;
      RECT  -4350.0 449100.0 -2550.0 450300.0 ;
      RECT  -13650.0 449100.0 -17250.0 450300.0 ;
      RECT  -4350.0 451800.0 -13650.0 452700.0 ;
      RECT  -13650.0 449100.0 -14850.0 450300.0 ;
      RECT  -13650.0 451500.0 -14850.0 452700.0 ;
      RECT  -13650.0 451500.0 -14850.0 452700.0 ;
      RECT  -13650.0 449100.0 -14850.0 450300.0 ;
      RECT  -4350.0 449100.0 -5550.0 450300.0 ;
      RECT  -4350.0 451500.0 -5550.0 452700.0 ;
      RECT  -4350.0 451500.0 -5550.0 452700.0 ;
      RECT  -4350.0 449100.0 -5550.0 450300.0 ;
      RECT  -14250.0 453900.0 -15450.0 455100.0 ;
      RECT  -4350.0 453900.0 -5550.0 455100.0 ;
      RECT  -9000.0 449700.0 -10200.0 450900.0 ;
      RECT  -9000.0 449700.0 -10200.0 450900.0 ;
      RECT  -9150.0 452250.0 -10050.0 453150.0 ;
      RECT  -16350.0 447300.0 -17250.0 456900.0 ;
      RECT  -2550.0 447300.0 -3450.0 456900.0 ;
      RECT  -10200.0 449700.0 -9000.0 450900.0 ;
      RECT  -18750.0 440700.0 -16800.0 439500.0 ;
      RECT  -30600.0 440700.0 -28650.0 439500.0 ;
      RECT  -29250.0 445500.0 -31050.0 444300.0 ;
      RECT  -19950.0 445500.0 -16350.0 444300.0 ;
      RECT  -29250.0 442800.0 -19950.0 441900.0 ;
      RECT  -19950.0 445500.0 -18750.0 444300.0 ;
      RECT  -19950.0 443100.0 -18750.0 441900.0 ;
      RECT  -19950.0 443100.0 -18750.0 441900.0 ;
      RECT  -19950.0 445500.0 -18750.0 444300.0 ;
      RECT  -29250.0 445500.0 -28050.0 444300.0 ;
      RECT  -29250.0 443100.0 -28050.0 441900.0 ;
      RECT  -29250.0 443100.0 -28050.0 441900.0 ;
      RECT  -29250.0 445500.0 -28050.0 444300.0 ;
      RECT  -19350.0 440700.0 -18150.0 439500.0 ;
      RECT  -29250.0 440700.0 -28050.0 439500.0 ;
      RECT  -24600.0 444900.0 -23400.0 443700.0 ;
      RECT  -24600.0 444900.0 -23400.0 443700.0 ;
      RECT  -24450.0 442350.0 -23550.0 441450.0 ;
      RECT  -17250.0 447300.0 -16350.0 437700.0 ;
      RECT  -31050.0 447300.0 -30150.0 437700.0 ;
      RECT  -24600.0 443700.0 -23400.0 444900.0 ;
      RECT  -18750.0 431100.0 -16800.0 429900.0 ;
      RECT  -30600.0 431100.0 -28650.0 429900.0 ;
      RECT  -29250.0 435900.0 -31050.0 434700.0 ;
      RECT  -19950.0 435900.0 -16350.0 434700.0 ;
      RECT  -29250.0 433200.0 -19950.0 432300.0 ;
      RECT  -19950.0 435900.0 -18750.0 434700.0 ;
      RECT  -19950.0 433500.0 -18750.0 432300.0 ;
      RECT  -19950.0 433500.0 -18750.0 432300.0 ;
      RECT  -19950.0 435900.0 -18750.0 434700.0 ;
      RECT  -29250.0 435900.0 -28050.0 434700.0 ;
      RECT  -29250.0 433500.0 -28050.0 432300.0 ;
      RECT  -29250.0 433500.0 -28050.0 432300.0 ;
      RECT  -29250.0 435900.0 -28050.0 434700.0 ;
      RECT  -19350.0 431100.0 -18150.0 429900.0 ;
      RECT  -29250.0 431100.0 -28050.0 429900.0 ;
      RECT  -24600.0 435300.0 -23400.0 434100.0 ;
      RECT  -24600.0 435300.0 -23400.0 434100.0 ;
      RECT  -24450.0 432750.0 -23550.0 431850.0 ;
      RECT  -17250.0 437700.0 -16350.0 428100.0 ;
      RECT  -31050.0 437700.0 -30150.0 428100.0 ;
      RECT  -24600.0 434100.0 -23400.0 435300.0 ;
      RECT  -18750.0 421500.0 -16800.0 420300.0 ;
      RECT  -30600.0 421500.0 -28650.0 420300.0 ;
      RECT  -29250.0 426300.0 -31050.0 425100.0 ;
      RECT  -19950.0 426300.0 -16350.0 425100.0 ;
      RECT  -29250.0 423600.0 -19950.0 422700.0 ;
      RECT  -19950.0 426300.0 -18750.0 425100.0 ;
      RECT  -19950.0 423900.0 -18750.0 422700.0 ;
      RECT  -19950.0 423900.0 -18750.0 422700.0 ;
      RECT  -19950.0 426300.0 -18750.0 425100.0 ;
      RECT  -29250.0 426300.0 -28050.0 425100.0 ;
      RECT  -29250.0 423900.0 -28050.0 422700.0 ;
      RECT  -29250.0 423900.0 -28050.0 422700.0 ;
      RECT  -29250.0 426300.0 -28050.0 425100.0 ;
      RECT  -19350.0 421500.0 -18150.0 420300.0 ;
      RECT  -29250.0 421500.0 -28050.0 420300.0 ;
      RECT  -24600.0 425700.0 -23400.0 424500.0 ;
      RECT  -24600.0 425700.0 -23400.0 424500.0 ;
      RECT  -24450.0 423150.0 -23550.0 422250.0 ;
      RECT  -17250.0 428100.0 -16350.0 418500.0 ;
      RECT  -31050.0 428100.0 -30150.0 418500.0 ;
      RECT  -24600.0 424500.0 -23400.0 425700.0 ;
      RECT  -18750.0 411900.0 -16800.0 410700.0 ;
      RECT  -30600.0 411900.0 -28650.0 410700.0 ;
      RECT  -29250.0 416700.0 -31050.0 415500.0 ;
      RECT  -19950.0 416700.0 -16350.0 415500.0 ;
      RECT  -29250.0 414000.0 -19950.0 413100.0 ;
      RECT  -19950.0 416700.0 -18750.0 415500.0 ;
      RECT  -19950.0 414300.0 -18750.0 413100.0 ;
      RECT  -19950.0 414300.0 -18750.0 413100.0 ;
      RECT  -19950.0 416700.0 -18750.0 415500.0 ;
      RECT  -29250.0 416700.0 -28050.0 415500.0 ;
      RECT  -29250.0 414300.0 -28050.0 413100.0 ;
      RECT  -29250.0 414300.0 -28050.0 413100.0 ;
      RECT  -29250.0 416700.0 -28050.0 415500.0 ;
      RECT  -19350.0 411900.0 -18150.0 410700.0 ;
      RECT  -29250.0 411900.0 -28050.0 410700.0 ;
      RECT  -24600.0 416100.0 -23400.0 414900.0 ;
      RECT  -24600.0 416100.0 -23400.0 414900.0 ;
      RECT  -24450.0 413550.0 -23550.0 412650.0 ;
      RECT  -17250.0 418500.0 -16350.0 408900.0 ;
      RECT  -31050.0 418500.0 -30150.0 408900.0 ;
      RECT  -24600.0 414900.0 -23400.0 416100.0 ;
      RECT  -18750.0 402300.0 -16800.0 401100.0 ;
      RECT  -30600.0 402300.0 -28650.0 401100.0 ;
      RECT  -29250.0 407100.0 -31050.0 405900.0 ;
      RECT  -19950.0 407100.0 -16350.0 405900.0 ;
      RECT  -29250.0 404400.0 -19950.0 403500.0 ;
      RECT  -19950.0 407100.0 -18750.0 405900.0 ;
      RECT  -19950.0 404700.0 -18750.0 403500.0 ;
      RECT  -19950.0 404700.0 -18750.0 403500.0 ;
      RECT  -19950.0 407100.0 -18750.0 405900.0 ;
      RECT  -29250.0 407100.0 -28050.0 405900.0 ;
      RECT  -29250.0 404700.0 -28050.0 403500.0 ;
      RECT  -29250.0 404700.0 -28050.0 403500.0 ;
      RECT  -29250.0 407100.0 -28050.0 405900.0 ;
      RECT  -19350.0 402300.0 -18150.0 401100.0 ;
      RECT  -29250.0 402300.0 -28050.0 401100.0 ;
      RECT  -24600.0 406500.0 -23400.0 405300.0 ;
      RECT  -24600.0 406500.0 -23400.0 405300.0 ;
      RECT  -24450.0 403950.0 -23550.0 403050.0 ;
      RECT  -17250.0 408900.0 -16350.0 399300.0 ;
      RECT  -31050.0 408900.0 -30150.0 399300.0 ;
      RECT  -24600.0 405300.0 -23400.0 406500.0 ;
      RECT  -18750.0 392700.0 -16800.0 391500.0 ;
      RECT  -30600.0 392700.0 -28650.0 391500.0 ;
      RECT  -29250.0 397500.0 -31050.0 396300.0 ;
      RECT  -19950.0 397500.0 -16350.0 396300.0 ;
      RECT  -29250.0 394800.0 -19950.0 393900.0 ;
      RECT  -19950.0 397500.0 -18750.0 396300.0 ;
      RECT  -19950.0 395100.0 -18750.0 393900.0 ;
      RECT  -19950.0 395100.0 -18750.0 393900.0 ;
      RECT  -19950.0 397500.0 -18750.0 396300.0 ;
      RECT  -29250.0 397500.0 -28050.0 396300.0 ;
      RECT  -29250.0 395100.0 -28050.0 393900.0 ;
      RECT  -29250.0 395100.0 -28050.0 393900.0 ;
      RECT  -29250.0 397500.0 -28050.0 396300.0 ;
      RECT  -19350.0 392700.0 -18150.0 391500.0 ;
      RECT  -29250.0 392700.0 -28050.0 391500.0 ;
      RECT  -24600.0 396900.0 -23400.0 395700.0 ;
      RECT  -24600.0 396900.0 -23400.0 395700.0 ;
      RECT  -24450.0 394350.0 -23550.0 393450.0 ;
      RECT  -17250.0 399300.0 -16350.0 389700.0 ;
      RECT  -31050.0 399300.0 -30150.0 389700.0 ;
      RECT  -24600.0 395700.0 -23400.0 396900.0 ;
      RECT  -10200.0 394500.0 -9000.0 395700.0 ;
      RECT  -10200.0 423300.0 -9000.0 424500.0 ;
      RECT  -10200.0 452100.0 -9000.0 453300.0 ;
      RECT  -24600.0 422100.0 -23400.0 423300.0 ;
      RECT  -10200.0 392100.0 -9000.0 393300.0 ;
      RECT  -24450.0 389700.0 -23550.0 393450.0 ;
      RECT  -17250.0 389700.0 -16350.0 456900.0 ;
      RECT  -31050.0 389700.0 -30150.0 456900.0 ;
      RECT  -3450.0 389700.0 -2550.0 456900.0 ;
      RECT  -36000.0 374700.0 -46200.0 360900.0 ;
      RECT  -36000.0 374700.0 -46200.0 388500.0 ;
      RECT  -36000.0 402300.0 -46200.0 388500.0 ;
      RECT  -36000.0 402300.0 -46200.0 416100.0 ;
      RECT  -36000.0 429900.0 -46200.0 416100.0 ;
      RECT  -35400.0 376200.0 -46800.0 377400.0 ;
      RECT  -35400.0 399600.0 -46800.0 400800.0 ;
      RECT  -35400.0 403800.0 -46800.0 405000.0 ;
      RECT  -35400.0 427200.0 -46800.0 428400.0 ;
      RECT  -35400.0 387900.0 -46800.0 388800.0 ;
      RECT  -35400.0 415500.0 -46800.0 416400.0 ;
      RECT  -30450.0 376200.0 -31650.0 377400.0 ;
      RECT  -30450.0 399600.0 -31650.0 400800.0 ;
      RECT  -30450.0 403800.0 -31650.0 405000.0 ;
      RECT  -30450.0 427200.0 -31650.0 428400.0 ;
      RECT  -30600.0 389700.0 -31800.0 390900.0 ;
      RECT  -30000.0 350100.0 -31200.0 351300.0 ;
      RECT  -36600.0 350700.0 -35400.0 351900.0 ;
      RECT  -46800.0 350700.0 -45600.0 351900.0 ;
      RECT  -23400.0 376500.0 -24600.0 377700.0 ;
      RECT  -33450.0 363000.0 -32250.0 364200.0 ;
      RECT  -33450.0 354900.0 -32250.0 356100.0 ;
      RECT  -40200.0 354900.0 -39000.0 356100.0 ;
      RECT  -9000.0 341700.0 -9900.0 392100.0 ;
      RECT  -23550.0 341700.0 -24450.0 355050.0 ;
      RECT  -48300.0 341700.0 -49200.0 432150.0 ;
      RECT  -16350.0 341700.0 -17250.0 389700.0 ;
      RECT  -30150.0 341700.0 -31050.0 351300.0 ;
      RECT  -2550.0 341700.0 -3450.0 389700.0 ;
      RECT  -8850.0 265050.0 -10050.0 263850.0 ;
      RECT  -8850.0 224100.0 -10050.0 222900.0 ;
      RECT  -18900.0 185250.0 -20100.0 184050.0 ;
      RECT  -22950.0 265050.0 -24150.0 263850.0 ;
      RECT  -25650.0 270450.0 -26850.0 269250.0 ;
      RECT  -22200.0 307800.0 -23400.0 306600.0 ;
      RECT  -24900.0 310800.0 -26100.0 309600.0 ;
      RECT  -10950.0 283950.0 -12150.0 282750.0 ;
      RECT  -9000.0 281250.0 -10200.0 280050.0 ;
      RECT  -7050.0 273150.0 -8250.0 271950.0 ;
      RECT  -38550.0 283950.0 -39750.0 282750.0 ;
      RECT  -36600.0 273150.0 -37800.0 271950.0 ;
      RECT  -34650.0 275850.0 -35850.0 274650.0 ;
      RECT  -22950.0 302100.0 -24150.0 303300.0 ;
      RECT  -22200.0 319200.0 -23400.0 320400.0 ;
      RECT  -36600.0 341700.0 -37800.0 342900.0 ;
      RECT  -23400.0 321900.0 -24600.0 323100.0 ;
      RECT  -2400.0 267750.0 -3600.0 266550.0 ;
      RECT  -16200.0 278550.0 -17400.0 277350.0 ;
      RECT  -30000.0 267750.0 -31200.0 266550.0 ;
      RECT  -43800.0 278550.0 -45000.0 277350.0 ;
      RECT  -9000.0 181800.0 -10200.0 185400.0 ;
      RECT  -16350.0 181800.0 -17250.0 182700.0 ;
      RECT  -2550.0 181800.0 -3450.0 182700.0 ;
   LAYER  metal2 ;
      RECT  109650.0 319800.0 110550.0 322500.0 ;
      RECT  106950.0 339600.0 107850.0 342300.0 ;
      RECT  101550.0 300000.0 102450.0 302700.0 ;
      RECT  98850.0 317100.0 99750.0 319800.0 ;
      RECT  104250.0 280650.0 105150.0 283350.0 ;
      RECT  96150.0 261750.0 97050.0 264450.0 ;
      RECT  6300.0 275250.0 7200.0 277950.0 ;
      RECT  -3000.0 266700.0 1800.0 267600.0 ;
      RECT  96150.0 0.0 97050.0 461850.0 ;
      RECT  98850.0 0.0 99750.0 461850.0 ;
      RECT  101550.0 0.0 102450.0 461850.0 ;
      RECT  104250.0 0.0 105150.0 461850.0 ;
      RECT  106950.0 0.0 107850.0 461850.0 ;
      RECT  109650.0 0.0 110550.0 461850.0 ;
      RECT  85350.0 47400.0 86250.0 209400.0 ;
      RECT  88050.0 47400.0 88950.0 209400.0 ;
      RECT  90750.0 47400.0 91650.0 209400.0 ;
      RECT  93450.0 47400.0 94350.0 209400.0 ;
      RECT  122550.0 432600.0 123450.0 433800.0 ;
      RECT  132750.0 432600.0 133650.0 433800.0 ;
      RECT  121050.0 15750.0 121950.0 16650.0 ;
      RECT  117900.0 15750.0 121500.0 16650.0 ;
      RECT  121050.0 16200.0 121950.0 18000.0 ;
      RECT  131250.0 15750.0 132150.0 16650.0 ;
      RECT  128100.0 15750.0 131700.0 16650.0 ;
      RECT  131250.0 16200.0 132150.0 18000.0 ;
      RECT  53400.0 430200.0 54300.0 432300.0 ;
      RECT  116400.0 209400.0 126600.0 223200.0 ;
      RECT  116400.0 237000.0 126600.0 223200.0 ;
      RECT  116400.0 237000.0 126600.0 250800.0 ;
      RECT  116400.0 264600.0 126600.0 250800.0 ;
      RECT  116400.0 264600.0 126600.0 278400.0 ;
      RECT  116400.0 292200.0 126600.0 278400.0 ;
      RECT  116400.0 292200.0 126600.0 306000.0 ;
      RECT  116400.0 319800.0 126600.0 306000.0 ;
      RECT  116400.0 319800.0 126600.0 333600.0 ;
      RECT  116400.0 347400.0 126600.0 333600.0 ;
      RECT  116400.0 347400.0 126600.0 361200.0 ;
      RECT  116400.0 375000.0 126600.0 361200.0 ;
      RECT  116400.0 375000.0 126600.0 388800.0 ;
      RECT  116400.0 402600.0 126600.0 388800.0 ;
      RECT  116400.0 402600.0 126600.0 416400.0 ;
      RECT  116400.0 430200.0 126600.0 416400.0 ;
      RECT  126600.0 209400.0 136800.0 223200.0 ;
      RECT  126600.0 237000.0 136800.0 223200.0 ;
      RECT  126600.0 237000.0 136800.0 250800.0 ;
      RECT  126600.0 264600.0 136800.0 250800.0 ;
      RECT  126600.0 264600.0 136800.0 278400.0 ;
      RECT  126600.0 292200.0 136800.0 278400.0 ;
      RECT  126600.0 292200.0 136800.0 306000.0 ;
      RECT  126600.0 319800.0 136800.0 306000.0 ;
      RECT  126600.0 319800.0 136800.0 333600.0 ;
      RECT  126600.0 347400.0 136800.0 333600.0 ;
      RECT  126600.0 347400.0 136800.0 361200.0 ;
      RECT  126600.0 375000.0 136800.0 361200.0 ;
      RECT  126600.0 375000.0 136800.0 388800.0 ;
      RECT  126600.0 402600.0 136800.0 388800.0 ;
      RECT  126600.0 402600.0 136800.0 416400.0 ;
      RECT  126600.0 430200.0 136800.0 416400.0 ;
      RECT  119400.0 210000.0 120600.0 433800.0 ;
      RECT  122400.0 208800.0 123600.0 432600.0 ;
      RECT  129600.0 210000.0 130800.0 433800.0 ;
      RECT  132600.0 208800.0 133800.0 432600.0 ;
      RECT  115800.0 208800.0 117000.0 432600.0 ;
      RECT  126000.0 208800.0 127200.0 432600.0 ;
      RECT  136200.0 208800.0 137400.0 432600.0 ;
      RECT  119400.0 436200.0 120600.0 437400.0 ;
      RECT  121800.0 436200.0 123450.0 437400.0 ;
      RECT  119400.0 443400.0 120600.0 444600.0 ;
      RECT  122550.0 443400.0 125400.0 444600.0 ;
      RECT  119400.0 436200.0 120600.0 437400.0 ;
      RECT  121800.0 436200.0 123000.0 437400.0 ;
      RECT  119400.0 443400.0 120600.0 444600.0 ;
      RECT  124200.0 443400.0 125400.0 444600.0 ;
      RECT  119550.0 433800.0 120450.0 450600.0 ;
      RECT  122550.0 433800.0 123450.0 450600.0 ;
      RECT  129600.0 436200.0 130800.0 437400.0 ;
      RECT  132000.0 436200.0 133650.0 437400.0 ;
      RECT  129600.0 443400.0 130800.0 444600.0 ;
      RECT  132750.0 443400.0 135600.0 444600.0 ;
      RECT  129600.0 436200.0 130800.0 437400.0 ;
      RECT  132000.0 436200.0 133200.0 437400.0 ;
      RECT  129600.0 443400.0 130800.0 444600.0 ;
      RECT  134400.0 443400.0 135600.0 444600.0 ;
      RECT  129750.0 433800.0 130650.0 450600.0 ;
      RECT  132750.0 433800.0 133650.0 450600.0 ;
      RECT  119550.0 433800.0 120450.0 450600.0 ;
      RECT  122550.0 433800.0 123450.0 450600.0 ;
      RECT  129750.0 433800.0 130650.0 450600.0 ;
      RECT  132750.0 433800.0 133650.0 450600.0 ;
      RECT  116400.0 160500.0 126600.0 209400.0 ;
      RECT  126600.0 160500.0 136800.0 209400.0 ;
      RECT  119400.0 160500.0 120600.0 173700.0 ;
      RECT  122400.0 160500.0 123600.0 173700.0 ;
      RECT  129600.0 160500.0 130800.0 173700.0 ;
      RECT  132600.0 160500.0 133800.0 173700.0 ;
      RECT  116400.0 99900.0 126600.0 160500.0 ;
      RECT  126600.0 99900.0 136800.0 160500.0 ;
      RECT  120900.0 99900.0 122100.0 102900.0 ;
      RECT  131100.0 99900.0 132300.0 102900.0 ;
      RECT  119400.0 158400.0 120600.0 160500.0 ;
      RECT  122400.0 153000.0 123600.0 160500.0 ;
      RECT  129600.0 158400.0 130800.0 160500.0 ;
      RECT  132600.0 153000.0 133800.0 160500.0 ;
      RECT  116400.0 39900.0 126600.0 99900.0 ;
      RECT  136800.0 39900.0 126600.0 99900.0 ;
      RECT  120900.0 97500.0 123600.0 98700.0 ;
      RECT  118200.0 95400.0 119400.0 99900.0 ;
      RECT  129600.0 97500.0 132300.0 98700.0 ;
      RECT  133800.0 95400.0 135000.0 99900.0 ;
      RECT  126000.0 39900.0 127200.0 99900.0 ;
      RECT  116400.0 39900.0 126600.0 18000.0 ;
      RECT  126600.0 39900.0 136800.0 18000.0 ;
      RECT  120900.0 24900.0 122100.0 18000.0 ;
      RECT  131100.0 24900.0 132300.0 18000.0 ;
      RECT  120900.0 39900.0 122100.0 38400.0 ;
      RECT  131100.0 39900.0 132300.0 38400.0 ;
      RECT  9900.0 99000.0 10800.0 430200.0 ;
      RECT  12000.0 99000.0 12900.0 430200.0 ;
      RECT  14100.0 99000.0 15000.0 430200.0 ;
      RECT  16200.0 99000.0 17100.0 430200.0 ;
      RECT  18300.0 99000.0 19200.0 430200.0 ;
      RECT  20400.0 99000.0 21300.0 430200.0 ;
      RECT  22500.0 99000.0 23400.0 430200.0 ;
      RECT  24600.0 99000.0 25500.0 430200.0 ;
      RECT  56700.0 99000.0 55800.0 152400.0 ;
      RECT  53700.0 99000.0 52800.0 152400.0 ;
      RECT  62700.0 99000.0 61800.0 152400.0 ;
      RECT  59700.0 99000.0 58800.0 152400.0 ;
      RECT  46350.0 106350.0 45450.0 107250.0 ;
      RECT  43950.0 106350.0 43050.0 107250.0 ;
      RECT  46350.0 106800.0 45450.0 109650.0 ;
      RECT  45900.0 106350.0 43500.0 107250.0 ;
      RECT  43950.0 102150.0 43050.0 106800.0 ;
      RECT  46500.0 109650.0 45300.0 110850.0 ;
      RECT  44100.0 100950.0 42900.0 102150.0 ;
      RECT  42900.0 106200.0 44100.0 107400.0 ;
      RECT  46350.0 119250.0 45450.0 118350.0 ;
      RECT  43950.0 119250.0 43050.0 118350.0 ;
      RECT  46350.0 118800.0 45450.0 115950.0 ;
      RECT  45900.0 119250.0 43500.0 118350.0 ;
      RECT  43950.0 123450.0 43050.0 118800.0 ;
      RECT  46500.0 115950.0 45300.0 114750.0 ;
      RECT  44100.0 124650.0 42900.0 123450.0 ;
      RECT  42900.0 119400.0 44100.0 118200.0 ;
      RECT  46350.0 133950.0 45450.0 134850.0 ;
      RECT  43950.0 133950.0 43050.0 134850.0 ;
      RECT  46350.0 134400.0 45450.0 137250.0 ;
      RECT  45900.0 133950.0 43500.0 134850.0 ;
      RECT  43950.0 129750.0 43050.0 134400.0 ;
      RECT  46500.0 137250.0 45300.0 138450.0 ;
      RECT  44100.0 128550.0 42900.0 129750.0 ;
      RECT  42900.0 133800.0 44100.0 135000.0 ;
      RECT  46350.0 146850.0 45450.0 145950.0 ;
      RECT  43950.0 146850.0 43050.0 145950.0 ;
      RECT  46350.0 146400.0 45450.0 143550.0 ;
      RECT  45900.0 146850.0 43500.0 145950.0 ;
      RECT  43950.0 151050.0 43050.0 146400.0 ;
      RECT  46500.0 143550.0 45300.0 142350.0 ;
      RECT  44100.0 152250.0 42900.0 151050.0 ;
      RECT  42900.0 147000.0 44100.0 145800.0 ;
      RECT  61650.0 109500.0 62850.0 110700.0 ;
      RECT  80250.0 105000.0 81450.0 106200.0 ;
      RECT  58650.0 123300.0 59850.0 124500.0 ;
      RECT  77250.0 119400.0 78450.0 120600.0 ;
      RECT  80250.0 128100.0 81450.0 129300.0 ;
      RECT  55650.0 128100.0 56850.0 129300.0 ;
      RECT  77250.0 141900.0 78450.0 143100.0 ;
      RECT  52650.0 141900.0 53850.0 143100.0 ;
      RECT  61650.0 106200.0 62850.0 107400.0 ;
      RECT  58650.0 103500.0 59850.0 104700.0 ;
      RECT  55650.0 118200.0 56850.0 119400.0 ;
      RECT  58650.0 120900.0 59850.0 122100.0 ;
      RECT  61650.0 133800.0 62850.0 135000.0 ;
      RECT  52650.0 131100.0 53850.0 132300.0 ;
      RECT  55650.0 145800.0 56850.0 147000.0 ;
      RECT  52650.0 148500.0 53850.0 149700.0 ;
      RECT  81300.0 99000.0 80400.0 152400.0 ;
      RECT  78300.0 99000.0 77400.0 152400.0 ;
      RECT  56700.0 154200.0 55800.0 207600.0 ;
      RECT  53700.0 154200.0 52800.0 207600.0 ;
      RECT  62700.0 154200.0 61800.0 207600.0 ;
      RECT  59700.0 154200.0 58800.0 207600.0 ;
      RECT  46350.0 161550.0 45450.0 162450.0 ;
      RECT  43950.0 161550.0 43050.0 162450.0 ;
      RECT  46350.0 162000.0 45450.0 164850.0 ;
      RECT  45900.0 161550.0 43500.0 162450.0 ;
      RECT  43950.0 157350.0 43050.0 162000.0 ;
      RECT  46500.0 164850.0 45300.0 166050.0 ;
      RECT  44100.0 156150.0 42900.0 157350.0 ;
      RECT  42900.0 161400.0 44100.0 162600.0 ;
      RECT  46350.0 174450.0 45450.0 173550.0 ;
      RECT  43950.0 174450.0 43050.0 173550.0 ;
      RECT  46350.0 174000.0 45450.0 171150.0 ;
      RECT  45900.0 174450.0 43500.0 173550.0 ;
      RECT  43950.0 178650.0 43050.0 174000.0 ;
      RECT  46500.0 171150.0 45300.0 169950.0 ;
      RECT  44100.0 179850.0 42900.0 178650.0 ;
      RECT  42900.0 174600.0 44100.0 173400.0 ;
      RECT  46350.0 189150.0 45450.0 190050.0 ;
      RECT  43950.0 189150.0 43050.0 190050.0 ;
      RECT  46350.0 189600.0 45450.0 192450.0 ;
      RECT  45900.0 189150.0 43500.0 190050.0 ;
      RECT  43950.0 184950.0 43050.0 189600.0 ;
      RECT  46500.0 192450.0 45300.0 193650.0 ;
      RECT  44100.0 183750.0 42900.0 184950.0 ;
      RECT  42900.0 189000.0 44100.0 190200.0 ;
      RECT  46350.0 202050.0 45450.0 201150.0 ;
      RECT  43950.0 202050.0 43050.0 201150.0 ;
      RECT  46350.0 201600.0 45450.0 198750.0 ;
      RECT  45900.0 202050.0 43500.0 201150.0 ;
      RECT  43950.0 206250.0 43050.0 201600.0 ;
      RECT  46500.0 198750.0 45300.0 197550.0 ;
      RECT  44100.0 207450.0 42900.0 206250.0 ;
      RECT  42900.0 202200.0 44100.0 201000.0 ;
      RECT  61650.0 164700.0 62850.0 165900.0 ;
      RECT  80250.0 160200.0 81450.0 161400.0 ;
      RECT  58650.0 178500.0 59850.0 179700.0 ;
      RECT  77250.0 174600.0 78450.0 175800.0 ;
      RECT  80250.0 183300.0 81450.0 184500.0 ;
      RECT  55650.0 183300.0 56850.0 184500.0 ;
      RECT  77250.0 197100.0 78450.0 198300.0 ;
      RECT  52650.0 197100.0 53850.0 198300.0 ;
      RECT  61650.0 161400.0 62850.0 162600.0 ;
      RECT  58650.0 158700.0 59850.0 159900.0 ;
      RECT  55650.0 173400.0 56850.0 174600.0 ;
      RECT  58650.0 176100.0 59850.0 177300.0 ;
      RECT  61650.0 189000.0 62850.0 190200.0 ;
      RECT  52650.0 186300.0 53850.0 187500.0 ;
      RECT  55650.0 201000.0 56850.0 202200.0 ;
      RECT  52650.0 203700.0 53850.0 204900.0 ;
      RECT  81300.0 154200.0 80400.0 207600.0 ;
      RECT  78300.0 154200.0 77400.0 207600.0 ;
      RECT  31050.0 216750.0 31950.0 217650.0 ;
      RECT  33450.0 216750.0 34350.0 217650.0 ;
      RECT  31050.0 217200.0 31950.0 220050.0 ;
      RECT  31500.0 216750.0 33900.0 217650.0 ;
      RECT  33450.0 212550.0 34350.0 217200.0 ;
      RECT  30900.0 220050.0 32100.0 221250.0 ;
      RECT  33300.0 211350.0 34500.0 212550.0 ;
      RECT  34500.0 216600.0 33300.0 217800.0 ;
      RECT  31050.0 229650.0 31950.0 228750.0 ;
      RECT  33450.0 229650.0 34350.0 228750.0 ;
      RECT  31050.0 229200.0 31950.0 226350.0 ;
      RECT  31500.0 229650.0 33900.0 228750.0 ;
      RECT  33450.0 233850.0 34350.0 229200.0 ;
      RECT  30900.0 226350.0 32100.0 225150.0 ;
      RECT  33300.0 235050.0 34500.0 233850.0 ;
      RECT  34500.0 229800.0 33300.0 228600.0 ;
      RECT  31050.0 244350.0 31950.0 245250.0 ;
      RECT  33450.0 244350.0 34350.0 245250.0 ;
      RECT  31050.0 244800.0 31950.0 247650.0 ;
      RECT  31500.0 244350.0 33900.0 245250.0 ;
      RECT  33450.0 240150.0 34350.0 244800.0 ;
      RECT  30900.0 247650.0 32100.0 248850.0 ;
      RECT  33300.0 238950.0 34500.0 240150.0 ;
      RECT  34500.0 244200.0 33300.0 245400.0 ;
      RECT  31050.0 257250.0 31950.0 256350.0 ;
      RECT  33450.0 257250.0 34350.0 256350.0 ;
      RECT  31050.0 256800.0 31950.0 253950.0 ;
      RECT  31500.0 257250.0 33900.0 256350.0 ;
      RECT  33450.0 261450.0 34350.0 256800.0 ;
      RECT  30900.0 253950.0 32100.0 252750.0 ;
      RECT  33300.0 262650.0 34500.0 261450.0 ;
      RECT  34500.0 257400.0 33300.0 256200.0 ;
      RECT  31050.0 271950.0 31950.0 272850.0 ;
      RECT  33450.0 271950.0 34350.0 272850.0 ;
      RECT  31050.0 272400.0 31950.0 275250.0 ;
      RECT  31500.0 271950.0 33900.0 272850.0 ;
      RECT  33450.0 267750.0 34350.0 272400.0 ;
      RECT  30900.0 275250.0 32100.0 276450.0 ;
      RECT  33300.0 266550.0 34500.0 267750.0 ;
      RECT  34500.0 271800.0 33300.0 273000.0 ;
      RECT  31050.0 284850.0 31950.0 283950.0 ;
      RECT  33450.0 284850.0 34350.0 283950.0 ;
      RECT  31050.0 284400.0 31950.0 281550.0 ;
      RECT  31500.0 284850.0 33900.0 283950.0 ;
      RECT  33450.0 289050.0 34350.0 284400.0 ;
      RECT  30900.0 281550.0 32100.0 280350.0 ;
      RECT  33300.0 290250.0 34500.0 289050.0 ;
      RECT  34500.0 285000.0 33300.0 283800.0 ;
      RECT  31050.0 299550.0 31950.0 300450.0 ;
      RECT  33450.0 299550.0 34350.0 300450.0 ;
      RECT  31050.0 300000.0 31950.0 302850.0 ;
      RECT  31500.0 299550.0 33900.0 300450.0 ;
      RECT  33450.0 295350.0 34350.0 300000.0 ;
      RECT  30900.0 302850.0 32100.0 304050.0 ;
      RECT  33300.0 294150.0 34500.0 295350.0 ;
      RECT  34500.0 299400.0 33300.0 300600.0 ;
      RECT  31050.0 312450.0 31950.0 311550.0 ;
      RECT  33450.0 312450.0 34350.0 311550.0 ;
      RECT  31050.0 312000.0 31950.0 309150.0 ;
      RECT  31500.0 312450.0 33900.0 311550.0 ;
      RECT  33450.0 316650.0 34350.0 312000.0 ;
      RECT  30900.0 309150.0 32100.0 307950.0 ;
      RECT  33300.0 317850.0 34500.0 316650.0 ;
      RECT  34500.0 312600.0 33300.0 311400.0 ;
      RECT  31050.0 327150.0 31950.0 328050.0 ;
      RECT  33450.0 327150.0 34350.0 328050.0 ;
      RECT  31050.0 327600.0 31950.0 330450.0 ;
      RECT  31500.0 327150.0 33900.0 328050.0 ;
      RECT  33450.0 322950.0 34350.0 327600.0 ;
      RECT  30900.0 330450.0 32100.0 331650.0 ;
      RECT  33300.0 321750.0 34500.0 322950.0 ;
      RECT  34500.0 327000.0 33300.0 328200.0 ;
      RECT  31050.0 340050.0 31950.0 339150.0 ;
      RECT  33450.0 340050.0 34350.0 339150.0 ;
      RECT  31050.0 339600.0 31950.0 336750.0 ;
      RECT  31500.0 340050.0 33900.0 339150.0 ;
      RECT  33450.0 344250.0 34350.0 339600.0 ;
      RECT  30900.0 336750.0 32100.0 335550.0 ;
      RECT  33300.0 345450.0 34500.0 344250.0 ;
      RECT  34500.0 340200.0 33300.0 339000.0 ;
      RECT  31050.0 354750.0 31950.0 355650.0 ;
      RECT  33450.0 354750.0 34350.0 355650.0 ;
      RECT  31050.0 355200.0 31950.0 358050.0 ;
      RECT  31500.0 354750.0 33900.0 355650.0 ;
      RECT  33450.0 350550.0 34350.0 355200.0 ;
      RECT  30900.0 358050.0 32100.0 359250.0 ;
      RECT  33300.0 349350.0 34500.0 350550.0 ;
      RECT  34500.0 354600.0 33300.0 355800.0 ;
      RECT  31050.0 367650.0 31950.0 366750.0 ;
      RECT  33450.0 367650.0 34350.0 366750.0 ;
      RECT  31050.0 367200.0 31950.0 364350.0 ;
      RECT  31500.0 367650.0 33900.0 366750.0 ;
      RECT  33450.0 371850.0 34350.0 367200.0 ;
      RECT  30900.0 364350.0 32100.0 363150.0 ;
      RECT  33300.0 373050.0 34500.0 371850.0 ;
      RECT  34500.0 367800.0 33300.0 366600.0 ;
      RECT  31050.0 382350.0 31950.0 383250.0 ;
      RECT  33450.0 382350.0 34350.0 383250.0 ;
      RECT  31050.0 382800.0 31950.0 385650.0 ;
      RECT  31500.0 382350.0 33900.0 383250.0 ;
      RECT  33450.0 378150.0 34350.0 382800.0 ;
      RECT  30900.0 385650.0 32100.0 386850.0 ;
      RECT  33300.0 376950.0 34500.0 378150.0 ;
      RECT  34500.0 382200.0 33300.0 383400.0 ;
      RECT  31050.0 395250.0 31950.0 394350.0 ;
      RECT  33450.0 395250.0 34350.0 394350.0 ;
      RECT  31050.0 394800.0 31950.0 391950.0 ;
      RECT  31500.0 395250.0 33900.0 394350.0 ;
      RECT  33450.0 399450.0 34350.0 394800.0 ;
      RECT  30900.0 391950.0 32100.0 390750.0 ;
      RECT  33300.0 400650.0 34500.0 399450.0 ;
      RECT  34500.0 395400.0 33300.0 394200.0 ;
      RECT  31050.0 409950.0 31950.0 410850.0 ;
      RECT  33450.0 409950.0 34350.0 410850.0 ;
      RECT  31050.0 410400.0 31950.0 413250.0 ;
      RECT  31500.0 409950.0 33900.0 410850.0 ;
      RECT  33450.0 405750.0 34350.0 410400.0 ;
      RECT  30900.0 413250.0 32100.0 414450.0 ;
      RECT  33300.0 404550.0 34500.0 405750.0 ;
      RECT  34500.0 409800.0 33300.0 411000.0 ;
      RECT  31050.0 422850.0 31950.0 421950.0 ;
      RECT  33450.0 422850.0 34350.0 421950.0 ;
      RECT  31050.0 422400.0 31950.0 419550.0 ;
      RECT  31500.0 422850.0 33900.0 421950.0 ;
      RECT  33450.0 427050.0 34350.0 422400.0 ;
      RECT  30900.0 419550.0 32100.0 418350.0 ;
      RECT  33300.0 428250.0 34500.0 427050.0 ;
      RECT  34500.0 423000.0 33300.0 421800.0 ;
      RECT  10950.0 105000.0 9750.0 106200.0 ;
      RECT  13050.0 119400.0 11850.0 120600.0 ;
      RECT  15150.0 132600.0 13950.0 133800.0 ;
      RECT  17250.0 147000.0 16050.0 148200.0 ;
      RECT  19350.0 160200.0 18150.0 161400.0 ;
      RECT  21450.0 174600.0 20250.0 175800.0 ;
      RECT  23550.0 187800.0 22350.0 189000.0 ;
      RECT  25650.0 202200.0 24450.0 203400.0 ;
      RECT  10950.0 216600.0 9750.0 217800.0 ;
      RECT  19350.0 213900.0 18150.0 215100.0 ;
      RECT  10950.0 228600.0 9750.0 229800.0 ;
      RECT  21450.0 231300.0 20250.0 232500.0 ;
      RECT  10950.0 244200.0 9750.0 245400.0 ;
      RECT  23550.0 241500.0 22350.0 242700.0 ;
      RECT  10950.0 256200.0 9750.0 257400.0 ;
      RECT  25650.0 258900.0 24450.0 260100.0 ;
      RECT  13050.0 271800.0 11850.0 273000.0 ;
      RECT  19350.0 269100.0 18150.0 270300.0 ;
      RECT  13050.0 283800.0 11850.0 285000.0 ;
      RECT  21450.0 286500.0 20250.0 287700.0 ;
      RECT  13050.0 299400.0 11850.0 300600.0 ;
      RECT  23550.0 296700.0 22350.0 297900.0 ;
      RECT  13050.0 311400.0 11850.0 312600.0 ;
      RECT  25650.0 314100.0 24450.0 315300.0 ;
      RECT  15150.0 327000.0 13950.0 328200.0 ;
      RECT  19350.0 324300.0 18150.0 325500.0 ;
      RECT  15150.0 339000.0 13950.0 340200.0 ;
      RECT  21450.0 341700.0 20250.0 342900.0 ;
      RECT  15150.0 354600.0 13950.0 355800.0 ;
      RECT  23550.0 351900.0 22350.0 353100.0 ;
      RECT  15150.0 366600.0 13950.0 367800.0 ;
      RECT  25650.0 369300.0 24450.0 370500.0 ;
      RECT  17250.0 382200.0 16050.0 383400.0 ;
      RECT  19350.0 379500.0 18150.0 380700.0 ;
      RECT  17250.0 394200.0 16050.0 395400.0 ;
      RECT  21450.0 396900.0 20250.0 398100.0 ;
      RECT  17250.0 409800.0 16050.0 411000.0 ;
      RECT  23550.0 407100.0 22350.0 408300.0 ;
      RECT  17250.0 421800.0 16050.0 423000.0 ;
      RECT  25650.0 424500.0 24450.0 425700.0 ;
      RECT  80400.0 99000.0 81300.0 152400.0 ;
      RECT  77400.0 99000.0 78300.0 152400.0 ;
      RECT  80400.0 154200.0 81300.0 207600.0 ;
      RECT  77400.0 154200.0 78300.0 207600.0 ;
      RECT  55350.0 214050.0 56250.0 214950.0 ;
      RECT  55350.0 213600.0 56250.0 214500.0 ;
      RECT  55800.0 214050.0 72000.0 214950.0 ;
      RECT  55350.0 231450.0 56250.0 232350.0 ;
      RECT  55350.0 231900.0 56250.0 232800.0 ;
      RECT  55800.0 231450.0 72000.0 232350.0 ;
      RECT  55350.0 241650.0 56250.0 242550.0 ;
      RECT  55350.0 241200.0 56250.0 242100.0 ;
      RECT  55800.0 241650.0 72000.0 242550.0 ;
      RECT  55350.0 259050.0 56250.0 259950.0 ;
      RECT  55350.0 259500.0 56250.0 260400.0 ;
      RECT  55800.0 259050.0 72000.0 259950.0 ;
      RECT  55350.0 269250.0 56250.0 270150.0 ;
      RECT  55350.0 268800.0 56250.0 269700.0 ;
      RECT  55800.0 269250.0 72000.0 270150.0 ;
      RECT  55350.0 286650.0 56250.0 287550.0 ;
      RECT  55350.0 287100.0 56250.0 288000.0 ;
      RECT  55800.0 286650.0 72000.0 287550.0 ;
      RECT  55350.0 296850.0 56250.0 297750.0 ;
      RECT  55350.0 296400.0 56250.0 297300.0 ;
      RECT  55800.0 296850.0 72000.0 297750.0 ;
      RECT  55350.0 314250.0 56250.0 315150.0 ;
      RECT  55350.0 314700.0 56250.0 315600.0 ;
      RECT  55800.0 314250.0 72000.0 315150.0 ;
      RECT  55350.0 324450.0 56250.0 325350.0 ;
      RECT  55350.0 324000.0 56250.0 324900.0 ;
      RECT  55800.0 324450.0 72000.0 325350.0 ;
      RECT  55350.0 341850.0 56250.0 342750.0 ;
      RECT  55350.0 342300.0 56250.0 343200.0 ;
      RECT  55800.0 341850.0 72000.0 342750.0 ;
      RECT  55350.0 352050.0 56250.0 352950.0 ;
      RECT  55350.0 351600.0 56250.0 352500.0 ;
      RECT  55800.0 352050.0 72000.0 352950.0 ;
      RECT  55350.0 369450.0 56250.0 370350.0 ;
      RECT  55350.0 369900.0 56250.0 370800.0 ;
      RECT  55800.0 369450.0 72000.0 370350.0 ;
      RECT  55350.0 379650.0 56250.0 380550.0 ;
      RECT  55350.0 379200.0 56250.0 380100.0 ;
      RECT  55800.0 379650.0 72000.0 380550.0 ;
      RECT  55350.0 397050.0 56250.0 397950.0 ;
      RECT  55350.0 397500.0 56250.0 398400.0 ;
      RECT  55800.0 397050.0 72000.0 397950.0 ;
      RECT  55350.0 407250.0 56250.0 408150.0 ;
      RECT  55350.0 406800.0 56250.0 407700.0 ;
      RECT  55800.0 407250.0 72000.0 408150.0 ;
      RECT  55350.0 424650.0 56250.0 425550.0 ;
      RECT  55350.0 425100.0 56250.0 426000.0 ;
      RECT  55800.0 424650.0 72000.0 425550.0 ;
      RECT  70950.0 216750.0 71850.0 217650.0 ;
      RECT  73350.0 216750.0 74250.0 217650.0 ;
      RECT  70950.0 217200.0 71850.0 220050.0 ;
      RECT  71400.0 216750.0 73800.0 217650.0 ;
      RECT  73350.0 212550.0 74250.0 217200.0 ;
      RECT  70800.0 220050.0 72000.0 221250.0 ;
      RECT  73200.0 211350.0 74400.0 212550.0 ;
      RECT  74400.0 216600.0 73200.0 217800.0 ;
      RECT  53250.0 215400.0 54450.0 216600.0 ;
      RECT  55200.0 213000.0 56400.0 214200.0 ;
      RECT  72000.0 213900.0 70800.0 215100.0 ;
      RECT  70950.0 229650.0 71850.0 228750.0 ;
      RECT  73350.0 229650.0 74250.0 228750.0 ;
      RECT  70950.0 229200.0 71850.0 226350.0 ;
      RECT  71400.0 229650.0 73800.0 228750.0 ;
      RECT  73350.0 233850.0 74250.0 229200.0 ;
      RECT  70800.0 226350.0 72000.0 225150.0 ;
      RECT  73200.0 235050.0 74400.0 233850.0 ;
      RECT  74400.0 229800.0 73200.0 228600.0 ;
      RECT  53250.0 229800.0 54450.0 231000.0 ;
      RECT  55200.0 232200.0 56400.0 233400.0 ;
      RECT  72000.0 231300.0 70800.0 232500.0 ;
      RECT  70950.0 244350.0 71850.0 245250.0 ;
      RECT  73350.0 244350.0 74250.0 245250.0 ;
      RECT  70950.0 244800.0 71850.0 247650.0 ;
      RECT  71400.0 244350.0 73800.0 245250.0 ;
      RECT  73350.0 240150.0 74250.0 244800.0 ;
      RECT  70800.0 247650.0 72000.0 248850.0 ;
      RECT  73200.0 238950.0 74400.0 240150.0 ;
      RECT  74400.0 244200.0 73200.0 245400.0 ;
      RECT  53250.0 243000.0 54450.0 244200.0 ;
      RECT  55200.0 240600.0 56400.0 241800.0 ;
      RECT  72000.0 241500.0 70800.0 242700.0 ;
      RECT  70950.0 257250.0 71850.0 256350.0 ;
      RECT  73350.0 257250.0 74250.0 256350.0 ;
      RECT  70950.0 256800.0 71850.0 253950.0 ;
      RECT  71400.0 257250.0 73800.0 256350.0 ;
      RECT  73350.0 261450.0 74250.0 256800.0 ;
      RECT  70800.0 253950.0 72000.0 252750.0 ;
      RECT  73200.0 262650.0 74400.0 261450.0 ;
      RECT  74400.0 257400.0 73200.0 256200.0 ;
      RECT  53250.0 257400.0 54450.0 258600.0 ;
      RECT  55200.0 259800.0 56400.0 261000.0 ;
      RECT  72000.0 258900.0 70800.0 260100.0 ;
      RECT  70950.0 271950.0 71850.0 272850.0 ;
      RECT  73350.0 271950.0 74250.0 272850.0 ;
      RECT  70950.0 272400.0 71850.0 275250.0 ;
      RECT  71400.0 271950.0 73800.0 272850.0 ;
      RECT  73350.0 267750.0 74250.0 272400.0 ;
      RECT  70800.0 275250.0 72000.0 276450.0 ;
      RECT  73200.0 266550.0 74400.0 267750.0 ;
      RECT  74400.0 271800.0 73200.0 273000.0 ;
      RECT  53250.0 270600.0 54450.0 271800.0 ;
      RECT  55200.0 268200.0 56400.0 269400.0 ;
      RECT  72000.0 269100.0 70800.0 270300.0 ;
      RECT  70950.0 284850.0 71850.0 283950.0 ;
      RECT  73350.0 284850.0 74250.0 283950.0 ;
      RECT  70950.0 284400.0 71850.0 281550.0 ;
      RECT  71400.0 284850.0 73800.0 283950.0 ;
      RECT  73350.0 289050.0 74250.0 284400.0 ;
      RECT  70800.0 281550.0 72000.0 280350.0 ;
      RECT  73200.0 290250.0 74400.0 289050.0 ;
      RECT  74400.0 285000.0 73200.0 283800.0 ;
      RECT  53250.0 285000.0 54450.0 286200.0 ;
      RECT  55200.0 287400.0 56400.0 288600.0 ;
      RECT  72000.0 286500.0 70800.0 287700.0 ;
      RECT  70950.0 299550.0 71850.0 300450.0 ;
      RECT  73350.0 299550.0 74250.0 300450.0 ;
      RECT  70950.0 300000.0 71850.0 302850.0 ;
      RECT  71400.0 299550.0 73800.0 300450.0 ;
      RECT  73350.0 295350.0 74250.0 300000.0 ;
      RECT  70800.0 302850.0 72000.0 304050.0 ;
      RECT  73200.0 294150.0 74400.0 295350.0 ;
      RECT  74400.0 299400.0 73200.0 300600.0 ;
      RECT  53250.0 298200.0 54450.0 299400.0 ;
      RECT  55200.0 295800.0 56400.0 297000.0 ;
      RECT  72000.0 296700.0 70800.0 297900.0 ;
      RECT  70950.0 312450.0 71850.0 311550.0 ;
      RECT  73350.0 312450.0 74250.0 311550.0 ;
      RECT  70950.0 312000.0 71850.0 309150.0 ;
      RECT  71400.0 312450.0 73800.0 311550.0 ;
      RECT  73350.0 316650.0 74250.0 312000.0 ;
      RECT  70800.0 309150.0 72000.0 307950.0 ;
      RECT  73200.0 317850.0 74400.0 316650.0 ;
      RECT  74400.0 312600.0 73200.0 311400.0 ;
      RECT  53250.0 312600.0 54450.0 313800.0 ;
      RECT  55200.0 315000.0 56400.0 316200.0 ;
      RECT  72000.0 314100.0 70800.0 315300.0 ;
      RECT  70950.0 327150.0 71850.0 328050.0 ;
      RECT  73350.0 327150.0 74250.0 328050.0 ;
      RECT  70950.0 327600.0 71850.0 330450.0 ;
      RECT  71400.0 327150.0 73800.0 328050.0 ;
      RECT  73350.0 322950.0 74250.0 327600.0 ;
      RECT  70800.0 330450.0 72000.0 331650.0 ;
      RECT  73200.0 321750.0 74400.0 322950.0 ;
      RECT  74400.0 327000.0 73200.0 328200.0 ;
      RECT  53250.0 325800.0 54450.0 327000.0 ;
      RECT  55200.0 323400.0 56400.0 324600.0 ;
      RECT  72000.0 324300.0 70800.0 325500.0 ;
      RECT  70950.0 340050.0 71850.0 339150.0 ;
      RECT  73350.0 340050.0 74250.0 339150.0 ;
      RECT  70950.0 339600.0 71850.0 336750.0 ;
      RECT  71400.0 340050.0 73800.0 339150.0 ;
      RECT  73350.0 344250.0 74250.0 339600.0 ;
      RECT  70800.0 336750.0 72000.0 335550.0 ;
      RECT  73200.0 345450.0 74400.0 344250.0 ;
      RECT  74400.0 340200.0 73200.0 339000.0 ;
      RECT  53250.0 340200.0 54450.0 341400.0 ;
      RECT  55200.0 342600.0 56400.0 343800.0 ;
      RECT  72000.0 341700.0 70800.0 342900.0 ;
      RECT  70950.0 354750.0 71850.0 355650.0 ;
      RECT  73350.0 354750.0 74250.0 355650.0 ;
      RECT  70950.0 355200.0 71850.0 358050.0 ;
      RECT  71400.0 354750.0 73800.0 355650.0 ;
      RECT  73350.0 350550.0 74250.0 355200.0 ;
      RECT  70800.0 358050.0 72000.0 359250.0 ;
      RECT  73200.0 349350.0 74400.0 350550.0 ;
      RECT  74400.0 354600.0 73200.0 355800.0 ;
      RECT  53250.0 353400.0 54450.0 354600.0 ;
      RECT  55200.0 351000.0 56400.0 352200.0 ;
      RECT  72000.0 351900.0 70800.0 353100.0 ;
      RECT  70950.0 367650.0 71850.0 366750.0 ;
      RECT  73350.0 367650.0 74250.0 366750.0 ;
      RECT  70950.0 367200.0 71850.0 364350.0 ;
      RECT  71400.0 367650.0 73800.0 366750.0 ;
      RECT  73350.0 371850.0 74250.0 367200.0 ;
      RECT  70800.0 364350.0 72000.0 363150.0 ;
      RECT  73200.0 373050.0 74400.0 371850.0 ;
      RECT  74400.0 367800.0 73200.0 366600.0 ;
      RECT  53250.0 367800.0 54450.0 369000.0 ;
      RECT  55200.0 370200.0 56400.0 371400.0 ;
      RECT  72000.0 369300.0 70800.0 370500.0 ;
      RECT  70950.0 382350.0 71850.0 383250.0 ;
      RECT  73350.0 382350.0 74250.0 383250.0 ;
      RECT  70950.0 382800.0 71850.0 385650.0 ;
      RECT  71400.0 382350.0 73800.0 383250.0 ;
      RECT  73350.0 378150.0 74250.0 382800.0 ;
      RECT  70800.0 385650.0 72000.0 386850.0 ;
      RECT  73200.0 376950.0 74400.0 378150.0 ;
      RECT  74400.0 382200.0 73200.0 383400.0 ;
      RECT  53250.0 381000.0 54450.0 382200.0 ;
      RECT  55200.0 378600.0 56400.0 379800.0 ;
      RECT  72000.0 379500.0 70800.0 380700.0 ;
      RECT  70950.0 395250.0 71850.0 394350.0 ;
      RECT  73350.0 395250.0 74250.0 394350.0 ;
      RECT  70950.0 394800.0 71850.0 391950.0 ;
      RECT  71400.0 395250.0 73800.0 394350.0 ;
      RECT  73350.0 399450.0 74250.0 394800.0 ;
      RECT  70800.0 391950.0 72000.0 390750.0 ;
      RECT  73200.0 400650.0 74400.0 399450.0 ;
      RECT  74400.0 395400.0 73200.0 394200.0 ;
      RECT  53250.0 395400.0 54450.0 396600.0 ;
      RECT  55200.0 397800.0 56400.0 399000.0 ;
      RECT  72000.0 396900.0 70800.0 398100.0 ;
      RECT  70950.0 409950.0 71850.0 410850.0 ;
      RECT  73350.0 409950.0 74250.0 410850.0 ;
      RECT  70950.0 410400.0 71850.0 413250.0 ;
      RECT  71400.0 409950.0 73800.0 410850.0 ;
      RECT  73350.0 405750.0 74250.0 410400.0 ;
      RECT  70800.0 413250.0 72000.0 414450.0 ;
      RECT  73200.0 404550.0 74400.0 405750.0 ;
      RECT  74400.0 409800.0 73200.0 411000.0 ;
      RECT  53250.0 408600.0 54450.0 409800.0 ;
      RECT  55200.0 406200.0 56400.0 407400.0 ;
      RECT  72000.0 407100.0 70800.0 408300.0 ;
      RECT  70950.0 422850.0 71850.0 421950.0 ;
      RECT  73350.0 422850.0 74250.0 421950.0 ;
      RECT  70950.0 422400.0 71850.0 419550.0 ;
      RECT  71400.0 422850.0 73800.0 421950.0 ;
      RECT  73350.0 427050.0 74250.0 422400.0 ;
      RECT  70800.0 419550.0 72000.0 418350.0 ;
      RECT  73200.0 428250.0 74400.0 427050.0 ;
      RECT  74400.0 423000.0 73200.0 421800.0 ;
      RECT  53250.0 423000.0 54450.0 424200.0 ;
      RECT  55200.0 425400.0 56400.0 426600.0 ;
      RECT  72000.0 424500.0 70800.0 425700.0 ;
      RECT  53400.0 209400.0 54300.0 430200.0 ;
      RECT  9900.0 93600.0 69900.0 83400.0 ;
      RECT  9900.0 73200.0 69900.0 83400.0 ;
      RECT  9900.0 73200.0 69900.0 63000.0 ;
      RECT  9900.0 52800.0 69900.0 63000.0 ;
      RECT  67500.0 89100.0 68700.0 86400.0 ;
      RECT  65400.0 91800.0 69900.0 90600.0 ;
      RECT  67500.0 80400.0 68700.0 77700.0 ;
      RECT  65400.0 76200.0 69900.0 75000.0 ;
      RECT  67500.0 68700.0 68700.0 66000.0 ;
      RECT  65400.0 71400.0 69900.0 70200.0 ;
      RECT  67500.0 60000.0 68700.0 57300.0 ;
      RECT  65400.0 55800.0 69900.0 54600.0 ;
      RECT  9900.0 84000.0 69900.0 82800.0 ;
      RECT  9900.0 63600.0 69900.0 62400.0 ;
      RECT  0.0 0.0 3600.0 3600.0 ;
      RECT  0.0 453300.0 3600.0 456900.0 ;
      RECT  139500.0 0.0 143100.0 3600.0 ;
      RECT  139500.0 453300.0 143100.0 456900.0 ;
      RECT  4950.0 4950.0 8550.0 8550.0 ;
      RECT  4950.0 458250.0 8550.0 461850.0 ;
      RECT  144450.0 4950.0 148050.0 8550.0 ;
      RECT  144450.0 458250.0 148050.0 461850.0 ;
      RECT  117450.0 15750.0 118650.0 16950.0 ;
      RECT  127650.0 15750.0 128850.0 16950.0 ;
      RECT  121200.0 300.0 122400.0 1500.0 ;
      RECT  131400.0 300.0 132600.0 1500.0 ;
      RECT  81300.0 101250.0 80100.0 102450.0 ;
      RECT  86400.0 101100.0 85200.0 102300.0 ;
      RECT  78300.0 115050.0 77100.0 116250.0 ;
      RECT  89100.0 114900.0 87900.0 116100.0 ;
      RECT  81300.0 156450.0 80100.0 157650.0 ;
      RECT  91800.0 156300.0 90600.0 157500.0 ;
      RECT  78300.0 170250.0 77100.0 171450.0 ;
      RECT  94500.0 170100.0 93300.0 171300.0 ;
      RECT  3600.0 98400.0 -5.3290705182e-12 99600.0 ;
      RECT  3600.0 126000.0 -5.3290705182e-12 127200.0 ;
      RECT  3600.0 153600.0 -5.3290705182e-12 154800.0 ;
      RECT  3600.0 181200.0 -5.3290705182e-12 182400.0 ;
      RECT  8550.0 112200.0 4950.0 113400.0 ;
      RECT  8550.0 139800.0 4950.0 141000.0 ;
      RECT  8550.0 167400.0 4950.0 168600.0 ;
      RECT  8550.0 195000.0 4950.0 196200.0 ;
      RECT  69300.0 87150.0 68100.0 88350.0 ;
      RECT  86400.0 87150.0 85200.0 88350.0 ;
      RECT  69300.0 78450.0 68100.0 79650.0 ;
      RECT  89100.0 78450.0 87900.0 79650.0 ;
      RECT  69300.0 66750.0 68100.0 67950.0 ;
      RECT  91800.0 66750.0 90600.0 67950.0 ;
      RECT  69300.0 58050.0 68100.0 59250.0 ;
      RECT  94500.0 58050.0 93300.0 59250.0 ;
      RECT  11100.0 82800.0 9900.0 84000.0 ;
      RECT  3600.0 82800.0 -5.3290705182e-12 84000.0 ;
      RECT  11100.0 62400.0 9900.0 63600.0 ;
      RECT  3600.0 62400.0 -5.3290705182e-12 63600.0 ;
      RECT  8550.0 50100.0 4950.0 51300.0 ;
      RECT  105300.0 42150.0 104100.0 43350.0 ;
      RECT  99900.0 37650.0 98700.0 38850.0 ;
      RECT  102600.0 35250.0 101400.0 36450.0 ;
      RECT  105300.0 438450.0 104100.0 439650.0 ;
      RECT  108000.0 106950.0 106800.0 108150.0 ;
      RECT  110700.0 205050.0 109500.0 206250.0 ;
      RECT  97200.0 95100.0 96000.0 96300.0 ;
      RECT  54450.0 431700.0 53250.0 432900.0 ;
      RECT  97200.0 431700.0 96000.0 432900.0 ;
      RECT  148050.0 449550.0 144450.0 450750.0 ;
      RECT  148050.0 177750.0 144450.0 178950.0 ;
      RECT  148050.0 109050.0 144450.0 110250.0 ;
      RECT  148050.0 96150.0 144450.0 97350.0 ;
      RECT  148050.0 19350.0 144450.0 20550.0 ;
      RECT  8550.0 222600.0 4950.0 223800.0 ;
      RECT  148050.0 222600.0 144450.0 223800.0 ;
      RECT  8550.0 250200.0 4950.0 251400.0 ;
      RECT  148050.0 250200.0 144450.0 251400.0 ;
      RECT  8550.0 277800.0 4950.0 279000.0 ;
      RECT  148050.0 277800.0 144450.0 279000.0 ;
      RECT  8550.0 305400.0 4950.0 306600.0 ;
      RECT  148050.0 305400.0 144450.0 306600.0 ;
      RECT  8550.0 333000.0 4950.0 334200.0 ;
      RECT  148050.0 333000.0 144450.0 334200.0 ;
      RECT  8550.0 360600.0 4950.0 361800.0 ;
      RECT  148050.0 360600.0 144450.0 361800.0 ;
      RECT  8550.0 388200.0 4950.0 389400.0 ;
      RECT  148050.0 388200.0 144450.0 389400.0 ;
      RECT  8550.0 415800.0 4950.0 417000.0 ;
      RECT  148050.0 415800.0 144450.0 417000.0 ;
      RECT  143100.0 33150.0 139500.0 34350.0 ;
      RECT  143100.0 202950.0 139500.0 204150.0 ;
      RECT  143100.0 104850.0 139500.0 106050.0 ;
      RECT  3600.0 208800.0 -5.3290705182e-12 210000.0 ;
      RECT  3600.0 236400.0 -5.3290705182e-12 237600.0 ;
      RECT  3600.0 264000.0 -5.3290705182e-12 265200.0 ;
      RECT  3600.0 291600.0 -5.3290705182e-12 292800.0 ;
      RECT  3600.0 319200.0 -5.3290705182e-12 320400.0 ;
      RECT  3600.0 346800.0 -5.3290705182e-12 348000.0 ;
      RECT  3600.0 374400.0 -5.3290705182e-12 375600.0 ;
      RECT  3600.0 402000.0 -5.3290705182e-12 403200.0 ;
      RECT  3600.0 429600.0 -5.3290705182e-12 430800.0 ;
      RECT  120900.0 0.0 121800.0 1800.0 ;
      RECT  131100.0 0.0 132000.0 1800.0 ;
      RECT  109650.0 0.0 110550.0 461850.0 ;
      RECT  106950.0 0.0 107850.0 461850.0 ;
      RECT  98850.0 0.0 99750.0 461850.0 ;
      RECT  101550.0 0.0 102450.0 461850.0 ;
      RECT  104250.0 0.0 105150.0 461850.0 ;
      RECT  96150.0 0.0 97050.0 461850.0 ;
      RECT  4950.0 0.0 8550.0 461850.0 ;
      RECT  144450.0 0.0 148050.0 461850.0 ;
      RECT  0.0 0.0 3600.0 461850.0 ;
      RECT  139500.0 0.0 143100.0 461850.0 ;
      RECT  -3000.0 269400.0 -52800.0 270300.0 ;
      RECT  -3000.0 272100.0 -52800.0 273000.0 ;
      RECT  -3000.0 274800.0 -52800.0 275700.0 ;
      RECT  -3000.0 280200.0 -52800.0 281100.0 ;
      RECT  -9450.0 223050.0 -16800.0 223950.0 ;
      RECT  -19050.0 184650.0 -19950.0 264450.0 ;
      RECT  -3000.0 266700.0 -5700.0 267600.0 ;
      RECT  -14100.0 277500.0 -16800.0 278400.0 ;
      RECT  -27900.0 266700.0 -30600.0 267600.0 ;
      RECT  -41700.0 277500.0 -44400.0 278400.0 ;
      RECT  -52800.0 181800.0 -42600.0 241800.0 ;
      RECT  -32400.0 181800.0 -42600.0 241800.0 ;
      RECT  -32400.0 181800.0 -22200.0 241800.0 ;
      RECT  -48300.0 239400.0 -45600.0 240600.0 ;
      RECT  -51000.0 237300.0 -49800.0 241800.0 ;
      RECT  -39600.0 239400.0 -36900.0 240600.0 ;
      RECT  -35400.0 237300.0 -34200.0 241800.0 ;
      RECT  -27900.0 239400.0 -25200.0 240600.0 ;
      RECT  -30600.0 237300.0 -29400.0 241800.0 ;
      RECT  -43200.0 181800.0 -42000.0 241800.0 ;
      RECT  -22800.0 181800.0 -21600.0 241800.0 ;
      RECT  -6150.0 297450.0 -13650.0 298350.0 ;
      RECT  -11100.0 292650.0 -12000.0 293550.0 ;
      RECT  -11100.0 297450.0 -12000.0 298350.0 ;
      RECT  -11550.0 292650.0 -13650.0 293550.0 ;
      RECT  -11100.0 293100.0 -12000.0 297900.0 ;
      RECT  -6150.0 297450.0 -11550.0 298350.0 ;
      RECT  -13650.0 292500.0 -14850.0 293700.0 ;
      RECT  -13650.0 297300.0 -14850.0 298500.0 ;
      RECT  -4950.0 297300.0 -6150.0 298500.0 ;
      RECT  -10950.0 297300.0 -12150.0 298500.0 ;
      RECT  -24000.0 295050.0 -23100.0 295950.0 ;
      RECT  -23550.0 295050.0 -20550.0 295950.0 ;
      RECT  -24000.0 295500.0 -23100.0 296400.0 ;
      RECT  -29100.0 295050.0 -28200.0 295950.0 ;
      RECT  -29100.0 293700.0 -28200.0 295500.0 ;
      RECT  -28650.0 295050.0 -23550.0 295950.0 ;
      RECT  -20550.0 294900.0 -19350.0 296100.0 ;
      RECT  -29250.0 293700.0 -28050.0 292500.0 ;
      RECT  -24150.0 297000.0 -22950.0 295800.0 ;
      RECT  -23250.0 309750.0 -22350.0 310650.0 ;
      RECT  -23250.0 312150.0 -22350.0 313050.0 ;
      RECT  -22800.0 309750.0 -19950.0 310650.0 ;
      RECT  -23250.0 310200.0 -22350.0 312600.0 ;
      RECT  -27450.0 312150.0 -22800.0 313050.0 ;
      RECT  -19950.0 309600.0 -18750.0 310800.0 ;
      RECT  -28650.0 312000.0 -27450.0 313200.0 ;
      RECT  -23400.0 313200.0 -22200.0 312000.0 ;
      RECT  -33750.0 307050.0 -41250.0 307950.0 ;
      RECT  -38700.0 302250.0 -39600.0 303150.0 ;
      RECT  -38700.0 307050.0 -39600.0 307950.0 ;
      RECT  -39150.0 302250.0 -41250.0 303150.0 ;
      RECT  -38700.0 302700.0 -39600.0 307500.0 ;
      RECT  -33750.0 307050.0 -39150.0 307950.0 ;
      RECT  -41250.0 302100.0 -42450.0 303300.0 ;
      RECT  -41250.0 306900.0 -42450.0 308100.0 ;
      RECT  -32550.0 306900.0 -33750.0 308100.0 ;
      RECT  -38550.0 306900.0 -39750.0 308100.0 ;
      RECT  -49800.0 242400.0 -51000.0 241200.0 ;
      RECT  -49800.0 281250.0 -51000.0 280050.0 ;
      RECT  -46350.0 241200.0 -47550.0 240000.0 ;
      RECT  -46350.0 270450.0 -47550.0 269250.0 ;
      RECT  -34200.0 242400.0 -35400.0 241200.0 ;
      RECT  -34200.0 273150.0 -35400.0 271950.0 ;
      RECT  -29400.0 242400.0 -30600.0 241200.0 ;
      RECT  -29400.0 275850.0 -30600.0 274650.0 ;
      RECT  -42000.0 242400.0 -43200.0 241200.0 ;
      RECT  -42000.0 267750.0 -43200.0 266550.0 ;
      RECT  -21600.0 242400.0 -22800.0 241200.0 ;
      RECT  -21600.0 267750.0 -22800.0 266550.0 ;
      RECT  -30150.0 351300.0 -31050.0 437100.0 ;
      RECT  -35550.0 351300.0 -36450.0 432300.0 ;
      RECT  -45750.0 351300.0 -46650.0 432300.0 ;
      RECT  -32400.0 355500.0 -33300.0 363600.0 ;
      RECT  -39150.0 355500.0 -40050.0 360300.0 ;
      RECT  -10050.0 395100.0 -9150.0 402300.0 ;
      RECT  -10050.0 402300.0 -9150.0 411900.0 ;
      RECT  -10050.0 411900.0 -9150.0 421500.0 ;
      RECT  -10050.0 423900.0 -9150.0 431100.0 ;
      RECT  -10050.0 431100.0 -9150.0 440700.0 ;
      RECT  -10050.0 440700.0 -9150.0 450300.0 ;
      RECT  -17250.0 452250.0 -16350.0 453150.0 ;
      RECT  -17250.0 443850.0 -16350.0 444750.0 ;
      RECT  -16800.0 452250.0 -9600.0 453150.0 ;
      RECT  -17250.0 444300.0 -16350.0 452700.0 ;
      RECT  -24000.0 443850.0 -16800.0 444750.0 ;
      RECT  -24450.0 434700.0 -23550.0 444300.0 ;
      RECT  -24450.0 425100.0 -23550.0 434700.0 ;
      RECT  -24450.0 415500.0 -23550.0 422700.0 ;
      RECT  -24450.0 405900.0 -23550.0 415500.0 ;
      RECT  -24450.0 396300.0 -23550.0 405900.0 ;
      RECT  -10200.0 401700.0 -9000.0 402900.0 ;
      RECT  -10200.0 411300.0 -9000.0 412500.0 ;
      RECT  -10200.0 420900.0 -9000.0 422100.0 ;
      RECT  -10200.0 430500.0 -9000.0 431700.0 ;
      RECT  -10200.0 440100.0 -9000.0 441300.0 ;
      RECT  -10200.0 449700.0 -9000.0 450900.0 ;
      RECT  -24600.0 443700.0 -23400.0 444900.0 ;
      RECT  -24600.0 434100.0 -23400.0 435300.0 ;
      RECT  -24600.0 424500.0 -23400.0 425700.0 ;
      RECT  -24600.0 414900.0 -23400.0 416100.0 ;
      RECT  -24600.0 405300.0 -23400.0 406500.0 ;
      RECT  -24600.0 395700.0 -23400.0 396900.0 ;
      RECT  -10200.0 394500.0 -9000.0 395700.0 ;
      RECT  -10200.0 423300.0 -9000.0 424500.0 ;
      RECT  -10200.0 452100.0 -9000.0 453300.0 ;
      RECT  -24600.0 422100.0 -23400.0 423300.0 ;
      RECT  -36000.0 374700.0 -46200.0 360900.0 ;
      RECT  -36000.0 374700.0 -46200.0 388500.0 ;
      RECT  -36000.0 402300.0 -46200.0 388500.0 ;
      RECT  -36000.0 402300.0 -46200.0 416100.0 ;
      RECT  -36000.0 429900.0 -46200.0 416100.0 ;
      RECT  -39000.0 375300.0 -40200.0 433500.0 ;
      RECT  -42000.0 374100.0 -43200.0 432300.0 ;
      RECT  -35400.0 374100.0 -36600.0 432300.0 ;
      RECT  -45600.0 374100.0 -46800.0 432300.0 ;
      RECT  -30450.0 376200.0 -31650.0 377400.0 ;
      RECT  -30450.0 399600.0 -31650.0 400800.0 ;
      RECT  -30450.0 403800.0 -31650.0 405000.0 ;
      RECT  -30450.0 427200.0 -31650.0 428400.0 ;
      RECT  -30600.0 389700.0 -31800.0 390900.0 ;
      RECT  -30000.0 350100.0 -31200.0 351300.0 ;
      RECT  -36600.0 350700.0 -35400.0 351900.0 ;
      RECT  -46800.0 350700.0 -45600.0 351900.0 ;
      RECT  -33450.0 363000.0 -32250.0 364200.0 ;
      RECT  -33450.0 354900.0 -32250.0 356100.0 ;
      RECT  -40200.0 354900.0 -39000.0 356100.0 ;
      RECT  -8850.0 265050.0 -10050.0 263850.0 ;
      RECT  -8850.0 224100.0 -10050.0 222900.0 ;
      RECT  -16200.0 224100.0 -17400.0 222900.0 ;
      RECT  -16200.0 283950.0 -17400.0 282750.0 ;
      RECT  -18900.0 185250.0 -20100.0 184050.0 ;
      RECT  -22950.0 265050.0 -24150.0 263850.0 ;
      RECT  -25650.0 270450.0 -26850.0 269250.0 ;
      RECT  -22200.0 307800.0 -23400.0 306600.0 ;
      RECT  -22200.0 307800.0 -23400.0 306600.0 ;
      RECT  -22200.0 283950.0 -23400.0 282750.0 ;
      RECT  -24900.0 310800.0 -26100.0 309600.0 ;
      RECT  -24900.0 310800.0 -26100.0 309600.0 ;
      RECT  -24900.0 281250.0 -26100.0 280050.0 ;
      RECT  -10950.0 283950.0 -12150.0 282750.0 ;
      RECT  -9000.0 281250.0 -10200.0 280050.0 ;
      RECT  -7050.0 273150.0 -8250.0 271950.0 ;
      RECT  -38550.0 283950.0 -39750.0 282750.0 ;
      RECT  -36600.0 273150.0 -37800.0 271950.0 ;
      RECT  -34650.0 275850.0 -35850.0 274650.0 ;
      RECT  -22950.0 302100.0 -24150.0 303300.0 ;
      RECT  -22200.0 319200.0 -23400.0 320400.0 ;
      RECT  -36600.0 341700.0 -37800.0 342900.0 ;
      RECT  -23400.0 321900.0 -24600.0 323100.0 ;
      RECT  -2400.0 267750.0 -3600.0 266550.0 ;
      RECT  -16200.0 278550.0 -17400.0 277350.0 ;
      RECT  -30000.0 267750.0 -31200.0 266550.0 ;
      RECT  -43800.0 278550.0 -45000.0 277350.0 ;
      RECT  -3000.0 322050.0 -24000.0 322950.0 ;
      RECT  -3000.0 341850.0 -37200.0 342750.0 ;
      RECT  -3000.0 302250.0 -23550.0 303150.0 ;
      RECT  -3000.0 319350.0 -22800.0 320250.0 ;
      RECT  -3000.0 282900.0 -52800.0 283800.0 ;
      RECT  -3000.0 264000.0 -52800.0 264900.0 ;
      RECT  -3000.0 277500.0 -52800.0 278400.0 ;
      RECT  -3000.0 266700.0 -52800.0 267600.0 ;
      RECT  110700.0 321900.0 109500.0 323100.0 ;
      RECT  -3300.0 322050.0 -4500.0 323250.0 ;
      RECT  108000.0 341700.0 106800.0 342900.0 ;
      RECT  -3300.0 341850.0 -4500.0 343050.0 ;
      RECT  102600.0 302100.0 101400.0 303300.0 ;
      RECT  -3300.0 302250.0 -4500.0 303450.0 ;
      RECT  99900.0 319200.0 98700.0 320400.0 ;
      RECT  -3300.0 319350.0 -4500.0 320550.0 ;
      RECT  105300.0 282750.0 104100.0 283950.0 ;
      RECT  -3300.0 282900.0 -4500.0 284100.0 ;
      RECT  97200.0 263850.0 96000.0 265050.0 ;
      RECT  -3300.0 264000.0 -4500.0 265200.0 ;
      RECT  7350.0 277350.0 6150.0 278550.0 ;
      RECT  -3300.0 277500.0 -4500.0 278700.0 ;
   LAYER  metal3 ;
      RECT  -3000.0 321750.0 110100.0 323250.0 ;
      RECT  -3000.0 341550.0 107400.0 343050.0 ;
      RECT  -3000.0 301950.0 102000.0 303450.0 ;
      RECT  -3000.0 319050.0 99300.0 320550.0 ;
      RECT  -3000.0 282600.0 104700.0 284100.0 ;
      RECT  -3000.0 263700.0 96600.0 265200.0 ;
      RECT  -3000.0 277200.0 6750.0 278700.0 ;
      RECT  117150.0 16200.0 118650.0 161400.0 ;
      RECT  127350.0 16200.0 128850.0 161400.0 ;
      RECT  120900.0 0.0 122400.0 39900.0 ;
      RECT  131100.0 0.0 132600.0 39900.0 ;
      RECT  117000.0 161400.0 118800.0 163200.0 ;
      RECT  127200.0 161400.0 129000.0 163200.0 ;
      RECT  120600.0 40800.0 122400.0 42600.0 ;
      RECT  130800.0 40800.0 132600.0 42600.0 ;
      RECT  10800.0 89400.0 12600.0 87600.0 ;
      RECT  10800.0 79200.0 12600.0 77400.0 ;
      RECT  10800.0 69000.0 12600.0 67200.0 ;
      RECT  10800.0 58800.0 12600.0 57000.0 ;
      RECT  117150.0 15450.0 118950.0 17250.0 ;
      RECT  127350.0 15450.0 129150.0 17250.0 ;
      RECT  120900.0 0.0 122700.0 1800.0 ;
      RECT  131100.0 0.0 132900.0 1800.0 ;
      RECT  0.0 87600.0 10800.0 89100.0 ;
      RECT  0.0 77400.0 10800.0 78900.0 ;
      RECT  0.0 67200.0 10800.0 68700.0 ;
      RECT  0.0 57000.0 10800.0 58500.0 ;
      RECT  -49650.0 241800.0 -51150.0 280650.0 ;
      RECT  -46200.0 240600.0 -47700.0 269850.0 ;
      RECT  -34050.0 241800.0 -35550.0 272550.0 ;
      RECT  -29250.0 241800.0 -30750.0 275250.0 ;
      RECT  -41850.0 241800.0 -43350.0 267150.0 ;
      RECT  -21450.0 241800.0 -22950.0 267150.0 ;
      RECT  -16050.0 223500.0 -17550.0 283350.0 ;
      RECT  -22050.0 283350.0 -23550.0 307200.0 ;
      RECT  -24750.0 280650.0 -26250.0 310200.0 ;
      RECT  -48600.0 182700.0 -46800.0 184500.0 ;
      RECT  -38400.0 182700.0 -36600.0 184500.0 ;
      RECT  -28200.0 182700.0 -26400.0 184500.0 ;
      RECT  -49500.0 242700.0 -51300.0 240900.0 ;
      RECT  -49500.0 281550.0 -51300.0 279750.0 ;
      RECT  -46050.0 241500.0 -47850.0 239700.0 ;
      RECT  -46050.0 270750.0 -47850.0 268950.0 ;
      RECT  -33900.0 242700.0 -35700.0 240900.0 ;
      RECT  -33900.0 273450.0 -35700.0 271650.0 ;
      RECT  -29100.0 242700.0 -30900.0 240900.0 ;
      RECT  -29100.0 276150.0 -30900.0 274350.0 ;
      RECT  -41700.0 242700.0 -43500.0 240900.0 ;
      RECT  -41700.0 268050.0 -43500.0 266250.0 ;
      RECT  -21300.0 242700.0 -23100.0 240900.0 ;
      RECT  -21300.0 268050.0 -23100.0 266250.0 ;
      RECT  -15900.0 224400.0 -17700.0 222600.0 ;
      RECT  -15900.0 284250.0 -17700.0 282450.0 ;
      RECT  -21900.0 308100.0 -23700.0 306300.0 ;
      RECT  -21900.0 284250.0 -23700.0 282450.0 ;
      RECT  -24600.0 311100.0 -26400.0 309300.0 ;
      RECT  -24600.0 281550.0 -26400.0 279750.0 ;
      RECT  -36600.0 182700.0 -38400.0 184500.0 ;
      RECT  -26400.0 182700.0 -28200.0 184500.0 ;
      RECT  -46800.0 182700.0 -48600.0 184500.0 ;
      RECT  111000.0 321600.0 109200.0 323400.0 ;
      RECT  -3000.0 321750.0 -4800.0 323550.0 ;
      RECT  108300.0 341400.0 106500.0 343200.0 ;
      RECT  -3000.0 341550.0 -4800.0 343350.0 ;
      RECT  102900.0 301800.0 101100.0 303600.0 ;
      RECT  -3000.0 301950.0 -4800.0 303750.0 ;
      RECT  100200.0 318900.0 98400.0 320700.0 ;
      RECT  -3000.0 319050.0 -4800.0 320850.0 ;
      RECT  105600.0 282450.0 103800.0 284250.0 ;
      RECT  -3000.0 282600.0 -4800.0 284400.0 ;
      RECT  97500.0 263550.0 95700.0 265350.0 ;
      RECT  -3000.0 263700.0 -4800.0 265500.0 ;
      RECT  7650.0 277050.0 5850.0 278850.0 ;
      RECT  -3000.0 277200.0 -4800.0 279000.0 ;
   END
   END    sram_2_16_1_scn3me_subm
END    LIBRARY
