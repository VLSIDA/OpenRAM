magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1296 -1277 1764 2731
<< nwell >>
rect -36 679 504 1471
<< poly >>
rect 114 225 144 1113
rect 214 225 244 1113
<< locali >>
rect 0 1397 468 1431
rect 62 1218 96 1397
rect 262 1218 296 1397
rect 366 1322 400 1397
rect 162 1168 196 1218
rect 162 1134 364 1168
rect 212 485 246 551
rect 112 237 146 303
rect 330 243 364 1134
rect 262 209 364 243
rect 262 158 296 209
rect 62 17 96 92
rect 366 17 400 92
rect 0 -17 468 17
use nmos_m1_w0_740_sactive_dli  nmos_m1_w0_740_sactive_dli_0
timestamp 1595931502
transform 1 0 154 0 1 51
box 0 -26 150 174
use pmos_m1_w1_120_sli_dli  pmos_m1_w1_120_sli_dli_1
timestamp 1595931502
transform 1 0 54 0 1 1139
box -59 -54 209 278
use pmos_m1_w1_120_sli_dli  pmos_m1_w1_120_sli_dli_0
timestamp 1595931502
transform 1 0 154 0 1 1139
box -59 -54 209 278
use contact_24  contact_24_0
timestamp 1595931502
transform 1 0 358 0 1 1281
box -59 -43 109 125
use contact_12  contact_12_1
timestamp 1595931502
transform 1 0 96 0 1 237
box 0 0 66 66
use contact_12  contact_12_0
timestamp 1595931502
transform 1 0 196 0 1 485
box 0 0 66 66
use nmos_m1_w0_740_sli_dactive  nmos_m1_w0_740_sli_dactive_0
timestamp 1595931502
transform 1 0 54 0 1 51
box 0 -26 150 174
use contact_25  contact_25_0
timestamp 1595931502
transform 1 0 358 0 1 51
box 0 0 50 82
<< labels >>
rlabel corelocali s 234 0 234 0 4 gnd
rlabel corelocali s 229 518 229 518 4 B
rlabel corelocali s 347 1151 347 1151 4 Z
rlabel corelocali s 129 270 129 270 4 A
rlabel corelocali s 234 1414 234 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 468 1414
<< end >>
