magic
tech gf180mcuD
magscale 1 10
timestamp 1694474583
<< nwell >>
rect 290 388 1009 1008
<< nmos >>
rect -174 728 -4 788
rect -174 618 -4 678
<< pmos >>
rect 380 758 721 818
rect 380 588 721 648
<< ndiff >>
rect -174 866 -4 888
rect -174 820 -112 866
rect -66 820 -4 866
rect -174 788 -4 820
rect -174 678 -4 728
rect -174 586 -4 618
rect -174 540 -112 586
rect -66 540 -4 586
rect -174 518 -4 540
<< pdiff >>
rect 380 896 721 918
rect 380 850 433 896
rect 668 850 721 896
rect 380 818 721 850
rect 380 726 721 758
rect 380 680 433 726
rect 668 680 721 726
rect 380 648 721 680
rect 380 556 721 588
rect 380 510 433 556
rect 668 510 721 556
rect 380 488 721 510
<< ndiffc >>
rect -112 820 -66 866
rect -112 540 -66 586
<< pdiffc >>
rect 433 850 668 896
rect 433 680 668 726
rect 433 510 668 556
<< psubdiff >>
rect -311 451 -204 468
rect -311 405 -271 451
rect -225 405 -204 451
rect -311 388 -204 405
<< nsubdiff >>
rect 787 535 867 572
rect 787 489 804 535
rect 850 489 867 535
rect 787 465 867 489
<< psubdiffcont >>
rect -271 405 -225 451
<< nsubdiffcont >>
rect 804 489 850 535
<< polysilicon >>
rect -297 801 -214 828
rect -297 755 -281 801
rect -235 788 -214 801
rect 46 788 380 818
rect -235 755 -174 788
rect -297 728 -174 755
rect -4 758 380 788
rect 721 758 771 818
rect -4 728 86 758
rect -297 662 -174 678
rect -297 616 -281 662
rect -235 618 -174 662
rect -4 648 86 678
rect -4 618 380 648
rect -235 616 -214 618
rect -297 578 -214 616
rect 46 588 380 618
rect 721 588 771 648
<< polycontact >>
rect -281 755 -235 801
rect -281 616 -235 662
<< metal1 >>
rect -174 866 66 868
rect -284 801 -232 853
rect -174 820 -112 866
rect -66 820 66 866
rect 422 850 433 896
rect 668 850 679 896
rect 518 844 530 850
rect 582 844 594 850
rect -174 818 66 820
rect -284 755 -281 801
rect -235 755 -232 801
rect -284 741 -232 755
rect 16 728 66 818
rect 781 728 827 896
rect 16 726 827 728
rect 16 680 433 726
rect 668 680 827 726
rect 16 678 827 680
rect -284 662 -232 676
rect -284 616 -281 662
rect -235 616 -232 662
rect -284 557 -232 616
rect -144 534 -112 586
rect -60 534 -37 586
rect 518 556 530 562
rect 582 556 594 562
rect -144 528 -37 534
rect 422 510 433 556
rect 668 510 679 556
rect 754 486 801 538
rect 853 486 865 538
rect -305 454 -206 464
rect -305 402 -274 454
rect -222 402 -206 454
rect -305 394 -206 402
<< via1 >>
rect 530 850 582 896
rect 530 844 582 850
rect -112 540 -66 586
rect -66 540 -60 586
rect -112 534 -60 540
rect 530 556 582 562
rect 530 510 582 556
rect 801 535 853 538
rect 801 489 804 535
rect 804 489 850 535
rect 850 489 853 535
rect 801 486 853 489
rect -274 451 -222 454
rect -274 405 -271 451
rect -271 405 -225 451
rect -225 405 -222 451
rect -274 402 -222 405
<< metal2 >>
rect -114 586 -58 948
rect -114 534 -112 586
rect -60 534 -58 586
rect -114 456 -58 534
rect -296 454 -58 456
rect -296 402 -274 454
rect -222 402 -58 454
rect 528 896 584 948
rect 528 844 530 896
rect 582 844 584 896
rect 528 562 584 844
rect 528 510 530 562
rect 582 540 584 562
rect 582 538 865 540
rect 582 510 801 538
rect 528 486 801 510
rect 853 486 865 538
rect 528 484 865 486
rect 528 436 584 484
rect -296 400 -58 402
<< labels >>
rlabel metal1 s -257 778 -257 778 4 B
rlabel metal1 s -257 639 -257 639 4 A
rlabel metal1 s 803 873 803 873 4 Y
rlabel metal2 s 556 461 556 461 4 VDD
rlabel metal2 s -85 484 -85 484 4 GND
<< properties >>
string FIXED_BBOX -384 388 1009 1009
<< end >>
