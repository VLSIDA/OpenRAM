magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1296 -1277 1772 2731
<< nwell >>
rect -36 679 512 1471
<< locali >>
rect 0 1397 476 1431
rect 64 648 98 714
rect 183 664 217 698
rect 0 -17 476 17
use pinv_9  pinv_9_0
timestamp 1595931502
transform 1 0 0 0 1 0
box -36 -17 512 1471
<< labels >>
rlabel corelocali s 238 0 238 0 4 gnd
rlabel corelocali s 200 681 200 681 4 Z
rlabel corelocali s 238 1414 238 1414 4 vdd
rlabel corelocali s 81 681 81 681 4 A
<< properties >>
string FIXED_BBOX 0 0 476 1414
<< end >>
