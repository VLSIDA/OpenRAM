magic
tech gf180mcuD
magscale 1 10
timestamp 1694492972
<< nwell >>
rect 675 -40 1355 640
<< nmos >>
rect 211 300 381 360
rect 211 190 381 250
<< pmos >>
rect 765 330 1106 390
rect 765 160 1106 220
<< ndiff >>
rect 211 438 381 460
rect 211 392 273 438
rect 319 392 381 438
rect 211 360 381 392
rect 211 250 381 300
rect 211 158 381 190
rect 211 112 273 158
rect 319 112 381 158
rect 211 90 381 112
<< pdiff >>
rect 765 468 1106 490
rect 765 422 818 468
rect 1052 422 1106 468
rect 765 390 1106 422
rect 765 298 1106 330
rect 765 252 818 298
rect 1052 252 1106 298
rect 765 220 1106 252
rect 765 128 1106 160
rect 765 82 818 128
rect 1052 82 1106 128
rect 765 60 1106 82
<< ndiffc >>
rect 273 392 319 438
rect 273 112 319 158
<< pdiffc >>
rect 818 422 1052 468
rect 818 252 1052 298
rect 818 82 1052 128
<< psubdiff >>
rect 74 23 181 40
rect 74 -23 114 23
rect 160 -23 181 23
rect 74 -40 181 -23
<< nsubdiff >>
rect 1172 107 1252 144
rect 1172 61 1189 107
rect 1235 61 1252 107
rect 1172 37 1252 61
<< psubdiffcont >>
rect 114 -23 160 23
<< nsubdiffcont >>
rect 1189 61 1235 107
<< polysilicon >>
rect 88 373 171 400
rect 88 327 104 373
rect 150 360 171 373
rect 431 360 765 390
rect 150 327 211 360
rect 88 300 211 327
rect 381 330 765 360
rect 1106 330 1156 390
rect 381 300 471 330
rect 88 234 211 250
rect 88 188 104 234
rect 150 190 211 234
rect 381 220 471 250
rect 381 190 765 220
rect 150 188 171 190
rect 88 150 171 188
rect 431 160 765 190
rect 1106 160 1156 220
<< polycontact >>
rect 104 327 150 373
rect 104 188 150 234
<< metal1 >>
rect 211 438 451 440
rect 101 373 153 425
rect 211 392 273 438
rect 319 392 451 438
rect 807 422 818 468
rect 1052 422 1064 468
rect 903 416 915 422
rect 967 416 979 422
rect 211 390 451 392
rect 101 327 104 373
rect 150 327 153 373
rect 101 313 153 327
rect 401 300 451 390
rect 1130 300 1182 463
rect 401 298 1182 300
rect 401 252 818 298
rect 1052 252 1182 298
rect 401 250 1182 252
rect 101 234 153 248
rect 101 188 104 234
rect 150 188 153 234
rect 101 129 153 188
rect 241 106 273 158
rect 325 106 348 158
rect 903 128 915 134
rect 967 128 979 134
rect 241 100 348 106
rect 807 82 818 128
rect 1052 82 1064 128
rect 1139 58 1186 110
rect 1238 58 1250 110
rect 80 26 179 36
rect 80 -26 111 26
rect 163 -26 179 26
rect 80 -34 179 -26
<< via1 >>
rect 915 422 967 468
rect 915 416 967 422
rect 273 112 319 158
rect 319 112 325 158
rect 273 106 325 112
rect 915 128 967 134
rect 915 82 967 128
rect 1186 107 1238 110
rect 1186 61 1189 107
rect 1189 61 1235 107
rect 1235 61 1238 107
rect 1186 58 1238 61
rect 111 23 163 26
rect 111 -23 114 23
rect 114 -23 160 23
rect 160 -23 163 23
rect 111 -26 163 -23
<< metal2 >>
rect 271 158 327 520
rect 271 106 273 158
rect 325 106 327 158
rect 271 28 327 106
rect 89 26 327 28
rect 89 -26 111 26
rect 163 -26 327 26
rect 913 468 969 520
rect 913 416 915 468
rect 967 416 969 468
rect 913 134 969 416
rect 913 82 915 134
rect 967 112 969 134
rect 967 110 1250 112
rect 967 82 1186 110
rect 913 58 1186 82
rect 1238 58 1250 110
rect 913 56 1250 58
rect 913 8 969 56
rect 89 -28 327 -26
<< labels >>
rlabel metal1 s 1156 439 1156 439 4 Y
rlabel metal1 s 127 211 127 211 4 B
rlabel metal1 s 127 350 127 350 4 A
rlabel metal2 s 941 33 941 33 4 VDD
rlabel metal2 s 300 56 300 56 4 GND
<< properties >>
string FIXED_BBOX -17 0 1373 522
<< end >>
