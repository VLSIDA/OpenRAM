magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1296 -1277 1664 2731
<< nwell >>
rect -36 679 404 1471
<< poly >>
rect 114 702 144 1113
rect 81 636 144 702
rect 114 149 144 636
<< locali >>
rect 0 1397 368 1431
rect 62 1218 96 1397
rect 266 1322 300 1397
rect 64 636 98 702
rect 162 686 196 1284
rect 162 652 213 686
rect 162 54 196 652
rect 62 17 96 54
rect 266 17 300 92
rect 0 -17 368 17
use pmos_m1_w1_120_sli_dli_da_p  pmos_m1_w1_120_sli_dli_da_p_0
timestamp 1595931502
transform 1 0 54 0 1 1139
box -59 -54 209 278
use contact_24  contact_24_0
timestamp 1595931502
transform 1 0 258 0 1 1281
box -59 -43 109 125
use nmos_m1_w0_360_sli_dli_da_p  nmos_m1_w0_360_sli_dli_da_p_0
timestamp 1595931502
transform 1 0 54 0 1 51
box 0 -26 150 98
use contact_12  contact_12_0
timestamp 1595931502
transform 1 0 48 0 1 636
box 0 0 66 66
use contact_25  contact_25_0
timestamp 1595931502
transform 1 0 258 0 1 51
box 0 0 50 82
<< labels >>
rlabel corelocali s 184 0 184 0 4 gnd
rlabel corelocali s 196 669 196 669 4 Z
rlabel corelocali s 184 1414 184 1414 4 vdd
rlabel corelocali s 81 669 81 669 4 A
<< properties >>
string FIXED_BBOX 0 0 368 1414
<< end >>
