VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 21695.0 by 42337.5 ;
END  MacroSite
MACRO sram_2_16_1_freepdk45
   CLASS BLOCK ;
   SIZE 21695.0 BY 42337.5 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN DATA[0]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  14837.5 0.0 14907.5 140.0 ;
      END
   END DATA[0]
   PIN DATA[1]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  15542.5 0.0 15612.5 140.0 ;
      END
   END DATA[1]
   PIN ADDR[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 7532.5 4655.0 7602.5 ;
      END
   END ADDR[0]
   PIN ADDR[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 6827.5 4655.0 6897.5 ;
      END
   END ADDR[1]
   PIN ADDR[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 6122.5 4655.0 6192.5 ;
      END
   END ADDR[2]
   PIN ADDR[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 5417.5 4655.0 5487.5 ;
      END
   END ADDR[3]
   PIN CSb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1187.5 19230.0 1257.5 19370.0 ;
      END
   END CSb
   PIN WEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1892.5 19230.0 1962.5 19370.0 ;
      END
   END WEb
   PIN OEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  482.5 19230.0 552.5 19370.0 ;
      END
   END OEb
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER metal1 ;
         RECT  3340.0 19230.0 3475.0 19420.0 ;
      END
   END clk
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal1 ;
         RECT  16125.0 0.0 16475.0 42337.5 ;
         LAYER metal1 ;
         RECT  4175.0 0.0 4525.0 42337.5 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal2 ;
         RECT  12427.5 0.0 12777.5 42337.5 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  4317.5 26935.0 4382.5 27140.0 ;
      RECT  8475.0 19685.0 8540.0 19750.0 ;
      RECT  8475.0 19412.5 8540.0 19477.5 ;
      RECT  8405.0 19685.0 8507.5 19750.0 ;
      RECT  8475.0 19445.0 8540.0 19717.5 ;
      RECT  8507.5 19412.5 8610.0 19477.5 ;
      RECT  12632.5 19685.0 12697.5 19750.0 ;
      RECT  12632.5 19197.5 12697.5 19262.5 ;
      RECT  10900.0 19685.0 12665.0 19750.0 ;
      RECT  12632.5 19230.0 12697.5 19717.5 ;
      RECT  12665.0 19197.5 14430.0 19262.5 ;
      RECT  8475.0 21120.0 8540.0 21185.0 ;
      RECT  8475.0 21392.5 8540.0 21457.5 ;
      RECT  8405.0 21120.0 8507.5 21185.0 ;
      RECT  8475.0 21152.5 8540.0 21425.0 ;
      RECT  8507.5 21392.5 8610.0 21457.5 ;
      RECT  12632.5 21120.0 12697.5 21185.0 ;
      RECT  12632.5 21607.5 12697.5 21672.5 ;
      RECT  10900.0 21120.0 12665.0 21185.0 ;
      RECT  12632.5 21152.5 12697.5 21640.0 ;
      RECT  12665.0 21607.5 14430.0 21672.5 ;
      RECT  8475.0 22375.0 8540.0 22440.0 ;
      RECT  8475.0 22102.5 8540.0 22167.5 ;
      RECT  8405.0 22375.0 8507.5 22440.0 ;
      RECT  8475.0 22135.0 8540.0 22407.5 ;
      RECT  8507.5 22102.5 8610.0 22167.5 ;
      RECT  12632.5 22375.0 12697.5 22440.0 ;
      RECT  12632.5 21887.5 12697.5 21952.5 ;
      RECT  10900.0 22375.0 12665.0 22440.0 ;
      RECT  12632.5 21920.0 12697.5 22407.5 ;
      RECT  12665.0 21887.5 14430.0 21952.5 ;
      RECT  8475.0 23810.0 8540.0 23875.0 ;
      RECT  8475.0 24082.5 8540.0 24147.5 ;
      RECT  8405.0 23810.0 8507.5 23875.0 ;
      RECT  8475.0 23842.5 8540.0 24115.0 ;
      RECT  8507.5 24082.5 8610.0 24147.5 ;
      RECT  12632.5 23810.0 12697.5 23875.0 ;
      RECT  12632.5 24297.5 12697.5 24362.5 ;
      RECT  10900.0 23810.0 12665.0 23875.0 ;
      RECT  12632.5 23842.5 12697.5 24330.0 ;
      RECT  12665.0 24297.5 14430.0 24362.5 ;
      RECT  8475.0 25065.0 8540.0 25130.0 ;
      RECT  8475.0 24792.5 8540.0 24857.5 ;
      RECT  8405.0 25065.0 8507.5 25130.0 ;
      RECT  8475.0 24825.0 8540.0 25097.5 ;
      RECT  8507.5 24792.5 8610.0 24857.5 ;
      RECT  12632.5 25065.0 12697.5 25130.0 ;
      RECT  12632.5 24577.5 12697.5 24642.5 ;
      RECT  10900.0 25065.0 12665.0 25130.0 ;
      RECT  12632.5 24610.0 12697.5 25097.5 ;
      RECT  12665.0 24577.5 14430.0 24642.5 ;
      RECT  8475.0 26500.0 8540.0 26565.0 ;
      RECT  8475.0 26772.5 8540.0 26837.5 ;
      RECT  8405.0 26500.0 8507.5 26565.0 ;
      RECT  8475.0 26532.5 8540.0 26805.0 ;
      RECT  8507.5 26772.5 8610.0 26837.5 ;
      RECT  12632.5 26500.0 12697.5 26565.0 ;
      RECT  12632.5 26987.5 12697.5 27052.5 ;
      RECT  10900.0 26500.0 12665.0 26565.0 ;
      RECT  12632.5 26532.5 12697.5 27020.0 ;
      RECT  12665.0 26987.5 14430.0 27052.5 ;
      RECT  8475.0 27755.0 8540.0 27820.0 ;
      RECT  8475.0 27482.5 8540.0 27547.5 ;
      RECT  8405.0 27755.0 8507.5 27820.0 ;
      RECT  8475.0 27515.0 8540.0 27787.5 ;
      RECT  8507.5 27482.5 8610.0 27547.5 ;
      RECT  12632.5 27755.0 12697.5 27820.0 ;
      RECT  12632.5 27267.5 12697.5 27332.5 ;
      RECT  10900.0 27755.0 12665.0 27820.0 ;
      RECT  12632.5 27300.0 12697.5 27787.5 ;
      RECT  12665.0 27267.5 14430.0 27332.5 ;
      RECT  8475.0 29190.0 8540.0 29255.0 ;
      RECT  8475.0 29462.5 8540.0 29527.5 ;
      RECT  8405.0 29190.0 8507.5 29255.0 ;
      RECT  8475.0 29222.5 8540.0 29495.0 ;
      RECT  8507.5 29462.5 8610.0 29527.5 ;
      RECT  12632.5 29190.0 12697.5 29255.0 ;
      RECT  12632.5 29677.5 12697.5 29742.5 ;
      RECT  10900.0 29190.0 12665.0 29255.0 ;
      RECT  12632.5 29222.5 12697.5 29710.0 ;
      RECT  12665.0 29677.5 14430.0 29742.5 ;
      RECT  8475.0 30445.0 8540.0 30510.0 ;
      RECT  8475.0 30172.5 8540.0 30237.5 ;
      RECT  8405.0 30445.0 8507.5 30510.0 ;
      RECT  8475.0 30205.0 8540.0 30477.5 ;
      RECT  8507.5 30172.5 8610.0 30237.5 ;
      RECT  12632.5 30445.0 12697.5 30510.0 ;
      RECT  12632.5 29957.5 12697.5 30022.5 ;
      RECT  10900.0 30445.0 12665.0 30510.0 ;
      RECT  12632.5 29990.0 12697.5 30477.5 ;
      RECT  12665.0 29957.5 14430.0 30022.5 ;
      RECT  8475.0 31880.0 8540.0 31945.0 ;
      RECT  8475.0 32152.5 8540.0 32217.5 ;
      RECT  8405.0 31880.0 8507.5 31945.0 ;
      RECT  8475.0 31912.5 8540.0 32185.0 ;
      RECT  8507.5 32152.5 8610.0 32217.5 ;
      RECT  12632.5 31880.0 12697.5 31945.0 ;
      RECT  12632.5 32367.5 12697.5 32432.5 ;
      RECT  10900.0 31880.0 12665.0 31945.0 ;
      RECT  12632.5 31912.5 12697.5 32400.0 ;
      RECT  12665.0 32367.5 14430.0 32432.5 ;
      RECT  8475.0 33135.0 8540.0 33200.0 ;
      RECT  8475.0 32862.5 8540.0 32927.5 ;
      RECT  8405.0 33135.0 8507.5 33200.0 ;
      RECT  8475.0 32895.0 8540.0 33167.5 ;
      RECT  8507.5 32862.5 8610.0 32927.5 ;
      RECT  12632.5 33135.0 12697.5 33200.0 ;
      RECT  12632.5 32647.5 12697.5 32712.5 ;
      RECT  10900.0 33135.0 12665.0 33200.0 ;
      RECT  12632.5 32680.0 12697.5 33167.5 ;
      RECT  12665.0 32647.5 14430.0 32712.5 ;
      RECT  8475.0 34570.0 8540.0 34635.0 ;
      RECT  8475.0 34842.5 8540.0 34907.5 ;
      RECT  8405.0 34570.0 8507.5 34635.0 ;
      RECT  8475.0 34602.5 8540.0 34875.0 ;
      RECT  8507.5 34842.5 8610.0 34907.5 ;
      RECT  12632.5 34570.0 12697.5 34635.0 ;
      RECT  12632.5 35057.5 12697.5 35122.5 ;
      RECT  10900.0 34570.0 12665.0 34635.0 ;
      RECT  12632.5 34602.5 12697.5 35090.0 ;
      RECT  12665.0 35057.5 14430.0 35122.5 ;
      RECT  8475.0 35825.0 8540.0 35890.0 ;
      RECT  8475.0 35552.5 8540.0 35617.5 ;
      RECT  8405.0 35825.0 8507.5 35890.0 ;
      RECT  8475.0 35585.0 8540.0 35857.5 ;
      RECT  8507.5 35552.5 8610.0 35617.5 ;
      RECT  12632.5 35825.0 12697.5 35890.0 ;
      RECT  12632.5 35337.5 12697.5 35402.5 ;
      RECT  10900.0 35825.0 12665.0 35890.0 ;
      RECT  12632.5 35370.0 12697.5 35857.5 ;
      RECT  12665.0 35337.5 14430.0 35402.5 ;
      RECT  8475.0 37260.0 8540.0 37325.0 ;
      RECT  8475.0 37532.5 8540.0 37597.5 ;
      RECT  8405.0 37260.0 8507.5 37325.0 ;
      RECT  8475.0 37292.5 8540.0 37565.0 ;
      RECT  8507.5 37532.5 8610.0 37597.5 ;
      RECT  12632.5 37260.0 12697.5 37325.0 ;
      RECT  12632.5 37747.5 12697.5 37812.5 ;
      RECT  10900.0 37260.0 12665.0 37325.0 ;
      RECT  12632.5 37292.5 12697.5 37780.0 ;
      RECT  12665.0 37747.5 14430.0 37812.5 ;
      RECT  8475.0 38515.0 8540.0 38580.0 ;
      RECT  8475.0 38242.5 8540.0 38307.5 ;
      RECT  8405.0 38515.0 8507.5 38580.0 ;
      RECT  8475.0 38275.0 8540.0 38547.5 ;
      RECT  8507.5 38242.5 8610.0 38307.5 ;
      RECT  12632.5 38515.0 12697.5 38580.0 ;
      RECT  12632.5 38027.5 12697.5 38092.5 ;
      RECT  10900.0 38515.0 12665.0 38580.0 ;
      RECT  12632.5 38060.0 12697.5 38547.5 ;
      RECT  12665.0 38027.5 14430.0 38092.5 ;
      RECT  8475.0 39950.0 8540.0 40015.0 ;
      RECT  8475.0 40222.5 8540.0 40287.5 ;
      RECT  8405.0 39950.0 8507.5 40015.0 ;
      RECT  8475.0 39982.5 8540.0 40255.0 ;
      RECT  8507.5 40222.5 8610.0 40287.5 ;
      RECT  12632.5 39950.0 12697.5 40015.0 ;
      RECT  12632.5 40437.5 12697.5 40502.5 ;
      RECT  10900.0 39950.0 12665.0 40015.0 ;
      RECT  12632.5 39982.5 12697.5 40470.0 ;
      RECT  12665.0 40437.5 14430.0 40502.5 ;
      RECT  9065.0 19057.5 14520.0 19122.5 ;
      RECT  9065.0 21747.5 14520.0 21812.5 ;
      RECT  9065.0 24437.5 14520.0 24502.5 ;
      RECT  9065.0 27127.5 14520.0 27192.5 ;
      RECT  9065.0 29817.5 14520.0 29882.5 ;
      RECT  9065.0 32507.5 14520.0 32572.5 ;
      RECT  9065.0 35197.5 14520.0 35262.5 ;
      RECT  9065.0 37887.5 14520.0 37952.5 ;
      RECT  9065.0 40577.5 14520.0 40642.5 ;
      RECT  4175.0 20402.5 16475.0 20467.5 ;
      RECT  4175.0 23092.5 16475.0 23157.5 ;
      RECT  4175.0 25782.5 16475.0 25847.5 ;
      RECT  4175.0 28472.5 16475.0 28537.5 ;
      RECT  4175.0 31162.5 16475.0 31227.5 ;
      RECT  4175.0 33852.5 16475.0 33917.5 ;
      RECT  4175.0 36542.5 16475.0 36607.5 ;
      RECT  4175.0 39232.5 16475.0 39297.5 ;
      RECT  11095.0 8502.5 11437.5 8567.5 ;
      RECT  10820.0 9847.5 11642.5 9912.5 ;
      RECT  11095.0 13882.5 11847.5 13947.5 ;
      RECT  10820.0 15227.5 12052.5 15292.5 ;
      RECT  11095.0 8297.5 11232.5 8362.5 ;
      RECT  11095.0 10987.5 11232.5 11052.5 ;
      RECT  11095.0 13677.5 11232.5 13742.5 ;
      RECT  11095.0 16367.5 11232.5 16432.5 ;
      RECT  4175.0 9642.5 11095.0 9707.5 ;
      RECT  4175.0 12332.5 11095.0 12397.5 ;
      RECT  4175.0 15022.5 11095.0 15087.5 ;
      RECT  4175.0 17712.5 11095.0 17777.5 ;
      RECT  11095.0 7535.0 11437.5 7600.0 ;
      RECT  11095.0 6830.0 11642.5 6895.0 ;
      RECT  11095.0 6125.0 11847.5 6190.0 ;
      RECT  11095.0 5420.0 12052.5 5485.0 ;
      RECT  11095.0 7887.5 12562.5 7952.5 ;
      RECT  11095.0 7182.5 12562.5 7247.5 ;
      RECT  11095.0 6477.5 12562.5 6542.5 ;
      RECT  11095.0 5772.5 12562.5 5837.5 ;
      RECT  11095.0 5067.5 12562.5 5132.5 ;
      RECT  7865.0 4862.5 7930.0 4927.5 ;
      RECT  7865.0 4895.0 7930.0 5100.0 ;
      RECT  4175.0 4862.5 7897.5 4927.5 ;
      RECT  10825.0 4862.5 10890.0 4927.5 ;
      RECT  10825.0 4895.0 10890.0 5100.0 ;
      RECT  4175.0 4862.5 10857.5 4927.5 ;
      RECT  5875.0 4862.5 5940.0 4927.5 ;
      RECT  5875.0 4895.0 5940.0 5100.0 ;
      RECT  4175.0 4862.5 5907.5 4927.5 ;
      RECT  8835.0 4862.5 8900.0 4927.5 ;
      RECT  8835.0 4895.0 8900.0 5100.0 ;
      RECT  4175.0 4862.5 8867.5 4927.5 ;
      RECT  13632.5 3795.0 14520.0 3860.0 ;
      RECT  13222.5 1610.0 14520.0 1675.0 ;
      RECT  13427.5 3157.5 14520.0 3222.5 ;
      RECT  13632.5 41587.5 14520.0 41652.5 ;
      RECT  13837.5 10297.5 14520.0 10362.5 ;
      RECT  14042.5 14322.5 14520.0 14387.5 ;
      RECT  4860.0 8092.5 4925.0 8157.5 ;
      RECT  4860.0 7920.0 4925.0 8125.0 ;
      RECT  4892.5 8092.5 13017.5 8157.5 ;
      RECT  8840.0 40782.5 13082.5 40847.5 ;
      RECT  14520.0 42272.5 16125.0 42337.5 ;
      RECT  14520.0 18895.0 16125.0 18960.0 ;
      RECT  14520.0 10427.5 16125.0 10492.5 ;
      RECT  14520.0 6800.0 16125.0 6865.0 ;
      RECT  14520.0 9760.0 16125.0 9825.0 ;
      RECT  14520.0 4810.0 16125.0 4875.0 ;
      RECT  14520.0 7770.0 16125.0 7835.0 ;
      RECT  14520.0 1740.0 16125.0 1805.0 ;
      RECT  12777.5 3027.5 14520.0 3092.5 ;
      RECT  12777.5 14452.5 14520.0 14517.5 ;
      RECT  12777.5 3955.0 14520.0 4020.0 ;
      RECT  12777.5 11230.0 14520.0 11295.0 ;
      RECT  14520.0 19090.0 15225.0 20435.0 ;
      RECT  14520.0 21780.0 15225.0 20435.0 ;
      RECT  14520.0 21780.0 15225.0 23125.0 ;
      RECT  14520.0 24470.0 15225.0 23125.0 ;
      RECT  14520.0 24470.0 15225.0 25815.0 ;
      RECT  14520.0 27160.0 15225.0 25815.0 ;
      RECT  14520.0 27160.0 15225.0 28505.0 ;
      RECT  14520.0 29850.0 15225.0 28505.0 ;
      RECT  14520.0 29850.0 15225.0 31195.0 ;
      RECT  14520.0 32540.0 15225.0 31195.0 ;
      RECT  14520.0 32540.0 15225.0 33885.0 ;
      RECT  14520.0 35230.0 15225.0 33885.0 ;
      RECT  14520.0 35230.0 15225.0 36575.0 ;
      RECT  14520.0 37920.0 15225.0 36575.0 ;
      RECT  14520.0 37920.0 15225.0 39265.0 ;
      RECT  14520.0 40610.0 15225.0 39265.0 ;
      RECT  15225.0 19090.0 15930.0 20435.0 ;
      RECT  15225.0 21780.0 15930.0 20435.0 ;
      RECT  15225.0 21780.0 15930.0 23125.0 ;
      RECT  15225.0 24470.0 15930.0 23125.0 ;
      RECT  15225.0 24470.0 15930.0 25815.0 ;
      RECT  15225.0 27160.0 15930.0 25815.0 ;
      RECT  15225.0 27160.0 15930.0 28505.0 ;
      RECT  15225.0 29850.0 15930.0 28505.0 ;
      RECT  15225.0 29850.0 15930.0 31195.0 ;
      RECT  15225.0 32540.0 15930.0 31195.0 ;
      RECT  15225.0 32540.0 15930.0 33885.0 ;
      RECT  15225.0 35230.0 15930.0 33885.0 ;
      RECT  15225.0 35230.0 15930.0 36575.0 ;
      RECT  15225.0 37920.0 15930.0 36575.0 ;
      RECT  15225.0 37920.0 15930.0 39265.0 ;
      RECT  15225.0 40610.0 15930.0 39265.0 ;
      RECT  14430.0 19197.5 16020.0 19262.5 ;
      RECT  14430.0 21607.5 16020.0 21672.5 ;
      RECT  14430.0 21887.5 16020.0 21952.5 ;
      RECT  14430.0 24297.5 16020.0 24362.5 ;
      RECT  14430.0 24577.5 16020.0 24642.5 ;
      RECT  14430.0 26987.5 16020.0 27052.5 ;
      RECT  14430.0 27267.5 16020.0 27332.5 ;
      RECT  14430.0 29677.5 16020.0 29742.5 ;
      RECT  14430.0 29957.5 16020.0 30022.5 ;
      RECT  14430.0 32367.5 16020.0 32432.5 ;
      RECT  14430.0 32647.5 16020.0 32712.5 ;
      RECT  14430.0 35057.5 16020.0 35122.5 ;
      RECT  14430.0 35337.5 16020.0 35402.5 ;
      RECT  14430.0 37747.5 16020.0 37812.5 ;
      RECT  14430.0 38027.5 16020.0 38092.5 ;
      RECT  14430.0 40437.5 16020.0 40502.5 ;
      RECT  14430.0 20402.5 16020.0 20467.5 ;
      RECT  14430.0 23092.5 16020.0 23157.5 ;
      RECT  14430.0 25782.5 16020.0 25847.5 ;
      RECT  14430.0 28472.5 16020.0 28537.5 ;
      RECT  14430.0 31162.5 16020.0 31227.5 ;
      RECT  14430.0 33852.5 16020.0 33917.5 ;
      RECT  14430.0 36542.5 16020.0 36607.5 ;
      RECT  14430.0 39232.5 16020.0 39297.5 ;
      RECT  14430.0 19057.5 16020.0 19122.5 ;
      RECT  14430.0 21747.5 16020.0 21812.5 ;
      RECT  14430.0 24437.5 16020.0 24502.5 ;
      RECT  14430.0 27127.5 16020.0 27192.5 ;
      RECT  14430.0 29817.5 16020.0 29882.5 ;
      RECT  14430.0 32507.5 16020.0 32572.5 ;
      RECT  14430.0 35197.5 16020.0 35262.5 ;
      RECT  14430.0 37887.5 16020.0 37952.5 ;
      RECT  14430.0 40577.5 16020.0 40642.5 ;
      RECT  14872.5 41822.5 14937.5 42337.5 ;
      RECT  14682.5 41292.5 14747.5 41427.5 ;
      RECT  14872.5 41292.5 14937.5 41427.5 ;
      RECT  14872.5 41292.5 14937.5 41427.5 ;
      RECT  14682.5 41292.5 14747.5 41427.5 ;
      RECT  14682.5 41822.5 14747.5 41957.5 ;
      RECT  14872.5 41822.5 14937.5 41957.5 ;
      RECT  14872.5 41822.5 14937.5 41957.5 ;
      RECT  14682.5 41822.5 14747.5 41957.5 ;
      RECT  14872.5 41822.5 14937.5 41957.5 ;
      RECT  15062.5 41822.5 15127.5 41957.5 ;
      RECT  15062.5 41822.5 15127.5 41957.5 ;
      RECT  14872.5 41822.5 14937.5 41957.5 ;
      RECT  14852.5 41587.5 14717.5 41652.5 ;
      RECT  14872.5 42135.0 14937.5 42270.0 ;
      RECT  14682.5 41292.5 14747.5 41427.5 ;
      RECT  14872.5 41292.5 14937.5 41427.5 ;
      RECT  14682.5 41822.5 14747.5 41957.5 ;
      RECT  15062.5 41822.5 15127.5 41957.5 ;
      RECT  14520.0 41587.5 15225.0 41652.5 ;
      RECT  14520.0 42272.5 15225.0 42337.5 ;
      RECT  15577.5 41822.5 15642.5 42337.5 ;
      RECT  15387.5 41292.5 15452.5 41427.5 ;
      RECT  15577.5 41292.5 15642.5 41427.5 ;
      RECT  15577.5 41292.5 15642.5 41427.5 ;
      RECT  15387.5 41292.5 15452.5 41427.5 ;
      RECT  15387.5 41822.5 15452.5 41957.5 ;
      RECT  15577.5 41822.5 15642.5 41957.5 ;
      RECT  15577.5 41822.5 15642.5 41957.5 ;
      RECT  15387.5 41822.5 15452.5 41957.5 ;
      RECT  15577.5 41822.5 15642.5 41957.5 ;
      RECT  15767.5 41822.5 15832.5 41957.5 ;
      RECT  15767.5 41822.5 15832.5 41957.5 ;
      RECT  15577.5 41822.5 15642.5 41957.5 ;
      RECT  15557.5 41587.5 15422.5 41652.5 ;
      RECT  15577.5 42135.0 15642.5 42270.0 ;
      RECT  15387.5 41292.5 15452.5 41427.5 ;
      RECT  15577.5 41292.5 15642.5 41427.5 ;
      RECT  15387.5 41822.5 15452.5 41957.5 ;
      RECT  15767.5 41822.5 15832.5 41957.5 ;
      RECT  15225.0 41587.5 15930.0 41652.5 ;
      RECT  15225.0 42272.5 15930.0 42337.5 ;
      RECT  14520.0 41587.5 15930.0 41652.5 ;
      RECT  14520.0 42272.5 15930.0 42337.5 ;
      RECT  14520.0 14205.0 15225.0 19090.0 ;
      RECT  15225.0 14205.0 15930.0 19090.0 ;
      RECT  14520.0 14322.5 15930.0 14387.5 ;
      RECT  14520.0 18895.0 15930.0 18960.0 ;
      RECT  14520.0 14452.5 15930.0 14517.5 ;
      RECT  14520.0 10030.0 15225.0 14205.0 ;
      RECT  15225.0 10030.0 15930.0 14205.0 ;
      RECT  14520.0 10297.5 15930.0 10362.5 ;
      RECT  14520.0 10427.5 15930.0 10492.5 ;
      RECT  14520.0 11230.0 15930.0 11295.0 ;
      RECT  14520.0 3590.0 15225.0 10030.0 ;
      RECT  15930.0 3590.0 15225.0 10030.0 ;
      RECT  14520.0 3795.0 15930.0 3860.0 ;
      RECT  14520.0 6800.0 15930.0 6865.0 ;
      RECT  14520.0 9760.0 15930.0 9825.0 ;
      RECT  14520.0 4810.0 15930.0 4875.0 ;
      RECT  14520.0 7770.0 15930.0 7835.0 ;
      RECT  14520.0 3955.0 15930.0 4020.0 ;
      RECT  14520.0 3590.0 15225.0 615.0 ;
      RECT  15225.0 3590.0 15930.0 615.0 ;
      RECT  14520.0 3222.5 15930.0 3157.5 ;
      RECT  14520.0 1675.0 15930.0 1610.0 ;
      RECT  14520.0 1805.0 15930.0 1740.0 ;
      RECT  14520.0 3092.5 15930.0 3027.5 ;
      RECT  7895.0 19697.5 7960.0 19762.5 ;
      RECT  7895.0 19685.0 7960.0 19750.0 ;
      RECT  7677.5 19697.5 7927.5 19762.5 ;
      RECT  7895.0 19717.5 7960.0 19730.0 ;
      RECT  7927.5 19685.0 8175.0 19750.0 ;
      RECT  7895.0 21107.5 7960.0 21172.5 ;
      RECT  7895.0 21120.0 7960.0 21185.0 ;
      RECT  7677.5 21107.5 7927.5 21172.5 ;
      RECT  7895.0 21140.0 7960.0 21152.5 ;
      RECT  7927.5 21120.0 8175.0 21185.0 ;
      RECT  7895.0 22387.5 7960.0 22452.5 ;
      RECT  7895.0 22375.0 7960.0 22440.0 ;
      RECT  7677.5 22387.5 7927.5 22452.5 ;
      RECT  7895.0 22407.5 7960.0 22420.0 ;
      RECT  7927.5 22375.0 8175.0 22440.0 ;
      RECT  7895.0 23797.5 7960.0 23862.5 ;
      RECT  7895.0 23810.0 7960.0 23875.0 ;
      RECT  7677.5 23797.5 7927.5 23862.5 ;
      RECT  7895.0 23830.0 7960.0 23842.5 ;
      RECT  7927.5 23810.0 8175.0 23875.0 ;
      RECT  7895.0 25077.5 7960.0 25142.5 ;
      RECT  7895.0 25065.0 7960.0 25130.0 ;
      RECT  7677.5 25077.5 7927.5 25142.5 ;
      RECT  7895.0 25097.5 7960.0 25110.0 ;
      RECT  7927.5 25065.0 8175.0 25130.0 ;
      RECT  7895.0 26487.5 7960.0 26552.5 ;
      RECT  7895.0 26500.0 7960.0 26565.0 ;
      RECT  7677.5 26487.5 7927.5 26552.5 ;
      RECT  7895.0 26520.0 7960.0 26532.5 ;
      RECT  7927.5 26500.0 8175.0 26565.0 ;
      RECT  7895.0 27767.5 7960.0 27832.5 ;
      RECT  7895.0 27755.0 7960.0 27820.0 ;
      RECT  7677.5 27767.5 7927.5 27832.5 ;
      RECT  7895.0 27787.5 7960.0 27800.0 ;
      RECT  7927.5 27755.0 8175.0 27820.0 ;
      RECT  7895.0 29177.5 7960.0 29242.5 ;
      RECT  7895.0 29190.0 7960.0 29255.0 ;
      RECT  7677.5 29177.5 7927.5 29242.5 ;
      RECT  7895.0 29210.0 7960.0 29222.5 ;
      RECT  7927.5 29190.0 8175.0 29255.0 ;
      RECT  7895.0 30457.5 7960.0 30522.5 ;
      RECT  7895.0 30445.0 7960.0 30510.0 ;
      RECT  7677.5 30457.5 7927.5 30522.5 ;
      RECT  7895.0 30477.5 7960.0 30490.0 ;
      RECT  7927.5 30445.0 8175.0 30510.0 ;
      RECT  7895.0 31867.5 7960.0 31932.5 ;
      RECT  7895.0 31880.0 7960.0 31945.0 ;
      RECT  7677.5 31867.5 7927.5 31932.5 ;
      RECT  7895.0 31900.0 7960.0 31912.5 ;
      RECT  7927.5 31880.0 8175.0 31945.0 ;
      RECT  7895.0 33147.5 7960.0 33212.5 ;
      RECT  7895.0 33135.0 7960.0 33200.0 ;
      RECT  7677.5 33147.5 7927.5 33212.5 ;
      RECT  7895.0 33167.5 7960.0 33180.0 ;
      RECT  7927.5 33135.0 8175.0 33200.0 ;
      RECT  7895.0 34557.5 7960.0 34622.5 ;
      RECT  7895.0 34570.0 7960.0 34635.0 ;
      RECT  7677.5 34557.5 7927.5 34622.5 ;
      RECT  7895.0 34590.0 7960.0 34602.5 ;
      RECT  7927.5 34570.0 8175.0 34635.0 ;
      RECT  7895.0 35837.5 7960.0 35902.5 ;
      RECT  7895.0 35825.0 7960.0 35890.0 ;
      RECT  7677.5 35837.5 7927.5 35902.5 ;
      RECT  7895.0 35857.5 7960.0 35870.0 ;
      RECT  7927.5 35825.0 8175.0 35890.0 ;
      RECT  7895.0 37247.5 7960.0 37312.5 ;
      RECT  7895.0 37260.0 7960.0 37325.0 ;
      RECT  7677.5 37247.5 7927.5 37312.5 ;
      RECT  7895.0 37280.0 7960.0 37292.5 ;
      RECT  7927.5 37260.0 8175.0 37325.0 ;
      RECT  7895.0 38527.5 7960.0 38592.5 ;
      RECT  7895.0 38515.0 7960.0 38580.0 ;
      RECT  7677.5 38527.5 7927.5 38592.5 ;
      RECT  7895.0 38547.5 7960.0 38560.0 ;
      RECT  7927.5 38515.0 8175.0 38580.0 ;
      RECT  7895.0 39937.5 7960.0 40002.5 ;
      RECT  7895.0 39950.0 7960.0 40015.0 ;
      RECT  7677.5 39937.5 7927.5 40002.5 ;
      RECT  7895.0 39970.0 7960.0 39982.5 ;
      RECT  7927.5 39950.0 8175.0 40015.0 ;
      RECT  5765.0 8925.0 7130.0 8990.0 ;
      RECT  5940.0 10360.0 7130.0 10425.0 ;
      RECT  6115.0 11615.0 7130.0 11680.0 ;
      RECT  6290.0 13050.0 7130.0 13115.0 ;
      RECT  6465.0 14305.0 7130.0 14370.0 ;
      RECT  6640.0 15740.0 7130.0 15805.0 ;
      RECT  6815.0 16995.0 7130.0 17060.0 ;
      RECT  6990.0 18430.0 7130.0 18495.0 ;
      RECT  5765.0 19697.5 7190.0 19762.5 ;
      RECT  6465.0 19482.5 7447.5 19547.5 ;
      RECT  5765.0 21107.5 7190.0 21172.5 ;
      RECT  6640.0 21322.5 7447.5 21387.5 ;
      RECT  5765.0 22387.5 7190.0 22452.5 ;
      RECT  6815.0 22172.5 7447.5 22237.5 ;
      RECT  5765.0 23797.5 7190.0 23862.5 ;
      RECT  6990.0 24012.5 7447.5 24077.5 ;
      RECT  5940.0 25077.5 7190.0 25142.5 ;
      RECT  6465.0 24862.5 7447.5 24927.5 ;
      RECT  5940.0 26487.5 7190.0 26552.5 ;
      RECT  6640.0 26702.5 7447.5 26767.5 ;
      RECT  5940.0 27767.5 7190.0 27832.5 ;
      RECT  6815.0 27552.5 7447.5 27617.5 ;
      RECT  5940.0 29177.5 7190.0 29242.5 ;
      RECT  6990.0 29392.5 7447.5 29457.5 ;
      RECT  6115.0 30457.5 7190.0 30522.5 ;
      RECT  6465.0 30242.5 7447.5 30307.5 ;
      RECT  6115.0 31867.5 7190.0 31932.5 ;
      RECT  6640.0 32082.5 7447.5 32147.5 ;
      RECT  6115.0 33147.5 7190.0 33212.5 ;
      RECT  6815.0 32932.5 7447.5 32997.5 ;
      RECT  6115.0 34557.5 7190.0 34622.5 ;
      RECT  6990.0 34772.5 7447.5 34837.5 ;
      RECT  6290.0 35837.5 7190.0 35902.5 ;
      RECT  6465.0 35622.5 7447.5 35687.5 ;
      RECT  6290.0 37247.5 7190.0 37312.5 ;
      RECT  6640.0 37462.5 7447.5 37527.5 ;
      RECT  6290.0 38527.5 7190.0 38592.5 ;
      RECT  6815.0 38312.5 7447.5 38377.5 ;
      RECT  6290.0 39937.5 7190.0 40002.5 ;
      RECT  6990.0 40152.5 7447.5 40217.5 ;
      RECT  9952.5 8925.0 9887.5 8990.0 ;
      RECT  9952.5 9447.5 9887.5 9512.5 ;
      RECT  10190.0 8925.0 9920.0 8990.0 ;
      RECT  9952.5 8957.5 9887.5 9480.0 ;
      RECT  9920.0 9447.5 9675.0 9512.5 ;
      RECT  11060.0 8925.0 10420.0 8990.0 ;
      RECT  9952.5 10360.0 9887.5 10425.0 ;
      RECT  9952.5 10792.5 9887.5 10857.5 ;
      RECT  10190.0 10360.0 9920.0 10425.0 ;
      RECT  9952.5 10392.5 9887.5 10825.0 ;
      RECT  9920.0 10792.5 9400.0 10857.5 ;
      RECT  10785.0 10360.0 10420.0 10425.0 ;
      RECT  11060.0 11122.5 9125.0 11187.5 ;
      RECT  10785.0 12467.5 8850.0 12532.5 ;
      RECT  9675.0 8937.5 8550.0 9002.5 ;
      RECT  9400.0 8722.5 8292.5 8787.5 ;
      RECT  9125.0 10347.5 8550.0 10412.5 ;
      RECT  9400.0 10562.5 8292.5 10627.5 ;
      RECT  9675.0 11627.5 8550.0 11692.5 ;
      RECT  8850.0 11412.5 8292.5 11477.5 ;
      RECT  9125.0 13037.5 8550.0 13102.5 ;
      RECT  8850.0 13252.5 8292.5 13317.5 ;
      RECT  7845.0 8937.5 7780.0 9002.5 ;
      RECT  7845.0 8925.0 7780.0 8990.0 ;
      RECT  8062.5 8937.5 7812.5 9002.5 ;
      RECT  7845.0 8957.5 7780.0 8970.0 ;
      RECT  7812.5 8925.0 7565.0 8990.0 ;
      RECT  7845.0 10347.5 7780.0 10412.5 ;
      RECT  7845.0 10360.0 7780.0 10425.0 ;
      RECT  8062.5 10347.5 7812.5 10412.5 ;
      RECT  7845.0 10380.0 7780.0 10392.5 ;
      RECT  7812.5 10360.0 7565.0 10425.0 ;
      RECT  7845.0 11627.5 7780.0 11692.5 ;
      RECT  7845.0 11615.0 7780.0 11680.0 ;
      RECT  8062.5 11627.5 7812.5 11692.5 ;
      RECT  7845.0 11647.5 7780.0 11660.0 ;
      RECT  7812.5 11615.0 7565.0 11680.0 ;
      RECT  7845.0 13037.5 7780.0 13102.5 ;
      RECT  7845.0 13050.0 7780.0 13115.0 ;
      RECT  8062.5 13037.5 7812.5 13102.5 ;
      RECT  7845.0 13070.0 7780.0 13082.5 ;
      RECT  7812.5 13050.0 7565.0 13115.0 ;
      RECT  10117.5 9490.0 10052.5 9675.0 ;
      RECT  10117.5 8330.0 10052.5 8515.0 ;
      RECT  10477.5 8447.5 10412.5 8297.5 ;
      RECT  10477.5 9332.5 10412.5 9707.5 ;
      RECT  10287.5 8447.5 10222.5 9332.5 ;
      RECT  10477.5 9332.5 10412.5 9467.5 ;
      RECT  10287.5 9332.5 10222.5 9467.5 ;
      RECT  10287.5 9332.5 10222.5 9467.5 ;
      RECT  10477.5 9332.5 10412.5 9467.5 ;
      RECT  10477.5 8447.5 10412.5 8582.5 ;
      RECT  10287.5 8447.5 10222.5 8582.5 ;
      RECT  10287.5 8447.5 10222.5 8582.5 ;
      RECT  10477.5 8447.5 10412.5 8582.5 ;
      RECT  10117.5 9422.5 10052.5 9557.5 ;
      RECT  10117.5 8447.5 10052.5 8582.5 ;
      RECT  10420.0 8890.0 10355.0 9025.0 ;
      RECT  10420.0 8890.0 10355.0 9025.0 ;
      RECT  10255.0 8925.0 10190.0 8990.0 ;
      RECT  10545.0 9642.5 9985.0 9707.5 ;
      RECT  10545.0 8297.5 9985.0 8362.5 ;
      RECT  10117.5 9860.0 10052.5 9675.0 ;
      RECT  10117.5 11020.0 10052.5 10835.0 ;
      RECT  10477.5 10902.5 10412.5 11052.5 ;
      RECT  10477.5 10017.5 10412.5 9642.5 ;
      RECT  10287.5 10902.5 10222.5 10017.5 ;
      RECT  10477.5 10017.5 10412.5 9882.5 ;
      RECT  10287.5 10017.5 10222.5 9882.5 ;
      RECT  10287.5 10017.5 10222.5 9882.5 ;
      RECT  10477.5 10017.5 10412.5 9882.5 ;
      RECT  10477.5 10902.5 10412.5 10767.5 ;
      RECT  10287.5 10902.5 10222.5 10767.5 ;
      RECT  10287.5 10902.5 10222.5 10767.5 ;
      RECT  10477.5 10902.5 10412.5 10767.5 ;
      RECT  10117.5 9927.5 10052.5 9792.5 ;
      RECT  10117.5 10902.5 10052.5 10767.5 ;
      RECT  10420.0 10460.0 10355.0 10325.0 ;
      RECT  10420.0 10460.0 10355.0 10325.0 ;
      RECT  10255.0 10425.0 10190.0 10360.0 ;
      RECT  10545.0 9707.5 9985.0 9642.5 ;
      RECT  10545.0 11052.5 9985.0 10987.5 ;
      RECT  7262.5 9490.0 7197.5 9675.0 ;
      RECT  7262.5 8330.0 7197.5 8515.0 ;
      RECT  7622.5 8447.5 7557.5 8297.5 ;
      RECT  7622.5 9332.5 7557.5 9707.5 ;
      RECT  7432.5 8447.5 7367.5 9332.5 ;
      RECT  7622.5 9332.5 7557.5 9467.5 ;
      RECT  7432.5 9332.5 7367.5 9467.5 ;
      RECT  7432.5 9332.5 7367.5 9467.5 ;
      RECT  7622.5 9332.5 7557.5 9467.5 ;
      RECT  7622.5 8447.5 7557.5 8582.5 ;
      RECT  7432.5 8447.5 7367.5 8582.5 ;
      RECT  7432.5 8447.5 7367.5 8582.5 ;
      RECT  7622.5 8447.5 7557.5 8582.5 ;
      RECT  7262.5 9422.5 7197.5 9557.5 ;
      RECT  7262.5 8447.5 7197.5 8582.5 ;
      RECT  7565.0 8890.0 7500.0 9025.0 ;
      RECT  7565.0 8890.0 7500.0 9025.0 ;
      RECT  7400.0 8925.0 7335.0 8990.0 ;
      RECT  7690.0 9642.5 7130.0 9707.5 ;
      RECT  7690.0 8297.5 7130.0 8362.5 ;
      RECT  7262.5 9860.0 7197.5 9675.0 ;
      RECT  7262.5 11020.0 7197.5 10835.0 ;
      RECT  7622.5 10902.5 7557.5 11052.5 ;
      RECT  7622.5 10017.5 7557.5 9642.5 ;
      RECT  7432.5 10902.5 7367.5 10017.5 ;
      RECT  7622.5 10017.5 7557.5 9882.5 ;
      RECT  7432.5 10017.5 7367.5 9882.5 ;
      RECT  7432.5 10017.5 7367.5 9882.5 ;
      RECT  7622.5 10017.5 7557.5 9882.5 ;
      RECT  7622.5 10902.5 7557.5 10767.5 ;
      RECT  7432.5 10902.5 7367.5 10767.5 ;
      RECT  7432.5 10902.5 7367.5 10767.5 ;
      RECT  7622.5 10902.5 7557.5 10767.5 ;
      RECT  7262.5 9927.5 7197.5 9792.5 ;
      RECT  7262.5 10902.5 7197.5 10767.5 ;
      RECT  7565.0 10460.0 7500.0 10325.0 ;
      RECT  7565.0 10460.0 7500.0 10325.0 ;
      RECT  7400.0 10425.0 7335.0 10360.0 ;
      RECT  7690.0 9707.5 7130.0 9642.5 ;
      RECT  7690.0 11052.5 7130.0 10987.5 ;
      RECT  7262.5 12180.0 7197.5 12365.0 ;
      RECT  7262.5 11020.0 7197.5 11205.0 ;
      RECT  7622.5 11137.5 7557.5 10987.5 ;
      RECT  7622.5 12022.5 7557.5 12397.5 ;
      RECT  7432.5 11137.5 7367.5 12022.5 ;
      RECT  7622.5 12022.5 7557.5 12157.5 ;
      RECT  7432.5 12022.5 7367.5 12157.5 ;
      RECT  7432.5 12022.5 7367.5 12157.5 ;
      RECT  7622.5 12022.5 7557.5 12157.5 ;
      RECT  7622.5 11137.5 7557.5 11272.5 ;
      RECT  7432.5 11137.5 7367.5 11272.5 ;
      RECT  7432.5 11137.5 7367.5 11272.5 ;
      RECT  7622.5 11137.5 7557.5 11272.5 ;
      RECT  7262.5 12112.5 7197.5 12247.5 ;
      RECT  7262.5 11137.5 7197.5 11272.5 ;
      RECT  7565.0 11580.0 7500.0 11715.0 ;
      RECT  7565.0 11580.0 7500.0 11715.0 ;
      RECT  7400.0 11615.0 7335.0 11680.0 ;
      RECT  7690.0 12332.5 7130.0 12397.5 ;
      RECT  7690.0 10987.5 7130.0 11052.5 ;
      RECT  7262.5 12550.0 7197.5 12365.0 ;
      RECT  7262.5 13710.0 7197.5 13525.0 ;
      RECT  7622.5 13592.5 7557.5 13742.5 ;
      RECT  7622.5 12707.5 7557.5 12332.5 ;
      RECT  7432.5 13592.5 7367.5 12707.5 ;
      RECT  7622.5 12707.5 7557.5 12572.5 ;
      RECT  7432.5 12707.5 7367.5 12572.5 ;
      RECT  7432.5 12707.5 7367.5 12572.5 ;
      RECT  7622.5 12707.5 7557.5 12572.5 ;
      RECT  7622.5 13592.5 7557.5 13457.5 ;
      RECT  7432.5 13592.5 7367.5 13457.5 ;
      RECT  7432.5 13592.5 7367.5 13457.5 ;
      RECT  7622.5 13592.5 7557.5 13457.5 ;
      RECT  7262.5 12617.5 7197.5 12482.5 ;
      RECT  7262.5 13592.5 7197.5 13457.5 ;
      RECT  7565.0 13150.0 7500.0 13015.0 ;
      RECT  7565.0 13150.0 7500.0 13015.0 ;
      RECT  7400.0 13115.0 7335.0 13050.0 ;
      RECT  7690.0 12397.5 7130.0 12332.5 ;
      RECT  7690.0 13742.5 7130.0 13677.5 ;
      RECT  8542.5 8492.5 8477.5 8297.5 ;
      RECT  8542.5 9332.5 8477.5 9707.5 ;
      RECT  8162.5 9332.5 8097.5 9707.5 ;
      RECT  7992.5 9490.0 7927.5 9675.0 ;
      RECT  7992.5 8330.0 7927.5 8515.0 ;
      RECT  8542.5 9332.5 8477.5 9467.5 ;
      RECT  8352.5 9332.5 8287.5 9467.5 ;
      RECT  8352.5 9332.5 8287.5 9467.5 ;
      RECT  8542.5 9332.5 8477.5 9467.5 ;
      RECT  8352.5 9332.5 8287.5 9467.5 ;
      RECT  8162.5 9332.5 8097.5 9467.5 ;
      RECT  8162.5 9332.5 8097.5 9467.5 ;
      RECT  8352.5 9332.5 8287.5 9467.5 ;
      RECT  8542.5 8492.5 8477.5 8627.5 ;
      RECT  8352.5 8492.5 8287.5 8627.5 ;
      RECT  8352.5 8492.5 8287.5 8627.5 ;
      RECT  8542.5 8492.5 8477.5 8627.5 ;
      RECT  8352.5 8492.5 8287.5 8627.5 ;
      RECT  8162.5 8492.5 8097.5 8627.5 ;
      RECT  8162.5 8492.5 8097.5 8627.5 ;
      RECT  8352.5 8492.5 8287.5 8627.5 ;
      RECT  7992.5 9422.5 7927.5 9557.5 ;
      RECT  7992.5 8447.5 7927.5 8582.5 ;
      RECT  8157.5 8722.5 8292.5 8787.5 ;
      RECT  8415.0 8937.5 8550.0 9002.5 ;
      RECT  8352.5 9332.5 8287.5 9467.5 ;
      RECT  8162.5 8492.5 8097.5 8627.5 ;
      RECT  8062.5 8937.5 8197.5 9002.5 ;
      RECT  8550.0 8937.5 8415.0 9002.5 ;
      RECT  8292.5 8722.5 8157.5 8787.5 ;
      RECT  8197.5 8937.5 8062.5 9002.5 ;
      RECT  8610.0 9642.5 7690.0 9707.5 ;
      RECT  8610.0 8297.5 7690.0 8362.5 ;
      RECT  8542.5 10857.5 8477.5 11052.5 ;
      RECT  8542.5 10017.5 8477.5 9642.5 ;
      RECT  8162.5 10017.5 8097.5 9642.5 ;
      RECT  7992.5 9860.0 7927.5 9675.0 ;
      RECT  7992.5 11020.0 7927.5 10835.0 ;
      RECT  8542.5 10017.5 8477.5 9882.5 ;
      RECT  8352.5 10017.5 8287.5 9882.5 ;
      RECT  8352.5 10017.5 8287.5 9882.5 ;
      RECT  8542.5 10017.5 8477.5 9882.5 ;
      RECT  8352.5 10017.5 8287.5 9882.5 ;
      RECT  8162.5 10017.5 8097.5 9882.5 ;
      RECT  8162.5 10017.5 8097.5 9882.5 ;
      RECT  8352.5 10017.5 8287.5 9882.5 ;
      RECT  8542.5 10857.5 8477.5 10722.5 ;
      RECT  8352.5 10857.5 8287.5 10722.5 ;
      RECT  8352.5 10857.5 8287.5 10722.5 ;
      RECT  8542.5 10857.5 8477.5 10722.5 ;
      RECT  8352.5 10857.5 8287.5 10722.5 ;
      RECT  8162.5 10857.5 8097.5 10722.5 ;
      RECT  8162.5 10857.5 8097.5 10722.5 ;
      RECT  8352.5 10857.5 8287.5 10722.5 ;
      RECT  7992.5 9927.5 7927.5 9792.5 ;
      RECT  7992.5 10902.5 7927.5 10767.5 ;
      RECT  8157.5 10627.5 8292.5 10562.5 ;
      RECT  8415.0 10412.5 8550.0 10347.5 ;
      RECT  8352.5 10017.5 8287.5 9882.5 ;
      RECT  8162.5 10857.5 8097.5 10722.5 ;
      RECT  8062.5 10412.5 8197.5 10347.5 ;
      RECT  8550.0 10412.5 8415.0 10347.5 ;
      RECT  8292.5 10627.5 8157.5 10562.5 ;
      RECT  8197.5 10412.5 8062.5 10347.5 ;
      RECT  8610.0 9707.5 7690.0 9642.5 ;
      RECT  8610.0 11052.5 7690.0 10987.5 ;
      RECT  8542.5 11182.5 8477.5 10987.5 ;
      RECT  8542.5 12022.5 8477.5 12397.5 ;
      RECT  8162.5 12022.5 8097.5 12397.5 ;
      RECT  7992.5 12180.0 7927.5 12365.0 ;
      RECT  7992.5 11020.0 7927.5 11205.0 ;
      RECT  8542.5 12022.5 8477.5 12157.5 ;
      RECT  8352.5 12022.5 8287.5 12157.5 ;
      RECT  8352.5 12022.5 8287.5 12157.5 ;
      RECT  8542.5 12022.5 8477.5 12157.5 ;
      RECT  8352.5 12022.5 8287.5 12157.5 ;
      RECT  8162.5 12022.5 8097.5 12157.5 ;
      RECT  8162.5 12022.5 8097.5 12157.5 ;
      RECT  8352.5 12022.5 8287.5 12157.5 ;
      RECT  8542.5 11182.5 8477.5 11317.5 ;
      RECT  8352.5 11182.5 8287.5 11317.5 ;
      RECT  8352.5 11182.5 8287.5 11317.5 ;
      RECT  8542.5 11182.5 8477.5 11317.5 ;
      RECT  8352.5 11182.5 8287.5 11317.5 ;
      RECT  8162.5 11182.5 8097.5 11317.5 ;
      RECT  8162.5 11182.5 8097.5 11317.5 ;
      RECT  8352.5 11182.5 8287.5 11317.5 ;
      RECT  7992.5 12112.5 7927.5 12247.5 ;
      RECT  7992.5 11137.5 7927.5 11272.5 ;
      RECT  8157.5 11412.5 8292.5 11477.5 ;
      RECT  8415.0 11627.5 8550.0 11692.5 ;
      RECT  8352.5 12022.5 8287.5 12157.5 ;
      RECT  8162.5 11182.5 8097.5 11317.5 ;
      RECT  8062.5 11627.5 8197.5 11692.5 ;
      RECT  8550.0 11627.5 8415.0 11692.5 ;
      RECT  8292.5 11412.5 8157.5 11477.5 ;
      RECT  8197.5 11627.5 8062.5 11692.5 ;
      RECT  8610.0 12332.5 7690.0 12397.5 ;
      RECT  8610.0 10987.5 7690.0 11052.5 ;
      RECT  8542.5 13547.5 8477.5 13742.5 ;
      RECT  8542.5 12707.5 8477.5 12332.5 ;
      RECT  8162.5 12707.5 8097.5 12332.5 ;
      RECT  7992.5 12550.0 7927.5 12365.0 ;
      RECT  7992.5 13710.0 7927.5 13525.0 ;
      RECT  8542.5 12707.5 8477.5 12572.5 ;
      RECT  8352.5 12707.5 8287.5 12572.5 ;
      RECT  8352.5 12707.5 8287.5 12572.5 ;
      RECT  8542.5 12707.5 8477.5 12572.5 ;
      RECT  8352.5 12707.5 8287.5 12572.5 ;
      RECT  8162.5 12707.5 8097.5 12572.5 ;
      RECT  8162.5 12707.5 8097.5 12572.5 ;
      RECT  8352.5 12707.5 8287.5 12572.5 ;
      RECT  8542.5 13547.5 8477.5 13412.5 ;
      RECT  8352.5 13547.5 8287.5 13412.5 ;
      RECT  8352.5 13547.5 8287.5 13412.5 ;
      RECT  8542.5 13547.5 8477.5 13412.5 ;
      RECT  8352.5 13547.5 8287.5 13412.5 ;
      RECT  8162.5 13547.5 8097.5 13412.5 ;
      RECT  8162.5 13547.5 8097.5 13412.5 ;
      RECT  8352.5 13547.5 8287.5 13412.5 ;
      RECT  7992.5 12617.5 7927.5 12482.5 ;
      RECT  7992.5 13592.5 7927.5 13457.5 ;
      RECT  8157.5 13317.5 8292.5 13252.5 ;
      RECT  8415.0 13102.5 8550.0 13037.5 ;
      RECT  8352.5 12707.5 8287.5 12572.5 ;
      RECT  8162.5 13547.5 8097.5 13412.5 ;
      RECT  8062.5 13102.5 8197.5 13037.5 ;
      RECT  8550.0 13102.5 8415.0 13037.5 ;
      RECT  8292.5 13317.5 8157.5 13252.5 ;
      RECT  8197.5 13102.5 8062.5 13037.5 ;
      RECT  8610.0 12397.5 7690.0 12332.5 ;
      RECT  8610.0 13742.5 7690.0 13677.5 ;
      RECT  9607.5 9447.5 9742.5 9512.5 ;
      RECT  10992.5 8925.0 11127.5 8990.0 ;
      RECT  9332.5 10792.5 9467.5 10857.5 ;
      RECT  10717.5 10360.0 10852.5 10425.0 ;
      RECT  10992.5 11122.5 11127.5 11187.5 ;
      RECT  9057.5 11122.5 9192.5 11187.5 ;
      RECT  10717.5 12467.5 10852.5 12532.5 ;
      RECT  8782.5 12467.5 8917.5 12532.5 ;
      RECT  9607.5 8937.5 9742.5 9002.5 ;
      RECT  9332.5 8722.5 9467.5 8787.5 ;
      RECT  9057.5 10347.5 9192.5 10412.5 ;
      RECT  9332.5 10562.5 9467.5 10627.5 ;
      RECT  9607.5 11627.5 9742.5 11692.5 ;
      RECT  8782.5 11412.5 8917.5 11477.5 ;
      RECT  9057.5 13037.5 9192.5 13102.5 ;
      RECT  8782.5 13252.5 8917.5 13317.5 ;
      RECT  7335.0 8925.0 7130.0 8990.0 ;
      RECT  7335.0 10360.0 7130.0 10425.0 ;
      RECT  7335.0 11615.0 7130.0 11680.0 ;
      RECT  7335.0 13050.0 7130.0 13115.0 ;
      RECT  11095.0 9642.5 7130.0 9707.5 ;
      RECT  11095.0 12332.5 7130.0 12397.5 ;
      RECT  11095.0 8297.5 7130.0 8362.5 ;
      RECT  11095.0 10987.5 7130.0 11052.5 ;
      RECT  11095.0 13677.5 7130.0 13742.5 ;
      RECT  9952.5 14305.0 9887.5 14370.0 ;
      RECT  9952.5 14827.5 9887.5 14892.5 ;
      RECT  10190.0 14305.0 9920.0 14370.0 ;
      RECT  9952.5 14337.5 9887.5 14860.0 ;
      RECT  9920.0 14827.5 9675.0 14892.5 ;
      RECT  11060.0 14305.0 10420.0 14370.0 ;
      RECT  9952.5 15740.0 9887.5 15805.0 ;
      RECT  9952.5 16172.5 9887.5 16237.5 ;
      RECT  10190.0 15740.0 9920.0 15805.0 ;
      RECT  9952.5 15772.5 9887.5 16205.0 ;
      RECT  9920.0 16172.5 9400.0 16237.5 ;
      RECT  10785.0 15740.0 10420.0 15805.0 ;
      RECT  11060.0 16502.5 9125.0 16567.5 ;
      RECT  10785.0 17847.5 8850.0 17912.5 ;
      RECT  9675.0 14317.5 8550.0 14382.5 ;
      RECT  9400.0 14102.5 8292.5 14167.5 ;
      RECT  9125.0 15727.5 8550.0 15792.5 ;
      RECT  9400.0 15942.5 8292.5 16007.5 ;
      RECT  9675.0 17007.5 8550.0 17072.5 ;
      RECT  8850.0 16792.5 8292.5 16857.5 ;
      RECT  9125.0 18417.5 8550.0 18482.5 ;
      RECT  8850.0 18632.5 8292.5 18697.5 ;
      RECT  7845.0 14317.5 7780.0 14382.5 ;
      RECT  7845.0 14305.0 7780.0 14370.0 ;
      RECT  8062.5 14317.5 7812.5 14382.5 ;
      RECT  7845.0 14337.5 7780.0 14350.0 ;
      RECT  7812.5 14305.0 7565.0 14370.0 ;
      RECT  7845.0 15727.5 7780.0 15792.5 ;
      RECT  7845.0 15740.0 7780.0 15805.0 ;
      RECT  8062.5 15727.5 7812.5 15792.5 ;
      RECT  7845.0 15760.0 7780.0 15772.5 ;
      RECT  7812.5 15740.0 7565.0 15805.0 ;
      RECT  7845.0 17007.5 7780.0 17072.5 ;
      RECT  7845.0 16995.0 7780.0 17060.0 ;
      RECT  8062.5 17007.5 7812.5 17072.5 ;
      RECT  7845.0 17027.5 7780.0 17040.0 ;
      RECT  7812.5 16995.0 7565.0 17060.0 ;
      RECT  7845.0 18417.5 7780.0 18482.5 ;
      RECT  7845.0 18430.0 7780.0 18495.0 ;
      RECT  8062.5 18417.5 7812.5 18482.5 ;
      RECT  7845.0 18450.0 7780.0 18462.5 ;
      RECT  7812.5 18430.0 7565.0 18495.0 ;
      RECT  10117.5 14870.0 10052.5 15055.0 ;
      RECT  10117.5 13710.0 10052.5 13895.0 ;
      RECT  10477.5 13827.5 10412.5 13677.5 ;
      RECT  10477.5 14712.5 10412.5 15087.5 ;
      RECT  10287.5 13827.5 10222.5 14712.5 ;
      RECT  10477.5 14712.5 10412.5 14847.5 ;
      RECT  10287.5 14712.5 10222.5 14847.5 ;
      RECT  10287.5 14712.5 10222.5 14847.5 ;
      RECT  10477.5 14712.5 10412.5 14847.5 ;
      RECT  10477.5 13827.5 10412.5 13962.5 ;
      RECT  10287.5 13827.5 10222.5 13962.5 ;
      RECT  10287.5 13827.5 10222.5 13962.5 ;
      RECT  10477.5 13827.5 10412.5 13962.5 ;
      RECT  10117.5 14802.5 10052.5 14937.5 ;
      RECT  10117.5 13827.5 10052.5 13962.5 ;
      RECT  10420.0 14270.0 10355.0 14405.0 ;
      RECT  10420.0 14270.0 10355.0 14405.0 ;
      RECT  10255.0 14305.0 10190.0 14370.0 ;
      RECT  10545.0 15022.5 9985.0 15087.5 ;
      RECT  10545.0 13677.5 9985.0 13742.5 ;
      RECT  10117.5 15240.0 10052.5 15055.0 ;
      RECT  10117.5 16400.0 10052.5 16215.0 ;
      RECT  10477.5 16282.5 10412.5 16432.5 ;
      RECT  10477.5 15397.5 10412.5 15022.5 ;
      RECT  10287.5 16282.5 10222.5 15397.5 ;
      RECT  10477.5 15397.5 10412.5 15262.5 ;
      RECT  10287.5 15397.5 10222.5 15262.5 ;
      RECT  10287.5 15397.5 10222.5 15262.5 ;
      RECT  10477.5 15397.5 10412.5 15262.5 ;
      RECT  10477.5 16282.5 10412.5 16147.5 ;
      RECT  10287.5 16282.5 10222.5 16147.5 ;
      RECT  10287.5 16282.5 10222.5 16147.5 ;
      RECT  10477.5 16282.5 10412.5 16147.5 ;
      RECT  10117.5 15307.5 10052.5 15172.5 ;
      RECT  10117.5 16282.5 10052.5 16147.5 ;
      RECT  10420.0 15840.0 10355.0 15705.0 ;
      RECT  10420.0 15840.0 10355.0 15705.0 ;
      RECT  10255.0 15805.0 10190.0 15740.0 ;
      RECT  10545.0 15087.5 9985.0 15022.5 ;
      RECT  10545.0 16432.5 9985.0 16367.5 ;
      RECT  7262.5 14870.0 7197.5 15055.0 ;
      RECT  7262.5 13710.0 7197.5 13895.0 ;
      RECT  7622.5 13827.5 7557.5 13677.5 ;
      RECT  7622.5 14712.5 7557.5 15087.5 ;
      RECT  7432.5 13827.5 7367.5 14712.5 ;
      RECT  7622.5 14712.5 7557.5 14847.5 ;
      RECT  7432.5 14712.5 7367.5 14847.5 ;
      RECT  7432.5 14712.5 7367.5 14847.5 ;
      RECT  7622.5 14712.5 7557.5 14847.5 ;
      RECT  7622.5 13827.5 7557.5 13962.5 ;
      RECT  7432.5 13827.5 7367.5 13962.5 ;
      RECT  7432.5 13827.5 7367.5 13962.5 ;
      RECT  7622.5 13827.5 7557.5 13962.5 ;
      RECT  7262.5 14802.5 7197.5 14937.5 ;
      RECT  7262.5 13827.5 7197.5 13962.5 ;
      RECT  7565.0 14270.0 7500.0 14405.0 ;
      RECT  7565.0 14270.0 7500.0 14405.0 ;
      RECT  7400.0 14305.0 7335.0 14370.0 ;
      RECT  7690.0 15022.5 7130.0 15087.5 ;
      RECT  7690.0 13677.5 7130.0 13742.5 ;
      RECT  7262.5 15240.0 7197.5 15055.0 ;
      RECT  7262.5 16400.0 7197.5 16215.0 ;
      RECT  7622.5 16282.5 7557.5 16432.5 ;
      RECT  7622.5 15397.5 7557.5 15022.5 ;
      RECT  7432.5 16282.5 7367.5 15397.5 ;
      RECT  7622.5 15397.5 7557.5 15262.5 ;
      RECT  7432.5 15397.5 7367.5 15262.5 ;
      RECT  7432.5 15397.5 7367.5 15262.5 ;
      RECT  7622.5 15397.5 7557.5 15262.5 ;
      RECT  7622.5 16282.5 7557.5 16147.5 ;
      RECT  7432.5 16282.5 7367.5 16147.5 ;
      RECT  7432.5 16282.5 7367.5 16147.5 ;
      RECT  7622.5 16282.5 7557.5 16147.5 ;
      RECT  7262.5 15307.5 7197.5 15172.5 ;
      RECT  7262.5 16282.5 7197.5 16147.5 ;
      RECT  7565.0 15840.0 7500.0 15705.0 ;
      RECT  7565.0 15840.0 7500.0 15705.0 ;
      RECT  7400.0 15805.0 7335.0 15740.0 ;
      RECT  7690.0 15087.5 7130.0 15022.5 ;
      RECT  7690.0 16432.5 7130.0 16367.5 ;
      RECT  7262.5 17560.0 7197.5 17745.0 ;
      RECT  7262.5 16400.0 7197.5 16585.0 ;
      RECT  7622.5 16517.5 7557.5 16367.5 ;
      RECT  7622.5 17402.5 7557.5 17777.5 ;
      RECT  7432.5 16517.5 7367.5 17402.5 ;
      RECT  7622.5 17402.5 7557.5 17537.5 ;
      RECT  7432.5 17402.5 7367.5 17537.5 ;
      RECT  7432.5 17402.5 7367.5 17537.5 ;
      RECT  7622.5 17402.5 7557.5 17537.5 ;
      RECT  7622.5 16517.5 7557.5 16652.5 ;
      RECT  7432.5 16517.5 7367.5 16652.5 ;
      RECT  7432.5 16517.5 7367.5 16652.5 ;
      RECT  7622.5 16517.5 7557.5 16652.5 ;
      RECT  7262.5 17492.5 7197.5 17627.5 ;
      RECT  7262.5 16517.5 7197.5 16652.5 ;
      RECT  7565.0 16960.0 7500.0 17095.0 ;
      RECT  7565.0 16960.0 7500.0 17095.0 ;
      RECT  7400.0 16995.0 7335.0 17060.0 ;
      RECT  7690.0 17712.5 7130.0 17777.5 ;
      RECT  7690.0 16367.5 7130.0 16432.5 ;
      RECT  7262.5 17930.0 7197.5 17745.0 ;
      RECT  7262.5 19090.0 7197.5 18905.0 ;
      RECT  7622.5 18972.5 7557.5 19122.5 ;
      RECT  7622.5 18087.5 7557.5 17712.5 ;
      RECT  7432.5 18972.5 7367.5 18087.5 ;
      RECT  7622.5 18087.5 7557.5 17952.5 ;
      RECT  7432.5 18087.5 7367.5 17952.5 ;
      RECT  7432.5 18087.5 7367.5 17952.5 ;
      RECT  7622.5 18087.5 7557.5 17952.5 ;
      RECT  7622.5 18972.5 7557.5 18837.5 ;
      RECT  7432.5 18972.5 7367.5 18837.5 ;
      RECT  7432.5 18972.5 7367.5 18837.5 ;
      RECT  7622.5 18972.5 7557.5 18837.5 ;
      RECT  7262.5 17997.5 7197.5 17862.5 ;
      RECT  7262.5 18972.5 7197.5 18837.5 ;
      RECT  7565.0 18530.0 7500.0 18395.0 ;
      RECT  7565.0 18530.0 7500.0 18395.0 ;
      RECT  7400.0 18495.0 7335.0 18430.0 ;
      RECT  7690.0 17777.5 7130.0 17712.5 ;
      RECT  7690.0 19122.5 7130.0 19057.5 ;
      RECT  8542.5 13872.5 8477.5 13677.5 ;
      RECT  8542.5 14712.5 8477.5 15087.5 ;
      RECT  8162.5 14712.5 8097.5 15087.5 ;
      RECT  7992.5 14870.0 7927.5 15055.0 ;
      RECT  7992.5 13710.0 7927.5 13895.0 ;
      RECT  8542.5 14712.5 8477.5 14847.5 ;
      RECT  8352.5 14712.5 8287.5 14847.5 ;
      RECT  8352.5 14712.5 8287.5 14847.5 ;
      RECT  8542.5 14712.5 8477.5 14847.5 ;
      RECT  8352.5 14712.5 8287.5 14847.5 ;
      RECT  8162.5 14712.5 8097.5 14847.5 ;
      RECT  8162.5 14712.5 8097.5 14847.5 ;
      RECT  8352.5 14712.5 8287.5 14847.5 ;
      RECT  8542.5 13872.5 8477.5 14007.5 ;
      RECT  8352.5 13872.5 8287.5 14007.5 ;
      RECT  8352.5 13872.5 8287.5 14007.5 ;
      RECT  8542.5 13872.5 8477.5 14007.5 ;
      RECT  8352.5 13872.5 8287.5 14007.5 ;
      RECT  8162.5 13872.5 8097.5 14007.5 ;
      RECT  8162.5 13872.5 8097.5 14007.5 ;
      RECT  8352.5 13872.5 8287.5 14007.5 ;
      RECT  7992.5 14802.5 7927.5 14937.5 ;
      RECT  7992.5 13827.5 7927.5 13962.5 ;
      RECT  8157.5 14102.5 8292.5 14167.5 ;
      RECT  8415.0 14317.5 8550.0 14382.5 ;
      RECT  8352.5 14712.5 8287.5 14847.5 ;
      RECT  8162.5 13872.5 8097.5 14007.5 ;
      RECT  8062.5 14317.5 8197.5 14382.5 ;
      RECT  8550.0 14317.5 8415.0 14382.5 ;
      RECT  8292.5 14102.5 8157.5 14167.5 ;
      RECT  8197.5 14317.5 8062.5 14382.5 ;
      RECT  8610.0 15022.5 7690.0 15087.5 ;
      RECT  8610.0 13677.5 7690.0 13742.5 ;
      RECT  8542.5 16237.5 8477.5 16432.5 ;
      RECT  8542.5 15397.5 8477.5 15022.5 ;
      RECT  8162.5 15397.5 8097.5 15022.5 ;
      RECT  7992.5 15240.0 7927.5 15055.0 ;
      RECT  7992.5 16400.0 7927.5 16215.0 ;
      RECT  8542.5 15397.5 8477.5 15262.5 ;
      RECT  8352.5 15397.5 8287.5 15262.5 ;
      RECT  8352.5 15397.5 8287.5 15262.5 ;
      RECT  8542.5 15397.5 8477.5 15262.5 ;
      RECT  8352.5 15397.5 8287.5 15262.5 ;
      RECT  8162.5 15397.5 8097.5 15262.5 ;
      RECT  8162.5 15397.5 8097.5 15262.5 ;
      RECT  8352.5 15397.5 8287.5 15262.5 ;
      RECT  8542.5 16237.5 8477.5 16102.5 ;
      RECT  8352.5 16237.5 8287.5 16102.5 ;
      RECT  8352.5 16237.5 8287.5 16102.5 ;
      RECT  8542.5 16237.5 8477.5 16102.5 ;
      RECT  8352.5 16237.5 8287.5 16102.5 ;
      RECT  8162.5 16237.5 8097.5 16102.5 ;
      RECT  8162.5 16237.5 8097.5 16102.5 ;
      RECT  8352.5 16237.5 8287.5 16102.5 ;
      RECT  7992.5 15307.5 7927.5 15172.5 ;
      RECT  7992.5 16282.5 7927.5 16147.5 ;
      RECT  8157.5 16007.5 8292.5 15942.5 ;
      RECT  8415.0 15792.5 8550.0 15727.5 ;
      RECT  8352.5 15397.5 8287.5 15262.5 ;
      RECT  8162.5 16237.5 8097.5 16102.5 ;
      RECT  8062.5 15792.5 8197.5 15727.5 ;
      RECT  8550.0 15792.5 8415.0 15727.5 ;
      RECT  8292.5 16007.5 8157.5 15942.5 ;
      RECT  8197.5 15792.5 8062.5 15727.5 ;
      RECT  8610.0 15087.5 7690.0 15022.5 ;
      RECT  8610.0 16432.5 7690.0 16367.5 ;
      RECT  8542.5 16562.5 8477.5 16367.5 ;
      RECT  8542.5 17402.5 8477.5 17777.5 ;
      RECT  8162.5 17402.5 8097.5 17777.5 ;
      RECT  7992.5 17560.0 7927.5 17745.0 ;
      RECT  7992.5 16400.0 7927.5 16585.0 ;
      RECT  8542.5 17402.5 8477.5 17537.5 ;
      RECT  8352.5 17402.5 8287.5 17537.5 ;
      RECT  8352.5 17402.5 8287.5 17537.5 ;
      RECT  8542.5 17402.5 8477.5 17537.5 ;
      RECT  8352.5 17402.5 8287.5 17537.5 ;
      RECT  8162.5 17402.5 8097.5 17537.5 ;
      RECT  8162.5 17402.5 8097.5 17537.5 ;
      RECT  8352.5 17402.5 8287.5 17537.5 ;
      RECT  8542.5 16562.5 8477.5 16697.5 ;
      RECT  8352.5 16562.5 8287.5 16697.5 ;
      RECT  8352.5 16562.5 8287.5 16697.5 ;
      RECT  8542.5 16562.5 8477.5 16697.5 ;
      RECT  8352.5 16562.5 8287.5 16697.5 ;
      RECT  8162.5 16562.5 8097.5 16697.5 ;
      RECT  8162.5 16562.5 8097.5 16697.5 ;
      RECT  8352.5 16562.5 8287.5 16697.5 ;
      RECT  7992.5 17492.5 7927.5 17627.5 ;
      RECT  7992.5 16517.5 7927.5 16652.5 ;
      RECT  8157.5 16792.5 8292.5 16857.5 ;
      RECT  8415.0 17007.5 8550.0 17072.5 ;
      RECT  8352.5 17402.5 8287.5 17537.5 ;
      RECT  8162.5 16562.5 8097.5 16697.5 ;
      RECT  8062.5 17007.5 8197.5 17072.5 ;
      RECT  8550.0 17007.5 8415.0 17072.5 ;
      RECT  8292.5 16792.5 8157.5 16857.5 ;
      RECT  8197.5 17007.5 8062.5 17072.5 ;
      RECT  8610.0 17712.5 7690.0 17777.5 ;
      RECT  8610.0 16367.5 7690.0 16432.5 ;
      RECT  8542.5 18927.5 8477.5 19122.5 ;
      RECT  8542.5 18087.5 8477.5 17712.5 ;
      RECT  8162.5 18087.5 8097.5 17712.5 ;
      RECT  7992.5 17930.0 7927.5 17745.0 ;
      RECT  7992.5 19090.0 7927.5 18905.0 ;
      RECT  8542.5 18087.5 8477.5 17952.5 ;
      RECT  8352.5 18087.5 8287.5 17952.5 ;
      RECT  8352.5 18087.5 8287.5 17952.5 ;
      RECT  8542.5 18087.5 8477.5 17952.5 ;
      RECT  8352.5 18087.5 8287.5 17952.5 ;
      RECT  8162.5 18087.5 8097.5 17952.5 ;
      RECT  8162.5 18087.5 8097.5 17952.5 ;
      RECT  8352.5 18087.5 8287.5 17952.5 ;
      RECT  8542.5 18927.5 8477.5 18792.5 ;
      RECT  8352.5 18927.5 8287.5 18792.5 ;
      RECT  8352.5 18927.5 8287.5 18792.5 ;
      RECT  8542.5 18927.5 8477.5 18792.5 ;
      RECT  8352.5 18927.5 8287.5 18792.5 ;
      RECT  8162.5 18927.5 8097.5 18792.5 ;
      RECT  8162.5 18927.5 8097.5 18792.5 ;
      RECT  8352.5 18927.5 8287.5 18792.5 ;
      RECT  7992.5 17997.5 7927.5 17862.5 ;
      RECT  7992.5 18972.5 7927.5 18837.5 ;
      RECT  8157.5 18697.5 8292.5 18632.5 ;
      RECT  8415.0 18482.5 8550.0 18417.5 ;
      RECT  8352.5 18087.5 8287.5 17952.5 ;
      RECT  8162.5 18927.5 8097.5 18792.5 ;
      RECT  8062.5 18482.5 8197.5 18417.5 ;
      RECT  8550.0 18482.5 8415.0 18417.5 ;
      RECT  8292.5 18697.5 8157.5 18632.5 ;
      RECT  8197.5 18482.5 8062.5 18417.5 ;
      RECT  8610.0 17777.5 7690.0 17712.5 ;
      RECT  8610.0 19122.5 7690.0 19057.5 ;
      RECT  9607.5 14827.5 9742.5 14892.5 ;
      RECT  10992.5 14305.0 11127.5 14370.0 ;
      RECT  9332.5 16172.5 9467.5 16237.5 ;
      RECT  10717.5 15740.0 10852.5 15805.0 ;
      RECT  10992.5 16502.5 11127.5 16567.5 ;
      RECT  9057.5 16502.5 9192.5 16567.5 ;
      RECT  10717.5 17847.5 10852.5 17912.5 ;
      RECT  8782.5 17847.5 8917.5 17912.5 ;
      RECT  9607.5 14317.5 9742.5 14382.5 ;
      RECT  9332.5 14102.5 9467.5 14167.5 ;
      RECT  9057.5 15727.5 9192.5 15792.5 ;
      RECT  9332.5 15942.5 9467.5 16007.5 ;
      RECT  9607.5 17007.5 9742.5 17072.5 ;
      RECT  8782.5 16792.5 8917.5 16857.5 ;
      RECT  9057.5 18417.5 9192.5 18482.5 ;
      RECT  8782.5 18632.5 8917.5 18697.5 ;
      RECT  7335.0 14305.0 7130.0 14370.0 ;
      RECT  7335.0 15740.0 7130.0 15805.0 ;
      RECT  7335.0 16995.0 7130.0 17060.0 ;
      RECT  7335.0 18430.0 7130.0 18495.0 ;
      RECT  11095.0 15022.5 7130.0 15087.5 ;
      RECT  11095.0 17712.5 7130.0 17777.5 ;
      RECT  11095.0 13677.5 7130.0 13742.5 ;
      RECT  11095.0 16367.5 7130.0 16432.5 ;
      RECT  11095.0 19057.5 7130.0 19122.5 ;
      RECT  7197.5 19252.5 7262.5 19057.5 ;
      RECT  7197.5 20092.5 7262.5 20467.5 ;
      RECT  7577.5 20092.5 7642.5 20467.5 ;
      RECT  7747.5 20250.0 7812.5 20435.0 ;
      RECT  7747.5 19090.0 7812.5 19275.0 ;
      RECT  7197.5 20092.5 7262.5 20227.5 ;
      RECT  7387.5 20092.5 7452.5 20227.5 ;
      RECT  7387.5 20092.5 7452.5 20227.5 ;
      RECT  7197.5 20092.5 7262.5 20227.5 ;
      RECT  7387.5 20092.5 7452.5 20227.5 ;
      RECT  7577.5 20092.5 7642.5 20227.5 ;
      RECT  7577.5 20092.5 7642.5 20227.5 ;
      RECT  7387.5 20092.5 7452.5 20227.5 ;
      RECT  7197.5 19252.5 7262.5 19387.5 ;
      RECT  7387.5 19252.5 7452.5 19387.5 ;
      RECT  7387.5 19252.5 7452.5 19387.5 ;
      RECT  7197.5 19252.5 7262.5 19387.5 ;
      RECT  7387.5 19252.5 7452.5 19387.5 ;
      RECT  7577.5 19252.5 7642.5 19387.5 ;
      RECT  7577.5 19252.5 7642.5 19387.5 ;
      RECT  7387.5 19252.5 7452.5 19387.5 ;
      RECT  7747.5 20182.5 7812.5 20317.5 ;
      RECT  7747.5 19207.5 7812.5 19342.5 ;
      RECT  7582.5 19482.5 7447.5 19547.5 ;
      RECT  7325.0 19697.5 7190.0 19762.5 ;
      RECT  7387.5 20092.5 7452.5 20227.5 ;
      RECT  7577.5 19252.5 7642.5 19387.5 ;
      RECT  7677.5 19697.5 7542.5 19762.5 ;
      RECT  7190.0 19697.5 7325.0 19762.5 ;
      RECT  7447.5 19482.5 7582.5 19547.5 ;
      RECT  7542.5 19697.5 7677.5 19762.5 ;
      RECT  7130.0 20402.5 8050.0 20467.5 ;
      RECT  7130.0 19057.5 8050.0 19122.5 ;
      RECT  7197.5 21617.5 7262.5 21812.5 ;
      RECT  7197.5 20777.5 7262.5 20402.5 ;
      RECT  7577.5 20777.5 7642.5 20402.5 ;
      RECT  7747.5 20620.0 7812.5 20435.0 ;
      RECT  7747.5 21780.0 7812.5 21595.0 ;
      RECT  7197.5 20777.5 7262.5 20642.5 ;
      RECT  7387.5 20777.5 7452.5 20642.5 ;
      RECT  7387.5 20777.5 7452.5 20642.5 ;
      RECT  7197.5 20777.5 7262.5 20642.5 ;
      RECT  7387.5 20777.5 7452.5 20642.5 ;
      RECT  7577.5 20777.5 7642.5 20642.5 ;
      RECT  7577.5 20777.5 7642.5 20642.5 ;
      RECT  7387.5 20777.5 7452.5 20642.5 ;
      RECT  7197.5 21617.5 7262.5 21482.5 ;
      RECT  7387.5 21617.5 7452.5 21482.5 ;
      RECT  7387.5 21617.5 7452.5 21482.5 ;
      RECT  7197.5 21617.5 7262.5 21482.5 ;
      RECT  7387.5 21617.5 7452.5 21482.5 ;
      RECT  7577.5 21617.5 7642.5 21482.5 ;
      RECT  7577.5 21617.5 7642.5 21482.5 ;
      RECT  7387.5 21617.5 7452.5 21482.5 ;
      RECT  7747.5 20687.5 7812.5 20552.5 ;
      RECT  7747.5 21662.5 7812.5 21527.5 ;
      RECT  7582.5 21387.5 7447.5 21322.5 ;
      RECT  7325.0 21172.5 7190.0 21107.5 ;
      RECT  7387.5 20777.5 7452.5 20642.5 ;
      RECT  7577.5 21617.5 7642.5 21482.5 ;
      RECT  7677.5 21172.5 7542.5 21107.5 ;
      RECT  7190.0 21172.5 7325.0 21107.5 ;
      RECT  7447.5 21387.5 7582.5 21322.5 ;
      RECT  7542.5 21172.5 7677.5 21107.5 ;
      RECT  7130.0 20467.5 8050.0 20402.5 ;
      RECT  7130.0 21812.5 8050.0 21747.5 ;
      RECT  7197.5 21942.5 7262.5 21747.5 ;
      RECT  7197.5 22782.5 7262.5 23157.5 ;
      RECT  7577.5 22782.5 7642.5 23157.5 ;
      RECT  7747.5 22940.0 7812.5 23125.0 ;
      RECT  7747.5 21780.0 7812.5 21965.0 ;
      RECT  7197.5 22782.5 7262.5 22917.5 ;
      RECT  7387.5 22782.5 7452.5 22917.5 ;
      RECT  7387.5 22782.5 7452.5 22917.5 ;
      RECT  7197.5 22782.5 7262.5 22917.5 ;
      RECT  7387.5 22782.5 7452.5 22917.5 ;
      RECT  7577.5 22782.5 7642.5 22917.5 ;
      RECT  7577.5 22782.5 7642.5 22917.5 ;
      RECT  7387.5 22782.5 7452.5 22917.5 ;
      RECT  7197.5 21942.5 7262.5 22077.5 ;
      RECT  7387.5 21942.5 7452.5 22077.5 ;
      RECT  7387.5 21942.5 7452.5 22077.5 ;
      RECT  7197.5 21942.5 7262.5 22077.5 ;
      RECT  7387.5 21942.5 7452.5 22077.5 ;
      RECT  7577.5 21942.5 7642.5 22077.5 ;
      RECT  7577.5 21942.5 7642.5 22077.5 ;
      RECT  7387.5 21942.5 7452.5 22077.5 ;
      RECT  7747.5 22872.5 7812.5 23007.5 ;
      RECT  7747.5 21897.5 7812.5 22032.5 ;
      RECT  7582.5 22172.5 7447.5 22237.5 ;
      RECT  7325.0 22387.5 7190.0 22452.5 ;
      RECT  7387.5 22782.5 7452.5 22917.5 ;
      RECT  7577.5 21942.5 7642.5 22077.5 ;
      RECT  7677.5 22387.5 7542.5 22452.5 ;
      RECT  7190.0 22387.5 7325.0 22452.5 ;
      RECT  7447.5 22172.5 7582.5 22237.5 ;
      RECT  7542.5 22387.5 7677.5 22452.5 ;
      RECT  7130.0 23092.5 8050.0 23157.5 ;
      RECT  7130.0 21747.5 8050.0 21812.5 ;
      RECT  7197.5 24307.5 7262.5 24502.5 ;
      RECT  7197.5 23467.5 7262.5 23092.5 ;
      RECT  7577.5 23467.5 7642.5 23092.5 ;
      RECT  7747.5 23310.0 7812.5 23125.0 ;
      RECT  7747.5 24470.0 7812.5 24285.0 ;
      RECT  7197.5 23467.5 7262.5 23332.5 ;
      RECT  7387.5 23467.5 7452.5 23332.5 ;
      RECT  7387.5 23467.5 7452.5 23332.5 ;
      RECT  7197.5 23467.5 7262.5 23332.5 ;
      RECT  7387.5 23467.5 7452.5 23332.5 ;
      RECT  7577.5 23467.5 7642.5 23332.5 ;
      RECT  7577.5 23467.5 7642.5 23332.5 ;
      RECT  7387.5 23467.5 7452.5 23332.5 ;
      RECT  7197.5 24307.5 7262.5 24172.5 ;
      RECT  7387.5 24307.5 7452.5 24172.5 ;
      RECT  7387.5 24307.5 7452.5 24172.5 ;
      RECT  7197.5 24307.5 7262.5 24172.5 ;
      RECT  7387.5 24307.5 7452.5 24172.5 ;
      RECT  7577.5 24307.5 7642.5 24172.5 ;
      RECT  7577.5 24307.5 7642.5 24172.5 ;
      RECT  7387.5 24307.5 7452.5 24172.5 ;
      RECT  7747.5 23377.5 7812.5 23242.5 ;
      RECT  7747.5 24352.5 7812.5 24217.5 ;
      RECT  7582.5 24077.5 7447.5 24012.5 ;
      RECT  7325.0 23862.5 7190.0 23797.5 ;
      RECT  7387.5 23467.5 7452.5 23332.5 ;
      RECT  7577.5 24307.5 7642.5 24172.5 ;
      RECT  7677.5 23862.5 7542.5 23797.5 ;
      RECT  7190.0 23862.5 7325.0 23797.5 ;
      RECT  7447.5 24077.5 7582.5 24012.5 ;
      RECT  7542.5 23862.5 7677.5 23797.5 ;
      RECT  7130.0 23157.5 8050.0 23092.5 ;
      RECT  7130.0 24502.5 8050.0 24437.5 ;
      RECT  7197.5 24632.5 7262.5 24437.5 ;
      RECT  7197.5 25472.5 7262.5 25847.5 ;
      RECT  7577.5 25472.5 7642.5 25847.5 ;
      RECT  7747.5 25630.0 7812.5 25815.0 ;
      RECT  7747.5 24470.0 7812.5 24655.0 ;
      RECT  7197.5 25472.5 7262.5 25607.5 ;
      RECT  7387.5 25472.5 7452.5 25607.5 ;
      RECT  7387.5 25472.5 7452.5 25607.5 ;
      RECT  7197.5 25472.5 7262.5 25607.5 ;
      RECT  7387.5 25472.5 7452.5 25607.5 ;
      RECT  7577.5 25472.5 7642.5 25607.5 ;
      RECT  7577.5 25472.5 7642.5 25607.5 ;
      RECT  7387.5 25472.5 7452.5 25607.5 ;
      RECT  7197.5 24632.5 7262.5 24767.5 ;
      RECT  7387.5 24632.5 7452.5 24767.5 ;
      RECT  7387.5 24632.5 7452.5 24767.5 ;
      RECT  7197.5 24632.5 7262.5 24767.5 ;
      RECT  7387.5 24632.5 7452.5 24767.5 ;
      RECT  7577.5 24632.5 7642.5 24767.5 ;
      RECT  7577.5 24632.5 7642.5 24767.5 ;
      RECT  7387.5 24632.5 7452.5 24767.5 ;
      RECT  7747.5 25562.5 7812.5 25697.5 ;
      RECT  7747.5 24587.5 7812.5 24722.5 ;
      RECT  7582.5 24862.5 7447.5 24927.5 ;
      RECT  7325.0 25077.5 7190.0 25142.5 ;
      RECT  7387.5 25472.5 7452.5 25607.5 ;
      RECT  7577.5 24632.5 7642.5 24767.5 ;
      RECT  7677.5 25077.5 7542.5 25142.5 ;
      RECT  7190.0 25077.5 7325.0 25142.5 ;
      RECT  7447.5 24862.5 7582.5 24927.5 ;
      RECT  7542.5 25077.5 7677.5 25142.5 ;
      RECT  7130.0 25782.5 8050.0 25847.5 ;
      RECT  7130.0 24437.5 8050.0 24502.5 ;
      RECT  7197.5 26997.5 7262.5 27192.5 ;
      RECT  7197.5 26157.5 7262.5 25782.5 ;
      RECT  7577.5 26157.5 7642.5 25782.5 ;
      RECT  7747.5 26000.0 7812.5 25815.0 ;
      RECT  7747.5 27160.0 7812.5 26975.0 ;
      RECT  7197.5 26157.5 7262.5 26022.5 ;
      RECT  7387.5 26157.5 7452.5 26022.5 ;
      RECT  7387.5 26157.5 7452.5 26022.5 ;
      RECT  7197.5 26157.5 7262.5 26022.5 ;
      RECT  7387.5 26157.5 7452.5 26022.5 ;
      RECT  7577.5 26157.5 7642.5 26022.5 ;
      RECT  7577.5 26157.5 7642.5 26022.5 ;
      RECT  7387.5 26157.5 7452.5 26022.5 ;
      RECT  7197.5 26997.5 7262.5 26862.5 ;
      RECT  7387.5 26997.5 7452.5 26862.5 ;
      RECT  7387.5 26997.5 7452.5 26862.5 ;
      RECT  7197.5 26997.5 7262.5 26862.5 ;
      RECT  7387.5 26997.5 7452.5 26862.5 ;
      RECT  7577.5 26997.5 7642.5 26862.5 ;
      RECT  7577.5 26997.5 7642.5 26862.5 ;
      RECT  7387.5 26997.5 7452.5 26862.5 ;
      RECT  7747.5 26067.5 7812.5 25932.5 ;
      RECT  7747.5 27042.5 7812.5 26907.5 ;
      RECT  7582.5 26767.5 7447.5 26702.5 ;
      RECT  7325.0 26552.5 7190.0 26487.5 ;
      RECT  7387.5 26157.5 7452.5 26022.5 ;
      RECT  7577.5 26997.5 7642.5 26862.5 ;
      RECT  7677.5 26552.5 7542.5 26487.5 ;
      RECT  7190.0 26552.5 7325.0 26487.5 ;
      RECT  7447.5 26767.5 7582.5 26702.5 ;
      RECT  7542.5 26552.5 7677.5 26487.5 ;
      RECT  7130.0 25847.5 8050.0 25782.5 ;
      RECT  7130.0 27192.5 8050.0 27127.5 ;
      RECT  7197.5 27322.5 7262.5 27127.5 ;
      RECT  7197.5 28162.5 7262.5 28537.5 ;
      RECT  7577.5 28162.5 7642.5 28537.5 ;
      RECT  7747.5 28320.0 7812.5 28505.0 ;
      RECT  7747.5 27160.0 7812.5 27345.0 ;
      RECT  7197.5 28162.5 7262.5 28297.5 ;
      RECT  7387.5 28162.5 7452.5 28297.5 ;
      RECT  7387.5 28162.5 7452.5 28297.5 ;
      RECT  7197.5 28162.5 7262.5 28297.5 ;
      RECT  7387.5 28162.5 7452.5 28297.5 ;
      RECT  7577.5 28162.5 7642.5 28297.5 ;
      RECT  7577.5 28162.5 7642.5 28297.5 ;
      RECT  7387.5 28162.5 7452.5 28297.5 ;
      RECT  7197.5 27322.5 7262.5 27457.5 ;
      RECT  7387.5 27322.5 7452.5 27457.5 ;
      RECT  7387.5 27322.5 7452.5 27457.5 ;
      RECT  7197.5 27322.5 7262.5 27457.5 ;
      RECT  7387.5 27322.5 7452.5 27457.5 ;
      RECT  7577.5 27322.5 7642.5 27457.5 ;
      RECT  7577.5 27322.5 7642.5 27457.5 ;
      RECT  7387.5 27322.5 7452.5 27457.5 ;
      RECT  7747.5 28252.5 7812.5 28387.5 ;
      RECT  7747.5 27277.5 7812.5 27412.5 ;
      RECT  7582.5 27552.5 7447.5 27617.5 ;
      RECT  7325.0 27767.5 7190.0 27832.5 ;
      RECT  7387.5 28162.5 7452.5 28297.5 ;
      RECT  7577.5 27322.5 7642.5 27457.5 ;
      RECT  7677.5 27767.5 7542.5 27832.5 ;
      RECT  7190.0 27767.5 7325.0 27832.5 ;
      RECT  7447.5 27552.5 7582.5 27617.5 ;
      RECT  7542.5 27767.5 7677.5 27832.5 ;
      RECT  7130.0 28472.5 8050.0 28537.5 ;
      RECT  7130.0 27127.5 8050.0 27192.5 ;
      RECT  7197.5 29687.5 7262.5 29882.5 ;
      RECT  7197.5 28847.5 7262.5 28472.5 ;
      RECT  7577.5 28847.5 7642.5 28472.5 ;
      RECT  7747.5 28690.0 7812.5 28505.0 ;
      RECT  7747.5 29850.0 7812.5 29665.0 ;
      RECT  7197.5 28847.5 7262.5 28712.5 ;
      RECT  7387.5 28847.5 7452.5 28712.5 ;
      RECT  7387.5 28847.5 7452.5 28712.5 ;
      RECT  7197.5 28847.5 7262.5 28712.5 ;
      RECT  7387.5 28847.5 7452.5 28712.5 ;
      RECT  7577.5 28847.5 7642.5 28712.5 ;
      RECT  7577.5 28847.5 7642.5 28712.5 ;
      RECT  7387.5 28847.5 7452.5 28712.5 ;
      RECT  7197.5 29687.5 7262.5 29552.5 ;
      RECT  7387.5 29687.5 7452.5 29552.5 ;
      RECT  7387.5 29687.5 7452.5 29552.5 ;
      RECT  7197.5 29687.5 7262.5 29552.5 ;
      RECT  7387.5 29687.5 7452.5 29552.5 ;
      RECT  7577.5 29687.5 7642.5 29552.5 ;
      RECT  7577.5 29687.5 7642.5 29552.5 ;
      RECT  7387.5 29687.5 7452.5 29552.5 ;
      RECT  7747.5 28757.5 7812.5 28622.5 ;
      RECT  7747.5 29732.5 7812.5 29597.5 ;
      RECT  7582.5 29457.5 7447.5 29392.5 ;
      RECT  7325.0 29242.5 7190.0 29177.5 ;
      RECT  7387.5 28847.5 7452.5 28712.5 ;
      RECT  7577.5 29687.5 7642.5 29552.5 ;
      RECT  7677.5 29242.5 7542.5 29177.5 ;
      RECT  7190.0 29242.5 7325.0 29177.5 ;
      RECT  7447.5 29457.5 7582.5 29392.5 ;
      RECT  7542.5 29242.5 7677.5 29177.5 ;
      RECT  7130.0 28537.5 8050.0 28472.5 ;
      RECT  7130.0 29882.5 8050.0 29817.5 ;
      RECT  7197.5 30012.5 7262.5 29817.5 ;
      RECT  7197.5 30852.5 7262.5 31227.5 ;
      RECT  7577.5 30852.5 7642.5 31227.5 ;
      RECT  7747.5 31010.0 7812.5 31195.0 ;
      RECT  7747.5 29850.0 7812.5 30035.0 ;
      RECT  7197.5 30852.5 7262.5 30987.5 ;
      RECT  7387.5 30852.5 7452.5 30987.5 ;
      RECT  7387.5 30852.5 7452.5 30987.5 ;
      RECT  7197.5 30852.5 7262.5 30987.5 ;
      RECT  7387.5 30852.5 7452.5 30987.5 ;
      RECT  7577.5 30852.5 7642.5 30987.5 ;
      RECT  7577.5 30852.5 7642.5 30987.5 ;
      RECT  7387.5 30852.5 7452.5 30987.5 ;
      RECT  7197.5 30012.5 7262.5 30147.5 ;
      RECT  7387.5 30012.5 7452.5 30147.5 ;
      RECT  7387.5 30012.5 7452.5 30147.5 ;
      RECT  7197.5 30012.5 7262.5 30147.5 ;
      RECT  7387.5 30012.5 7452.5 30147.5 ;
      RECT  7577.5 30012.5 7642.5 30147.5 ;
      RECT  7577.5 30012.5 7642.5 30147.5 ;
      RECT  7387.5 30012.5 7452.5 30147.5 ;
      RECT  7747.5 30942.5 7812.5 31077.5 ;
      RECT  7747.5 29967.5 7812.5 30102.5 ;
      RECT  7582.5 30242.5 7447.5 30307.5 ;
      RECT  7325.0 30457.5 7190.0 30522.5 ;
      RECT  7387.5 30852.5 7452.5 30987.5 ;
      RECT  7577.5 30012.5 7642.5 30147.5 ;
      RECT  7677.5 30457.5 7542.5 30522.5 ;
      RECT  7190.0 30457.5 7325.0 30522.5 ;
      RECT  7447.5 30242.5 7582.5 30307.5 ;
      RECT  7542.5 30457.5 7677.5 30522.5 ;
      RECT  7130.0 31162.5 8050.0 31227.5 ;
      RECT  7130.0 29817.5 8050.0 29882.5 ;
      RECT  7197.5 32377.5 7262.5 32572.5 ;
      RECT  7197.5 31537.5 7262.5 31162.5 ;
      RECT  7577.5 31537.5 7642.5 31162.5 ;
      RECT  7747.5 31380.0 7812.5 31195.0 ;
      RECT  7747.5 32540.0 7812.5 32355.0 ;
      RECT  7197.5 31537.5 7262.5 31402.5 ;
      RECT  7387.5 31537.5 7452.5 31402.5 ;
      RECT  7387.5 31537.5 7452.5 31402.5 ;
      RECT  7197.5 31537.5 7262.5 31402.5 ;
      RECT  7387.5 31537.5 7452.5 31402.5 ;
      RECT  7577.5 31537.5 7642.5 31402.5 ;
      RECT  7577.5 31537.5 7642.5 31402.5 ;
      RECT  7387.5 31537.5 7452.5 31402.5 ;
      RECT  7197.5 32377.5 7262.5 32242.5 ;
      RECT  7387.5 32377.5 7452.5 32242.5 ;
      RECT  7387.5 32377.5 7452.5 32242.5 ;
      RECT  7197.5 32377.5 7262.5 32242.5 ;
      RECT  7387.5 32377.5 7452.5 32242.5 ;
      RECT  7577.5 32377.5 7642.5 32242.5 ;
      RECT  7577.5 32377.5 7642.5 32242.5 ;
      RECT  7387.5 32377.5 7452.5 32242.5 ;
      RECT  7747.5 31447.5 7812.5 31312.5 ;
      RECT  7747.5 32422.5 7812.5 32287.5 ;
      RECT  7582.5 32147.5 7447.5 32082.5 ;
      RECT  7325.0 31932.5 7190.0 31867.5 ;
      RECT  7387.5 31537.5 7452.5 31402.5 ;
      RECT  7577.5 32377.5 7642.5 32242.5 ;
      RECT  7677.5 31932.5 7542.5 31867.5 ;
      RECT  7190.0 31932.5 7325.0 31867.5 ;
      RECT  7447.5 32147.5 7582.5 32082.5 ;
      RECT  7542.5 31932.5 7677.5 31867.5 ;
      RECT  7130.0 31227.5 8050.0 31162.5 ;
      RECT  7130.0 32572.5 8050.0 32507.5 ;
      RECT  7197.5 32702.5 7262.5 32507.5 ;
      RECT  7197.5 33542.5 7262.5 33917.5 ;
      RECT  7577.5 33542.5 7642.5 33917.5 ;
      RECT  7747.5 33700.0 7812.5 33885.0 ;
      RECT  7747.5 32540.0 7812.5 32725.0 ;
      RECT  7197.5 33542.5 7262.5 33677.5 ;
      RECT  7387.5 33542.5 7452.5 33677.5 ;
      RECT  7387.5 33542.5 7452.5 33677.5 ;
      RECT  7197.5 33542.5 7262.5 33677.5 ;
      RECT  7387.5 33542.5 7452.5 33677.5 ;
      RECT  7577.5 33542.5 7642.5 33677.5 ;
      RECT  7577.5 33542.5 7642.5 33677.5 ;
      RECT  7387.5 33542.5 7452.5 33677.5 ;
      RECT  7197.5 32702.5 7262.5 32837.5 ;
      RECT  7387.5 32702.5 7452.5 32837.5 ;
      RECT  7387.5 32702.5 7452.5 32837.5 ;
      RECT  7197.5 32702.5 7262.5 32837.5 ;
      RECT  7387.5 32702.5 7452.5 32837.5 ;
      RECT  7577.5 32702.5 7642.5 32837.5 ;
      RECT  7577.5 32702.5 7642.5 32837.5 ;
      RECT  7387.5 32702.5 7452.5 32837.5 ;
      RECT  7747.5 33632.5 7812.5 33767.5 ;
      RECT  7747.5 32657.5 7812.5 32792.5 ;
      RECT  7582.5 32932.5 7447.5 32997.5 ;
      RECT  7325.0 33147.5 7190.0 33212.5 ;
      RECT  7387.5 33542.5 7452.5 33677.5 ;
      RECT  7577.5 32702.5 7642.5 32837.5 ;
      RECT  7677.5 33147.5 7542.5 33212.5 ;
      RECT  7190.0 33147.5 7325.0 33212.5 ;
      RECT  7447.5 32932.5 7582.5 32997.5 ;
      RECT  7542.5 33147.5 7677.5 33212.5 ;
      RECT  7130.0 33852.5 8050.0 33917.5 ;
      RECT  7130.0 32507.5 8050.0 32572.5 ;
      RECT  7197.5 35067.5 7262.5 35262.5 ;
      RECT  7197.5 34227.5 7262.5 33852.5 ;
      RECT  7577.5 34227.5 7642.5 33852.5 ;
      RECT  7747.5 34070.0 7812.5 33885.0 ;
      RECT  7747.5 35230.0 7812.5 35045.0 ;
      RECT  7197.5 34227.5 7262.5 34092.5 ;
      RECT  7387.5 34227.5 7452.5 34092.5 ;
      RECT  7387.5 34227.5 7452.5 34092.5 ;
      RECT  7197.5 34227.5 7262.5 34092.5 ;
      RECT  7387.5 34227.5 7452.5 34092.5 ;
      RECT  7577.5 34227.5 7642.5 34092.5 ;
      RECT  7577.5 34227.5 7642.5 34092.5 ;
      RECT  7387.5 34227.5 7452.5 34092.5 ;
      RECT  7197.5 35067.5 7262.5 34932.5 ;
      RECT  7387.5 35067.5 7452.5 34932.5 ;
      RECT  7387.5 35067.5 7452.5 34932.5 ;
      RECT  7197.5 35067.5 7262.5 34932.5 ;
      RECT  7387.5 35067.5 7452.5 34932.5 ;
      RECT  7577.5 35067.5 7642.5 34932.5 ;
      RECT  7577.5 35067.5 7642.5 34932.5 ;
      RECT  7387.5 35067.5 7452.5 34932.5 ;
      RECT  7747.5 34137.5 7812.5 34002.5 ;
      RECT  7747.5 35112.5 7812.5 34977.5 ;
      RECT  7582.5 34837.5 7447.5 34772.5 ;
      RECT  7325.0 34622.5 7190.0 34557.5 ;
      RECT  7387.5 34227.5 7452.5 34092.5 ;
      RECT  7577.5 35067.5 7642.5 34932.5 ;
      RECT  7677.5 34622.5 7542.5 34557.5 ;
      RECT  7190.0 34622.5 7325.0 34557.5 ;
      RECT  7447.5 34837.5 7582.5 34772.5 ;
      RECT  7542.5 34622.5 7677.5 34557.5 ;
      RECT  7130.0 33917.5 8050.0 33852.5 ;
      RECT  7130.0 35262.5 8050.0 35197.5 ;
      RECT  7197.5 35392.5 7262.5 35197.5 ;
      RECT  7197.5 36232.5 7262.5 36607.5 ;
      RECT  7577.5 36232.5 7642.5 36607.5 ;
      RECT  7747.5 36390.0 7812.5 36575.0 ;
      RECT  7747.5 35230.0 7812.5 35415.0 ;
      RECT  7197.5 36232.5 7262.5 36367.5 ;
      RECT  7387.5 36232.5 7452.5 36367.5 ;
      RECT  7387.5 36232.5 7452.5 36367.5 ;
      RECT  7197.5 36232.5 7262.5 36367.5 ;
      RECT  7387.5 36232.5 7452.5 36367.5 ;
      RECT  7577.5 36232.5 7642.5 36367.5 ;
      RECT  7577.5 36232.5 7642.5 36367.5 ;
      RECT  7387.5 36232.5 7452.5 36367.5 ;
      RECT  7197.5 35392.5 7262.5 35527.5 ;
      RECT  7387.5 35392.5 7452.5 35527.5 ;
      RECT  7387.5 35392.5 7452.5 35527.5 ;
      RECT  7197.5 35392.5 7262.5 35527.5 ;
      RECT  7387.5 35392.5 7452.5 35527.5 ;
      RECT  7577.5 35392.5 7642.5 35527.5 ;
      RECT  7577.5 35392.5 7642.5 35527.5 ;
      RECT  7387.5 35392.5 7452.5 35527.5 ;
      RECT  7747.5 36322.5 7812.5 36457.5 ;
      RECT  7747.5 35347.5 7812.5 35482.5 ;
      RECT  7582.5 35622.5 7447.5 35687.5 ;
      RECT  7325.0 35837.5 7190.0 35902.5 ;
      RECT  7387.5 36232.5 7452.5 36367.5 ;
      RECT  7577.5 35392.5 7642.5 35527.5 ;
      RECT  7677.5 35837.5 7542.5 35902.5 ;
      RECT  7190.0 35837.5 7325.0 35902.5 ;
      RECT  7447.5 35622.5 7582.5 35687.5 ;
      RECT  7542.5 35837.5 7677.5 35902.5 ;
      RECT  7130.0 36542.5 8050.0 36607.5 ;
      RECT  7130.0 35197.5 8050.0 35262.5 ;
      RECT  7197.5 37757.5 7262.5 37952.5 ;
      RECT  7197.5 36917.5 7262.5 36542.5 ;
      RECT  7577.5 36917.5 7642.5 36542.5 ;
      RECT  7747.5 36760.0 7812.5 36575.0 ;
      RECT  7747.5 37920.0 7812.5 37735.0 ;
      RECT  7197.5 36917.5 7262.5 36782.5 ;
      RECT  7387.5 36917.5 7452.5 36782.5 ;
      RECT  7387.5 36917.5 7452.5 36782.5 ;
      RECT  7197.5 36917.5 7262.5 36782.5 ;
      RECT  7387.5 36917.5 7452.5 36782.5 ;
      RECT  7577.5 36917.5 7642.5 36782.5 ;
      RECT  7577.5 36917.5 7642.5 36782.5 ;
      RECT  7387.5 36917.5 7452.5 36782.5 ;
      RECT  7197.5 37757.5 7262.5 37622.5 ;
      RECT  7387.5 37757.5 7452.5 37622.5 ;
      RECT  7387.5 37757.5 7452.5 37622.5 ;
      RECT  7197.5 37757.5 7262.5 37622.5 ;
      RECT  7387.5 37757.5 7452.5 37622.5 ;
      RECT  7577.5 37757.5 7642.5 37622.5 ;
      RECT  7577.5 37757.5 7642.5 37622.5 ;
      RECT  7387.5 37757.5 7452.5 37622.5 ;
      RECT  7747.5 36827.5 7812.5 36692.5 ;
      RECT  7747.5 37802.5 7812.5 37667.5 ;
      RECT  7582.5 37527.5 7447.5 37462.5 ;
      RECT  7325.0 37312.5 7190.0 37247.5 ;
      RECT  7387.5 36917.5 7452.5 36782.5 ;
      RECT  7577.5 37757.5 7642.5 37622.5 ;
      RECT  7677.5 37312.5 7542.5 37247.5 ;
      RECT  7190.0 37312.5 7325.0 37247.5 ;
      RECT  7447.5 37527.5 7582.5 37462.5 ;
      RECT  7542.5 37312.5 7677.5 37247.5 ;
      RECT  7130.0 36607.5 8050.0 36542.5 ;
      RECT  7130.0 37952.5 8050.0 37887.5 ;
      RECT  7197.5 38082.5 7262.5 37887.5 ;
      RECT  7197.5 38922.5 7262.5 39297.5 ;
      RECT  7577.5 38922.5 7642.5 39297.5 ;
      RECT  7747.5 39080.0 7812.5 39265.0 ;
      RECT  7747.5 37920.0 7812.5 38105.0 ;
      RECT  7197.5 38922.5 7262.5 39057.5 ;
      RECT  7387.5 38922.5 7452.5 39057.5 ;
      RECT  7387.5 38922.5 7452.5 39057.5 ;
      RECT  7197.5 38922.5 7262.5 39057.5 ;
      RECT  7387.5 38922.5 7452.5 39057.5 ;
      RECT  7577.5 38922.5 7642.5 39057.5 ;
      RECT  7577.5 38922.5 7642.5 39057.5 ;
      RECT  7387.5 38922.5 7452.5 39057.5 ;
      RECT  7197.5 38082.5 7262.5 38217.5 ;
      RECT  7387.5 38082.5 7452.5 38217.5 ;
      RECT  7387.5 38082.5 7452.5 38217.5 ;
      RECT  7197.5 38082.5 7262.5 38217.5 ;
      RECT  7387.5 38082.5 7452.5 38217.5 ;
      RECT  7577.5 38082.5 7642.5 38217.5 ;
      RECT  7577.5 38082.5 7642.5 38217.5 ;
      RECT  7387.5 38082.5 7452.5 38217.5 ;
      RECT  7747.5 39012.5 7812.5 39147.5 ;
      RECT  7747.5 38037.5 7812.5 38172.5 ;
      RECT  7582.5 38312.5 7447.5 38377.5 ;
      RECT  7325.0 38527.5 7190.0 38592.5 ;
      RECT  7387.5 38922.5 7452.5 39057.5 ;
      RECT  7577.5 38082.5 7642.5 38217.5 ;
      RECT  7677.5 38527.5 7542.5 38592.5 ;
      RECT  7190.0 38527.5 7325.0 38592.5 ;
      RECT  7447.5 38312.5 7582.5 38377.5 ;
      RECT  7542.5 38527.5 7677.5 38592.5 ;
      RECT  7130.0 39232.5 8050.0 39297.5 ;
      RECT  7130.0 37887.5 8050.0 37952.5 ;
      RECT  7197.5 40447.5 7262.5 40642.5 ;
      RECT  7197.5 39607.5 7262.5 39232.5 ;
      RECT  7577.5 39607.5 7642.5 39232.5 ;
      RECT  7747.5 39450.0 7812.5 39265.0 ;
      RECT  7747.5 40610.0 7812.5 40425.0 ;
      RECT  7197.5 39607.5 7262.5 39472.5 ;
      RECT  7387.5 39607.5 7452.5 39472.5 ;
      RECT  7387.5 39607.5 7452.5 39472.5 ;
      RECT  7197.5 39607.5 7262.5 39472.5 ;
      RECT  7387.5 39607.5 7452.5 39472.5 ;
      RECT  7577.5 39607.5 7642.5 39472.5 ;
      RECT  7577.5 39607.5 7642.5 39472.5 ;
      RECT  7387.5 39607.5 7452.5 39472.5 ;
      RECT  7197.5 40447.5 7262.5 40312.5 ;
      RECT  7387.5 40447.5 7452.5 40312.5 ;
      RECT  7387.5 40447.5 7452.5 40312.5 ;
      RECT  7197.5 40447.5 7262.5 40312.5 ;
      RECT  7387.5 40447.5 7452.5 40312.5 ;
      RECT  7577.5 40447.5 7642.5 40312.5 ;
      RECT  7577.5 40447.5 7642.5 40312.5 ;
      RECT  7387.5 40447.5 7452.5 40312.5 ;
      RECT  7747.5 39517.5 7812.5 39382.5 ;
      RECT  7747.5 40492.5 7812.5 40357.5 ;
      RECT  7582.5 40217.5 7447.5 40152.5 ;
      RECT  7325.0 40002.5 7190.0 39937.5 ;
      RECT  7387.5 39607.5 7452.5 39472.5 ;
      RECT  7577.5 40447.5 7642.5 40312.5 ;
      RECT  7677.5 40002.5 7542.5 39937.5 ;
      RECT  7190.0 40002.5 7325.0 39937.5 ;
      RECT  7447.5 40217.5 7582.5 40152.5 ;
      RECT  7542.5 40002.5 7677.5 39937.5 ;
      RECT  7130.0 39297.5 8050.0 39232.5 ;
      RECT  7130.0 40642.5 8050.0 40577.5 ;
      RECT  8477.5 20250.0 8542.5 20435.0 ;
      RECT  8477.5 19090.0 8542.5 19275.0 ;
      RECT  8117.5 19207.5 8182.5 19057.5 ;
      RECT  8117.5 20092.5 8182.5 20467.5 ;
      RECT  8307.5 19207.5 8372.5 20092.5 ;
      RECT  8117.5 20092.5 8182.5 20227.5 ;
      RECT  8307.5 20092.5 8372.5 20227.5 ;
      RECT  8307.5 20092.5 8372.5 20227.5 ;
      RECT  8117.5 20092.5 8182.5 20227.5 ;
      RECT  8117.5 19207.5 8182.5 19342.5 ;
      RECT  8307.5 19207.5 8372.5 19342.5 ;
      RECT  8307.5 19207.5 8372.5 19342.5 ;
      RECT  8117.5 19207.5 8182.5 19342.5 ;
      RECT  8477.5 20182.5 8542.5 20317.5 ;
      RECT  8477.5 19207.5 8542.5 19342.5 ;
      RECT  8175.0 19650.0 8240.0 19785.0 ;
      RECT  8175.0 19650.0 8240.0 19785.0 ;
      RECT  8340.0 19685.0 8405.0 19750.0 ;
      RECT  8050.0 20402.5 8610.0 20467.5 ;
      RECT  8050.0 19057.5 8610.0 19122.5 ;
      RECT  8477.5 20620.0 8542.5 20435.0 ;
      RECT  8477.5 21780.0 8542.5 21595.0 ;
      RECT  8117.5 21662.5 8182.5 21812.5 ;
      RECT  8117.5 20777.5 8182.5 20402.5 ;
      RECT  8307.5 21662.5 8372.5 20777.5 ;
      RECT  8117.5 20777.5 8182.5 20642.5 ;
      RECT  8307.5 20777.5 8372.5 20642.5 ;
      RECT  8307.5 20777.5 8372.5 20642.5 ;
      RECT  8117.5 20777.5 8182.5 20642.5 ;
      RECT  8117.5 21662.5 8182.5 21527.5 ;
      RECT  8307.5 21662.5 8372.5 21527.5 ;
      RECT  8307.5 21662.5 8372.5 21527.5 ;
      RECT  8117.5 21662.5 8182.5 21527.5 ;
      RECT  8477.5 20687.5 8542.5 20552.5 ;
      RECT  8477.5 21662.5 8542.5 21527.5 ;
      RECT  8175.0 21220.0 8240.0 21085.0 ;
      RECT  8175.0 21220.0 8240.0 21085.0 ;
      RECT  8340.0 21185.0 8405.0 21120.0 ;
      RECT  8050.0 20467.5 8610.0 20402.5 ;
      RECT  8050.0 21812.5 8610.0 21747.5 ;
      RECT  8477.5 22940.0 8542.5 23125.0 ;
      RECT  8477.5 21780.0 8542.5 21965.0 ;
      RECT  8117.5 21897.5 8182.5 21747.5 ;
      RECT  8117.5 22782.5 8182.5 23157.5 ;
      RECT  8307.5 21897.5 8372.5 22782.5 ;
      RECT  8117.5 22782.5 8182.5 22917.5 ;
      RECT  8307.5 22782.5 8372.5 22917.5 ;
      RECT  8307.5 22782.5 8372.5 22917.5 ;
      RECT  8117.5 22782.5 8182.5 22917.5 ;
      RECT  8117.5 21897.5 8182.5 22032.5 ;
      RECT  8307.5 21897.5 8372.5 22032.5 ;
      RECT  8307.5 21897.5 8372.5 22032.5 ;
      RECT  8117.5 21897.5 8182.5 22032.5 ;
      RECT  8477.5 22872.5 8542.5 23007.5 ;
      RECT  8477.5 21897.5 8542.5 22032.5 ;
      RECT  8175.0 22340.0 8240.0 22475.0 ;
      RECT  8175.0 22340.0 8240.0 22475.0 ;
      RECT  8340.0 22375.0 8405.0 22440.0 ;
      RECT  8050.0 23092.5 8610.0 23157.5 ;
      RECT  8050.0 21747.5 8610.0 21812.5 ;
      RECT  8477.5 23310.0 8542.5 23125.0 ;
      RECT  8477.5 24470.0 8542.5 24285.0 ;
      RECT  8117.5 24352.5 8182.5 24502.5 ;
      RECT  8117.5 23467.5 8182.5 23092.5 ;
      RECT  8307.5 24352.5 8372.5 23467.5 ;
      RECT  8117.5 23467.5 8182.5 23332.5 ;
      RECT  8307.5 23467.5 8372.5 23332.5 ;
      RECT  8307.5 23467.5 8372.5 23332.5 ;
      RECT  8117.5 23467.5 8182.5 23332.5 ;
      RECT  8117.5 24352.5 8182.5 24217.5 ;
      RECT  8307.5 24352.5 8372.5 24217.5 ;
      RECT  8307.5 24352.5 8372.5 24217.5 ;
      RECT  8117.5 24352.5 8182.5 24217.5 ;
      RECT  8477.5 23377.5 8542.5 23242.5 ;
      RECT  8477.5 24352.5 8542.5 24217.5 ;
      RECT  8175.0 23910.0 8240.0 23775.0 ;
      RECT  8175.0 23910.0 8240.0 23775.0 ;
      RECT  8340.0 23875.0 8405.0 23810.0 ;
      RECT  8050.0 23157.5 8610.0 23092.5 ;
      RECT  8050.0 24502.5 8610.0 24437.5 ;
      RECT  8477.5 25630.0 8542.5 25815.0 ;
      RECT  8477.5 24470.0 8542.5 24655.0 ;
      RECT  8117.5 24587.5 8182.5 24437.5 ;
      RECT  8117.5 25472.5 8182.5 25847.5 ;
      RECT  8307.5 24587.5 8372.5 25472.5 ;
      RECT  8117.5 25472.5 8182.5 25607.5 ;
      RECT  8307.5 25472.5 8372.5 25607.5 ;
      RECT  8307.5 25472.5 8372.5 25607.5 ;
      RECT  8117.5 25472.5 8182.5 25607.5 ;
      RECT  8117.5 24587.5 8182.5 24722.5 ;
      RECT  8307.5 24587.5 8372.5 24722.5 ;
      RECT  8307.5 24587.5 8372.5 24722.5 ;
      RECT  8117.5 24587.5 8182.5 24722.5 ;
      RECT  8477.5 25562.5 8542.5 25697.5 ;
      RECT  8477.5 24587.5 8542.5 24722.5 ;
      RECT  8175.0 25030.0 8240.0 25165.0 ;
      RECT  8175.0 25030.0 8240.0 25165.0 ;
      RECT  8340.0 25065.0 8405.0 25130.0 ;
      RECT  8050.0 25782.5 8610.0 25847.5 ;
      RECT  8050.0 24437.5 8610.0 24502.5 ;
      RECT  8477.5 26000.0 8542.5 25815.0 ;
      RECT  8477.5 27160.0 8542.5 26975.0 ;
      RECT  8117.5 27042.5 8182.5 27192.5 ;
      RECT  8117.5 26157.5 8182.5 25782.5 ;
      RECT  8307.5 27042.5 8372.5 26157.5 ;
      RECT  8117.5 26157.5 8182.5 26022.5 ;
      RECT  8307.5 26157.5 8372.5 26022.5 ;
      RECT  8307.5 26157.5 8372.5 26022.5 ;
      RECT  8117.5 26157.5 8182.5 26022.5 ;
      RECT  8117.5 27042.5 8182.5 26907.5 ;
      RECT  8307.5 27042.5 8372.5 26907.5 ;
      RECT  8307.5 27042.5 8372.5 26907.5 ;
      RECT  8117.5 27042.5 8182.5 26907.5 ;
      RECT  8477.5 26067.5 8542.5 25932.5 ;
      RECT  8477.5 27042.5 8542.5 26907.5 ;
      RECT  8175.0 26600.0 8240.0 26465.0 ;
      RECT  8175.0 26600.0 8240.0 26465.0 ;
      RECT  8340.0 26565.0 8405.0 26500.0 ;
      RECT  8050.0 25847.5 8610.0 25782.5 ;
      RECT  8050.0 27192.5 8610.0 27127.5 ;
      RECT  8477.5 28320.0 8542.5 28505.0 ;
      RECT  8477.5 27160.0 8542.5 27345.0 ;
      RECT  8117.5 27277.5 8182.5 27127.5 ;
      RECT  8117.5 28162.5 8182.5 28537.5 ;
      RECT  8307.5 27277.5 8372.5 28162.5 ;
      RECT  8117.5 28162.5 8182.5 28297.5 ;
      RECT  8307.5 28162.5 8372.5 28297.5 ;
      RECT  8307.5 28162.5 8372.5 28297.5 ;
      RECT  8117.5 28162.5 8182.5 28297.5 ;
      RECT  8117.5 27277.5 8182.5 27412.5 ;
      RECT  8307.5 27277.5 8372.5 27412.5 ;
      RECT  8307.5 27277.5 8372.5 27412.5 ;
      RECT  8117.5 27277.5 8182.5 27412.5 ;
      RECT  8477.5 28252.5 8542.5 28387.5 ;
      RECT  8477.5 27277.5 8542.5 27412.5 ;
      RECT  8175.0 27720.0 8240.0 27855.0 ;
      RECT  8175.0 27720.0 8240.0 27855.0 ;
      RECT  8340.0 27755.0 8405.0 27820.0 ;
      RECT  8050.0 28472.5 8610.0 28537.5 ;
      RECT  8050.0 27127.5 8610.0 27192.5 ;
      RECT  8477.5 28690.0 8542.5 28505.0 ;
      RECT  8477.5 29850.0 8542.5 29665.0 ;
      RECT  8117.5 29732.5 8182.5 29882.5 ;
      RECT  8117.5 28847.5 8182.5 28472.5 ;
      RECT  8307.5 29732.5 8372.5 28847.5 ;
      RECT  8117.5 28847.5 8182.5 28712.5 ;
      RECT  8307.5 28847.5 8372.5 28712.5 ;
      RECT  8307.5 28847.5 8372.5 28712.5 ;
      RECT  8117.5 28847.5 8182.5 28712.5 ;
      RECT  8117.5 29732.5 8182.5 29597.5 ;
      RECT  8307.5 29732.5 8372.5 29597.5 ;
      RECT  8307.5 29732.5 8372.5 29597.5 ;
      RECT  8117.5 29732.5 8182.5 29597.5 ;
      RECT  8477.5 28757.5 8542.5 28622.5 ;
      RECT  8477.5 29732.5 8542.5 29597.5 ;
      RECT  8175.0 29290.0 8240.0 29155.0 ;
      RECT  8175.0 29290.0 8240.0 29155.0 ;
      RECT  8340.0 29255.0 8405.0 29190.0 ;
      RECT  8050.0 28537.5 8610.0 28472.5 ;
      RECT  8050.0 29882.5 8610.0 29817.5 ;
      RECT  8477.5 31010.0 8542.5 31195.0 ;
      RECT  8477.5 29850.0 8542.5 30035.0 ;
      RECT  8117.5 29967.5 8182.5 29817.5 ;
      RECT  8117.5 30852.5 8182.5 31227.5 ;
      RECT  8307.5 29967.5 8372.5 30852.5 ;
      RECT  8117.5 30852.5 8182.5 30987.5 ;
      RECT  8307.5 30852.5 8372.5 30987.5 ;
      RECT  8307.5 30852.5 8372.5 30987.5 ;
      RECT  8117.5 30852.5 8182.5 30987.5 ;
      RECT  8117.5 29967.5 8182.5 30102.5 ;
      RECT  8307.5 29967.5 8372.5 30102.5 ;
      RECT  8307.5 29967.5 8372.5 30102.5 ;
      RECT  8117.5 29967.5 8182.5 30102.5 ;
      RECT  8477.5 30942.5 8542.5 31077.5 ;
      RECT  8477.5 29967.5 8542.5 30102.5 ;
      RECT  8175.0 30410.0 8240.0 30545.0 ;
      RECT  8175.0 30410.0 8240.0 30545.0 ;
      RECT  8340.0 30445.0 8405.0 30510.0 ;
      RECT  8050.0 31162.5 8610.0 31227.5 ;
      RECT  8050.0 29817.5 8610.0 29882.5 ;
      RECT  8477.5 31380.0 8542.5 31195.0 ;
      RECT  8477.5 32540.0 8542.5 32355.0 ;
      RECT  8117.5 32422.5 8182.5 32572.5 ;
      RECT  8117.5 31537.5 8182.5 31162.5 ;
      RECT  8307.5 32422.5 8372.5 31537.5 ;
      RECT  8117.5 31537.5 8182.5 31402.5 ;
      RECT  8307.5 31537.5 8372.5 31402.5 ;
      RECT  8307.5 31537.5 8372.5 31402.5 ;
      RECT  8117.5 31537.5 8182.5 31402.5 ;
      RECT  8117.5 32422.5 8182.5 32287.5 ;
      RECT  8307.5 32422.5 8372.5 32287.5 ;
      RECT  8307.5 32422.5 8372.5 32287.5 ;
      RECT  8117.5 32422.5 8182.5 32287.5 ;
      RECT  8477.5 31447.5 8542.5 31312.5 ;
      RECT  8477.5 32422.5 8542.5 32287.5 ;
      RECT  8175.0 31980.0 8240.0 31845.0 ;
      RECT  8175.0 31980.0 8240.0 31845.0 ;
      RECT  8340.0 31945.0 8405.0 31880.0 ;
      RECT  8050.0 31227.5 8610.0 31162.5 ;
      RECT  8050.0 32572.5 8610.0 32507.5 ;
      RECT  8477.5 33700.0 8542.5 33885.0 ;
      RECT  8477.5 32540.0 8542.5 32725.0 ;
      RECT  8117.5 32657.5 8182.5 32507.5 ;
      RECT  8117.5 33542.5 8182.5 33917.5 ;
      RECT  8307.5 32657.5 8372.5 33542.5 ;
      RECT  8117.5 33542.5 8182.5 33677.5 ;
      RECT  8307.5 33542.5 8372.5 33677.5 ;
      RECT  8307.5 33542.5 8372.5 33677.5 ;
      RECT  8117.5 33542.5 8182.5 33677.5 ;
      RECT  8117.5 32657.5 8182.5 32792.5 ;
      RECT  8307.5 32657.5 8372.5 32792.5 ;
      RECT  8307.5 32657.5 8372.5 32792.5 ;
      RECT  8117.5 32657.5 8182.5 32792.5 ;
      RECT  8477.5 33632.5 8542.5 33767.5 ;
      RECT  8477.5 32657.5 8542.5 32792.5 ;
      RECT  8175.0 33100.0 8240.0 33235.0 ;
      RECT  8175.0 33100.0 8240.0 33235.0 ;
      RECT  8340.0 33135.0 8405.0 33200.0 ;
      RECT  8050.0 33852.5 8610.0 33917.5 ;
      RECT  8050.0 32507.5 8610.0 32572.5 ;
      RECT  8477.5 34070.0 8542.5 33885.0 ;
      RECT  8477.5 35230.0 8542.5 35045.0 ;
      RECT  8117.5 35112.5 8182.5 35262.5 ;
      RECT  8117.5 34227.5 8182.5 33852.5 ;
      RECT  8307.5 35112.5 8372.5 34227.5 ;
      RECT  8117.5 34227.5 8182.5 34092.5 ;
      RECT  8307.5 34227.5 8372.5 34092.5 ;
      RECT  8307.5 34227.5 8372.5 34092.5 ;
      RECT  8117.5 34227.5 8182.5 34092.5 ;
      RECT  8117.5 35112.5 8182.5 34977.5 ;
      RECT  8307.5 35112.5 8372.5 34977.5 ;
      RECT  8307.5 35112.5 8372.5 34977.5 ;
      RECT  8117.5 35112.5 8182.5 34977.5 ;
      RECT  8477.5 34137.5 8542.5 34002.5 ;
      RECT  8477.5 35112.5 8542.5 34977.5 ;
      RECT  8175.0 34670.0 8240.0 34535.0 ;
      RECT  8175.0 34670.0 8240.0 34535.0 ;
      RECT  8340.0 34635.0 8405.0 34570.0 ;
      RECT  8050.0 33917.5 8610.0 33852.5 ;
      RECT  8050.0 35262.5 8610.0 35197.5 ;
      RECT  8477.5 36390.0 8542.5 36575.0 ;
      RECT  8477.5 35230.0 8542.5 35415.0 ;
      RECT  8117.5 35347.5 8182.5 35197.5 ;
      RECT  8117.5 36232.5 8182.5 36607.5 ;
      RECT  8307.5 35347.5 8372.5 36232.5 ;
      RECT  8117.5 36232.5 8182.5 36367.5 ;
      RECT  8307.5 36232.5 8372.5 36367.5 ;
      RECT  8307.5 36232.5 8372.5 36367.5 ;
      RECT  8117.5 36232.5 8182.5 36367.5 ;
      RECT  8117.5 35347.5 8182.5 35482.5 ;
      RECT  8307.5 35347.5 8372.5 35482.5 ;
      RECT  8307.5 35347.5 8372.5 35482.5 ;
      RECT  8117.5 35347.5 8182.5 35482.5 ;
      RECT  8477.5 36322.5 8542.5 36457.5 ;
      RECT  8477.5 35347.5 8542.5 35482.5 ;
      RECT  8175.0 35790.0 8240.0 35925.0 ;
      RECT  8175.0 35790.0 8240.0 35925.0 ;
      RECT  8340.0 35825.0 8405.0 35890.0 ;
      RECT  8050.0 36542.5 8610.0 36607.5 ;
      RECT  8050.0 35197.5 8610.0 35262.5 ;
      RECT  8477.5 36760.0 8542.5 36575.0 ;
      RECT  8477.5 37920.0 8542.5 37735.0 ;
      RECT  8117.5 37802.5 8182.5 37952.5 ;
      RECT  8117.5 36917.5 8182.5 36542.5 ;
      RECT  8307.5 37802.5 8372.5 36917.5 ;
      RECT  8117.5 36917.5 8182.5 36782.5 ;
      RECT  8307.5 36917.5 8372.5 36782.5 ;
      RECT  8307.5 36917.5 8372.5 36782.5 ;
      RECT  8117.5 36917.5 8182.5 36782.5 ;
      RECT  8117.5 37802.5 8182.5 37667.5 ;
      RECT  8307.5 37802.5 8372.5 37667.5 ;
      RECT  8307.5 37802.5 8372.5 37667.5 ;
      RECT  8117.5 37802.5 8182.5 37667.5 ;
      RECT  8477.5 36827.5 8542.5 36692.5 ;
      RECT  8477.5 37802.5 8542.5 37667.5 ;
      RECT  8175.0 37360.0 8240.0 37225.0 ;
      RECT  8175.0 37360.0 8240.0 37225.0 ;
      RECT  8340.0 37325.0 8405.0 37260.0 ;
      RECT  8050.0 36607.5 8610.0 36542.5 ;
      RECT  8050.0 37952.5 8610.0 37887.5 ;
      RECT  8477.5 39080.0 8542.5 39265.0 ;
      RECT  8477.5 37920.0 8542.5 38105.0 ;
      RECT  8117.5 38037.5 8182.5 37887.5 ;
      RECT  8117.5 38922.5 8182.5 39297.5 ;
      RECT  8307.5 38037.5 8372.5 38922.5 ;
      RECT  8117.5 38922.5 8182.5 39057.5 ;
      RECT  8307.5 38922.5 8372.5 39057.5 ;
      RECT  8307.5 38922.5 8372.5 39057.5 ;
      RECT  8117.5 38922.5 8182.5 39057.5 ;
      RECT  8117.5 38037.5 8182.5 38172.5 ;
      RECT  8307.5 38037.5 8372.5 38172.5 ;
      RECT  8307.5 38037.5 8372.5 38172.5 ;
      RECT  8117.5 38037.5 8182.5 38172.5 ;
      RECT  8477.5 39012.5 8542.5 39147.5 ;
      RECT  8477.5 38037.5 8542.5 38172.5 ;
      RECT  8175.0 38480.0 8240.0 38615.0 ;
      RECT  8175.0 38480.0 8240.0 38615.0 ;
      RECT  8340.0 38515.0 8405.0 38580.0 ;
      RECT  8050.0 39232.5 8610.0 39297.5 ;
      RECT  8050.0 37887.5 8610.0 37952.5 ;
      RECT  8477.5 39450.0 8542.5 39265.0 ;
      RECT  8477.5 40610.0 8542.5 40425.0 ;
      RECT  8117.5 40492.5 8182.5 40642.5 ;
      RECT  8117.5 39607.5 8182.5 39232.5 ;
      RECT  8307.5 40492.5 8372.5 39607.5 ;
      RECT  8117.5 39607.5 8182.5 39472.5 ;
      RECT  8307.5 39607.5 8372.5 39472.5 ;
      RECT  8307.5 39607.5 8372.5 39472.5 ;
      RECT  8117.5 39607.5 8182.5 39472.5 ;
      RECT  8117.5 40492.5 8182.5 40357.5 ;
      RECT  8307.5 40492.5 8372.5 40357.5 ;
      RECT  8307.5 40492.5 8372.5 40357.5 ;
      RECT  8117.5 40492.5 8182.5 40357.5 ;
      RECT  8477.5 39517.5 8542.5 39382.5 ;
      RECT  8477.5 40492.5 8542.5 40357.5 ;
      RECT  8175.0 40050.0 8240.0 39915.0 ;
      RECT  8175.0 40050.0 8240.0 39915.0 ;
      RECT  8340.0 40015.0 8405.0 39950.0 ;
      RECT  8050.0 39297.5 8610.0 39232.5 ;
      RECT  8050.0 40642.5 8610.0 40577.5 ;
      RECT  5832.5 8925.0 5697.5 8990.0 ;
      RECT  6007.5 10360.0 5872.5 10425.0 ;
      RECT  6182.5 11615.0 6047.5 11680.0 ;
      RECT  6357.5 13050.0 6222.5 13115.0 ;
      RECT  6532.5 14305.0 6397.5 14370.0 ;
      RECT  6707.5 15740.0 6572.5 15805.0 ;
      RECT  6882.5 16995.0 6747.5 17060.0 ;
      RECT  7057.5 18430.0 6922.5 18495.0 ;
      RECT  5832.5 19697.5 5697.5 19762.5 ;
      RECT  6532.5 19482.5 6397.5 19547.5 ;
      RECT  5832.5 21107.5 5697.5 21172.5 ;
      RECT  6707.5 21322.5 6572.5 21387.5 ;
      RECT  5832.5 22387.5 5697.5 22452.5 ;
      RECT  6882.5 22172.5 6747.5 22237.5 ;
      RECT  5832.5 23797.5 5697.5 23862.5 ;
      RECT  7057.5 24012.5 6922.5 24077.5 ;
      RECT  6007.5 25077.5 5872.5 25142.5 ;
      RECT  6532.5 24862.5 6397.5 24927.5 ;
      RECT  6007.5 26487.5 5872.5 26552.5 ;
      RECT  6707.5 26702.5 6572.5 26767.5 ;
      RECT  6007.5 27767.5 5872.5 27832.5 ;
      RECT  6882.5 27552.5 6747.5 27617.5 ;
      RECT  6007.5 29177.5 5872.5 29242.5 ;
      RECT  7057.5 29392.5 6922.5 29457.5 ;
      RECT  6182.5 30457.5 6047.5 30522.5 ;
      RECT  6532.5 30242.5 6397.5 30307.5 ;
      RECT  6182.5 31867.5 6047.5 31932.5 ;
      RECT  6707.5 32082.5 6572.5 32147.5 ;
      RECT  6182.5 33147.5 6047.5 33212.5 ;
      RECT  6882.5 32932.5 6747.5 32997.5 ;
      RECT  6182.5 34557.5 6047.5 34622.5 ;
      RECT  7057.5 34772.5 6922.5 34837.5 ;
      RECT  6357.5 35837.5 6222.5 35902.5 ;
      RECT  6532.5 35622.5 6397.5 35687.5 ;
      RECT  6357.5 37247.5 6222.5 37312.5 ;
      RECT  6707.5 37462.5 6572.5 37527.5 ;
      RECT  6357.5 38527.5 6222.5 38592.5 ;
      RECT  6882.5 38312.5 6747.5 38377.5 ;
      RECT  6357.5 39937.5 6222.5 40002.5 ;
      RECT  7057.5 40152.5 6922.5 40217.5 ;
      RECT  8340.0 19685.0 8405.0 19750.0 ;
      RECT  8340.0 21120.0 8405.0 21185.0 ;
      RECT  8340.0 22375.0 8405.0 22440.0 ;
      RECT  8340.0 23810.0 8405.0 23875.0 ;
      RECT  8340.0 25065.0 8405.0 25130.0 ;
      RECT  8340.0 26500.0 8405.0 26565.0 ;
      RECT  8340.0 27755.0 8405.0 27820.0 ;
      RECT  8340.0 29190.0 8405.0 29255.0 ;
      RECT  8340.0 30445.0 8405.0 30510.0 ;
      RECT  8340.0 31880.0 8405.0 31945.0 ;
      RECT  8340.0 33135.0 8405.0 33200.0 ;
      RECT  8340.0 34570.0 8405.0 34635.0 ;
      RECT  8340.0 35825.0 8405.0 35890.0 ;
      RECT  8340.0 37260.0 8405.0 37325.0 ;
      RECT  8340.0 38515.0 8405.0 38580.0 ;
      RECT  8340.0 39950.0 8405.0 40015.0 ;
      RECT  5730.0 9642.5 11095.0 9707.5 ;
      RECT  5730.0 12332.5 11095.0 12397.5 ;
      RECT  5730.0 15022.5 11095.0 15087.5 ;
      RECT  5730.0 17712.5 11095.0 17777.5 ;
      RECT  5730.0 20402.5 11095.0 20467.5 ;
      RECT  5730.0 23092.5 11095.0 23157.5 ;
      RECT  5730.0 25782.5 11095.0 25847.5 ;
      RECT  5730.0 28472.5 11095.0 28537.5 ;
      RECT  5730.0 31162.5 11095.0 31227.5 ;
      RECT  5730.0 33852.5 11095.0 33917.5 ;
      RECT  5730.0 36542.5 11095.0 36607.5 ;
      RECT  5730.0 39232.5 11095.0 39297.5 ;
      RECT  5730.0 8297.5 11095.0 8362.5 ;
      RECT  5730.0 10987.5 11095.0 11052.5 ;
      RECT  5730.0 13677.5 11095.0 13742.5 ;
      RECT  5730.0 16367.5 11095.0 16432.5 ;
      RECT  5730.0 19057.5 11095.0 19122.5 ;
      RECT  5730.0 21747.5 11095.0 21812.5 ;
      RECT  5730.0 24437.5 11095.0 24502.5 ;
      RECT  5730.0 27127.5 11095.0 27192.5 ;
      RECT  5730.0 29817.5 11095.0 29882.5 ;
      RECT  5730.0 32507.5 11095.0 32572.5 ;
      RECT  5730.0 35197.5 11095.0 35262.5 ;
      RECT  5730.0 37887.5 11095.0 37952.5 ;
      RECT  5730.0 40577.5 11095.0 40642.5 ;
      RECT  8840.0 19685.0 9190.0 19750.0 ;
      RECT  9355.0 19697.5 9420.0 19762.5 ;
      RECT  9355.0 19685.0 9420.0 19750.0 ;
      RECT  9355.0 19730.0 9420.0 19750.0 ;
      RECT  9387.5 19697.5 9685.0 19762.5 ;
      RECT  9685.0 19697.5 9820.0 19762.5 ;
      RECT  10390.0 19697.5 10455.0 19762.5 ;
      RECT  10390.0 19685.0 10455.0 19750.0 ;
      RECT  10172.5 19697.5 10422.5 19762.5 ;
      RECT  10390.0 19717.5 10455.0 19730.0 ;
      RECT  10422.5 19685.0 10670.0 19750.0 ;
      RECT  8840.0 21120.0 9190.0 21185.0 ;
      RECT  9355.0 21107.5 9420.0 21172.5 ;
      RECT  9355.0 21120.0 9420.0 21185.0 ;
      RECT  9355.0 21140.0 9420.0 21185.0 ;
      RECT  9387.5 21107.5 9685.0 21172.5 ;
      RECT  9685.0 21107.5 9820.0 21172.5 ;
      RECT  10390.0 21107.5 10455.0 21172.5 ;
      RECT  10390.0 21120.0 10455.0 21185.0 ;
      RECT  10172.5 21107.5 10422.5 21172.5 ;
      RECT  10390.0 21140.0 10455.0 21152.5 ;
      RECT  10422.5 21120.0 10670.0 21185.0 ;
      RECT  8840.0 22375.0 9190.0 22440.0 ;
      RECT  9355.0 22387.5 9420.0 22452.5 ;
      RECT  9355.0 22375.0 9420.0 22440.0 ;
      RECT  9355.0 22420.0 9420.0 22440.0 ;
      RECT  9387.5 22387.5 9685.0 22452.5 ;
      RECT  9685.0 22387.5 9820.0 22452.5 ;
      RECT  10390.0 22387.5 10455.0 22452.5 ;
      RECT  10390.0 22375.0 10455.0 22440.0 ;
      RECT  10172.5 22387.5 10422.5 22452.5 ;
      RECT  10390.0 22407.5 10455.0 22420.0 ;
      RECT  10422.5 22375.0 10670.0 22440.0 ;
      RECT  8840.0 23810.0 9190.0 23875.0 ;
      RECT  9355.0 23797.5 9420.0 23862.5 ;
      RECT  9355.0 23810.0 9420.0 23875.0 ;
      RECT  9355.0 23830.0 9420.0 23875.0 ;
      RECT  9387.5 23797.5 9685.0 23862.5 ;
      RECT  9685.0 23797.5 9820.0 23862.5 ;
      RECT  10390.0 23797.5 10455.0 23862.5 ;
      RECT  10390.0 23810.0 10455.0 23875.0 ;
      RECT  10172.5 23797.5 10422.5 23862.5 ;
      RECT  10390.0 23830.0 10455.0 23842.5 ;
      RECT  10422.5 23810.0 10670.0 23875.0 ;
      RECT  8840.0 25065.0 9190.0 25130.0 ;
      RECT  9355.0 25077.5 9420.0 25142.5 ;
      RECT  9355.0 25065.0 9420.0 25130.0 ;
      RECT  9355.0 25110.0 9420.0 25130.0 ;
      RECT  9387.5 25077.5 9685.0 25142.5 ;
      RECT  9685.0 25077.5 9820.0 25142.5 ;
      RECT  10390.0 25077.5 10455.0 25142.5 ;
      RECT  10390.0 25065.0 10455.0 25130.0 ;
      RECT  10172.5 25077.5 10422.5 25142.5 ;
      RECT  10390.0 25097.5 10455.0 25110.0 ;
      RECT  10422.5 25065.0 10670.0 25130.0 ;
      RECT  8840.0 26500.0 9190.0 26565.0 ;
      RECT  9355.0 26487.5 9420.0 26552.5 ;
      RECT  9355.0 26500.0 9420.0 26565.0 ;
      RECT  9355.0 26520.0 9420.0 26565.0 ;
      RECT  9387.5 26487.5 9685.0 26552.5 ;
      RECT  9685.0 26487.5 9820.0 26552.5 ;
      RECT  10390.0 26487.5 10455.0 26552.5 ;
      RECT  10390.0 26500.0 10455.0 26565.0 ;
      RECT  10172.5 26487.5 10422.5 26552.5 ;
      RECT  10390.0 26520.0 10455.0 26532.5 ;
      RECT  10422.5 26500.0 10670.0 26565.0 ;
      RECT  8840.0 27755.0 9190.0 27820.0 ;
      RECT  9355.0 27767.5 9420.0 27832.5 ;
      RECT  9355.0 27755.0 9420.0 27820.0 ;
      RECT  9355.0 27800.0 9420.0 27820.0 ;
      RECT  9387.5 27767.5 9685.0 27832.5 ;
      RECT  9685.0 27767.5 9820.0 27832.5 ;
      RECT  10390.0 27767.5 10455.0 27832.5 ;
      RECT  10390.0 27755.0 10455.0 27820.0 ;
      RECT  10172.5 27767.5 10422.5 27832.5 ;
      RECT  10390.0 27787.5 10455.0 27800.0 ;
      RECT  10422.5 27755.0 10670.0 27820.0 ;
      RECT  8840.0 29190.0 9190.0 29255.0 ;
      RECT  9355.0 29177.5 9420.0 29242.5 ;
      RECT  9355.0 29190.0 9420.0 29255.0 ;
      RECT  9355.0 29210.0 9420.0 29255.0 ;
      RECT  9387.5 29177.5 9685.0 29242.5 ;
      RECT  9685.0 29177.5 9820.0 29242.5 ;
      RECT  10390.0 29177.5 10455.0 29242.5 ;
      RECT  10390.0 29190.0 10455.0 29255.0 ;
      RECT  10172.5 29177.5 10422.5 29242.5 ;
      RECT  10390.0 29210.0 10455.0 29222.5 ;
      RECT  10422.5 29190.0 10670.0 29255.0 ;
      RECT  8840.0 30445.0 9190.0 30510.0 ;
      RECT  9355.0 30457.5 9420.0 30522.5 ;
      RECT  9355.0 30445.0 9420.0 30510.0 ;
      RECT  9355.0 30490.0 9420.0 30510.0 ;
      RECT  9387.5 30457.5 9685.0 30522.5 ;
      RECT  9685.0 30457.5 9820.0 30522.5 ;
      RECT  10390.0 30457.5 10455.0 30522.5 ;
      RECT  10390.0 30445.0 10455.0 30510.0 ;
      RECT  10172.5 30457.5 10422.5 30522.5 ;
      RECT  10390.0 30477.5 10455.0 30490.0 ;
      RECT  10422.5 30445.0 10670.0 30510.0 ;
      RECT  8840.0 31880.0 9190.0 31945.0 ;
      RECT  9355.0 31867.5 9420.0 31932.5 ;
      RECT  9355.0 31880.0 9420.0 31945.0 ;
      RECT  9355.0 31900.0 9420.0 31945.0 ;
      RECT  9387.5 31867.5 9685.0 31932.5 ;
      RECT  9685.0 31867.5 9820.0 31932.5 ;
      RECT  10390.0 31867.5 10455.0 31932.5 ;
      RECT  10390.0 31880.0 10455.0 31945.0 ;
      RECT  10172.5 31867.5 10422.5 31932.5 ;
      RECT  10390.0 31900.0 10455.0 31912.5 ;
      RECT  10422.5 31880.0 10670.0 31945.0 ;
      RECT  8840.0 33135.0 9190.0 33200.0 ;
      RECT  9355.0 33147.5 9420.0 33212.5 ;
      RECT  9355.0 33135.0 9420.0 33200.0 ;
      RECT  9355.0 33180.0 9420.0 33200.0 ;
      RECT  9387.5 33147.5 9685.0 33212.5 ;
      RECT  9685.0 33147.5 9820.0 33212.5 ;
      RECT  10390.0 33147.5 10455.0 33212.5 ;
      RECT  10390.0 33135.0 10455.0 33200.0 ;
      RECT  10172.5 33147.5 10422.5 33212.5 ;
      RECT  10390.0 33167.5 10455.0 33180.0 ;
      RECT  10422.5 33135.0 10670.0 33200.0 ;
      RECT  8840.0 34570.0 9190.0 34635.0 ;
      RECT  9355.0 34557.5 9420.0 34622.5 ;
      RECT  9355.0 34570.0 9420.0 34635.0 ;
      RECT  9355.0 34590.0 9420.0 34635.0 ;
      RECT  9387.5 34557.5 9685.0 34622.5 ;
      RECT  9685.0 34557.5 9820.0 34622.5 ;
      RECT  10390.0 34557.5 10455.0 34622.5 ;
      RECT  10390.0 34570.0 10455.0 34635.0 ;
      RECT  10172.5 34557.5 10422.5 34622.5 ;
      RECT  10390.0 34590.0 10455.0 34602.5 ;
      RECT  10422.5 34570.0 10670.0 34635.0 ;
      RECT  8840.0 35825.0 9190.0 35890.0 ;
      RECT  9355.0 35837.5 9420.0 35902.5 ;
      RECT  9355.0 35825.0 9420.0 35890.0 ;
      RECT  9355.0 35870.0 9420.0 35890.0 ;
      RECT  9387.5 35837.5 9685.0 35902.5 ;
      RECT  9685.0 35837.5 9820.0 35902.5 ;
      RECT  10390.0 35837.5 10455.0 35902.5 ;
      RECT  10390.0 35825.0 10455.0 35890.0 ;
      RECT  10172.5 35837.5 10422.5 35902.5 ;
      RECT  10390.0 35857.5 10455.0 35870.0 ;
      RECT  10422.5 35825.0 10670.0 35890.0 ;
      RECT  8840.0 37260.0 9190.0 37325.0 ;
      RECT  9355.0 37247.5 9420.0 37312.5 ;
      RECT  9355.0 37260.0 9420.0 37325.0 ;
      RECT  9355.0 37280.0 9420.0 37325.0 ;
      RECT  9387.5 37247.5 9685.0 37312.5 ;
      RECT  9685.0 37247.5 9820.0 37312.5 ;
      RECT  10390.0 37247.5 10455.0 37312.5 ;
      RECT  10390.0 37260.0 10455.0 37325.0 ;
      RECT  10172.5 37247.5 10422.5 37312.5 ;
      RECT  10390.0 37280.0 10455.0 37292.5 ;
      RECT  10422.5 37260.0 10670.0 37325.0 ;
      RECT  8840.0 38515.0 9190.0 38580.0 ;
      RECT  9355.0 38527.5 9420.0 38592.5 ;
      RECT  9355.0 38515.0 9420.0 38580.0 ;
      RECT  9355.0 38560.0 9420.0 38580.0 ;
      RECT  9387.5 38527.5 9685.0 38592.5 ;
      RECT  9685.0 38527.5 9820.0 38592.5 ;
      RECT  10390.0 38527.5 10455.0 38592.5 ;
      RECT  10390.0 38515.0 10455.0 38580.0 ;
      RECT  10172.5 38527.5 10422.5 38592.5 ;
      RECT  10390.0 38547.5 10455.0 38560.0 ;
      RECT  10422.5 38515.0 10670.0 38580.0 ;
      RECT  8840.0 39950.0 9190.0 40015.0 ;
      RECT  9355.0 39937.5 9420.0 40002.5 ;
      RECT  9355.0 39950.0 9420.0 40015.0 ;
      RECT  9355.0 39970.0 9420.0 40015.0 ;
      RECT  9387.5 39937.5 9685.0 40002.5 ;
      RECT  9685.0 39937.5 9820.0 40002.5 ;
      RECT  10390.0 39937.5 10455.0 40002.5 ;
      RECT  10390.0 39950.0 10455.0 40015.0 ;
      RECT  10172.5 39937.5 10422.5 40002.5 ;
      RECT  10390.0 39970.0 10455.0 39982.5 ;
      RECT  10422.5 39950.0 10670.0 40015.0 ;
      RECT  9492.5 20250.0 9557.5 20435.0 ;
      RECT  9492.5 19090.0 9557.5 19275.0 ;
      RECT  9132.5 19207.5 9197.5 19057.5 ;
      RECT  9132.5 20092.5 9197.5 20467.5 ;
      RECT  9322.5 19207.5 9387.5 20092.5 ;
      RECT  9132.5 20092.5 9197.5 20227.5 ;
      RECT  9322.5 20092.5 9387.5 20227.5 ;
      RECT  9322.5 20092.5 9387.5 20227.5 ;
      RECT  9132.5 20092.5 9197.5 20227.5 ;
      RECT  9132.5 19207.5 9197.5 19342.5 ;
      RECT  9322.5 19207.5 9387.5 19342.5 ;
      RECT  9322.5 19207.5 9387.5 19342.5 ;
      RECT  9132.5 19207.5 9197.5 19342.5 ;
      RECT  9492.5 20182.5 9557.5 20317.5 ;
      RECT  9492.5 19207.5 9557.5 19342.5 ;
      RECT  9190.0 19650.0 9255.0 19785.0 ;
      RECT  9190.0 19650.0 9255.0 19785.0 ;
      RECT  9355.0 19685.0 9420.0 19750.0 ;
      RECT  9065.0 20402.5 9625.0 20467.5 ;
      RECT  9065.0 19057.5 9625.0 19122.5 ;
      RECT  9692.5 19252.5 9757.5 19057.5 ;
      RECT  9692.5 20092.5 9757.5 20467.5 ;
      RECT  10072.5 20092.5 10137.5 20467.5 ;
      RECT  10242.5 20250.0 10307.5 20435.0 ;
      RECT  10242.5 19090.0 10307.5 19275.0 ;
      RECT  9692.5 20092.5 9757.5 20227.5 ;
      RECT  9882.5 20092.5 9947.5 20227.5 ;
      RECT  9882.5 20092.5 9947.5 20227.5 ;
      RECT  9692.5 20092.5 9757.5 20227.5 ;
      RECT  9882.5 20092.5 9947.5 20227.5 ;
      RECT  10072.5 20092.5 10137.5 20227.5 ;
      RECT  10072.5 20092.5 10137.5 20227.5 ;
      RECT  9882.5 20092.5 9947.5 20227.5 ;
      RECT  9692.5 19252.5 9757.5 19387.5 ;
      RECT  9882.5 19252.5 9947.5 19387.5 ;
      RECT  9882.5 19252.5 9947.5 19387.5 ;
      RECT  9692.5 19252.5 9757.5 19387.5 ;
      RECT  9882.5 19252.5 9947.5 19387.5 ;
      RECT  10072.5 19252.5 10137.5 19387.5 ;
      RECT  10072.5 19252.5 10137.5 19387.5 ;
      RECT  9882.5 19252.5 9947.5 19387.5 ;
      RECT  10242.5 20182.5 10307.5 20317.5 ;
      RECT  10242.5 19207.5 10307.5 19342.5 ;
      RECT  10077.5 19482.5 9942.5 19547.5 ;
      RECT  9820.0 19697.5 9685.0 19762.5 ;
      RECT  9882.5 20092.5 9947.5 20227.5 ;
      RECT  10072.5 19252.5 10137.5 19387.5 ;
      RECT  10172.5 19697.5 10037.5 19762.5 ;
      RECT  9685.0 19697.5 9820.0 19762.5 ;
      RECT  9942.5 19482.5 10077.5 19547.5 ;
      RECT  10037.5 19697.5 10172.5 19762.5 ;
      RECT  9625.0 20402.5 10545.0 20467.5 ;
      RECT  9625.0 19057.5 10545.0 19122.5 ;
      RECT  10972.5 20250.0 11037.5 20435.0 ;
      RECT  10972.5 19090.0 11037.5 19275.0 ;
      RECT  10612.5 19207.5 10677.5 19057.5 ;
      RECT  10612.5 20092.5 10677.5 20467.5 ;
      RECT  10802.5 19207.5 10867.5 20092.5 ;
      RECT  10612.5 20092.5 10677.5 20227.5 ;
      RECT  10802.5 20092.5 10867.5 20227.5 ;
      RECT  10802.5 20092.5 10867.5 20227.5 ;
      RECT  10612.5 20092.5 10677.5 20227.5 ;
      RECT  10612.5 19207.5 10677.5 19342.5 ;
      RECT  10802.5 19207.5 10867.5 19342.5 ;
      RECT  10802.5 19207.5 10867.5 19342.5 ;
      RECT  10612.5 19207.5 10677.5 19342.5 ;
      RECT  10972.5 20182.5 11037.5 20317.5 ;
      RECT  10972.5 19207.5 11037.5 19342.5 ;
      RECT  10670.0 19650.0 10735.0 19785.0 ;
      RECT  10670.0 19650.0 10735.0 19785.0 ;
      RECT  10835.0 19685.0 10900.0 19750.0 ;
      RECT  10545.0 20402.5 11105.0 20467.5 ;
      RECT  10545.0 19057.5 11105.0 19122.5 ;
      RECT  8807.5 19650.0 8872.5 19785.0 ;
      RECT  8947.5 19377.5 9012.5 19512.5 ;
      RECT  9942.5 19482.5 9807.5 19547.5 ;
      RECT  9492.5 20620.0 9557.5 20435.0 ;
      RECT  9492.5 21780.0 9557.5 21595.0 ;
      RECT  9132.5 21662.5 9197.5 21812.5 ;
      RECT  9132.5 20777.5 9197.5 20402.5 ;
      RECT  9322.5 21662.5 9387.5 20777.5 ;
      RECT  9132.5 20777.5 9197.5 20642.5 ;
      RECT  9322.5 20777.5 9387.5 20642.5 ;
      RECT  9322.5 20777.5 9387.5 20642.5 ;
      RECT  9132.5 20777.5 9197.5 20642.5 ;
      RECT  9132.5 21662.5 9197.5 21527.5 ;
      RECT  9322.5 21662.5 9387.5 21527.5 ;
      RECT  9322.5 21662.5 9387.5 21527.5 ;
      RECT  9132.5 21662.5 9197.5 21527.5 ;
      RECT  9492.5 20687.5 9557.5 20552.5 ;
      RECT  9492.5 21662.5 9557.5 21527.5 ;
      RECT  9190.0 21220.0 9255.0 21085.0 ;
      RECT  9190.0 21220.0 9255.0 21085.0 ;
      RECT  9355.0 21185.0 9420.0 21120.0 ;
      RECT  9065.0 20467.5 9625.0 20402.5 ;
      RECT  9065.0 21812.5 9625.0 21747.5 ;
      RECT  9692.5 21617.5 9757.5 21812.5 ;
      RECT  9692.5 20777.5 9757.5 20402.5 ;
      RECT  10072.5 20777.5 10137.5 20402.5 ;
      RECT  10242.5 20620.0 10307.5 20435.0 ;
      RECT  10242.5 21780.0 10307.5 21595.0 ;
      RECT  9692.5 20777.5 9757.5 20642.5 ;
      RECT  9882.5 20777.5 9947.5 20642.5 ;
      RECT  9882.5 20777.5 9947.5 20642.5 ;
      RECT  9692.5 20777.5 9757.5 20642.5 ;
      RECT  9882.5 20777.5 9947.5 20642.5 ;
      RECT  10072.5 20777.5 10137.5 20642.5 ;
      RECT  10072.5 20777.5 10137.5 20642.5 ;
      RECT  9882.5 20777.5 9947.5 20642.5 ;
      RECT  9692.5 21617.5 9757.5 21482.5 ;
      RECT  9882.5 21617.5 9947.5 21482.5 ;
      RECT  9882.5 21617.5 9947.5 21482.5 ;
      RECT  9692.5 21617.5 9757.5 21482.5 ;
      RECT  9882.5 21617.5 9947.5 21482.5 ;
      RECT  10072.5 21617.5 10137.5 21482.5 ;
      RECT  10072.5 21617.5 10137.5 21482.5 ;
      RECT  9882.5 21617.5 9947.5 21482.5 ;
      RECT  10242.5 20687.5 10307.5 20552.5 ;
      RECT  10242.5 21662.5 10307.5 21527.5 ;
      RECT  10077.5 21387.5 9942.5 21322.5 ;
      RECT  9820.0 21172.5 9685.0 21107.5 ;
      RECT  9882.5 20777.5 9947.5 20642.5 ;
      RECT  10072.5 21617.5 10137.5 21482.5 ;
      RECT  10172.5 21172.5 10037.5 21107.5 ;
      RECT  9685.0 21172.5 9820.0 21107.5 ;
      RECT  9942.5 21387.5 10077.5 21322.5 ;
      RECT  10037.5 21172.5 10172.5 21107.5 ;
      RECT  9625.0 20467.5 10545.0 20402.5 ;
      RECT  9625.0 21812.5 10545.0 21747.5 ;
      RECT  10972.5 20620.0 11037.5 20435.0 ;
      RECT  10972.5 21780.0 11037.5 21595.0 ;
      RECT  10612.5 21662.5 10677.5 21812.5 ;
      RECT  10612.5 20777.5 10677.5 20402.5 ;
      RECT  10802.5 21662.5 10867.5 20777.5 ;
      RECT  10612.5 20777.5 10677.5 20642.5 ;
      RECT  10802.5 20777.5 10867.5 20642.5 ;
      RECT  10802.5 20777.5 10867.5 20642.5 ;
      RECT  10612.5 20777.5 10677.5 20642.5 ;
      RECT  10612.5 21662.5 10677.5 21527.5 ;
      RECT  10802.5 21662.5 10867.5 21527.5 ;
      RECT  10802.5 21662.5 10867.5 21527.5 ;
      RECT  10612.5 21662.5 10677.5 21527.5 ;
      RECT  10972.5 20687.5 11037.5 20552.5 ;
      RECT  10972.5 21662.5 11037.5 21527.5 ;
      RECT  10670.0 21220.0 10735.0 21085.0 ;
      RECT  10670.0 21220.0 10735.0 21085.0 ;
      RECT  10835.0 21185.0 10900.0 21120.0 ;
      RECT  10545.0 20467.5 11105.0 20402.5 ;
      RECT  10545.0 21812.5 11105.0 21747.5 ;
      RECT  8807.5 21085.0 8872.5 21220.0 ;
      RECT  8947.5 21357.5 9012.5 21492.5 ;
      RECT  9942.5 21322.5 9807.5 21387.5 ;
      RECT  9492.5 22940.0 9557.5 23125.0 ;
      RECT  9492.5 21780.0 9557.5 21965.0 ;
      RECT  9132.5 21897.5 9197.5 21747.5 ;
      RECT  9132.5 22782.5 9197.5 23157.5 ;
      RECT  9322.5 21897.5 9387.5 22782.5 ;
      RECT  9132.5 22782.5 9197.5 22917.5 ;
      RECT  9322.5 22782.5 9387.5 22917.5 ;
      RECT  9322.5 22782.5 9387.5 22917.5 ;
      RECT  9132.5 22782.5 9197.5 22917.5 ;
      RECT  9132.5 21897.5 9197.5 22032.5 ;
      RECT  9322.5 21897.5 9387.5 22032.5 ;
      RECT  9322.5 21897.5 9387.5 22032.5 ;
      RECT  9132.5 21897.5 9197.5 22032.5 ;
      RECT  9492.5 22872.5 9557.5 23007.5 ;
      RECT  9492.5 21897.5 9557.5 22032.5 ;
      RECT  9190.0 22340.0 9255.0 22475.0 ;
      RECT  9190.0 22340.0 9255.0 22475.0 ;
      RECT  9355.0 22375.0 9420.0 22440.0 ;
      RECT  9065.0 23092.5 9625.0 23157.5 ;
      RECT  9065.0 21747.5 9625.0 21812.5 ;
      RECT  9692.5 21942.5 9757.5 21747.5 ;
      RECT  9692.5 22782.5 9757.5 23157.5 ;
      RECT  10072.5 22782.5 10137.5 23157.5 ;
      RECT  10242.5 22940.0 10307.5 23125.0 ;
      RECT  10242.5 21780.0 10307.5 21965.0 ;
      RECT  9692.5 22782.5 9757.5 22917.5 ;
      RECT  9882.5 22782.5 9947.5 22917.5 ;
      RECT  9882.5 22782.5 9947.5 22917.5 ;
      RECT  9692.5 22782.5 9757.5 22917.5 ;
      RECT  9882.5 22782.5 9947.5 22917.5 ;
      RECT  10072.5 22782.5 10137.5 22917.5 ;
      RECT  10072.5 22782.5 10137.5 22917.5 ;
      RECT  9882.5 22782.5 9947.5 22917.5 ;
      RECT  9692.5 21942.5 9757.5 22077.5 ;
      RECT  9882.5 21942.5 9947.5 22077.5 ;
      RECT  9882.5 21942.5 9947.5 22077.5 ;
      RECT  9692.5 21942.5 9757.5 22077.5 ;
      RECT  9882.5 21942.5 9947.5 22077.5 ;
      RECT  10072.5 21942.5 10137.5 22077.5 ;
      RECT  10072.5 21942.5 10137.5 22077.5 ;
      RECT  9882.5 21942.5 9947.5 22077.5 ;
      RECT  10242.5 22872.5 10307.5 23007.5 ;
      RECT  10242.5 21897.5 10307.5 22032.5 ;
      RECT  10077.5 22172.5 9942.5 22237.5 ;
      RECT  9820.0 22387.5 9685.0 22452.5 ;
      RECT  9882.5 22782.5 9947.5 22917.5 ;
      RECT  10072.5 21942.5 10137.5 22077.5 ;
      RECT  10172.5 22387.5 10037.5 22452.5 ;
      RECT  9685.0 22387.5 9820.0 22452.5 ;
      RECT  9942.5 22172.5 10077.5 22237.5 ;
      RECT  10037.5 22387.5 10172.5 22452.5 ;
      RECT  9625.0 23092.5 10545.0 23157.5 ;
      RECT  9625.0 21747.5 10545.0 21812.5 ;
      RECT  10972.5 22940.0 11037.5 23125.0 ;
      RECT  10972.5 21780.0 11037.5 21965.0 ;
      RECT  10612.5 21897.5 10677.5 21747.5 ;
      RECT  10612.5 22782.5 10677.5 23157.5 ;
      RECT  10802.5 21897.5 10867.5 22782.5 ;
      RECT  10612.5 22782.5 10677.5 22917.5 ;
      RECT  10802.5 22782.5 10867.5 22917.5 ;
      RECT  10802.5 22782.5 10867.5 22917.5 ;
      RECT  10612.5 22782.5 10677.5 22917.5 ;
      RECT  10612.5 21897.5 10677.5 22032.5 ;
      RECT  10802.5 21897.5 10867.5 22032.5 ;
      RECT  10802.5 21897.5 10867.5 22032.5 ;
      RECT  10612.5 21897.5 10677.5 22032.5 ;
      RECT  10972.5 22872.5 11037.5 23007.5 ;
      RECT  10972.5 21897.5 11037.5 22032.5 ;
      RECT  10670.0 22340.0 10735.0 22475.0 ;
      RECT  10670.0 22340.0 10735.0 22475.0 ;
      RECT  10835.0 22375.0 10900.0 22440.0 ;
      RECT  10545.0 23092.5 11105.0 23157.5 ;
      RECT  10545.0 21747.5 11105.0 21812.5 ;
      RECT  8807.5 22340.0 8872.5 22475.0 ;
      RECT  8947.5 22067.5 9012.5 22202.5 ;
      RECT  9942.5 22172.5 9807.5 22237.5 ;
      RECT  9492.5 23310.0 9557.5 23125.0 ;
      RECT  9492.5 24470.0 9557.5 24285.0 ;
      RECT  9132.5 24352.5 9197.5 24502.5 ;
      RECT  9132.5 23467.5 9197.5 23092.5 ;
      RECT  9322.5 24352.5 9387.5 23467.5 ;
      RECT  9132.5 23467.5 9197.5 23332.5 ;
      RECT  9322.5 23467.5 9387.5 23332.5 ;
      RECT  9322.5 23467.5 9387.5 23332.5 ;
      RECT  9132.5 23467.5 9197.5 23332.5 ;
      RECT  9132.5 24352.5 9197.5 24217.5 ;
      RECT  9322.5 24352.5 9387.5 24217.5 ;
      RECT  9322.5 24352.5 9387.5 24217.5 ;
      RECT  9132.5 24352.5 9197.5 24217.5 ;
      RECT  9492.5 23377.5 9557.5 23242.5 ;
      RECT  9492.5 24352.5 9557.5 24217.5 ;
      RECT  9190.0 23910.0 9255.0 23775.0 ;
      RECT  9190.0 23910.0 9255.0 23775.0 ;
      RECT  9355.0 23875.0 9420.0 23810.0 ;
      RECT  9065.0 23157.5 9625.0 23092.5 ;
      RECT  9065.0 24502.5 9625.0 24437.5 ;
      RECT  9692.5 24307.5 9757.5 24502.5 ;
      RECT  9692.5 23467.5 9757.5 23092.5 ;
      RECT  10072.5 23467.5 10137.5 23092.5 ;
      RECT  10242.5 23310.0 10307.5 23125.0 ;
      RECT  10242.5 24470.0 10307.5 24285.0 ;
      RECT  9692.5 23467.5 9757.5 23332.5 ;
      RECT  9882.5 23467.5 9947.5 23332.5 ;
      RECT  9882.5 23467.5 9947.5 23332.5 ;
      RECT  9692.5 23467.5 9757.5 23332.5 ;
      RECT  9882.5 23467.5 9947.5 23332.5 ;
      RECT  10072.5 23467.5 10137.5 23332.5 ;
      RECT  10072.5 23467.5 10137.5 23332.5 ;
      RECT  9882.5 23467.5 9947.5 23332.5 ;
      RECT  9692.5 24307.5 9757.5 24172.5 ;
      RECT  9882.5 24307.5 9947.5 24172.5 ;
      RECT  9882.5 24307.5 9947.5 24172.5 ;
      RECT  9692.5 24307.5 9757.5 24172.5 ;
      RECT  9882.5 24307.5 9947.5 24172.5 ;
      RECT  10072.5 24307.5 10137.5 24172.5 ;
      RECT  10072.5 24307.5 10137.5 24172.5 ;
      RECT  9882.5 24307.5 9947.5 24172.5 ;
      RECT  10242.5 23377.5 10307.5 23242.5 ;
      RECT  10242.5 24352.5 10307.5 24217.5 ;
      RECT  10077.5 24077.5 9942.5 24012.5 ;
      RECT  9820.0 23862.5 9685.0 23797.5 ;
      RECT  9882.5 23467.5 9947.5 23332.5 ;
      RECT  10072.5 24307.5 10137.5 24172.5 ;
      RECT  10172.5 23862.5 10037.5 23797.5 ;
      RECT  9685.0 23862.5 9820.0 23797.5 ;
      RECT  9942.5 24077.5 10077.5 24012.5 ;
      RECT  10037.5 23862.5 10172.5 23797.5 ;
      RECT  9625.0 23157.5 10545.0 23092.5 ;
      RECT  9625.0 24502.5 10545.0 24437.5 ;
      RECT  10972.5 23310.0 11037.5 23125.0 ;
      RECT  10972.5 24470.0 11037.5 24285.0 ;
      RECT  10612.5 24352.5 10677.5 24502.5 ;
      RECT  10612.5 23467.5 10677.5 23092.5 ;
      RECT  10802.5 24352.5 10867.5 23467.5 ;
      RECT  10612.5 23467.5 10677.5 23332.5 ;
      RECT  10802.5 23467.5 10867.5 23332.5 ;
      RECT  10802.5 23467.5 10867.5 23332.5 ;
      RECT  10612.5 23467.5 10677.5 23332.5 ;
      RECT  10612.5 24352.5 10677.5 24217.5 ;
      RECT  10802.5 24352.5 10867.5 24217.5 ;
      RECT  10802.5 24352.5 10867.5 24217.5 ;
      RECT  10612.5 24352.5 10677.5 24217.5 ;
      RECT  10972.5 23377.5 11037.5 23242.5 ;
      RECT  10972.5 24352.5 11037.5 24217.5 ;
      RECT  10670.0 23910.0 10735.0 23775.0 ;
      RECT  10670.0 23910.0 10735.0 23775.0 ;
      RECT  10835.0 23875.0 10900.0 23810.0 ;
      RECT  10545.0 23157.5 11105.0 23092.5 ;
      RECT  10545.0 24502.5 11105.0 24437.5 ;
      RECT  8807.5 23775.0 8872.5 23910.0 ;
      RECT  8947.5 24047.5 9012.5 24182.5 ;
      RECT  9942.5 24012.5 9807.5 24077.5 ;
      RECT  9492.5 25630.0 9557.5 25815.0 ;
      RECT  9492.5 24470.0 9557.5 24655.0 ;
      RECT  9132.5 24587.5 9197.5 24437.5 ;
      RECT  9132.5 25472.5 9197.5 25847.5 ;
      RECT  9322.5 24587.5 9387.5 25472.5 ;
      RECT  9132.5 25472.5 9197.5 25607.5 ;
      RECT  9322.5 25472.5 9387.5 25607.5 ;
      RECT  9322.5 25472.5 9387.5 25607.5 ;
      RECT  9132.5 25472.5 9197.5 25607.5 ;
      RECT  9132.5 24587.5 9197.5 24722.5 ;
      RECT  9322.5 24587.5 9387.5 24722.5 ;
      RECT  9322.5 24587.5 9387.5 24722.5 ;
      RECT  9132.5 24587.5 9197.5 24722.5 ;
      RECT  9492.5 25562.5 9557.5 25697.5 ;
      RECT  9492.5 24587.5 9557.5 24722.5 ;
      RECT  9190.0 25030.0 9255.0 25165.0 ;
      RECT  9190.0 25030.0 9255.0 25165.0 ;
      RECT  9355.0 25065.0 9420.0 25130.0 ;
      RECT  9065.0 25782.5 9625.0 25847.5 ;
      RECT  9065.0 24437.5 9625.0 24502.5 ;
      RECT  9692.5 24632.5 9757.5 24437.5 ;
      RECT  9692.5 25472.5 9757.5 25847.5 ;
      RECT  10072.5 25472.5 10137.5 25847.5 ;
      RECT  10242.5 25630.0 10307.5 25815.0 ;
      RECT  10242.5 24470.0 10307.5 24655.0 ;
      RECT  9692.5 25472.5 9757.5 25607.5 ;
      RECT  9882.5 25472.5 9947.5 25607.5 ;
      RECT  9882.5 25472.5 9947.5 25607.5 ;
      RECT  9692.5 25472.5 9757.5 25607.5 ;
      RECT  9882.5 25472.5 9947.5 25607.5 ;
      RECT  10072.5 25472.5 10137.5 25607.5 ;
      RECT  10072.5 25472.5 10137.5 25607.5 ;
      RECT  9882.5 25472.5 9947.5 25607.5 ;
      RECT  9692.5 24632.5 9757.5 24767.5 ;
      RECT  9882.5 24632.5 9947.5 24767.5 ;
      RECT  9882.5 24632.5 9947.5 24767.5 ;
      RECT  9692.5 24632.5 9757.5 24767.5 ;
      RECT  9882.5 24632.5 9947.5 24767.5 ;
      RECT  10072.5 24632.5 10137.5 24767.5 ;
      RECT  10072.5 24632.5 10137.5 24767.5 ;
      RECT  9882.5 24632.5 9947.5 24767.5 ;
      RECT  10242.5 25562.5 10307.5 25697.5 ;
      RECT  10242.5 24587.5 10307.5 24722.5 ;
      RECT  10077.5 24862.5 9942.5 24927.5 ;
      RECT  9820.0 25077.5 9685.0 25142.5 ;
      RECT  9882.5 25472.5 9947.5 25607.5 ;
      RECT  10072.5 24632.5 10137.5 24767.5 ;
      RECT  10172.5 25077.5 10037.5 25142.5 ;
      RECT  9685.0 25077.5 9820.0 25142.5 ;
      RECT  9942.5 24862.5 10077.5 24927.5 ;
      RECT  10037.5 25077.5 10172.5 25142.5 ;
      RECT  9625.0 25782.5 10545.0 25847.5 ;
      RECT  9625.0 24437.5 10545.0 24502.5 ;
      RECT  10972.5 25630.0 11037.5 25815.0 ;
      RECT  10972.5 24470.0 11037.5 24655.0 ;
      RECT  10612.5 24587.5 10677.5 24437.5 ;
      RECT  10612.5 25472.5 10677.5 25847.5 ;
      RECT  10802.5 24587.5 10867.5 25472.5 ;
      RECT  10612.5 25472.5 10677.5 25607.5 ;
      RECT  10802.5 25472.5 10867.5 25607.5 ;
      RECT  10802.5 25472.5 10867.5 25607.5 ;
      RECT  10612.5 25472.5 10677.5 25607.5 ;
      RECT  10612.5 24587.5 10677.5 24722.5 ;
      RECT  10802.5 24587.5 10867.5 24722.5 ;
      RECT  10802.5 24587.5 10867.5 24722.5 ;
      RECT  10612.5 24587.5 10677.5 24722.5 ;
      RECT  10972.5 25562.5 11037.5 25697.5 ;
      RECT  10972.5 24587.5 11037.5 24722.5 ;
      RECT  10670.0 25030.0 10735.0 25165.0 ;
      RECT  10670.0 25030.0 10735.0 25165.0 ;
      RECT  10835.0 25065.0 10900.0 25130.0 ;
      RECT  10545.0 25782.5 11105.0 25847.5 ;
      RECT  10545.0 24437.5 11105.0 24502.5 ;
      RECT  8807.5 25030.0 8872.5 25165.0 ;
      RECT  8947.5 24757.5 9012.5 24892.5 ;
      RECT  9942.5 24862.5 9807.5 24927.5 ;
      RECT  9492.5 26000.0 9557.5 25815.0 ;
      RECT  9492.5 27160.0 9557.5 26975.0 ;
      RECT  9132.5 27042.5 9197.5 27192.5 ;
      RECT  9132.5 26157.5 9197.5 25782.5 ;
      RECT  9322.5 27042.5 9387.5 26157.5 ;
      RECT  9132.5 26157.5 9197.5 26022.5 ;
      RECT  9322.5 26157.5 9387.5 26022.5 ;
      RECT  9322.5 26157.5 9387.5 26022.5 ;
      RECT  9132.5 26157.5 9197.5 26022.5 ;
      RECT  9132.5 27042.5 9197.5 26907.5 ;
      RECT  9322.5 27042.5 9387.5 26907.5 ;
      RECT  9322.5 27042.5 9387.5 26907.5 ;
      RECT  9132.5 27042.5 9197.5 26907.5 ;
      RECT  9492.5 26067.5 9557.5 25932.5 ;
      RECT  9492.5 27042.5 9557.5 26907.5 ;
      RECT  9190.0 26600.0 9255.0 26465.0 ;
      RECT  9190.0 26600.0 9255.0 26465.0 ;
      RECT  9355.0 26565.0 9420.0 26500.0 ;
      RECT  9065.0 25847.5 9625.0 25782.5 ;
      RECT  9065.0 27192.5 9625.0 27127.5 ;
      RECT  9692.5 26997.5 9757.5 27192.5 ;
      RECT  9692.5 26157.5 9757.5 25782.5 ;
      RECT  10072.5 26157.5 10137.5 25782.5 ;
      RECT  10242.5 26000.0 10307.5 25815.0 ;
      RECT  10242.5 27160.0 10307.5 26975.0 ;
      RECT  9692.5 26157.5 9757.5 26022.5 ;
      RECT  9882.5 26157.5 9947.5 26022.5 ;
      RECT  9882.5 26157.5 9947.5 26022.5 ;
      RECT  9692.5 26157.5 9757.5 26022.5 ;
      RECT  9882.5 26157.5 9947.5 26022.5 ;
      RECT  10072.5 26157.5 10137.5 26022.5 ;
      RECT  10072.5 26157.5 10137.5 26022.5 ;
      RECT  9882.5 26157.5 9947.5 26022.5 ;
      RECT  9692.5 26997.5 9757.5 26862.5 ;
      RECT  9882.5 26997.5 9947.5 26862.5 ;
      RECT  9882.5 26997.5 9947.5 26862.5 ;
      RECT  9692.5 26997.5 9757.5 26862.5 ;
      RECT  9882.5 26997.5 9947.5 26862.5 ;
      RECT  10072.5 26997.5 10137.5 26862.5 ;
      RECT  10072.5 26997.5 10137.5 26862.5 ;
      RECT  9882.5 26997.5 9947.5 26862.5 ;
      RECT  10242.5 26067.5 10307.5 25932.5 ;
      RECT  10242.5 27042.5 10307.5 26907.5 ;
      RECT  10077.5 26767.5 9942.5 26702.5 ;
      RECT  9820.0 26552.5 9685.0 26487.5 ;
      RECT  9882.5 26157.5 9947.5 26022.5 ;
      RECT  10072.5 26997.5 10137.5 26862.5 ;
      RECT  10172.5 26552.5 10037.5 26487.5 ;
      RECT  9685.0 26552.5 9820.0 26487.5 ;
      RECT  9942.5 26767.5 10077.5 26702.5 ;
      RECT  10037.5 26552.5 10172.5 26487.5 ;
      RECT  9625.0 25847.5 10545.0 25782.5 ;
      RECT  9625.0 27192.5 10545.0 27127.5 ;
      RECT  10972.5 26000.0 11037.5 25815.0 ;
      RECT  10972.5 27160.0 11037.5 26975.0 ;
      RECT  10612.5 27042.5 10677.5 27192.5 ;
      RECT  10612.5 26157.5 10677.5 25782.5 ;
      RECT  10802.5 27042.5 10867.5 26157.5 ;
      RECT  10612.5 26157.5 10677.5 26022.5 ;
      RECT  10802.5 26157.5 10867.5 26022.5 ;
      RECT  10802.5 26157.5 10867.5 26022.5 ;
      RECT  10612.5 26157.5 10677.5 26022.5 ;
      RECT  10612.5 27042.5 10677.5 26907.5 ;
      RECT  10802.5 27042.5 10867.5 26907.5 ;
      RECT  10802.5 27042.5 10867.5 26907.5 ;
      RECT  10612.5 27042.5 10677.5 26907.5 ;
      RECT  10972.5 26067.5 11037.5 25932.5 ;
      RECT  10972.5 27042.5 11037.5 26907.5 ;
      RECT  10670.0 26600.0 10735.0 26465.0 ;
      RECT  10670.0 26600.0 10735.0 26465.0 ;
      RECT  10835.0 26565.0 10900.0 26500.0 ;
      RECT  10545.0 25847.5 11105.0 25782.5 ;
      RECT  10545.0 27192.5 11105.0 27127.5 ;
      RECT  8807.5 26465.0 8872.5 26600.0 ;
      RECT  8947.5 26737.5 9012.5 26872.5 ;
      RECT  9942.5 26702.5 9807.5 26767.5 ;
      RECT  9492.5 28320.0 9557.5 28505.0 ;
      RECT  9492.5 27160.0 9557.5 27345.0 ;
      RECT  9132.5 27277.5 9197.5 27127.5 ;
      RECT  9132.5 28162.5 9197.5 28537.5 ;
      RECT  9322.5 27277.5 9387.5 28162.5 ;
      RECT  9132.5 28162.5 9197.5 28297.5 ;
      RECT  9322.5 28162.5 9387.5 28297.5 ;
      RECT  9322.5 28162.5 9387.5 28297.5 ;
      RECT  9132.5 28162.5 9197.5 28297.5 ;
      RECT  9132.5 27277.5 9197.5 27412.5 ;
      RECT  9322.5 27277.5 9387.5 27412.5 ;
      RECT  9322.5 27277.5 9387.5 27412.5 ;
      RECT  9132.5 27277.5 9197.5 27412.5 ;
      RECT  9492.5 28252.5 9557.5 28387.5 ;
      RECT  9492.5 27277.5 9557.5 27412.5 ;
      RECT  9190.0 27720.0 9255.0 27855.0 ;
      RECT  9190.0 27720.0 9255.0 27855.0 ;
      RECT  9355.0 27755.0 9420.0 27820.0 ;
      RECT  9065.0 28472.5 9625.0 28537.5 ;
      RECT  9065.0 27127.5 9625.0 27192.5 ;
      RECT  9692.5 27322.5 9757.5 27127.5 ;
      RECT  9692.5 28162.5 9757.5 28537.5 ;
      RECT  10072.5 28162.5 10137.5 28537.5 ;
      RECT  10242.5 28320.0 10307.5 28505.0 ;
      RECT  10242.5 27160.0 10307.5 27345.0 ;
      RECT  9692.5 28162.5 9757.5 28297.5 ;
      RECT  9882.5 28162.5 9947.5 28297.5 ;
      RECT  9882.5 28162.5 9947.5 28297.5 ;
      RECT  9692.5 28162.5 9757.5 28297.5 ;
      RECT  9882.5 28162.5 9947.5 28297.5 ;
      RECT  10072.5 28162.5 10137.5 28297.5 ;
      RECT  10072.5 28162.5 10137.5 28297.5 ;
      RECT  9882.5 28162.5 9947.5 28297.5 ;
      RECT  9692.5 27322.5 9757.5 27457.5 ;
      RECT  9882.5 27322.5 9947.5 27457.5 ;
      RECT  9882.5 27322.5 9947.5 27457.5 ;
      RECT  9692.5 27322.5 9757.5 27457.5 ;
      RECT  9882.5 27322.5 9947.5 27457.5 ;
      RECT  10072.5 27322.5 10137.5 27457.5 ;
      RECT  10072.5 27322.5 10137.5 27457.5 ;
      RECT  9882.5 27322.5 9947.5 27457.5 ;
      RECT  10242.5 28252.5 10307.5 28387.5 ;
      RECT  10242.5 27277.5 10307.5 27412.5 ;
      RECT  10077.5 27552.5 9942.5 27617.5 ;
      RECT  9820.0 27767.5 9685.0 27832.5 ;
      RECT  9882.5 28162.5 9947.5 28297.5 ;
      RECT  10072.5 27322.5 10137.5 27457.5 ;
      RECT  10172.5 27767.5 10037.5 27832.5 ;
      RECT  9685.0 27767.5 9820.0 27832.5 ;
      RECT  9942.5 27552.5 10077.5 27617.5 ;
      RECT  10037.5 27767.5 10172.5 27832.5 ;
      RECT  9625.0 28472.5 10545.0 28537.5 ;
      RECT  9625.0 27127.5 10545.0 27192.5 ;
      RECT  10972.5 28320.0 11037.5 28505.0 ;
      RECT  10972.5 27160.0 11037.5 27345.0 ;
      RECT  10612.5 27277.5 10677.5 27127.5 ;
      RECT  10612.5 28162.5 10677.5 28537.5 ;
      RECT  10802.5 27277.5 10867.5 28162.5 ;
      RECT  10612.5 28162.5 10677.5 28297.5 ;
      RECT  10802.5 28162.5 10867.5 28297.5 ;
      RECT  10802.5 28162.5 10867.5 28297.5 ;
      RECT  10612.5 28162.5 10677.5 28297.5 ;
      RECT  10612.5 27277.5 10677.5 27412.5 ;
      RECT  10802.5 27277.5 10867.5 27412.5 ;
      RECT  10802.5 27277.5 10867.5 27412.5 ;
      RECT  10612.5 27277.5 10677.5 27412.5 ;
      RECT  10972.5 28252.5 11037.5 28387.5 ;
      RECT  10972.5 27277.5 11037.5 27412.5 ;
      RECT  10670.0 27720.0 10735.0 27855.0 ;
      RECT  10670.0 27720.0 10735.0 27855.0 ;
      RECT  10835.0 27755.0 10900.0 27820.0 ;
      RECT  10545.0 28472.5 11105.0 28537.5 ;
      RECT  10545.0 27127.5 11105.0 27192.5 ;
      RECT  8807.5 27720.0 8872.5 27855.0 ;
      RECT  8947.5 27447.5 9012.5 27582.5 ;
      RECT  9942.5 27552.5 9807.5 27617.5 ;
      RECT  9492.5 28690.0 9557.5 28505.0 ;
      RECT  9492.5 29850.0 9557.5 29665.0 ;
      RECT  9132.5 29732.5 9197.5 29882.5 ;
      RECT  9132.5 28847.5 9197.5 28472.5 ;
      RECT  9322.5 29732.5 9387.5 28847.5 ;
      RECT  9132.5 28847.5 9197.5 28712.5 ;
      RECT  9322.5 28847.5 9387.5 28712.5 ;
      RECT  9322.5 28847.5 9387.5 28712.5 ;
      RECT  9132.5 28847.5 9197.5 28712.5 ;
      RECT  9132.5 29732.5 9197.5 29597.5 ;
      RECT  9322.5 29732.5 9387.5 29597.5 ;
      RECT  9322.5 29732.5 9387.5 29597.5 ;
      RECT  9132.5 29732.5 9197.5 29597.5 ;
      RECT  9492.5 28757.5 9557.5 28622.5 ;
      RECT  9492.5 29732.5 9557.5 29597.5 ;
      RECT  9190.0 29290.0 9255.0 29155.0 ;
      RECT  9190.0 29290.0 9255.0 29155.0 ;
      RECT  9355.0 29255.0 9420.0 29190.0 ;
      RECT  9065.0 28537.5 9625.0 28472.5 ;
      RECT  9065.0 29882.5 9625.0 29817.5 ;
      RECT  9692.5 29687.5 9757.5 29882.5 ;
      RECT  9692.5 28847.5 9757.5 28472.5 ;
      RECT  10072.5 28847.5 10137.5 28472.5 ;
      RECT  10242.5 28690.0 10307.5 28505.0 ;
      RECT  10242.5 29850.0 10307.5 29665.0 ;
      RECT  9692.5 28847.5 9757.5 28712.5 ;
      RECT  9882.5 28847.5 9947.5 28712.5 ;
      RECT  9882.5 28847.5 9947.5 28712.5 ;
      RECT  9692.5 28847.5 9757.5 28712.5 ;
      RECT  9882.5 28847.5 9947.5 28712.5 ;
      RECT  10072.5 28847.5 10137.5 28712.5 ;
      RECT  10072.5 28847.5 10137.5 28712.5 ;
      RECT  9882.5 28847.5 9947.5 28712.5 ;
      RECT  9692.5 29687.5 9757.5 29552.5 ;
      RECT  9882.5 29687.5 9947.5 29552.5 ;
      RECT  9882.5 29687.5 9947.5 29552.5 ;
      RECT  9692.5 29687.5 9757.5 29552.5 ;
      RECT  9882.5 29687.5 9947.5 29552.5 ;
      RECT  10072.5 29687.5 10137.5 29552.5 ;
      RECT  10072.5 29687.5 10137.5 29552.5 ;
      RECT  9882.5 29687.5 9947.5 29552.5 ;
      RECT  10242.5 28757.5 10307.5 28622.5 ;
      RECT  10242.5 29732.5 10307.5 29597.5 ;
      RECT  10077.5 29457.5 9942.5 29392.5 ;
      RECT  9820.0 29242.5 9685.0 29177.5 ;
      RECT  9882.5 28847.5 9947.5 28712.5 ;
      RECT  10072.5 29687.5 10137.5 29552.5 ;
      RECT  10172.5 29242.5 10037.5 29177.5 ;
      RECT  9685.0 29242.5 9820.0 29177.5 ;
      RECT  9942.5 29457.5 10077.5 29392.5 ;
      RECT  10037.5 29242.5 10172.5 29177.5 ;
      RECT  9625.0 28537.5 10545.0 28472.5 ;
      RECT  9625.0 29882.5 10545.0 29817.5 ;
      RECT  10972.5 28690.0 11037.5 28505.0 ;
      RECT  10972.5 29850.0 11037.5 29665.0 ;
      RECT  10612.5 29732.5 10677.5 29882.5 ;
      RECT  10612.5 28847.5 10677.5 28472.5 ;
      RECT  10802.5 29732.5 10867.5 28847.5 ;
      RECT  10612.5 28847.5 10677.5 28712.5 ;
      RECT  10802.5 28847.5 10867.5 28712.5 ;
      RECT  10802.5 28847.5 10867.5 28712.5 ;
      RECT  10612.5 28847.5 10677.5 28712.5 ;
      RECT  10612.5 29732.5 10677.5 29597.5 ;
      RECT  10802.5 29732.5 10867.5 29597.5 ;
      RECT  10802.5 29732.5 10867.5 29597.5 ;
      RECT  10612.5 29732.5 10677.5 29597.5 ;
      RECT  10972.5 28757.5 11037.5 28622.5 ;
      RECT  10972.5 29732.5 11037.5 29597.5 ;
      RECT  10670.0 29290.0 10735.0 29155.0 ;
      RECT  10670.0 29290.0 10735.0 29155.0 ;
      RECT  10835.0 29255.0 10900.0 29190.0 ;
      RECT  10545.0 28537.5 11105.0 28472.5 ;
      RECT  10545.0 29882.5 11105.0 29817.5 ;
      RECT  8807.5 29155.0 8872.5 29290.0 ;
      RECT  8947.5 29427.5 9012.5 29562.5 ;
      RECT  9942.5 29392.5 9807.5 29457.5 ;
      RECT  9492.5 31010.0 9557.5 31195.0 ;
      RECT  9492.5 29850.0 9557.5 30035.0 ;
      RECT  9132.5 29967.5 9197.5 29817.5 ;
      RECT  9132.5 30852.5 9197.5 31227.5 ;
      RECT  9322.5 29967.5 9387.5 30852.5 ;
      RECT  9132.5 30852.5 9197.5 30987.5 ;
      RECT  9322.5 30852.5 9387.5 30987.5 ;
      RECT  9322.5 30852.5 9387.5 30987.5 ;
      RECT  9132.5 30852.5 9197.5 30987.5 ;
      RECT  9132.5 29967.5 9197.5 30102.5 ;
      RECT  9322.5 29967.5 9387.5 30102.5 ;
      RECT  9322.5 29967.5 9387.5 30102.5 ;
      RECT  9132.5 29967.5 9197.5 30102.5 ;
      RECT  9492.5 30942.5 9557.5 31077.5 ;
      RECT  9492.5 29967.5 9557.5 30102.5 ;
      RECT  9190.0 30410.0 9255.0 30545.0 ;
      RECT  9190.0 30410.0 9255.0 30545.0 ;
      RECT  9355.0 30445.0 9420.0 30510.0 ;
      RECT  9065.0 31162.5 9625.0 31227.5 ;
      RECT  9065.0 29817.5 9625.0 29882.5 ;
      RECT  9692.5 30012.5 9757.5 29817.5 ;
      RECT  9692.5 30852.5 9757.5 31227.5 ;
      RECT  10072.5 30852.5 10137.5 31227.5 ;
      RECT  10242.5 31010.0 10307.5 31195.0 ;
      RECT  10242.5 29850.0 10307.5 30035.0 ;
      RECT  9692.5 30852.5 9757.5 30987.5 ;
      RECT  9882.5 30852.5 9947.5 30987.5 ;
      RECT  9882.5 30852.5 9947.5 30987.5 ;
      RECT  9692.5 30852.5 9757.5 30987.5 ;
      RECT  9882.5 30852.5 9947.5 30987.5 ;
      RECT  10072.5 30852.5 10137.5 30987.5 ;
      RECT  10072.5 30852.5 10137.5 30987.5 ;
      RECT  9882.5 30852.5 9947.5 30987.5 ;
      RECT  9692.5 30012.5 9757.5 30147.5 ;
      RECT  9882.5 30012.5 9947.5 30147.5 ;
      RECT  9882.5 30012.5 9947.5 30147.5 ;
      RECT  9692.5 30012.5 9757.5 30147.5 ;
      RECT  9882.5 30012.5 9947.5 30147.5 ;
      RECT  10072.5 30012.5 10137.5 30147.5 ;
      RECT  10072.5 30012.5 10137.5 30147.5 ;
      RECT  9882.5 30012.5 9947.5 30147.5 ;
      RECT  10242.5 30942.5 10307.5 31077.5 ;
      RECT  10242.5 29967.5 10307.5 30102.5 ;
      RECT  10077.5 30242.5 9942.5 30307.5 ;
      RECT  9820.0 30457.5 9685.0 30522.5 ;
      RECT  9882.5 30852.5 9947.5 30987.5 ;
      RECT  10072.5 30012.5 10137.5 30147.5 ;
      RECT  10172.5 30457.5 10037.5 30522.5 ;
      RECT  9685.0 30457.5 9820.0 30522.5 ;
      RECT  9942.5 30242.5 10077.5 30307.5 ;
      RECT  10037.5 30457.5 10172.5 30522.5 ;
      RECT  9625.0 31162.5 10545.0 31227.5 ;
      RECT  9625.0 29817.5 10545.0 29882.5 ;
      RECT  10972.5 31010.0 11037.5 31195.0 ;
      RECT  10972.5 29850.0 11037.5 30035.0 ;
      RECT  10612.5 29967.5 10677.5 29817.5 ;
      RECT  10612.5 30852.5 10677.5 31227.5 ;
      RECT  10802.5 29967.5 10867.5 30852.5 ;
      RECT  10612.5 30852.5 10677.5 30987.5 ;
      RECT  10802.5 30852.5 10867.5 30987.5 ;
      RECT  10802.5 30852.5 10867.5 30987.5 ;
      RECT  10612.5 30852.5 10677.5 30987.5 ;
      RECT  10612.5 29967.5 10677.5 30102.5 ;
      RECT  10802.5 29967.5 10867.5 30102.5 ;
      RECT  10802.5 29967.5 10867.5 30102.5 ;
      RECT  10612.5 29967.5 10677.5 30102.5 ;
      RECT  10972.5 30942.5 11037.5 31077.5 ;
      RECT  10972.5 29967.5 11037.5 30102.5 ;
      RECT  10670.0 30410.0 10735.0 30545.0 ;
      RECT  10670.0 30410.0 10735.0 30545.0 ;
      RECT  10835.0 30445.0 10900.0 30510.0 ;
      RECT  10545.0 31162.5 11105.0 31227.5 ;
      RECT  10545.0 29817.5 11105.0 29882.5 ;
      RECT  8807.5 30410.0 8872.5 30545.0 ;
      RECT  8947.5 30137.5 9012.5 30272.5 ;
      RECT  9942.5 30242.5 9807.5 30307.5 ;
      RECT  9492.5 31380.0 9557.5 31195.0 ;
      RECT  9492.5 32540.0 9557.5 32355.0 ;
      RECT  9132.5 32422.5 9197.5 32572.5 ;
      RECT  9132.5 31537.5 9197.5 31162.5 ;
      RECT  9322.5 32422.5 9387.5 31537.5 ;
      RECT  9132.5 31537.5 9197.5 31402.5 ;
      RECT  9322.5 31537.5 9387.5 31402.5 ;
      RECT  9322.5 31537.5 9387.5 31402.5 ;
      RECT  9132.5 31537.5 9197.5 31402.5 ;
      RECT  9132.5 32422.5 9197.5 32287.5 ;
      RECT  9322.5 32422.5 9387.5 32287.5 ;
      RECT  9322.5 32422.5 9387.5 32287.5 ;
      RECT  9132.5 32422.5 9197.5 32287.5 ;
      RECT  9492.5 31447.5 9557.5 31312.5 ;
      RECT  9492.5 32422.5 9557.5 32287.5 ;
      RECT  9190.0 31980.0 9255.0 31845.0 ;
      RECT  9190.0 31980.0 9255.0 31845.0 ;
      RECT  9355.0 31945.0 9420.0 31880.0 ;
      RECT  9065.0 31227.5 9625.0 31162.5 ;
      RECT  9065.0 32572.5 9625.0 32507.5 ;
      RECT  9692.5 32377.5 9757.5 32572.5 ;
      RECT  9692.5 31537.5 9757.5 31162.5 ;
      RECT  10072.5 31537.5 10137.5 31162.5 ;
      RECT  10242.5 31380.0 10307.5 31195.0 ;
      RECT  10242.5 32540.0 10307.5 32355.0 ;
      RECT  9692.5 31537.5 9757.5 31402.5 ;
      RECT  9882.5 31537.5 9947.5 31402.5 ;
      RECT  9882.5 31537.5 9947.5 31402.5 ;
      RECT  9692.5 31537.5 9757.5 31402.5 ;
      RECT  9882.5 31537.5 9947.5 31402.5 ;
      RECT  10072.5 31537.5 10137.5 31402.5 ;
      RECT  10072.5 31537.5 10137.5 31402.5 ;
      RECT  9882.5 31537.5 9947.5 31402.5 ;
      RECT  9692.5 32377.5 9757.5 32242.5 ;
      RECT  9882.5 32377.5 9947.5 32242.5 ;
      RECT  9882.5 32377.5 9947.5 32242.5 ;
      RECT  9692.5 32377.5 9757.5 32242.5 ;
      RECT  9882.5 32377.5 9947.5 32242.5 ;
      RECT  10072.5 32377.5 10137.5 32242.5 ;
      RECT  10072.5 32377.5 10137.5 32242.5 ;
      RECT  9882.5 32377.5 9947.5 32242.5 ;
      RECT  10242.5 31447.5 10307.5 31312.5 ;
      RECT  10242.5 32422.5 10307.5 32287.5 ;
      RECT  10077.5 32147.5 9942.5 32082.5 ;
      RECT  9820.0 31932.5 9685.0 31867.5 ;
      RECT  9882.5 31537.5 9947.5 31402.5 ;
      RECT  10072.5 32377.5 10137.5 32242.5 ;
      RECT  10172.5 31932.5 10037.5 31867.5 ;
      RECT  9685.0 31932.5 9820.0 31867.5 ;
      RECT  9942.5 32147.5 10077.5 32082.5 ;
      RECT  10037.5 31932.5 10172.5 31867.5 ;
      RECT  9625.0 31227.5 10545.0 31162.5 ;
      RECT  9625.0 32572.5 10545.0 32507.5 ;
      RECT  10972.5 31380.0 11037.5 31195.0 ;
      RECT  10972.5 32540.0 11037.5 32355.0 ;
      RECT  10612.5 32422.5 10677.5 32572.5 ;
      RECT  10612.5 31537.5 10677.5 31162.5 ;
      RECT  10802.5 32422.5 10867.5 31537.5 ;
      RECT  10612.5 31537.5 10677.5 31402.5 ;
      RECT  10802.5 31537.5 10867.5 31402.5 ;
      RECT  10802.5 31537.5 10867.5 31402.5 ;
      RECT  10612.5 31537.5 10677.5 31402.5 ;
      RECT  10612.5 32422.5 10677.5 32287.5 ;
      RECT  10802.5 32422.5 10867.5 32287.5 ;
      RECT  10802.5 32422.5 10867.5 32287.5 ;
      RECT  10612.5 32422.5 10677.5 32287.5 ;
      RECT  10972.5 31447.5 11037.5 31312.5 ;
      RECT  10972.5 32422.5 11037.5 32287.5 ;
      RECT  10670.0 31980.0 10735.0 31845.0 ;
      RECT  10670.0 31980.0 10735.0 31845.0 ;
      RECT  10835.0 31945.0 10900.0 31880.0 ;
      RECT  10545.0 31227.5 11105.0 31162.5 ;
      RECT  10545.0 32572.5 11105.0 32507.5 ;
      RECT  8807.5 31845.0 8872.5 31980.0 ;
      RECT  8947.5 32117.5 9012.5 32252.5 ;
      RECT  9942.5 32082.5 9807.5 32147.5 ;
      RECT  9492.5 33700.0 9557.5 33885.0 ;
      RECT  9492.5 32540.0 9557.5 32725.0 ;
      RECT  9132.5 32657.5 9197.5 32507.5 ;
      RECT  9132.5 33542.5 9197.5 33917.5 ;
      RECT  9322.5 32657.5 9387.5 33542.5 ;
      RECT  9132.5 33542.5 9197.5 33677.5 ;
      RECT  9322.5 33542.5 9387.5 33677.5 ;
      RECT  9322.5 33542.5 9387.5 33677.5 ;
      RECT  9132.5 33542.5 9197.5 33677.5 ;
      RECT  9132.5 32657.5 9197.5 32792.5 ;
      RECT  9322.5 32657.5 9387.5 32792.5 ;
      RECT  9322.5 32657.5 9387.5 32792.5 ;
      RECT  9132.5 32657.5 9197.5 32792.5 ;
      RECT  9492.5 33632.5 9557.5 33767.5 ;
      RECT  9492.5 32657.5 9557.5 32792.5 ;
      RECT  9190.0 33100.0 9255.0 33235.0 ;
      RECT  9190.0 33100.0 9255.0 33235.0 ;
      RECT  9355.0 33135.0 9420.0 33200.0 ;
      RECT  9065.0 33852.5 9625.0 33917.5 ;
      RECT  9065.0 32507.5 9625.0 32572.5 ;
      RECT  9692.5 32702.5 9757.5 32507.5 ;
      RECT  9692.5 33542.5 9757.5 33917.5 ;
      RECT  10072.5 33542.5 10137.5 33917.5 ;
      RECT  10242.5 33700.0 10307.5 33885.0 ;
      RECT  10242.5 32540.0 10307.5 32725.0 ;
      RECT  9692.5 33542.5 9757.5 33677.5 ;
      RECT  9882.5 33542.5 9947.5 33677.5 ;
      RECT  9882.5 33542.5 9947.5 33677.5 ;
      RECT  9692.5 33542.5 9757.5 33677.5 ;
      RECT  9882.5 33542.5 9947.5 33677.5 ;
      RECT  10072.5 33542.5 10137.5 33677.5 ;
      RECT  10072.5 33542.5 10137.5 33677.5 ;
      RECT  9882.5 33542.5 9947.5 33677.5 ;
      RECT  9692.5 32702.5 9757.5 32837.5 ;
      RECT  9882.5 32702.5 9947.5 32837.5 ;
      RECT  9882.5 32702.5 9947.5 32837.5 ;
      RECT  9692.5 32702.5 9757.5 32837.5 ;
      RECT  9882.5 32702.5 9947.5 32837.5 ;
      RECT  10072.5 32702.5 10137.5 32837.5 ;
      RECT  10072.5 32702.5 10137.5 32837.5 ;
      RECT  9882.5 32702.5 9947.5 32837.5 ;
      RECT  10242.5 33632.5 10307.5 33767.5 ;
      RECT  10242.5 32657.5 10307.5 32792.5 ;
      RECT  10077.5 32932.5 9942.5 32997.5 ;
      RECT  9820.0 33147.5 9685.0 33212.5 ;
      RECT  9882.5 33542.5 9947.5 33677.5 ;
      RECT  10072.5 32702.5 10137.5 32837.5 ;
      RECT  10172.5 33147.5 10037.5 33212.5 ;
      RECT  9685.0 33147.5 9820.0 33212.5 ;
      RECT  9942.5 32932.5 10077.5 32997.5 ;
      RECT  10037.5 33147.5 10172.5 33212.5 ;
      RECT  9625.0 33852.5 10545.0 33917.5 ;
      RECT  9625.0 32507.5 10545.0 32572.5 ;
      RECT  10972.5 33700.0 11037.5 33885.0 ;
      RECT  10972.5 32540.0 11037.5 32725.0 ;
      RECT  10612.5 32657.5 10677.5 32507.5 ;
      RECT  10612.5 33542.5 10677.5 33917.5 ;
      RECT  10802.5 32657.5 10867.5 33542.5 ;
      RECT  10612.5 33542.5 10677.5 33677.5 ;
      RECT  10802.5 33542.5 10867.5 33677.5 ;
      RECT  10802.5 33542.5 10867.5 33677.5 ;
      RECT  10612.5 33542.5 10677.5 33677.5 ;
      RECT  10612.5 32657.5 10677.5 32792.5 ;
      RECT  10802.5 32657.5 10867.5 32792.5 ;
      RECT  10802.5 32657.5 10867.5 32792.5 ;
      RECT  10612.5 32657.5 10677.5 32792.5 ;
      RECT  10972.5 33632.5 11037.5 33767.5 ;
      RECT  10972.5 32657.5 11037.5 32792.5 ;
      RECT  10670.0 33100.0 10735.0 33235.0 ;
      RECT  10670.0 33100.0 10735.0 33235.0 ;
      RECT  10835.0 33135.0 10900.0 33200.0 ;
      RECT  10545.0 33852.5 11105.0 33917.5 ;
      RECT  10545.0 32507.5 11105.0 32572.5 ;
      RECT  8807.5 33100.0 8872.5 33235.0 ;
      RECT  8947.5 32827.5 9012.5 32962.5 ;
      RECT  9942.5 32932.5 9807.5 32997.5 ;
      RECT  9492.5 34070.0 9557.5 33885.0 ;
      RECT  9492.5 35230.0 9557.5 35045.0 ;
      RECT  9132.5 35112.5 9197.5 35262.5 ;
      RECT  9132.5 34227.5 9197.5 33852.5 ;
      RECT  9322.5 35112.5 9387.5 34227.5 ;
      RECT  9132.5 34227.5 9197.5 34092.5 ;
      RECT  9322.5 34227.5 9387.5 34092.5 ;
      RECT  9322.5 34227.5 9387.5 34092.5 ;
      RECT  9132.5 34227.5 9197.5 34092.5 ;
      RECT  9132.5 35112.5 9197.5 34977.5 ;
      RECT  9322.5 35112.5 9387.5 34977.5 ;
      RECT  9322.5 35112.5 9387.5 34977.5 ;
      RECT  9132.5 35112.5 9197.5 34977.5 ;
      RECT  9492.5 34137.5 9557.5 34002.5 ;
      RECT  9492.5 35112.5 9557.5 34977.5 ;
      RECT  9190.0 34670.0 9255.0 34535.0 ;
      RECT  9190.0 34670.0 9255.0 34535.0 ;
      RECT  9355.0 34635.0 9420.0 34570.0 ;
      RECT  9065.0 33917.5 9625.0 33852.5 ;
      RECT  9065.0 35262.5 9625.0 35197.5 ;
      RECT  9692.5 35067.5 9757.5 35262.5 ;
      RECT  9692.5 34227.5 9757.5 33852.5 ;
      RECT  10072.5 34227.5 10137.5 33852.5 ;
      RECT  10242.5 34070.0 10307.5 33885.0 ;
      RECT  10242.5 35230.0 10307.5 35045.0 ;
      RECT  9692.5 34227.5 9757.5 34092.5 ;
      RECT  9882.5 34227.5 9947.5 34092.5 ;
      RECT  9882.5 34227.5 9947.5 34092.5 ;
      RECT  9692.5 34227.5 9757.5 34092.5 ;
      RECT  9882.5 34227.5 9947.5 34092.5 ;
      RECT  10072.5 34227.5 10137.5 34092.5 ;
      RECT  10072.5 34227.5 10137.5 34092.5 ;
      RECT  9882.5 34227.5 9947.5 34092.5 ;
      RECT  9692.5 35067.5 9757.5 34932.5 ;
      RECT  9882.5 35067.5 9947.5 34932.5 ;
      RECT  9882.5 35067.5 9947.5 34932.5 ;
      RECT  9692.5 35067.5 9757.5 34932.5 ;
      RECT  9882.5 35067.5 9947.5 34932.5 ;
      RECT  10072.5 35067.5 10137.5 34932.5 ;
      RECT  10072.5 35067.5 10137.5 34932.5 ;
      RECT  9882.5 35067.5 9947.5 34932.5 ;
      RECT  10242.5 34137.5 10307.5 34002.5 ;
      RECT  10242.5 35112.5 10307.5 34977.5 ;
      RECT  10077.5 34837.5 9942.5 34772.5 ;
      RECT  9820.0 34622.5 9685.0 34557.5 ;
      RECT  9882.5 34227.5 9947.5 34092.5 ;
      RECT  10072.5 35067.5 10137.5 34932.5 ;
      RECT  10172.5 34622.5 10037.5 34557.5 ;
      RECT  9685.0 34622.5 9820.0 34557.5 ;
      RECT  9942.5 34837.5 10077.5 34772.5 ;
      RECT  10037.5 34622.5 10172.5 34557.5 ;
      RECT  9625.0 33917.5 10545.0 33852.5 ;
      RECT  9625.0 35262.5 10545.0 35197.5 ;
      RECT  10972.5 34070.0 11037.5 33885.0 ;
      RECT  10972.5 35230.0 11037.5 35045.0 ;
      RECT  10612.5 35112.5 10677.5 35262.5 ;
      RECT  10612.5 34227.5 10677.5 33852.5 ;
      RECT  10802.5 35112.5 10867.5 34227.5 ;
      RECT  10612.5 34227.5 10677.5 34092.5 ;
      RECT  10802.5 34227.5 10867.5 34092.5 ;
      RECT  10802.5 34227.5 10867.5 34092.5 ;
      RECT  10612.5 34227.5 10677.5 34092.5 ;
      RECT  10612.5 35112.5 10677.5 34977.5 ;
      RECT  10802.5 35112.5 10867.5 34977.5 ;
      RECT  10802.5 35112.5 10867.5 34977.5 ;
      RECT  10612.5 35112.5 10677.5 34977.5 ;
      RECT  10972.5 34137.5 11037.5 34002.5 ;
      RECT  10972.5 35112.5 11037.5 34977.5 ;
      RECT  10670.0 34670.0 10735.0 34535.0 ;
      RECT  10670.0 34670.0 10735.0 34535.0 ;
      RECT  10835.0 34635.0 10900.0 34570.0 ;
      RECT  10545.0 33917.5 11105.0 33852.5 ;
      RECT  10545.0 35262.5 11105.0 35197.5 ;
      RECT  8807.5 34535.0 8872.5 34670.0 ;
      RECT  8947.5 34807.5 9012.5 34942.5 ;
      RECT  9942.5 34772.5 9807.5 34837.5 ;
      RECT  9492.5 36390.0 9557.5 36575.0 ;
      RECT  9492.5 35230.0 9557.5 35415.0 ;
      RECT  9132.5 35347.5 9197.5 35197.5 ;
      RECT  9132.5 36232.5 9197.5 36607.5 ;
      RECT  9322.5 35347.5 9387.5 36232.5 ;
      RECT  9132.5 36232.5 9197.5 36367.5 ;
      RECT  9322.5 36232.5 9387.5 36367.5 ;
      RECT  9322.5 36232.5 9387.5 36367.5 ;
      RECT  9132.5 36232.5 9197.5 36367.5 ;
      RECT  9132.5 35347.5 9197.5 35482.5 ;
      RECT  9322.5 35347.5 9387.5 35482.5 ;
      RECT  9322.5 35347.5 9387.5 35482.5 ;
      RECT  9132.5 35347.5 9197.5 35482.5 ;
      RECT  9492.5 36322.5 9557.5 36457.5 ;
      RECT  9492.5 35347.5 9557.5 35482.5 ;
      RECT  9190.0 35790.0 9255.0 35925.0 ;
      RECT  9190.0 35790.0 9255.0 35925.0 ;
      RECT  9355.0 35825.0 9420.0 35890.0 ;
      RECT  9065.0 36542.5 9625.0 36607.5 ;
      RECT  9065.0 35197.5 9625.0 35262.5 ;
      RECT  9692.5 35392.5 9757.5 35197.5 ;
      RECT  9692.5 36232.5 9757.5 36607.5 ;
      RECT  10072.5 36232.5 10137.5 36607.5 ;
      RECT  10242.5 36390.0 10307.5 36575.0 ;
      RECT  10242.5 35230.0 10307.5 35415.0 ;
      RECT  9692.5 36232.5 9757.5 36367.5 ;
      RECT  9882.5 36232.5 9947.5 36367.5 ;
      RECT  9882.5 36232.5 9947.5 36367.5 ;
      RECT  9692.5 36232.5 9757.5 36367.5 ;
      RECT  9882.5 36232.5 9947.5 36367.5 ;
      RECT  10072.5 36232.5 10137.5 36367.5 ;
      RECT  10072.5 36232.5 10137.5 36367.5 ;
      RECT  9882.5 36232.5 9947.5 36367.5 ;
      RECT  9692.5 35392.5 9757.5 35527.5 ;
      RECT  9882.5 35392.5 9947.5 35527.5 ;
      RECT  9882.5 35392.5 9947.5 35527.5 ;
      RECT  9692.5 35392.5 9757.5 35527.5 ;
      RECT  9882.5 35392.5 9947.5 35527.5 ;
      RECT  10072.5 35392.5 10137.5 35527.5 ;
      RECT  10072.5 35392.5 10137.5 35527.5 ;
      RECT  9882.5 35392.5 9947.5 35527.5 ;
      RECT  10242.5 36322.5 10307.5 36457.5 ;
      RECT  10242.5 35347.5 10307.5 35482.5 ;
      RECT  10077.5 35622.5 9942.5 35687.5 ;
      RECT  9820.0 35837.5 9685.0 35902.5 ;
      RECT  9882.5 36232.5 9947.5 36367.5 ;
      RECT  10072.5 35392.5 10137.5 35527.5 ;
      RECT  10172.5 35837.5 10037.5 35902.5 ;
      RECT  9685.0 35837.5 9820.0 35902.5 ;
      RECT  9942.5 35622.5 10077.5 35687.5 ;
      RECT  10037.5 35837.5 10172.5 35902.5 ;
      RECT  9625.0 36542.5 10545.0 36607.5 ;
      RECT  9625.0 35197.5 10545.0 35262.5 ;
      RECT  10972.5 36390.0 11037.5 36575.0 ;
      RECT  10972.5 35230.0 11037.5 35415.0 ;
      RECT  10612.5 35347.5 10677.5 35197.5 ;
      RECT  10612.5 36232.5 10677.5 36607.5 ;
      RECT  10802.5 35347.5 10867.5 36232.5 ;
      RECT  10612.5 36232.5 10677.5 36367.5 ;
      RECT  10802.5 36232.5 10867.5 36367.5 ;
      RECT  10802.5 36232.5 10867.5 36367.5 ;
      RECT  10612.5 36232.5 10677.5 36367.5 ;
      RECT  10612.5 35347.5 10677.5 35482.5 ;
      RECT  10802.5 35347.5 10867.5 35482.5 ;
      RECT  10802.5 35347.5 10867.5 35482.5 ;
      RECT  10612.5 35347.5 10677.5 35482.5 ;
      RECT  10972.5 36322.5 11037.5 36457.5 ;
      RECT  10972.5 35347.5 11037.5 35482.5 ;
      RECT  10670.0 35790.0 10735.0 35925.0 ;
      RECT  10670.0 35790.0 10735.0 35925.0 ;
      RECT  10835.0 35825.0 10900.0 35890.0 ;
      RECT  10545.0 36542.5 11105.0 36607.5 ;
      RECT  10545.0 35197.5 11105.0 35262.5 ;
      RECT  8807.5 35790.0 8872.5 35925.0 ;
      RECT  8947.5 35517.5 9012.5 35652.5 ;
      RECT  9942.5 35622.5 9807.5 35687.5 ;
      RECT  9492.5 36760.0 9557.5 36575.0 ;
      RECT  9492.5 37920.0 9557.5 37735.0 ;
      RECT  9132.5 37802.5 9197.5 37952.5 ;
      RECT  9132.5 36917.5 9197.5 36542.5 ;
      RECT  9322.5 37802.5 9387.5 36917.5 ;
      RECT  9132.5 36917.5 9197.5 36782.5 ;
      RECT  9322.5 36917.5 9387.5 36782.5 ;
      RECT  9322.5 36917.5 9387.5 36782.5 ;
      RECT  9132.5 36917.5 9197.5 36782.5 ;
      RECT  9132.5 37802.5 9197.5 37667.5 ;
      RECT  9322.5 37802.5 9387.5 37667.5 ;
      RECT  9322.5 37802.5 9387.5 37667.5 ;
      RECT  9132.5 37802.5 9197.5 37667.5 ;
      RECT  9492.5 36827.5 9557.5 36692.5 ;
      RECT  9492.5 37802.5 9557.5 37667.5 ;
      RECT  9190.0 37360.0 9255.0 37225.0 ;
      RECT  9190.0 37360.0 9255.0 37225.0 ;
      RECT  9355.0 37325.0 9420.0 37260.0 ;
      RECT  9065.0 36607.5 9625.0 36542.5 ;
      RECT  9065.0 37952.5 9625.0 37887.5 ;
      RECT  9692.5 37757.5 9757.5 37952.5 ;
      RECT  9692.5 36917.5 9757.5 36542.5 ;
      RECT  10072.5 36917.5 10137.5 36542.5 ;
      RECT  10242.5 36760.0 10307.5 36575.0 ;
      RECT  10242.5 37920.0 10307.5 37735.0 ;
      RECT  9692.5 36917.5 9757.5 36782.5 ;
      RECT  9882.5 36917.5 9947.5 36782.5 ;
      RECT  9882.5 36917.5 9947.5 36782.5 ;
      RECT  9692.5 36917.5 9757.5 36782.5 ;
      RECT  9882.5 36917.5 9947.5 36782.5 ;
      RECT  10072.5 36917.5 10137.5 36782.5 ;
      RECT  10072.5 36917.5 10137.5 36782.5 ;
      RECT  9882.5 36917.5 9947.5 36782.5 ;
      RECT  9692.5 37757.5 9757.5 37622.5 ;
      RECT  9882.5 37757.5 9947.5 37622.5 ;
      RECT  9882.5 37757.5 9947.5 37622.5 ;
      RECT  9692.5 37757.5 9757.5 37622.5 ;
      RECT  9882.5 37757.5 9947.5 37622.5 ;
      RECT  10072.5 37757.5 10137.5 37622.5 ;
      RECT  10072.5 37757.5 10137.5 37622.5 ;
      RECT  9882.5 37757.5 9947.5 37622.5 ;
      RECT  10242.5 36827.5 10307.5 36692.5 ;
      RECT  10242.5 37802.5 10307.5 37667.5 ;
      RECT  10077.5 37527.5 9942.5 37462.5 ;
      RECT  9820.0 37312.5 9685.0 37247.5 ;
      RECT  9882.5 36917.5 9947.5 36782.5 ;
      RECT  10072.5 37757.5 10137.5 37622.5 ;
      RECT  10172.5 37312.5 10037.5 37247.5 ;
      RECT  9685.0 37312.5 9820.0 37247.5 ;
      RECT  9942.5 37527.5 10077.5 37462.5 ;
      RECT  10037.5 37312.5 10172.5 37247.5 ;
      RECT  9625.0 36607.5 10545.0 36542.5 ;
      RECT  9625.0 37952.5 10545.0 37887.5 ;
      RECT  10972.5 36760.0 11037.5 36575.0 ;
      RECT  10972.5 37920.0 11037.5 37735.0 ;
      RECT  10612.5 37802.5 10677.5 37952.5 ;
      RECT  10612.5 36917.5 10677.5 36542.5 ;
      RECT  10802.5 37802.5 10867.5 36917.5 ;
      RECT  10612.5 36917.5 10677.5 36782.5 ;
      RECT  10802.5 36917.5 10867.5 36782.5 ;
      RECT  10802.5 36917.5 10867.5 36782.5 ;
      RECT  10612.5 36917.5 10677.5 36782.5 ;
      RECT  10612.5 37802.5 10677.5 37667.5 ;
      RECT  10802.5 37802.5 10867.5 37667.5 ;
      RECT  10802.5 37802.5 10867.5 37667.5 ;
      RECT  10612.5 37802.5 10677.5 37667.5 ;
      RECT  10972.5 36827.5 11037.5 36692.5 ;
      RECT  10972.5 37802.5 11037.5 37667.5 ;
      RECT  10670.0 37360.0 10735.0 37225.0 ;
      RECT  10670.0 37360.0 10735.0 37225.0 ;
      RECT  10835.0 37325.0 10900.0 37260.0 ;
      RECT  10545.0 36607.5 11105.0 36542.5 ;
      RECT  10545.0 37952.5 11105.0 37887.5 ;
      RECT  8807.5 37225.0 8872.5 37360.0 ;
      RECT  8947.5 37497.5 9012.5 37632.5 ;
      RECT  9942.5 37462.5 9807.5 37527.5 ;
      RECT  9492.5 39080.0 9557.5 39265.0 ;
      RECT  9492.5 37920.0 9557.5 38105.0 ;
      RECT  9132.5 38037.5 9197.5 37887.5 ;
      RECT  9132.5 38922.5 9197.5 39297.5 ;
      RECT  9322.5 38037.5 9387.5 38922.5 ;
      RECT  9132.5 38922.5 9197.5 39057.5 ;
      RECT  9322.5 38922.5 9387.5 39057.5 ;
      RECT  9322.5 38922.5 9387.5 39057.5 ;
      RECT  9132.5 38922.5 9197.5 39057.5 ;
      RECT  9132.5 38037.5 9197.5 38172.5 ;
      RECT  9322.5 38037.5 9387.5 38172.5 ;
      RECT  9322.5 38037.5 9387.5 38172.5 ;
      RECT  9132.5 38037.5 9197.5 38172.5 ;
      RECT  9492.5 39012.5 9557.5 39147.5 ;
      RECT  9492.5 38037.5 9557.5 38172.5 ;
      RECT  9190.0 38480.0 9255.0 38615.0 ;
      RECT  9190.0 38480.0 9255.0 38615.0 ;
      RECT  9355.0 38515.0 9420.0 38580.0 ;
      RECT  9065.0 39232.5 9625.0 39297.5 ;
      RECT  9065.0 37887.5 9625.0 37952.5 ;
      RECT  9692.5 38082.5 9757.5 37887.5 ;
      RECT  9692.5 38922.5 9757.5 39297.5 ;
      RECT  10072.5 38922.5 10137.5 39297.5 ;
      RECT  10242.5 39080.0 10307.5 39265.0 ;
      RECT  10242.5 37920.0 10307.5 38105.0 ;
      RECT  9692.5 38922.5 9757.5 39057.5 ;
      RECT  9882.5 38922.5 9947.5 39057.5 ;
      RECT  9882.5 38922.5 9947.5 39057.5 ;
      RECT  9692.5 38922.5 9757.5 39057.5 ;
      RECT  9882.5 38922.5 9947.5 39057.5 ;
      RECT  10072.5 38922.5 10137.5 39057.5 ;
      RECT  10072.5 38922.5 10137.5 39057.5 ;
      RECT  9882.5 38922.5 9947.5 39057.5 ;
      RECT  9692.5 38082.5 9757.5 38217.5 ;
      RECT  9882.5 38082.5 9947.5 38217.5 ;
      RECT  9882.5 38082.5 9947.5 38217.5 ;
      RECT  9692.5 38082.5 9757.5 38217.5 ;
      RECT  9882.5 38082.5 9947.5 38217.5 ;
      RECT  10072.5 38082.5 10137.5 38217.5 ;
      RECT  10072.5 38082.5 10137.5 38217.5 ;
      RECT  9882.5 38082.5 9947.5 38217.5 ;
      RECT  10242.5 39012.5 10307.5 39147.5 ;
      RECT  10242.5 38037.5 10307.5 38172.5 ;
      RECT  10077.5 38312.5 9942.5 38377.5 ;
      RECT  9820.0 38527.5 9685.0 38592.5 ;
      RECT  9882.5 38922.5 9947.5 39057.5 ;
      RECT  10072.5 38082.5 10137.5 38217.5 ;
      RECT  10172.5 38527.5 10037.5 38592.5 ;
      RECT  9685.0 38527.5 9820.0 38592.5 ;
      RECT  9942.5 38312.5 10077.5 38377.5 ;
      RECT  10037.5 38527.5 10172.5 38592.5 ;
      RECT  9625.0 39232.5 10545.0 39297.5 ;
      RECT  9625.0 37887.5 10545.0 37952.5 ;
      RECT  10972.5 39080.0 11037.5 39265.0 ;
      RECT  10972.5 37920.0 11037.5 38105.0 ;
      RECT  10612.5 38037.5 10677.5 37887.5 ;
      RECT  10612.5 38922.5 10677.5 39297.5 ;
      RECT  10802.5 38037.5 10867.5 38922.5 ;
      RECT  10612.5 38922.5 10677.5 39057.5 ;
      RECT  10802.5 38922.5 10867.5 39057.5 ;
      RECT  10802.5 38922.5 10867.5 39057.5 ;
      RECT  10612.5 38922.5 10677.5 39057.5 ;
      RECT  10612.5 38037.5 10677.5 38172.5 ;
      RECT  10802.5 38037.5 10867.5 38172.5 ;
      RECT  10802.5 38037.5 10867.5 38172.5 ;
      RECT  10612.5 38037.5 10677.5 38172.5 ;
      RECT  10972.5 39012.5 11037.5 39147.5 ;
      RECT  10972.5 38037.5 11037.5 38172.5 ;
      RECT  10670.0 38480.0 10735.0 38615.0 ;
      RECT  10670.0 38480.0 10735.0 38615.0 ;
      RECT  10835.0 38515.0 10900.0 38580.0 ;
      RECT  10545.0 39232.5 11105.0 39297.5 ;
      RECT  10545.0 37887.5 11105.0 37952.5 ;
      RECT  8807.5 38480.0 8872.5 38615.0 ;
      RECT  8947.5 38207.5 9012.5 38342.5 ;
      RECT  9942.5 38312.5 9807.5 38377.5 ;
      RECT  9492.5 39450.0 9557.5 39265.0 ;
      RECT  9492.5 40610.0 9557.5 40425.0 ;
      RECT  9132.5 40492.5 9197.5 40642.5 ;
      RECT  9132.5 39607.5 9197.5 39232.5 ;
      RECT  9322.5 40492.5 9387.5 39607.5 ;
      RECT  9132.5 39607.5 9197.5 39472.5 ;
      RECT  9322.5 39607.5 9387.5 39472.5 ;
      RECT  9322.5 39607.5 9387.5 39472.5 ;
      RECT  9132.5 39607.5 9197.5 39472.5 ;
      RECT  9132.5 40492.5 9197.5 40357.5 ;
      RECT  9322.5 40492.5 9387.5 40357.5 ;
      RECT  9322.5 40492.5 9387.5 40357.5 ;
      RECT  9132.5 40492.5 9197.5 40357.5 ;
      RECT  9492.5 39517.5 9557.5 39382.5 ;
      RECT  9492.5 40492.5 9557.5 40357.5 ;
      RECT  9190.0 40050.0 9255.0 39915.0 ;
      RECT  9190.0 40050.0 9255.0 39915.0 ;
      RECT  9355.0 40015.0 9420.0 39950.0 ;
      RECT  9065.0 39297.5 9625.0 39232.5 ;
      RECT  9065.0 40642.5 9625.0 40577.5 ;
      RECT  9692.5 40447.5 9757.5 40642.5 ;
      RECT  9692.5 39607.5 9757.5 39232.5 ;
      RECT  10072.5 39607.5 10137.5 39232.5 ;
      RECT  10242.5 39450.0 10307.5 39265.0 ;
      RECT  10242.5 40610.0 10307.5 40425.0 ;
      RECT  9692.5 39607.5 9757.5 39472.5 ;
      RECT  9882.5 39607.5 9947.5 39472.5 ;
      RECT  9882.5 39607.5 9947.5 39472.5 ;
      RECT  9692.5 39607.5 9757.5 39472.5 ;
      RECT  9882.5 39607.5 9947.5 39472.5 ;
      RECT  10072.5 39607.5 10137.5 39472.5 ;
      RECT  10072.5 39607.5 10137.5 39472.5 ;
      RECT  9882.5 39607.5 9947.5 39472.5 ;
      RECT  9692.5 40447.5 9757.5 40312.5 ;
      RECT  9882.5 40447.5 9947.5 40312.5 ;
      RECT  9882.5 40447.5 9947.5 40312.5 ;
      RECT  9692.5 40447.5 9757.5 40312.5 ;
      RECT  9882.5 40447.5 9947.5 40312.5 ;
      RECT  10072.5 40447.5 10137.5 40312.5 ;
      RECT  10072.5 40447.5 10137.5 40312.5 ;
      RECT  9882.5 40447.5 9947.5 40312.5 ;
      RECT  10242.5 39517.5 10307.5 39382.5 ;
      RECT  10242.5 40492.5 10307.5 40357.5 ;
      RECT  10077.5 40217.5 9942.5 40152.5 ;
      RECT  9820.0 40002.5 9685.0 39937.5 ;
      RECT  9882.5 39607.5 9947.5 39472.5 ;
      RECT  10072.5 40447.5 10137.5 40312.5 ;
      RECT  10172.5 40002.5 10037.5 39937.5 ;
      RECT  9685.0 40002.5 9820.0 39937.5 ;
      RECT  9942.5 40217.5 10077.5 40152.5 ;
      RECT  10037.5 40002.5 10172.5 39937.5 ;
      RECT  9625.0 39297.5 10545.0 39232.5 ;
      RECT  9625.0 40642.5 10545.0 40577.5 ;
      RECT  10972.5 39450.0 11037.5 39265.0 ;
      RECT  10972.5 40610.0 11037.5 40425.0 ;
      RECT  10612.5 40492.5 10677.5 40642.5 ;
      RECT  10612.5 39607.5 10677.5 39232.5 ;
      RECT  10802.5 40492.5 10867.5 39607.5 ;
      RECT  10612.5 39607.5 10677.5 39472.5 ;
      RECT  10802.5 39607.5 10867.5 39472.5 ;
      RECT  10802.5 39607.5 10867.5 39472.5 ;
      RECT  10612.5 39607.5 10677.5 39472.5 ;
      RECT  10612.5 40492.5 10677.5 40357.5 ;
      RECT  10802.5 40492.5 10867.5 40357.5 ;
      RECT  10802.5 40492.5 10867.5 40357.5 ;
      RECT  10612.5 40492.5 10677.5 40357.5 ;
      RECT  10972.5 39517.5 11037.5 39382.5 ;
      RECT  10972.5 40492.5 11037.5 40357.5 ;
      RECT  10670.0 40050.0 10735.0 39915.0 ;
      RECT  10670.0 40050.0 10735.0 39915.0 ;
      RECT  10835.0 40015.0 10900.0 39950.0 ;
      RECT  10545.0 39297.5 11105.0 39232.5 ;
      RECT  10545.0 40642.5 11105.0 40577.5 ;
      RECT  8807.5 39915.0 8872.5 40050.0 ;
      RECT  8947.5 40187.5 9012.5 40322.5 ;
      RECT  9942.5 40152.5 9807.5 40217.5 ;
      RECT  8610.0 19412.5 8980.0 19477.5 ;
      RECT  8610.0 21392.5 8980.0 21457.5 ;
      RECT  8610.0 22102.5 8980.0 22167.5 ;
      RECT  8610.0 24082.5 8980.0 24147.5 ;
      RECT  8610.0 24792.5 8980.0 24857.5 ;
      RECT  8610.0 26772.5 8980.0 26837.5 ;
      RECT  8610.0 27482.5 8980.0 27547.5 ;
      RECT  8610.0 29462.5 8980.0 29527.5 ;
      RECT  8610.0 30172.5 8980.0 30237.5 ;
      RECT  8610.0 32152.5 8980.0 32217.5 ;
      RECT  8610.0 32862.5 8980.0 32927.5 ;
      RECT  8610.0 34842.5 8980.0 34907.5 ;
      RECT  8610.0 35552.5 8980.0 35617.5 ;
      RECT  8610.0 37532.5 8980.0 37597.5 ;
      RECT  8610.0 38242.5 8980.0 38307.5 ;
      RECT  8610.0 40222.5 8980.0 40287.5 ;
      RECT  10835.0 19685.0 10900.0 19750.0 ;
      RECT  10835.0 21120.0 10900.0 21185.0 ;
      RECT  10835.0 22375.0 10900.0 22440.0 ;
      RECT  10835.0 23810.0 10900.0 23875.0 ;
      RECT  10835.0 25065.0 10900.0 25130.0 ;
      RECT  10835.0 26500.0 10900.0 26565.0 ;
      RECT  10835.0 27755.0 10900.0 27820.0 ;
      RECT  10835.0 29190.0 10900.0 29255.0 ;
      RECT  10835.0 30445.0 10900.0 30510.0 ;
      RECT  10835.0 31880.0 10900.0 31945.0 ;
      RECT  10835.0 33135.0 10900.0 33200.0 ;
      RECT  10835.0 34570.0 10900.0 34635.0 ;
      RECT  10835.0 35825.0 10900.0 35890.0 ;
      RECT  10835.0 37260.0 10900.0 37325.0 ;
      RECT  10835.0 38515.0 10900.0 38580.0 ;
      RECT  10835.0 39950.0 10900.0 40015.0 ;
      RECT  8610.0 20402.5 9065.0 20467.5 ;
      RECT  8610.0 23092.5 9065.0 23157.5 ;
      RECT  8610.0 25782.5 9065.0 25847.5 ;
      RECT  8610.0 28472.5 9065.0 28537.5 ;
      RECT  8610.0 31162.5 9065.0 31227.5 ;
      RECT  8610.0 33852.5 9065.0 33917.5 ;
      RECT  8610.0 36542.5 9065.0 36607.5 ;
      RECT  8610.0 39232.5 9065.0 39297.5 ;
      RECT  8610.0 19057.5 9065.0 19122.5 ;
      RECT  8610.0 21747.5 9065.0 21812.5 ;
      RECT  8610.0 24437.5 9065.0 24502.5 ;
      RECT  8610.0 27127.5 9065.0 27192.5 ;
      RECT  8610.0 29817.5 9065.0 29882.5 ;
      RECT  8610.0 32507.5 9065.0 32572.5 ;
      RECT  8610.0 35197.5 9065.0 35262.5 ;
      RECT  8610.0 37887.5 9065.0 37952.5 ;
      RECT  8610.0 40577.5 9065.0 40642.5 ;
      RECT  4655.0 7920.0 11095.0 7215.0 ;
      RECT  4655.0 6510.0 11095.0 7215.0 ;
      RECT  4655.0 6510.0 11095.0 5805.0 ;
      RECT  4655.0 5100.0 11095.0 5805.0 ;
      RECT  4860.0 7920.0 4925.0 5100.0 ;
      RECT  7865.0 7920.0 7930.0 5100.0 ;
      RECT  10825.0 7920.0 10890.0 5100.0 ;
      RECT  5875.0 7920.0 5940.0 5100.0 ;
      RECT  8835.0 7920.0 8900.0 5100.0 ;
      RECT  5020.0 7920.0 5085.0 5100.0 ;
      RECT  12427.5 19122.5 12562.5 19057.5 ;
      RECT  12427.5 21812.5 12562.5 21747.5 ;
      RECT  12427.5 24502.5 12562.5 24437.5 ;
      RECT  12427.5 27192.5 12562.5 27127.5 ;
      RECT  12427.5 29882.5 12562.5 29817.5 ;
      RECT  12427.5 32572.5 12562.5 32507.5 ;
      RECT  12427.5 35262.5 12562.5 35197.5 ;
      RECT  12427.5 37952.5 12562.5 37887.5 ;
      RECT  12427.5 40642.5 12562.5 40577.5 ;
      RECT  11095.0 8502.5 10960.0 8567.5 ;
      RECT  11505.0 8502.5 11370.0 8567.5 ;
      RECT  10820.0 9847.5 10685.0 9912.5 ;
      RECT  11710.0 9847.5 11575.0 9912.5 ;
      RECT  11095.0 13882.5 10960.0 13947.5 ;
      RECT  11915.0 13882.5 11780.0 13947.5 ;
      RECT  10820.0 15227.5 10685.0 15292.5 ;
      RECT  12120.0 15227.5 11985.0 15292.5 ;
      RECT  11300.0 8297.5 11165.0 8362.5 ;
      RECT  11300.0 10987.5 11165.0 11052.5 ;
      RECT  11300.0 13677.5 11165.0 13742.5 ;
      RECT  11300.0 16367.5 11165.0 16432.5 ;
      RECT  11162.5 7535.0 11027.5 7600.0 ;
      RECT  11505.0 7535.0 11370.0 7600.0 ;
      RECT  11162.5 6830.0 11027.5 6895.0 ;
      RECT  11710.0 6830.0 11575.0 6895.0 ;
      RECT  11162.5 6125.0 11027.5 6190.0 ;
      RECT  11915.0 6125.0 11780.0 6190.0 ;
      RECT  11162.5 5420.0 11027.5 5485.0 ;
      RECT  12120.0 5420.0 11985.0 5485.0 ;
      RECT  11230.0 7887.5 11095.0 7952.5 ;
      RECT  12562.5 7887.5 12427.5 7952.5 ;
      RECT  11230.0 7182.5 11095.0 7247.5 ;
      RECT  12562.5 7182.5 12427.5 7247.5 ;
      RECT  11230.0 6477.5 11095.0 6542.5 ;
      RECT  12562.5 6477.5 12427.5 6542.5 ;
      RECT  11230.0 5772.5 11095.0 5837.5 ;
      RECT  12562.5 5772.5 12427.5 5837.5 ;
      RECT  11230.0 5067.5 11095.0 5132.5 ;
      RECT  12562.5 5067.5 12427.5 5132.5 ;
      RECT  13700.0 3795.0 13565.0 3860.0 ;
      RECT  13290.0 1610.0 13155.0 1675.0 ;
      RECT  13495.0 3157.5 13360.0 3222.5 ;
      RECT  13700.0 41587.5 13565.0 41652.5 ;
      RECT  13905.0 10297.5 13770.0 10362.5 ;
      RECT  14110.0 14322.5 13975.0 14387.5 ;
      RECT  13085.0 8092.5 12950.0 8157.5 ;
      RECT  8907.5 40782.5 8772.5 40847.5 ;
      RECT  13085.0 40782.5 12950.0 40847.5 ;
      RECT  12777.5 3027.5 12642.5 3092.5 ;
      RECT  12777.5 14452.5 12642.5 14517.5 ;
      RECT  12777.5 3955.0 12642.5 4020.0 ;
      RECT  12777.5 11230.0 12642.5 11295.0 ;
      RECT  16125.0 0.0 16475.0 42337.5 ;
      RECT  4175.0 0.0 4525.0 42337.5 ;
      RECT  3455.0 19520.0 3390.0 19585.0 ;
      RECT  3422.5 19520.0 3407.5 19585.0 ;
      RECT  3455.0 19552.5 3390.0 20137.5 ;
      RECT  3455.0 20682.5 3390.0 21077.5 ;
      RECT  3455.0 22002.5 3390.0 22587.5 ;
      RECT  2657.5 22440.0 2280.0 22505.0 ;
      RECT  2657.5 25400.0 2280.0 25465.0 ;
      RECT  2657.5 20450.0 2280.0 20515.0 ;
      RECT  2657.5 23410.0 2280.0 23475.0 ;
      RECT  3440.0 19520.0 3375.0 19585.0 ;
      RECT  3455.0 20650.0 3390.0 20715.0 ;
      RECT  2005.0 31335.0 1940.0 32100.0 ;
      RECT  3455.0 24685.0 3390.0 26115.0 ;
      RECT  2485.0 19435.0 2280.0 19500.0 ;
      RECT  1962.5 26115.0 1897.5 28052.5 ;
      RECT  1747.5 26525.0 1682.5 28310.0 ;
      RECT  3380.0 27550.0 3315.0 28120.0 ;
      RECT  3520.0 27345.0 3455.0 28310.0 ;
      RECT  3660.0 26730.0 3595.0 28500.0 ;
      RECT  3380.0 29060.0 3315.0 29125.0 ;
      RECT  3380.0 28595.0 3315.0 29092.5 ;
      RECT  3407.5 29060.0 3347.5 29125.0 ;
      RECT  3475.0 29225.0 3410.0 29290.0 ;
      RECT  3442.5 29225.0 3407.5 29290.0 ;
      RECT  3475.0 29257.5 3410.0 32797.5 ;
      RECT  690.0 27550.0 625.0 28680.0 ;
      RECT  830.0 26730.0 765.0 28870.0 ;
      RECT  970.0 26935.0 905.0 29060.0 ;
      RECT  690.0 29620.0 625.0 29685.0 ;
      RECT  690.0 29155.0 625.0 29652.5 ;
      RECT  717.5 29620.0 657.5 29685.0 ;
      RECT  750.0 29817.5 685.0 30212.5 ;
      RECT  750.0 30377.5 685.0 30772.5 ;
      RECT  2005.0 31302.5 1940.0 31367.5 ;
      RECT  1972.5 31302.5 1940.0 31367.5 ;
      RECT  2005.0 31210.0 1940.0 31335.0 ;
      RECT  2005.0 30617.5 1940.0 31012.5 ;
      RECT  1962.5 28475.0 1897.5 28845.0 ;
      RECT  2017.5 29550.0 1952.5 29990.0 ;
      RECT  750.0 30937.5 685.0 31175.0 ;
      RECT  2005.0 30215.0 1940.0 30452.5 ;
      RECT  4067.5 19230.0 4002.5 31335.0 ;
      RECT  4067.5 26320.0 4002.5 27925.0 ;
      RECT  2722.5 19230.0 2657.5 31335.0 ;
      RECT  2722.5 27140.0 2657.5 27925.0 ;
      RECT  1377.5 27925.0 1312.5 31335.0 ;
      RECT  1377.5 26320.0 1312.5 27925.0 ;
      RECT  32.5 27925.0 -32.5 31335.0 ;
      RECT  32.5 27140.0 -32.5 27925.0 ;
      RECT  32.5 31302.5 -32.5 31367.5 ;
      RECT  32.5 31130.0 -32.5 31335.0 ;
      RECT  8.881784197e-13 31302.5 -45.0 31367.5 ;
      RECT  165.0 19230.0 870.0 25670.0 ;
      RECT  1575.0 19230.0 870.0 25670.0 ;
      RECT  1575.0 19230.0 2280.0 25670.0 ;
      RECT  165.0 19435.0 2280.0 19500.0 ;
      RECT  165.0 22440.0 2280.0 22505.0 ;
      RECT  165.0 25400.0 2280.0 25465.0 ;
      RECT  165.0 20450.0 2280.0 20515.0 ;
      RECT  165.0 23410.0 2280.0 23475.0 ;
      RECT  165.0 19595.0 2280.0 19660.0 ;
      RECT  2875.0 19847.5 2690.0 19912.5 ;
      RECT  4035.0 19847.5 3850.0 19912.5 ;
      RECT  2832.5 19297.5 2657.5 19742.5 ;
      RECT  3917.5 19487.5 3032.5 19552.5 ;
      RECT  2965.0 19297.5 2800.0 19362.5 ;
      RECT  2965.0 19677.5 2800.0 19742.5 ;
      RECT  3032.5 19297.5 2897.5 19362.5 ;
      RECT  3032.5 19677.5 2897.5 19742.5 ;
      RECT  3032.5 19487.5 2897.5 19552.5 ;
      RECT  3032.5 19487.5 2897.5 19552.5 ;
      RECT  2832.5 19297.5 2767.5 19742.5 ;
      RECT  4015.0 19297.5 3850.0 19362.5 ;
      RECT  4015.0 19677.5 3850.0 19742.5 ;
      RECT  3917.5 19297.5 3782.5 19362.5 ;
      RECT  3917.5 19677.5 3782.5 19742.5 ;
      RECT  3917.5 19487.5 3782.5 19552.5 ;
      RECT  3917.5 19487.5 3782.5 19552.5 ;
      RECT  4047.5 19297.5 3982.5 19742.5 ;
      RECT  2942.5 19847.5 2807.5 19912.5 ;
      RECT  3917.5 19847.5 3782.5 19912.5 ;
      RECT  3475.0 19355.0 3340.0 19420.0 ;
      RECT  3475.0 19355.0 3340.0 19420.0 ;
      RECT  3440.0 19520.0 3375.0 19585.0 ;
      RECT  2722.5 19230.0 2657.5 19980.0 ;
      RECT  4067.5 19230.0 4002.5 19980.0 ;
      RECT  2875.0 20787.5 2690.0 20852.5 ;
      RECT  4035.0 20787.5 3850.0 20852.5 ;
      RECT  2877.5 20047.5 2657.5 20492.5 ;
      RECT  3702.5 20617.5 3207.5 20682.5 ;
      RECT  3010.0 20047.5 2845.0 20112.5 ;
      RECT  3010.0 20427.5 2845.0 20492.5 ;
      RECT  3175.0 20237.5 3010.0 20302.5 ;
      RECT  3175.0 20617.5 3010.0 20682.5 ;
      RECT  3077.5 20047.5 2942.5 20112.5 ;
      RECT  3077.5 20427.5 2942.5 20492.5 ;
      RECT  3077.5 20237.5 2942.5 20302.5 ;
      RECT  3077.5 20617.5 2942.5 20682.5 ;
      RECT  3207.5 20237.5 3142.5 20682.5 ;
      RECT  2877.5 20047.5 2812.5 20492.5 ;
      RECT  4000.0 20047.5 3835.0 20112.5 ;
      RECT  4000.0 20427.5 3835.0 20492.5 ;
      RECT  3835.0 20237.5 3670.0 20302.5 ;
      RECT  3835.0 20617.5 3670.0 20682.5 ;
      RECT  3902.5 20047.5 3767.5 20112.5 ;
      RECT  3902.5 20427.5 3767.5 20492.5 ;
      RECT  3902.5 20237.5 3767.5 20302.5 ;
      RECT  3902.5 20617.5 3767.5 20682.5 ;
      RECT  3702.5 20237.5 3637.5 20682.5 ;
      RECT  4032.5 20047.5 3967.5 20492.5 ;
      RECT  2942.5 20787.5 2807.5 20852.5 ;
      RECT  3917.5 20787.5 3782.5 20852.5 ;
      RECT  3490.0 20105.0 3355.0 20170.0 ;
      RECT  3490.0 20105.0 3355.0 20170.0 ;
      RECT  3455.0 20650.0 3390.0 20715.0 ;
      RECT  2722.5 19980.0 2657.5 20920.0 ;
      RECT  4067.5 19980.0 4002.5 20920.0 ;
      RECT  2875.0 22297.5 2690.0 22362.5 ;
      RECT  4035.0 22297.5 3850.0 22362.5 ;
      RECT  2877.5 20987.5 2657.5 22192.5 ;
      RECT  3702.5 21937.5 3207.5 22002.5 ;
      RECT  3010.0 20987.5 2845.0 21052.5 ;
      RECT  3010.0 21367.5 2845.0 21432.5 ;
      RECT  3010.0 21747.5 2845.0 21812.5 ;
      RECT  3010.0 22127.5 2845.0 22192.5 ;
      RECT  3175.0 21177.5 3010.0 21242.5 ;
      RECT  3175.0 21557.5 3010.0 21622.5 ;
      RECT  3175.0 21937.5 3010.0 22002.5 ;
      RECT  3077.5 20987.5 2942.5 21052.5 ;
      RECT  3077.5 21367.5 2942.5 21432.5 ;
      RECT  3077.5 21747.5 2942.5 21812.5 ;
      RECT  3077.5 22127.5 2942.5 22192.5 ;
      RECT  3077.5 21177.5 2942.5 21242.5 ;
      RECT  3077.5 21557.5 2942.5 21622.5 ;
      RECT  3077.5 21937.5 2942.5 22002.5 ;
      RECT  3207.5 21177.5 3142.5 22002.5 ;
      RECT  2877.5 20987.5 2812.5 22192.5 ;
      RECT  4000.0 20987.5 3835.0 21052.5 ;
      RECT  4000.0 21367.5 3835.0 21432.5 ;
      RECT  4000.0 21747.5 3835.0 21812.5 ;
      RECT  4000.0 22127.5 3835.0 22192.5 ;
      RECT  3835.0 21177.5 3670.0 21242.5 ;
      RECT  3835.0 21557.5 3670.0 21622.5 ;
      RECT  3835.0 21937.5 3670.0 22002.5 ;
      RECT  3902.5 20987.5 3767.5 21052.5 ;
      RECT  3902.5 21367.5 3767.5 21432.5 ;
      RECT  3902.5 21747.5 3767.5 21812.5 ;
      RECT  3902.5 22127.5 3767.5 22192.5 ;
      RECT  3902.5 21177.5 3767.5 21242.5 ;
      RECT  3902.5 21557.5 3767.5 21622.5 ;
      RECT  3902.5 21937.5 3767.5 22002.5 ;
      RECT  3702.5 21177.5 3637.5 22002.5 ;
      RECT  4032.5 20987.5 3967.5 22192.5 ;
      RECT  2942.5 22297.5 2807.5 22362.5 ;
      RECT  3917.5 22297.5 3782.5 22362.5 ;
      RECT  3490.0 21045.0 3355.0 21110.0 ;
      RECT  3490.0 21045.0 3355.0 21110.0 ;
      RECT  3455.0 21970.0 3390.0 22035.0 ;
      RECT  2722.5 20920.0 2657.5 22430.0 ;
      RECT  4067.5 20920.0 4002.5 22430.0 ;
      RECT  2875.0 24947.5 2690.0 25012.5 ;
      RECT  4035.0 24947.5 3850.0 25012.5 ;
      RECT  2877.5 22497.5 2657.5 24842.5 ;
      RECT  3702.5 24587.5 3207.5 24652.5 ;
      RECT  3010.0 22497.5 2845.0 22562.5 ;
      RECT  3010.0 22877.5 2845.0 22942.5 ;
      RECT  3010.0 23257.5 2845.0 23322.5 ;
      RECT  3010.0 23637.5 2845.0 23702.5 ;
      RECT  3010.0 24017.5 2845.0 24082.5 ;
      RECT  3010.0 24397.5 2845.0 24462.5 ;
      RECT  3010.0 24777.5 2845.0 24842.5 ;
      RECT  3175.0 22687.5 3010.0 22752.5 ;
      RECT  3175.0 23067.5 3010.0 23132.5 ;
      RECT  3175.0 23447.5 3010.0 23512.5 ;
      RECT  3175.0 23827.5 3010.0 23892.5 ;
      RECT  3175.0 24207.5 3010.0 24272.5 ;
      RECT  3175.0 24587.5 3010.0 24652.5 ;
      RECT  3077.5 22497.5 2942.5 22562.5 ;
      RECT  3077.5 22877.5 2942.5 22942.5 ;
      RECT  3077.5 23257.5 2942.5 23322.5 ;
      RECT  3077.5 23637.5 2942.5 23702.5 ;
      RECT  3077.5 24017.5 2942.5 24082.5 ;
      RECT  3077.5 24397.5 2942.5 24462.5 ;
      RECT  3077.5 24777.5 2942.5 24842.5 ;
      RECT  3077.5 22687.5 2942.5 22752.5 ;
      RECT  3077.5 23067.5 2942.5 23132.5 ;
      RECT  3077.5 23447.5 2942.5 23512.5 ;
      RECT  3077.5 23827.5 2942.5 23892.5 ;
      RECT  3077.5 24207.5 2942.5 24272.5 ;
      RECT  3077.5 24587.5 2942.5 24652.5 ;
      RECT  3207.5 22687.5 3142.5 24652.5 ;
      RECT  2877.5 22497.5 2812.5 24842.5 ;
      RECT  4000.0 22497.5 3835.0 22562.5 ;
      RECT  4000.0 22877.5 3835.0 22942.5 ;
      RECT  4000.0 23257.5 3835.0 23322.5 ;
      RECT  4000.0 23637.5 3835.0 23702.5 ;
      RECT  4000.0 24017.5 3835.0 24082.5 ;
      RECT  4000.0 24397.5 3835.0 24462.5 ;
      RECT  4000.0 24777.5 3835.0 24842.5 ;
      RECT  3835.0 22687.5 3670.0 22752.5 ;
      RECT  3835.0 23067.5 3670.0 23132.5 ;
      RECT  3835.0 23447.5 3670.0 23512.5 ;
      RECT  3835.0 23827.5 3670.0 23892.5 ;
      RECT  3835.0 24207.5 3670.0 24272.5 ;
      RECT  3835.0 24587.5 3670.0 24652.5 ;
      RECT  3902.5 22497.5 3767.5 22562.5 ;
      RECT  3902.5 22877.5 3767.5 22942.5 ;
      RECT  3902.5 23257.5 3767.5 23322.5 ;
      RECT  3902.5 23637.5 3767.5 23702.5 ;
      RECT  3902.5 24017.5 3767.5 24082.5 ;
      RECT  3902.5 24397.5 3767.5 24462.5 ;
      RECT  3902.5 24777.5 3767.5 24842.5 ;
      RECT  3902.5 22687.5 3767.5 22752.5 ;
      RECT  3902.5 23067.5 3767.5 23132.5 ;
      RECT  3902.5 23447.5 3767.5 23512.5 ;
      RECT  3902.5 23827.5 3767.5 23892.5 ;
      RECT  3902.5 24207.5 3767.5 24272.5 ;
      RECT  3902.5 24587.5 3767.5 24652.5 ;
      RECT  3702.5 22687.5 3637.5 24652.5 ;
      RECT  4032.5 22497.5 3967.5 24842.5 ;
      RECT  2942.5 24947.5 2807.5 25012.5 ;
      RECT  3917.5 24947.5 3782.5 25012.5 ;
      RECT  3490.0 22555.0 3355.0 22620.0 ;
      RECT  3490.0 22555.0 3355.0 22620.0 ;
      RECT  3455.0 24620.0 3390.0 24685.0 ;
      RECT  2722.5 22430.0 2657.5 25080.0 ;
      RECT  4067.5 22430.0 4002.5 25080.0 ;
      RECT  3872.5 27992.5 4067.5 28057.5 ;
      RECT  3032.5 27992.5 2657.5 28057.5 ;
      RECT  3032.5 28372.5 2657.5 28437.5 ;
      RECT  2875.0 28732.5 2690.0 28797.5 ;
      RECT  4035.0 28732.5 3850.0 28797.5 ;
      RECT  3032.5 27992.5 2897.5 28057.5 ;
      RECT  3032.5 28182.5 2897.5 28247.5 ;
      RECT  3032.5 28182.5 2897.5 28247.5 ;
      RECT  3032.5 27992.5 2897.5 28057.5 ;
      RECT  3032.5 28182.5 2897.5 28247.5 ;
      RECT  3032.5 28372.5 2897.5 28437.5 ;
      RECT  3032.5 28372.5 2897.5 28437.5 ;
      RECT  3032.5 28182.5 2897.5 28247.5 ;
      RECT  3032.5 28372.5 2897.5 28437.5 ;
      RECT  3032.5 28562.5 2897.5 28627.5 ;
      RECT  3032.5 28562.5 2897.5 28627.5 ;
      RECT  3032.5 28372.5 2897.5 28437.5 ;
      RECT  3872.5 27992.5 3737.5 28057.5 ;
      RECT  3872.5 28182.5 3737.5 28247.5 ;
      RECT  3872.5 28182.5 3737.5 28247.5 ;
      RECT  3872.5 27992.5 3737.5 28057.5 ;
      RECT  3872.5 28182.5 3737.5 28247.5 ;
      RECT  3872.5 28372.5 3737.5 28437.5 ;
      RECT  3872.5 28372.5 3737.5 28437.5 ;
      RECT  3872.5 28182.5 3737.5 28247.5 ;
      RECT  3872.5 28372.5 3737.5 28437.5 ;
      RECT  3872.5 28562.5 3737.5 28627.5 ;
      RECT  3872.5 28562.5 3737.5 28627.5 ;
      RECT  3872.5 28372.5 3737.5 28437.5 ;
      RECT  2942.5 28732.5 2807.5 28797.5 ;
      RECT  3917.5 28732.5 3782.5 28797.5 ;
      RECT  3660.0 28567.5 3595.0 28432.5 ;
      RECT  3520.0 28377.5 3455.0 28242.5 ;
      RECT  3380.0 28187.5 3315.0 28052.5 ;
      RECT  3032.5 28182.5 2897.5 28247.5 ;
      RECT  3032.5 28562.5 2897.5 28627.5 ;
      RECT  3872.5 28562.5 3737.5 28627.5 ;
      RECT  3415.0 28562.5 3280.0 28627.5 ;
      RECT  3380.0 28052.5 3315.0 28187.5 ;
      RECT  3520.0 28242.5 3455.0 28377.5 ;
      RECT  3660.0 28432.5 3595.0 28567.5 ;
      RECT  3415.0 28562.5 3280.0 28627.5 ;
      RECT  2722.5 27925.0 2657.5 28935.0 ;
      RECT  4067.5 27925.0 4002.5 28935.0 ;
      RECT  2875.0 29362.5 2690.0 29427.5 ;
      RECT  4035.0 29362.5 3850.0 29427.5 ;
      RECT  3917.5 29002.5 4067.5 29067.5 ;
      RECT  3032.5 29002.5 2657.5 29067.5 ;
      RECT  3917.5 29192.5 3032.5 29257.5 ;
      RECT  3032.5 29002.5 2897.5 29067.5 ;
      RECT  3032.5 29192.5 2897.5 29257.5 ;
      RECT  3032.5 29192.5 2897.5 29257.5 ;
      RECT  3032.5 29002.5 2897.5 29067.5 ;
      RECT  3917.5 29002.5 3782.5 29067.5 ;
      RECT  3917.5 29192.5 3782.5 29257.5 ;
      RECT  3917.5 29192.5 3782.5 29257.5 ;
      RECT  3917.5 29002.5 3782.5 29067.5 ;
      RECT  2942.5 29362.5 2807.5 29427.5 ;
      RECT  3917.5 29362.5 3782.5 29427.5 ;
      RECT  3475.0 29060.0 3340.0 29125.0 ;
      RECT  3475.0 29060.0 3340.0 29125.0 ;
      RECT  3440.0 29225.0 3375.0 29290.0 ;
      RECT  2722.5 28935.0 2657.5 29495.0 ;
      RECT  4067.5 28935.0 4002.5 29495.0 ;
      RECT  1462.5 27992.5 1312.5 28057.5 ;
      RECT  1462.5 28372.5 1312.5 28437.5 ;
      RECT  2280.0 27992.5 2722.5 28057.5 ;
      RECT  2505.0 28542.5 2690.0 28607.5 ;
      RECT  1345.0 28542.5 1530.0 28607.5 ;
      RECT  2280.0 27992.5 2415.0 28057.5 ;
      RECT  2280.0 28182.5 2415.0 28247.5 ;
      RECT  2280.0 28182.5 2415.0 28247.5 ;
      RECT  2280.0 27992.5 2415.0 28057.5 ;
      RECT  2280.0 28182.5 2415.0 28247.5 ;
      RECT  2280.0 28372.5 2415.0 28437.5 ;
      RECT  2280.0 28372.5 2415.0 28437.5 ;
      RECT  2280.0 28182.5 2415.0 28247.5 ;
      RECT  1462.5 27992.5 1597.5 28057.5 ;
      RECT  1462.5 28182.5 1597.5 28247.5 ;
      RECT  1462.5 28182.5 1597.5 28247.5 ;
      RECT  1462.5 27992.5 1597.5 28057.5 ;
      RECT  1462.5 28182.5 1597.5 28247.5 ;
      RECT  1462.5 28372.5 1597.5 28437.5 ;
      RECT  1462.5 28372.5 1597.5 28437.5 ;
      RECT  1462.5 28182.5 1597.5 28247.5 ;
      RECT  2437.5 28542.5 2572.5 28607.5 ;
      RECT  1462.5 28542.5 1597.5 28607.5 ;
      RECT  1682.5 28377.5 1747.5 28242.5 ;
      RECT  1897.5 28120.0 1962.5 27985.0 ;
      RECT  2280.0 28372.5 2415.0 28437.5 ;
      RECT  1497.5 28282.5 1562.5 28147.5 ;
      RECT  1897.5 28542.5 1962.5 28407.5 ;
      RECT  1897.5 27985.0 1962.5 28120.0 ;
      RECT  1682.5 28242.5 1747.5 28377.5 ;
      RECT  1897.5 28407.5 1962.5 28542.5 ;
      RECT  2657.5 27925.0 2722.5 28845.0 ;
      RECT  1312.5 27925.0 1377.5 28845.0 ;
      RECT  1507.5 29137.5 1312.5 29202.5 ;
      RECT  2347.5 29137.5 2722.5 29202.5 ;
      RECT  2347.5 29517.5 2722.5 29582.5 ;
      RECT  2505.0 29687.5 2690.0 29752.5 ;
      RECT  1345.0 29687.5 1530.0 29752.5 ;
      RECT  2347.5 29137.5 2482.5 29202.5 ;
      RECT  2347.5 29327.5 2482.5 29392.5 ;
      RECT  2347.5 29327.5 2482.5 29392.5 ;
      RECT  2347.5 29137.5 2482.5 29202.5 ;
      RECT  2347.5 29327.5 2482.5 29392.5 ;
      RECT  2347.5 29517.5 2482.5 29582.5 ;
      RECT  2347.5 29517.5 2482.5 29582.5 ;
      RECT  2347.5 29327.5 2482.5 29392.5 ;
      RECT  1507.5 29137.5 1642.5 29202.5 ;
      RECT  1507.5 29327.5 1642.5 29392.5 ;
      RECT  1507.5 29327.5 1642.5 29392.5 ;
      RECT  1507.5 29137.5 1642.5 29202.5 ;
      RECT  1507.5 29327.5 1642.5 29392.5 ;
      RECT  1507.5 29517.5 1642.5 29582.5 ;
      RECT  1507.5 29517.5 1642.5 29582.5 ;
      RECT  1507.5 29327.5 1642.5 29392.5 ;
      RECT  2437.5 29687.5 2572.5 29752.5 ;
      RECT  1462.5 29687.5 1597.5 29752.5 ;
      RECT  1737.5 29522.5 1802.5 29387.5 ;
      RECT  1952.5 29265.0 2017.5 29130.0 ;
      RECT  2347.5 29327.5 2482.5 29392.5 ;
      RECT  1507.5 29517.5 1642.5 29582.5 ;
      RECT  1952.5 29617.5 2017.5 29482.5 ;
      RECT  1952.5 29130.0 2017.5 29265.0 ;
      RECT  1737.5 29387.5 1802.5 29522.5 ;
      RECT  1952.5 29482.5 2017.5 29617.5 ;
      RECT  2657.5 29070.0 2722.5 29990.0 ;
      RECT  1312.5 29070.0 1377.5 29990.0 ;
      RECT  2505.0 30347.5 2690.0 30282.5 ;
      RECT  1345.0 30347.5 1530.0 30282.5 ;
      RECT  1462.5 30707.5 1312.5 30642.5 ;
      RECT  2347.5 30707.5 2722.5 30642.5 ;
      RECT  1462.5 30517.5 2347.5 30452.5 ;
      RECT  2347.5 30707.5 2482.5 30642.5 ;
      RECT  2347.5 30517.5 2482.5 30452.5 ;
      RECT  2347.5 30517.5 2482.5 30452.5 ;
      RECT  2347.5 30707.5 2482.5 30642.5 ;
      RECT  1462.5 30707.5 1597.5 30642.5 ;
      RECT  1462.5 30517.5 1597.5 30452.5 ;
      RECT  1462.5 30517.5 1597.5 30452.5 ;
      RECT  1462.5 30707.5 1597.5 30642.5 ;
      RECT  2437.5 30347.5 2572.5 30282.5 ;
      RECT  1462.5 30347.5 1597.5 30282.5 ;
      RECT  1905.0 30650.0 2040.0 30585.0 ;
      RECT  1905.0 30650.0 2040.0 30585.0 ;
      RECT  1940.0 30485.0 2005.0 30420.0 ;
      RECT  2657.5 30775.0 2722.5 30215.0 ;
      RECT  1312.5 30775.0 1377.5 30215.0 ;
      RECT  2505.0 30907.5 2690.0 30842.5 ;
      RECT  1345.0 30907.5 1530.0 30842.5 ;
      RECT  1462.5 31267.5 1312.5 31202.5 ;
      RECT  2347.5 31267.5 2722.5 31202.5 ;
      RECT  1462.5 31077.5 2347.5 31012.5 ;
      RECT  2347.5 31267.5 2482.5 31202.5 ;
      RECT  2347.5 31077.5 2482.5 31012.5 ;
      RECT  2347.5 31077.5 2482.5 31012.5 ;
      RECT  2347.5 31267.5 2482.5 31202.5 ;
      RECT  1462.5 31267.5 1597.5 31202.5 ;
      RECT  1462.5 31077.5 1597.5 31012.5 ;
      RECT  1462.5 31077.5 1597.5 31012.5 ;
      RECT  1462.5 31267.5 1597.5 31202.5 ;
      RECT  2437.5 30907.5 2572.5 30842.5 ;
      RECT  1462.5 30907.5 1597.5 30842.5 ;
      RECT  1905.0 31210.0 2040.0 31145.0 ;
      RECT  1905.0 31210.0 2040.0 31145.0 ;
      RECT  1940.0 31045.0 2005.0 30980.0 ;
      RECT  2657.5 31335.0 2722.5 30775.0 ;
      RECT  1312.5 31335.0 1377.5 30775.0 ;
      RECT  1182.5 28552.5 1377.5 28617.5 ;
      RECT  342.5 28552.5 -32.5 28617.5 ;
      RECT  342.5 28932.5 -32.5 28997.5 ;
      RECT  185.0 29292.5 8.881784197e-13 29357.5 ;
      RECT  1345.0 29292.5 1160.0 29357.5 ;
      RECT  342.5 28552.5 207.5 28617.5 ;
      RECT  342.5 28742.5 207.5 28807.5 ;
      RECT  342.5 28742.5 207.5 28807.5 ;
      RECT  342.5 28552.5 207.5 28617.5 ;
      RECT  342.5 28742.5 207.5 28807.5 ;
      RECT  342.5 28932.5 207.5 28997.5 ;
      RECT  342.5 28932.5 207.5 28997.5 ;
      RECT  342.5 28742.5 207.5 28807.5 ;
      RECT  342.5 28932.5 207.5 28997.5 ;
      RECT  342.5 29122.5 207.5 29187.5 ;
      RECT  342.5 29122.5 207.5 29187.5 ;
      RECT  342.5 28932.5 207.5 28997.5 ;
      RECT  1182.5 28552.5 1047.5 28617.5 ;
      RECT  1182.5 28742.5 1047.5 28807.5 ;
      RECT  1182.5 28742.5 1047.5 28807.5 ;
      RECT  1182.5 28552.5 1047.5 28617.5 ;
      RECT  1182.5 28742.5 1047.5 28807.5 ;
      RECT  1182.5 28932.5 1047.5 28997.5 ;
      RECT  1182.5 28932.5 1047.5 28997.5 ;
      RECT  1182.5 28742.5 1047.5 28807.5 ;
      RECT  1182.5 28932.5 1047.5 28997.5 ;
      RECT  1182.5 29122.5 1047.5 29187.5 ;
      RECT  1182.5 29122.5 1047.5 29187.5 ;
      RECT  1182.5 28932.5 1047.5 28997.5 ;
      RECT  252.5 29292.5 117.5 29357.5 ;
      RECT  1227.5 29292.5 1092.5 29357.5 ;
      RECT  970.0 29127.5 905.0 28992.5 ;
      RECT  830.0 28937.5 765.0 28802.5 ;
      RECT  690.0 28747.5 625.0 28612.5 ;
      RECT  342.5 28742.5 207.5 28807.5 ;
      RECT  342.5 29122.5 207.5 29187.5 ;
      RECT  1182.5 29122.5 1047.5 29187.5 ;
      RECT  725.0 29122.5 590.0 29187.5 ;
      RECT  690.0 28612.5 625.0 28747.5 ;
      RECT  830.0 28802.5 765.0 28937.5 ;
      RECT  970.0 28992.5 905.0 29127.5 ;
      RECT  725.0 29122.5 590.0 29187.5 ;
      RECT  32.5 28485.0 -32.5 29495.0 ;
      RECT  1377.5 28485.0 1312.5 29495.0 ;
      RECT  185.0 29922.5 8.881784197e-13 29987.5 ;
      RECT  1345.0 29922.5 1160.0 29987.5 ;
      RECT  1227.5 29562.5 1377.5 29627.5 ;
      RECT  342.5 29562.5 -32.5 29627.5 ;
      RECT  1227.5 29752.5 342.5 29817.5 ;
      RECT  342.5 29562.5 207.5 29627.5 ;
      RECT  342.5 29752.5 207.5 29817.5 ;
      RECT  342.5 29752.5 207.5 29817.5 ;
      RECT  342.5 29562.5 207.5 29627.5 ;
      RECT  1227.5 29562.5 1092.5 29627.5 ;
      RECT  1227.5 29752.5 1092.5 29817.5 ;
      RECT  1227.5 29752.5 1092.5 29817.5 ;
      RECT  1227.5 29562.5 1092.5 29627.5 ;
      RECT  252.5 29922.5 117.5 29987.5 ;
      RECT  1227.5 29922.5 1092.5 29987.5 ;
      RECT  785.0 29620.0 650.0 29685.0 ;
      RECT  785.0 29620.0 650.0 29685.0 ;
      RECT  750.0 29785.0 685.0 29850.0 ;
      RECT  32.5 29495.0 -32.5 30055.0 ;
      RECT  1377.5 29495.0 1312.5 30055.0 ;
      RECT  185.0 30482.5 8.881784197e-13 30547.5 ;
      RECT  1345.0 30482.5 1160.0 30547.5 ;
      RECT  1227.5 30122.5 1377.5 30187.5 ;
      RECT  342.5 30122.5 -32.5 30187.5 ;
      RECT  1227.5 30312.5 342.5 30377.5 ;
      RECT  342.5 30122.5 207.5 30187.5 ;
      RECT  342.5 30312.5 207.5 30377.5 ;
      RECT  342.5 30312.5 207.5 30377.5 ;
      RECT  342.5 30122.5 207.5 30187.5 ;
      RECT  1227.5 30122.5 1092.5 30187.5 ;
      RECT  1227.5 30312.5 1092.5 30377.5 ;
      RECT  1227.5 30312.5 1092.5 30377.5 ;
      RECT  1227.5 30122.5 1092.5 30187.5 ;
      RECT  252.5 30482.5 117.5 30547.5 ;
      RECT  1227.5 30482.5 1092.5 30547.5 ;
      RECT  785.0 30180.0 650.0 30245.0 ;
      RECT  785.0 30180.0 650.0 30245.0 ;
      RECT  750.0 30345.0 685.0 30410.0 ;
      RECT  32.5 30055.0 -32.5 30615.0 ;
      RECT  1377.5 30055.0 1312.5 30615.0 ;
      RECT  185.0 31042.5 8.881784197e-13 31107.5 ;
      RECT  1345.0 31042.5 1160.0 31107.5 ;
      RECT  1227.5 30682.5 1377.5 30747.5 ;
      RECT  342.5 30682.5 -32.5 30747.5 ;
      RECT  1227.5 30872.5 342.5 30937.5 ;
      RECT  342.5 30682.5 207.5 30747.5 ;
      RECT  342.5 30872.5 207.5 30937.5 ;
      RECT  342.5 30872.5 207.5 30937.5 ;
      RECT  342.5 30682.5 207.5 30747.5 ;
      RECT  1227.5 30682.5 1092.5 30747.5 ;
      RECT  1227.5 30872.5 1092.5 30937.5 ;
      RECT  1227.5 30872.5 1092.5 30937.5 ;
      RECT  1227.5 30682.5 1092.5 30747.5 ;
      RECT  252.5 31042.5 117.5 31107.5 ;
      RECT  1227.5 31042.5 1092.5 31107.5 ;
      RECT  785.0 30740.0 650.0 30805.0 ;
      RECT  785.0 30740.0 650.0 30805.0 ;
      RECT  750.0 30905.0 685.0 30970.0 ;
      RECT  32.5 30615.0 -32.5 31175.0 ;
      RECT  1377.5 30615.0 1312.5 31175.0 ;
      RECT  1312.5 33907.5 1025.0 33972.5 ;
      RECT  1312.5 36317.5 1025.0 36382.5 ;
      RECT  1377.5 31862.5 935.0 31927.5 ;
      RECT  935.0 31862.5 230.0 31927.5 ;
      RECT  20.0 35112.5 935.0 35177.5 ;
      RECT  20.0 32422.5 935.0 32487.5 ;
      RECT  2005.0 33435.0 1940.0 34135.0 ;
      RECT  2005.0 33627.5 1940.0 33692.5 ;
      RECT  2005.0 33435.0 1940.0 33660.0 ;
      RECT  1972.5 33627.5 1025.0 33692.5 ;
      RECT  2690.0 33497.5 2465.0 33562.5 ;
      RECT  2430.0 32627.5 2365.0 32692.5 ;
      RECT  2005.0 32627.5 1940.0 32692.5 ;
      RECT  2430.0 32660.0 2365.0 33307.5 ;
      RECT  2397.5 32627.5 1972.5 32692.5 ;
      RECT  2005.0 32330.0 1940.0 32660.0 ;
      RECT  1972.5 32627.5 1172.5 32692.5 ;
      RECT  1172.5 32030.0 750.0 32095.0 ;
      RECT  2040.0 32265.0 1905.0 32330.0 ;
      RECT  2005.0 34135.0 1940.0 34340.0 ;
      RECT  2505.0 32027.5 2690.0 31962.5 ;
      RECT  1345.0 32027.5 1530.0 31962.5 ;
      RECT  1462.5 32387.5 1312.5 32322.5 ;
      RECT  2347.5 32387.5 2722.5 32322.5 ;
      RECT  1462.5 32197.5 2347.5 32132.5 ;
      RECT  2347.5 32387.5 2482.5 32322.5 ;
      RECT  2347.5 32197.5 2482.5 32132.5 ;
      RECT  2347.5 32197.5 2482.5 32132.5 ;
      RECT  2347.5 32387.5 2482.5 32322.5 ;
      RECT  1462.5 32387.5 1597.5 32322.5 ;
      RECT  1462.5 32197.5 1597.5 32132.5 ;
      RECT  1462.5 32197.5 1597.5 32132.5 ;
      RECT  1462.5 32387.5 1597.5 32322.5 ;
      RECT  2437.5 32027.5 2572.5 31962.5 ;
      RECT  1462.5 32027.5 1597.5 31962.5 ;
      RECT  1905.0 32330.0 2040.0 32265.0 ;
      RECT  1905.0 32330.0 2040.0 32265.0 ;
      RECT  1940.0 32165.0 2005.0 32100.0 ;
      RECT  2657.5 32455.0 2722.5 31895.0 ;
      RECT  1312.5 32455.0 1377.5 31895.0 ;
      RECT  2330.0 33307.5 2465.0 33372.5 ;
      RECT  2330.0 33497.5 2465.0 33562.5 ;
      RECT  2330.0 33497.5 2465.0 33562.5 ;
      RECT  2330.0 33307.5 2465.0 33372.5 ;
      RECT  1312.5 35352.5 1377.5 35417.5 ;
      RECT  4002.5 35352.5 4067.5 35417.5 ;
      RECT  1312.5 35255.0 1377.5 35385.0 ;
      RECT  1345.0 35352.5 4035.0 35417.5 ;
      RECT  4002.5 35255.0 4067.5 35385.0 ;
      RECT  2875.0 34562.5 2690.0 34627.5 ;
      RECT  4035.0 34562.5 3850.0 34627.5 ;
      RECT  3917.5 34202.5 4067.5 34267.5 ;
      RECT  3032.5 34202.5 2657.5 34267.5 ;
      RECT  3917.5 34392.5 3032.5 34457.5 ;
      RECT  3032.5 34202.5 2897.5 34267.5 ;
      RECT  3032.5 34392.5 2897.5 34457.5 ;
      RECT  3032.5 34392.5 2897.5 34457.5 ;
      RECT  3032.5 34202.5 2897.5 34267.5 ;
      RECT  3917.5 34202.5 3782.5 34267.5 ;
      RECT  3917.5 34392.5 3782.5 34457.5 ;
      RECT  3917.5 34392.5 3782.5 34457.5 ;
      RECT  3917.5 34202.5 3782.5 34267.5 ;
      RECT  2942.5 34562.5 2807.5 34627.5 ;
      RECT  3917.5 34562.5 3782.5 34627.5 ;
      RECT  3475.0 34260.0 3340.0 34325.0 ;
      RECT  3475.0 34260.0 3340.0 34325.0 ;
      RECT  3440.0 34425.0 3375.0 34490.0 ;
      RECT  2722.5 34135.0 2657.5 34695.0 ;
      RECT  4067.5 34135.0 4002.5 34695.0 ;
      RECT  2875.0 35122.5 2690.0 35187.5 ;
      RECT  4035.0 35122.5 3850.0 35187.5 ;
      RECT  3917.5 34762.5 4067.5 34827.5 ;
      RECT  3032.5 34762.5 2657.5 34827.5 ;
      RECT  3917.5 34952.5 3032.5 35017.5 ;
      RECT  3032.5 34762.5 2897.5 34827.5 ;
      RECT  3032.5 34952.5 2897.5 35017.5 ;
      RECT  3032.5 34952.5 2897.5 35017.5 ;
      RECT  3032.5 34762.5 2897.5 34827.5 ;
      RECT  3917.5 34762.5 3782.5 34827.5 ;
      RECT  3917.5 34952.5 3782.5 35017.5 ;
      RECT  3917.5 34952.5 3782.5 35017.5 ;
      RECT  3917.5 34762.5 3782.5 34827.5 ;
      RECT  2942.5 35122.5 2807.5 35187.5 ;
      RECT  3917.5 35122.5 3782.5 35187.5 ;
      RECT  3475.0 34820.0 3340.0 34885.0 ;
      RECT  3475.0 34820.0 3340.0 34885.0 ;
      RECT  3440.0 34985.0 3375.0 35050.0 ;
      RECT  2722.5 34695.0 2657.5 35255.0 ;
      RECT  4067.5 34695.0 4002.5 35255.0 ;
      RECT  3340.0 34820.0 3475.0 34885.0 ;
      RECT  2505.0 34827.5 2690.0 34762.5 ;
      RECT  1345.0 34827.5 1530.0 34762.5 ;
      RECT  1462.5 35187.5 1312.5 35122.5 ;
      RECT  2347.5 35187.5 2722.5 35122.5 ;
      RECT  1462.5 34997.5 2347.5 34932.5 ;
      RECT  2347.5 35187.5 2482.5 35122.5 ;
      RECT  2347.5 34997.5 2482.5 34932.5 ;
      RECT  2347.5 34997.5 2482.5 34932.5 ;
      RECT  2347.5 35187.5 2482.5 35122.5 ;
      RECT  1462.5 35187.5 1597.5 35122.5 ;
      RECT  1462.5 34997.5 1597.5 34932.5 ;
      RECT  1462.5 34997.5 1597.5 34932.5 ;
      RECT  1462.5 35187.5 1597.5 35122.5 ;
      RECT  2437.5 34827.5 2572.5 34762.5 ;
      RECT  1462.5 34827.5 1597.5 34762.5 ;
      RECT  1905.0 35130.0 2040.0 35065.0 ;
      RECT  1905.0 35130.0 2040.0 35065.0 ;
      RECT  1940.0 34965.0 2005.0 34900.0 ;
      RECT  2657.5 35255.0 2722.5 34695.0 ;
      RECT  1312.5 35255.0 1377.5 34695.0 ;
      RECT  1905.0 35065.0 2040.0 35130.0 ;
      RECT  2505.0 34267.5 2690.0 34202.5 ;
      RECT  1345.0 34267.5 1530.0 34202.5 ;
      RECT  1462.5 34627.5 1312.5 34562.5 ;
      RECT  2347.5 34627.5 2722.5 34562.5 ;
      RECT  1462.5 34437.5 2347.5 34372.5 ;
      RECT  2347.5 34627.5 2482.5 34562.5 ;
      RECT  2347.5 34437.5 2482.5 34372.5 ;
      RECT  2347.5 34437.5 2482.5 34372.5 ;
      RECT  2347.5 34627.5 2482.5 34562.5 ;
      RECT  1462.5 34627.5 1597.5 34562.5 ;
      RECT  1462.5 34437.5 1597.5 34372.5 ;
      RECT  1462.5 34437.5 1597.5 34372.5 ;
      RECT  1462.5 34627.5 1597.5 34562.5 ;
      RECT  2437.5 34267.5 2572.5 34202.5 ;
      RECT  1462.5 34267.5 1597.5 34202.5 ;
      RECT  1905.0 34570.0 2040.0 34505.0 ;
      RECT  1905.0 34570.0 2040.0 34505.0 ;
      RECT  1940.0 34405.0 2005.0 34340.0 ;
      RECT  2657.5 34695.0 2722.5 34135.0 ;
      RECT  1312.5 34695.0 1377.5 34135.0 ;
      RECT  1905.0 34505.0 2040.0 34570.0 ;
      RECT  3340.0 34425.0 3475.0 34490.0 ;
      RECT  3340.0 34985.0 3475.0 35050.0 ;
      RECT  1905.0 34900.0 2040.0 34965.0 ;
      RECT  3340.0 34260.0 3475.0 34325.0 ;
      RECT  1940.0 34135.0 2005.0 34340.0 ;
      RECT  2657.5 34135.0 2722.5 35255.0 ;
      RECT  1312.5 34135.0 1377.5 35255.0 ;
      RECT  4002.5 34135.0 4067.5 35255.0 ;
      RECT  935.0 33800.0 225.0 32455.0 ;
      RECT  935.0 33800.0 230.0 35145.0 ;
      RECT  935.0 36490.0 230.0 35145.0 ;
      RECT  1025.0 33907.5 140.0 33972.5 ;
      RECT  1025.0 36317.5 140.0 36382.5 ;
      RECT  1025.0 35112.5 140.0 35177.5 ;
      RECT  1025.0 33767.5 140.0 33832.5 ;
      RECT  1025.0 36457.5 140.0 36522.5 ;
      RECT  1345.0 33872.5 1280.0 34007.5 ;
      RECT  1345.0 36282.5 1280.0 36417.5 ;
      RECT  1342.5 34135.0 1277.5 34270.0 ;
      RECT  1377.5 31760.0 1312.5 31895.0 ;
      RECT  867.5 31862.5 1002.5 31927.5 ;
      RECT  162.5 31862.5 297.5 31927.5 ;
      RECT  2005.0 33367.5 1940.0 33502.5 ;
      RECT  1105.0 32627.5 1240.0 32692.5 ;
      RECT  1105.0 32030.0 1240.0 32095.0 ;
      RECT  682.5 32030.0 817.5 32095.0 ;
      RECT  3475.0 31335.0 3410.0 34260.0 ;
      RECT  2005.0 31335.0 1940.0 32100.0 ;
      RECT  20.0 31335.0 -45.0 36577.5 ;
      RECT  2722.5 31335.0 2657.5 34135.0 ;
      RECT  1377.5 31335.0 1312.5 31895.0 ;
      RECT  4067.5 31335.0 4002.5 34135.0 ;
      RECT  3455.0 26182.5 3390.0 26047.5 ;
      RECT  3455.0 22102.5 3390.0 21967.5 ;
      RECT  2517.5 19535.0 2452.5 19400.0 ;
      RECT  1962.5 26182.5 1897.5 26047.5 ;
      RECT  1747.5 26592.5 1682.5 26457.5 ;
      RECT  2017.5 29130.0 1952.5 28995.0 ;
      RECT  1802.5 29387.5 1737.5 29252.5 ;
      RECT  3380.0 27617.5 3315.0 27482.5 ;
      RECT  3520.0 27412.5 3455.0 27277.5 ;
      RECT  3660.0 26797.5 3595.0 26662.5 ;
      RECT  690.0 27617.5 625.0 27482.5 ;
      RECT  830.0 26797.5 765.0 26662.5 ;
      RECT  970.0 27002.5 905.0 26867.5 ;
      RECT  1997.5 28812.5 1862.5 28877.5 ;
      RECT  2052.5 29957.5 1917.5 30022.5 ;
      RECT  785.0 31142.5 650.0 31207.5 ;
      RECT  2040.0 30182.5 1905.0 30247.5 ;
      RECT  4067.5 26387.5 4002.5 26252.5 ;
      RECT  2722.5 27207.5 2657.5 27072.5 ;
      RECT  1377.5 26387.5 1312.5 26252.5 ;
      RECT  32.5 27207.5 -32.5 27072.5 ;
      RECT  3475.0 19230.0 3340.0 19420.0 ;
      RECT  2722.5 19230.0 2657.5 19295.0 ;
      RECT  4067.5 19230.0 4002.5 19295.0 ;
      RECT  4417.5 27107.5 4282.5 27172.5 ;
   LAYER  metal2 ;
      RECT  14007.5 30010.0 14077.5 30215.0 ;
      RECT  13802.5 30970.0 13872.5 31175.0 ;
      RECT  13392.5 28640.0 13462.5 28845.0 ;
      RECT  13187.5 29785.0 13257.5 29990.0 ;
      RECT  13597.5 27345.0 13667.5 27550.0 ;
      RECT  12982.5 25910.0 13052.5 26115.0 ;
      RECT  4035.0 27105.0 4350.0 27175.0 ;
      RECT  12567.5 26115.0 12637.5 26320.0 ;
      RECT  12982.5 0.0 13052.5 42337.5 ;
      RECT  13187.5 0.0 13257.5 42337.5 ;
      RECT  13392.5 0.0 13462.5 42337.5 ;
      RECT  13597.5 0.0 13667.5 42337.5 ;
      RECT  13802.5 0.0 13872.5 42337.5 ;
      RECT  14007.5 0.0 14077.5 42337.5 ;
      RECT  11402.5 4690.0 11472.5 19090.0 ;
      RECT  11607.5 4690.0 11677.5 19090.0 ;
      RECT  11812.5 4690.0 11882.5 19090.0 ;
      RECT  12017.5 4690.0 12087.5 19090.0 ;
      RECT  14670.0 40765.0 14740.0 41170.0 ;
      RECT  15005.0 40765.0 15075.0 41170.0 ;
      RECT  15375.0 40765.0 15445.0 41170.0 ;
      RECT  15710.0 40765.0 15780.0 41170.0 ;
      RECT  14837.5 440.0 14907.5 510.0 ;
      RECT  14662.5 440.0 14872.5 510.0 ;
      RECT  14837.5 475.0 14907.5 615.0 ;
      RECT  15542.5 440.0 15612.5 510.0 ;
      RECT  15367.5 440.0 15577.5 510.0 ;
      RECT  15542.5 475.0 15612.5 615.0 ;
      RECT  8805.0 40610.0 8875.0 40815.0 ;
      RECT  14520.0 19090.0 15225.0 20435.0 ;
      RECT  14520.0 21780.0 15225.0 20435.0 ;
      RECT  14520.0 21780.0 15225.0 23125.0 ;
      RECT  14520.0 24470.0 15225.0 23125.0 ;
      RECT  14520.0 24470.0 15225.0 25815.0 ;
      RECT  14520.0 27160.0 15225.0 25815.0 ;
      RECT  14520.0 27160.0 15225.0 28505.0 ;
      RECT  14520.0 29850.0 15225.0 28505.0 ;
      RECT  14520.0 29850.0 15225.0 31195.0 ;
      RECT  14520.0 32540.0 15225.0 31195.0 ;
      RECT  14520.0 32540.0 15225.0 33885.0 ;
      RECT  14520.0 35230.0 15225.0 33885.0 ;
      RECT  14520.0 35230.0 15225.0 36575.0 ;
      RECT  14520.0 37920.0 15225.0 36575.0 ;
      RECT  14520.0 37920.0 15225.0 39265.0 ;
      RECT  14520.0 40610.0 15225.0 39265.0 ;
      RECT  15225.0 19090.0 15930.0 20435.0 ;
      RECT  15225.0 21780.0 15930.0 20435.0 ;
      RECT  15225.0 21780.0 15930.0 23125.0 ;
      RECT  15225.0 24470.0 15930.0 23125.0 ;
      RECT  15225.0 24470.0 15930.0 25815.0 ;
      RECT  15225.0 27160.0 15930.0 25815.0 ;
      RECT  15225.0 27160.0 15930.0 28505.0 ;
      RECT  15225.0 29850.0 15930.0 28505.0 ;
      RECT  15225.0 29850.0 15930.0 31195.0 ;
      RECT  15225.0 32540.0 15930.0 31195.0 ;
      RECT  15225.0 32540.0 15930.0 33885.0 ;
      RECT  15225.0 35230.0 15930.0 33885.0 ;
      RECT  15225.0 35230.0 15930.0 36575.0 ;
      RECT  15225.0 37920.0 15930.0 36575.0 ;
      RECT  15225.0 37920.0 15930.0 39265.0 ;
      RECT  15225.0 40610.0 15930.0 39265.0 ;
      RECT  14670.0 18990.0 14740.0 40765.0 ;
      RECT  15005.0 18990.0 15075.0 40765.0 ;
      RECT  15375.0 18990.0 15445.0 40765.0 ;
      RECT  15710.0 18990.0 15780.0 40765.0 ;
      RECT  14485.0 18990.0 14555.0 40765.0 ;
      RECT  15190.0 18990.0 15260.0 40765.0 ;
      RECT  15895.0 18990.0 15965.0 40765.0 ;
      RECT  14670.0 41292.5 14747.5 41427.5 ;
      RECT  14872.5 41292.5 15075.0 41427.5 ;
      RECT  14670.0 41822.5 14747.5 41957.5 ;
      RECT  15005.0 41822.5 15127.5 41957.5 ;
      RECT  14680.0 41292.5 14750.0 41427.5 ;
      RECT  14870.0 41292.5 14940.0 41427.5 ;
      RECT  14680.0 41822.5 14750.0 41957.5 ;
      RECT  15060.0 41822.5 15130.0 41957.5 ;
      RECT  14670.0 41170.0 14740.0 42337.5 ;
      RECT  15005.0 41170.0 15075.0 42337.5 ;
      RECT  15375.0 41292.5 15452.5 41427.5 ;
      RECT  15577.5 41292.5 15780.0 41427.5 ;
      RECT  15375.0 41822.5 15452.5 41957.5 ;
      RECT  15710.0 41822.5 15832.5 41957.5 ;
      RECT  15385.0 41292.5 15455.0 41427.5 ;
      RECT  15575.0 41292.5 15645.0 41427.5 ;
      RECT  15385.0 41822.5 15455.0 41957.5 ;
      RECT  15765.0 41822.5 15835.0 41957.5 ;
      RECT  15375.0 41170.0 15445.0 42337.5 ;
      RECT  15710.0 41170.0 15780.0 42337.5 ;
      RECT  14670.0 41170.0 14740.0 42337.5 ;
      RECT  15005.0 41170.0 15075.0 42337.5 ;
      RECT  15375.0 41170.0 15445.0 42337.5 ;
      RECT  15710.0 41170.0 15780.0 42337.5 ;
      RECT  14520.0 14205.0 15225.0 19090.0 ;
      RECT  15225.0 14205.0 15930.0 19090.0 ;
      RECT  14670.0 14205.0 14740.0 19090.0 ;
      RECT  15005.0 14205.0 15075.0 18290.0 ;
      RECT  15375.0 14205.0 15445.0 19090.0 ;
      RECT  15710.0 14205.0 15780.0 18290.0 ;
      RECT  14520.0 10030.0 15225.0 14205.0 ;
      RECT  15225.0 10030.0 15930.0 14205.0 ;
      RECT  14837.5 10030.0 14907.5 10170.0 ;
      RECT  15542.5 10030.0 15612.5 10170.0 ;
      RECT  14670.0 13905.0 14740.0 14205.0 ;
      RECT  15005.0 11765.0 15075.0 14205.0 ;
      RECT  15375.0 13905.0 15445.0 14205.0 ;
      RECT  15710.0 11765.0 15780.0 14205.0 ;
      RECT  14520.0 3590.0 15225.0 10030.0 ;
      RECT  15930.0 3590.0 15225.0 10030.0 ;
      RECT  14837.5 3590.0 14907.5 3735.0 ;
      RECT  15542.5 3590.0 15612.5 3735.0 ;
      RECT  14837.5 9760.0 14907.5 10030.0 ;
      RECT  14682.5 9342.5 14752.5 10030.0 ;
      RECT  15542.5 9760.0 15612.5 10030.0 ;
      RECT  15697.5 9342.5 15767.5 10030.0 ;
      RECT  14485.0 3590.0 14555.0 10030.0 ;
      RECT  15190.0 3590.0 15260.0 10030.0 ;
      RECT  15895.0 3590.0 15965.0 10030.0 ;
      RECT  14520.0 3590.0 15225.0 615.0 ;
      RECT  15225.0 3590.0 15930.0 615.0 ;
      RECT  14837.5 855.0 14907.5 615.0 ;
      RECT  15542.5 855.0 15612.5 615.0 ;
      RECT  14837.5 3590.0 14907.5 3240.0 ;
      RECT  15542.5 3590.0 15612.5 3240.0 ;
      RECT  5730.0 8330.0 5800.0 40610.0 ;
      RECT  5905.0 8330.0 5975.0 40610.0 ;
      RECT  6080.0 8330.0 6150.0 40610.0 ;
      RECT  6255.0 8330.0 6325.0 40610.0 ;
      RECT  6430.0 8330.0 6500.0 40610.0 ;
      RECT  6605.0 8330.0 6675.0 40610.0 ;
      RECT  6780.0 8330.0 6850.0 40610.0 ;
      RECT  6955.0 8330.0 7025.0 40610.0 ;
      RECT  9160.0 8330.0 9090.0 13570.0 ;
      RECT  8885.0 8330.0 8815.0 13570.0 ;
      RECT  9710.0 8330.0 9640.0 13570.0 ;
      RECT  9435.0 8330.0 9365.0 13570.0 ;
      RECT  8355.0 8935.0 8285.0 9005.0 ;
      RECT  8165.0 8935.0 8095.0 9005.0 ;
      RECT  8355.0 8970.0 8285.0 9332.5 ;
      RECT  8320.0 8935.0 8130.0 9005.0 ;
      RECT  8165.0 8627.5 8095.0 8970.0 ;
      RECT  8355.0 9332.5 8285.0 9467.5 ;
      RECT  8165.0 8492.5 8095.0 8627.5 ;
      RECT  8062.5 8935.0 8197.5 9005.0 ;
      RECT  8355.0 10415.0 8285.0 10345.0 ;
      RECT  8165.0 10415.0 8095.0 10345.0 ;
      RECT  8355.0 10380.0 8285.0 10017.5 ;
      RECT  8320.0 10415.0 8130.0 10345.0 ;
      RECT  8165.0 10722.5 8095.0 10380.0 ;
      RECT  8355.0 10017.5 8285.0 9882.5 ;
      RECT  8165.0 10857.5 8095.0 10722.5 ;
      RECT  8062.5 10415.0 8197.5 10345.0 ;
      RECT  8355.0 11625.0 8285.0 11695.0 ;
      RECT  8165.0 11625.0 8095.0 11695.0 ;
      RECT  8355.0 11660.0 8285.0 12022.5 ;
      RECT  8320.0 11625.0 8130.0 11695.0 ;
      RECT  8165.0 11317.5 8095.0 11660.0 ;
      RECT  8355.0 12022.5 8285.0 12157.5 ;
      RECT  8165.0 11182.5 8095.0 11317.5 ;
      RECT  8062.5 11625.0 8197.5 11695.0 ;
      RECT  8355.0 13105.0 8285.0 13035.0 ;
      RECT  8165.0 13105.0 8095.0 13035.0 ;
      RECT  8355.0 13070.0 8285.0 12707.5 ;
      RECT  8320.0 13105.0 8130.0 13035.0 ;
      RECT  8165.0 13412.5 8095.0 13070.0 ;
      RECT  8355.0 12707.5 8285.0 12572.5 ;
      RECT  8165.0 13547.5 8095.0 13412.5 ;
      RECT  8062.5 13105.0 8197.5 13035.0 ;
      RECT  9607.5 9445.0 9742.5 9515.0 ;
      RECT  10992.5 8922.5 11127.5 8992.5 ;
      RECT  9332.5 10790.0 9467.5 10860.0 ;
      RECT  10717.5 10357.5 10852.5 10427.5 ;
      RECT  10992.5 11120.0 11127.5 11190.0 ;
      RECT  9057.5 11120.0 9192.5 11190.0 ;
      RECT  10717.5 12465.0 10852.5 12535.0 ;
      RECT  8782.5 12465.0 8917.5 12535.0 ;
      RECT  9607.5 8935.0 9742.5 9005.0 ;
      RECT  9332.5 8720.0 9467.5 8790.0 ;
      RECT  9057.5 10345.0 9192.5 10415.0 ;
      RECT  9332.5 10560.0 9467.5 10630.0 ;
      RECT  9607.5 11625.0 9742.5 11695.0 ;
      RECT  8782.5 11410.0 8917.5 11480.0 ;
      RECT  9057.5 13035.0 9192.5 13105.0 ;
      RECT  8782.5 13250.0 8917.5 13320.0 ;
      RECT  11095.0 8330.0 11025.0 13570.0 ;
      RECT  10820.0 8330.0 10750.0 13570.0 ;
      RECT  9160.0 13710.0 9090.0 18950.0 ;
      RECT  8885.0 13710.0 8815.0 18950.0 ;
      RECT  9710.0 13710.0 9640.0 18950.0 ;
      RECT  9435.0 13710.0 9365.0 18950.0 ;
      RECT  8355.0 14315.0 8285.0 14385.0 ;
      RECT  8165.0 14315.0 8095.0 14385.0 ;
      RECT  8355.0 14350.0 8285.0 14712.5 ;
      RECT  8320.0 14315.0 8130.0 14385.0 ;
      RECT  8165.0 14007.5 8095.0 14350.0 ;
      RECT  8355.0 14712.5 8285.0 14847.5 ;
      RECT  8165.0 13872.5 8095.0 14007.5 ;
      RECT  8062.5 14315.0 8197.5 14385.0 ;
      RECT  8355.0 15795.0 8285.0 15725.0 ;
      RECT  8165.0 15795.0 8095.0 15725.0 ;
      RECT  8355.0 15760.0 8285.0 15397.5 ;
      RECT  8320.0 15795.0 8130.0 15725.0 ;
      RECT  8165.0 16102.5 8095.0 15760.0 ;
      RECT  8355.0 15397.5 8285.0 15262.5 ;
      RECT  8165.0 16237.5 8095.0 16102.5 ;
      RECT  8062.5 15795.0 8197.5 15725.0 ;
      RECT  8355.0 17005.0 8285.0 17075.0 ;
      RECT  8165.0 17005.0 8095.0 17075.0 ;
      RECT  8355.0 17040.0 8285.0 17402.5 ;
      RECT  8320.0 17005.0 8130.0 17075.0 ;
      RECT  8165.0 16697.5 8095.0 17040.0 ;
      RECT  8355.0 17402.5 8285.0 17537.5 ;
      RECT  8165.0 16562.5 8095.0 16697.5 ;
      RECT  8062.5 17005.0 8197.5 17075.0 ;
      RECT  8355.0 18485.0 8285.0 18415.0 ;
      RECT  8165.0 18485.0 8095.0 18415.0 ;
      RECT  8355.0 18450.0 8285.0 18087.5 ;
      RECT  8320.0 18485.0 8130.0 18415.0 ;
      RECT  8165.0 18792.5 8095.0 18450.0 ;
      RECT  8355.0 18087.5 8285.0 17952.5 ;
      RECT  8165.0 18927.5 8095.0 18792.5 ;
      RECT  8062.5 18485.0 8197.5 18415.0 ;
      RECT  9607.5 14825.0 9742.5 14895.0 ;
      RECT  10992.5 14302.5 11127.5 14372.5 ;
      RECT  9332.5 16170.0 9467.5 16240.0 ;
      RECT  10717.5 15737.5 10852.5 15807.5 ;
      RECT  10992.5 16500.0 11127.5 16570.0 ;
      RECT  9057.5 16500.0 9192.5 16570.0 ;
      RECT  10717.5 17845.0 10852.5 17915.0 ;
      RECT  8782.5 17845.0 8917.5 17915.0 ;
      RECT  9607.5 14315.0 9742.5 14385.0 ;
      RECT  9332.5 14100.0 9467.5 14170.0 ;
      RECT  9057.5 15725.0 9192.5 15795.0 ;
      RECT  9332.5 15940.0 9467.5 16010.0 ;
      RECT  9607.5 17005.0 9742.5 17075.0 ;
      RECT  8782.5 16790.0 8917.5 16860.0 ;
      RECT  9057.5 18415.0 9192.5 18485.0 ;
      RECT  8782.5 18630.0 8917.5 18700.0 ;
      RECT  11095.0 13710.0 11025.0 18950.0 ;
      RECT  10820.0 13710.0 10750.0 18950.0 ;
      RECT  7385.0 19695.0 7455.0 19765.0 ;
      RECT  7575.0 19695.0 7645.0 19765.0 ;
      RECT  7385.0 19730.0 7455.0 20092.5 ;
      RECT  7420.0 19695.0 7610.0 19765.0 ;
      RECT  7575.0 19387.5 7645.0 19730.0 ;
      RECT  7385.0 20092.5 7455.0 20227.5 ;
      RECT  7575.0 19252.5 7645.0 19387.5 ;
      RECT  7677.5 19695.0 7542.5 19765.0 ;
      RECT  7385.0 21175.0 7455.0 21105.0 ;
      RECT  7575.0 21175.0 7645.0 21105.0 ;
      RECT  7385.0 21140.0 7455.0 20777.5 ;
      RECT  7420.0 21175.0 7610.0 21105.0 ;
      RECT  7575.0 21482.5 7645.0 21140.0 ;
      RECT  7385.0 20777.5 7455.0 20642.5 ;
      RECT  7575.0 21617.5 7645.0 21482.5 ;
      RECT  7677.5 21175.0 7542.5 21105.0 ;
      RECT  7385.0 22385.0 7455.0 22455.0 ;
      RECT  7575.0 22385.0 7645.0 22455.0 ;
      RECT  7385.0 22420.0 7455.0 22782.5 ;
      RECT  7420.0 22385.0 7610.0 22455.0 ;
      RECT  7575.0 22077.5 7645.0 22420.0 ;
      RECT  7385.0 22782.5 7455.0 22917.5 ;
      RECT  7575.0 21942.5 7645.0 22077.5 ;
      RECT  7677.5 22385.0 7542.5 22455.0 ;
      RECT  7385.0 23865.0 7455.0 23795.0 ;
      RECT  7575.0 23865.0 7645.0 23795.0 ;
      RECT  7385.0 23830.0 7455.0 23467.5 ;
      RECT  7420.0 23865.0 7610.0 23795.0 ;
      RECT  7575.0 24172.5 7645.0 23830.0 ;
      RECT  7385.0 23467.5 7455.0 23332.5 ;
      RECT  7575.0 24307.5 7645.0 24172.5 ;
      RECT  7677.5 23865.0 7542.5 23795.0 ;
      RECT  7385.0 25075.0 7455.0 25145.0 ;
      RECT  7575.0 25075.0 7645.0 25145.0 ;
      RECT  7385.0 25110.0 7455.0 25472.5 ;
      RECT  7420.0 25075.0 7610.0 25145.0 ;
      RECT  7575.0 24767.5 7645.0 25110.0 ;
      RECT  7385.0 25472.5 7455.0 25607.5 ;
      RECT  7575.0 24632.5 7645.0 24767.5 ;
      RECT  7677.5 25075.0 7542.5 25145.0 ;
      RECT  7385.0 26555.0 7455.0 26485.0 ;
      RECT  7575.0 26555.0 7645.0 26485.0 ;
      RECT  7385.0 26520.0 7455.0 26157.5 ;
      RECT  7420.0 26555.0 7610.0 26485.0 ;
      RECT  7575.0 26862.5 7645.0 26520.0 ;
      RECT  7385.0 26157.5 7455.0 26022.5 ;
      RECT  7575.0 26997.5 7645.0 26862.5 ;
      RECT  7677.5 26555.0 7542.5 26485.0 ;
      RECT  7385.0 27765.0 7455.0 27835.0 ;
      RECT  7575.0 27765.0 7645.0 27835.0 ;
      RECT  7385.0 27800.0 7455.0 28162.5 ;
      RECT  7420.0 27765.0 7610.0 27835.0 ;
      RECT  7575.0 27457.5 7645.0 27800.0 ;
      RECT  7385.0 28162.5 7455.0 28297.5 ;
      RECT  7575.0 27322.5 7645.0 27457.5 ;
      RECT  7677.5 27765.0 7542.5 27835.0 ;
      RECT  7385.0 29245.0 7455.0 29175.0 ;
      RECT  7575.0 29245.0 7645.0 29175.0 ;
      RECT  7385.0 29210.0 7455.0 28847.5 ;
      RECT  7420.0 29245.0 7610.0 29175.0 ;
      RECT  7575.0 29552.5 7645.0 29210.0 ;
      RECT  7385.0 28847.5 7455.0 28712.5 ;
      RECT  7575.0 29687.5 7645.0 29552.5 ;
      RECT  7677.5 29245.0 7542.5 29175.0 ;
      RECT  7385.0 30455.0 7455.0 30525.0 ;
      RECT  7575.0 30455.0 7645.0 30525.0 ;
      RECT  7385.0 30490.0 7455.0 30852.5 ;
      RECT  7420.0 30455.0 7610.0 30525.0 ;
      RECT  7575.0 30147.5 7645.0 30490.0 ;
      RECT  7385.0 30852.5 7455.0 30987.5 ;
      RECT  7575.0 30012.5 7645.0 30147.5 ;
      RECT  7677.5 30455.0 7542.5 30525.0 ;
      RECT  7385.0 31935.0 7455.0 31865.0 ;
      RECT  7575.0 31935.0 7645.0 31865.0 ;
      RECT  7385.0 31900.0 7455.0 31537.5 ;
      RECT  7420.0 31935.0 7610.0 31865.0 ;
      RECT  7575.0 32242.5 7645.0 31900.0 ;
      RECT  7385.0 31537.5 7455.0 31402.5 ;
      RECT  7575.0 32377.5 7645.0 32242.5 ;
      RECT  7677.5 31935.0 7542.5 31865.0 ;
      RECT  7385.0 33145.0 7455.0 33215.0 ;
      RECT  7575.0 33145.0 7645.0 33215.0 ;
      RECT  7385.0 33180.0 7455.0 33542.5 ;
      RECT  7420.0 33145.0 7610.0 33215.0 ;
      RECT  7575.0 32837.5 7645.0 33180.0 ;
      RECT  7385.0 33542.5 7455.0 33677.5 ;
      RECT  7575.0 32702.5 7645.0 32837.5 ;
      RECT  7677.5 33145.0 7542.5 33215.0 ;
      RECT  7385.0 34625.0 7455.0 34555.0 ;
      RECT  7575.0 34625.0 7645.0 34555.0 ;
      RECT  7385.0 34590.0 7455.0 34227.5 ;
      RECT  7420.0 34625.0 7610.0 34555.0 ;
      RECT  7575.0 34932.5 7645.0 34590.0 ;
      RECT  7385.0 34227.5 7455.0 34092.5 ;
      RECT  7575.0 35067.5 7645.0 34932.5 ;
      RECT  7677.5 34625.0 7542.5 34555.0 ;
      RECT  7385.0 35835.0 7455.0 35905.0 ;
      RECT  7575.0 35835.0 7645.0 35905.0 ;
      RECT  7385.0 35870.0 7455.0 36232.5 ;
      RECT  7420.0 35835.0 7610.0 35905.0 ;
      RECT  7575.0 35527.5 7645.0 35870.0 ;
      RECT  7385.0 36232.5 7455.0 36367.5 ;
      RECT  7575.0 35392.5 7645.0 35527.5 ;
      RECT  7677.5 35835.0 7542.5 35905.0 ;
      RECT  7385.0 37315.0 7455.0 37245.0 ;
      RECT  7575.0 37315.0 7645.0 37245.0 ;
      RECT  7385.0 37280.0 7455.0 36917.5 ;
      RECT  7420.0 37315.0 7610.0 37245.0 ;
      RECT  7575.0 37622.5 7645.0 37280.0 ;
      RECT  7385.0 36917.5 7455.0 36782.5 ;
      RECT  7575.0 37757.5 7645.0 37622.5 ;
      RECT  7677.5 37315.0 7542.5 37245.0 ;
      RECT  7385.0 38525.0 7455.0 38595.0 ;
      RECT  7575.0 38525.0 7645.0 38595.0 ;
      RECT  7385.0 38560.0 7455.0 38922.5 ;
      RECT  7420.0 38525.0 7610.0 38595.0 ;
      RECT  7575.0 38217.5 7645.0 38560.0 ;
      RECT  7385.0 38922.5 7455.0 39057.5 ;
      RECT  7575.0 38082.5 7645.0 38217.5 ;
      RECT  7677.5 38525.0 7542.5 38595.0 ;
      RECT  7385.0 40005.0 7455.0 39935.0 ;
      RECT  7575.0 40005.0 7645.0 39935.0 ;
      RECT  7385.0 39970.0 7455.0 39607.5 ;
      RECT  7420.0 40005.0 7610.0 39935.0 ;
      RECT  7575.0 40312.5 7645.0 39970.0 ;
      RECT  7385.0 39607.5 7455.0 39472.5 ;
      RECT  7575.0 40447.5 7645.0 40312.5 ;
      RECT  7677.5 40005.0 7542.5 39935.0 ;
      RECT  5832.5 8922.5 5697.5 8992.5 ;
      RECT  6007.5 10357.5 5872.5 10427.5 ;
      RECT  6182.5 11612.5 6047.5 11682.5 ;
      RECT  6357.5 13047.5 6222.5 13117.5 ;
      RECT  6532.5 14302.5 6397.5 14372.5 ;
      RECT  6707.5 15737.5 6572.5 15807.5 ;
      RECT  6882.5 16992.5 6747.5 17062.5 ;
      RECT  7057.5 18427.5 6922.5 18497.5 ;
      RECT  5832.5 19695.0 5697.5 19765.0 ;
      RECT  6532.5 19480.0 6397.5 19550.0 ;
      RECT  5832.5 21105.0 5697.5 21175.0 ;
      RECT  6707.5 21320.0 6572.5 21390.0 ;
      RECT  5832.5 22385.0 5697.5 22455.0 ;
      RECT  6882.5 22170.0 6747.5 22240.0 ;
      RECT  5832.5 23795.0 5697.5 23865.0 ;
      RECT  7057.5 24010.0 6922.5 24080.0 ;
      RECT  6007.5 25075.0 5872.5 25145.0 ;
      RECT  6532.5 24860.0 6397.5 24930.0 ;
      RECT  6007.5 26485.0 5872.5 26555.0 ;
      RECT  6707.5 26700.0 6572.5 26770.0 ;
      RECT  6007.5 27765.0 5872.5 27835.0 ;
      RECT  6882.5 27550.0 6747.5 27620.0 ;
      RECT  6007.5 29175.0 5872.5 29245.0 ;
      RECT  7057.5 29390.0 6922.5 29460.0 ;
      RECT  6182.5 30455.0 6047.5 30525.0 ;
      RECT  6532.5 30240.0 6397.5 30310.0 ;
      RECT  6182.5 31865.0 6047.5 31935.0 ;
      RECT  6707.5 32080.0 6572.5 32150.0 ;
      RECT  6182.5 33145.0 6047.5 33215.0 ;
      RECT  6882.5 32930.0 6747.5 33000.0 ;
      RECT  6182.5 34555.0 6047.5 34625.0 ;
      RECT  7057.5 34770.0 6922.5 34840.0 ;
      RECT  6357.5 35835.0 6222.5 35905.0 ;
      RECT  6532.5 35620.0 6397.5 35690.0 ;
      RECT  6357.5 37245.0 6222.5 37315.0 ;
      RECT  6707.5 37460.0 6572.5 37530.0 ;
      RECT  6357.5 38525.0 6222.5 38595.0 ;
      RECT  6882.5 38310.0 6747.5 38380.0 ;
      RECT  6357.5 39935.0 6222.5 40005.0 ;
      RECT  7057.5 40150.0 6922.5 40220.0 ;
      RECT  11025.0 8330.0 11095.0 13570.0 ;
      RECT  10750.0 8330.0 10820.0 13570.0 ;
      RECT  11025.0 13710.0 11095.0 18950.0 ;
      RECT  10750.0 13710.0 10820.0 18950.0 ;
      RECT  8945.0 19480.0 9015.0 19550.0 ;
      RECT  8945.0 19445.0 9015.0 19515.0 ;
      RECT  8980.0 19480.0 9942.5 19550.0 ;
      RECT  8945.0 21320.0 9015.0 21390.0 ;
      RECT  8945.0 21355.0 9015.0 21425.0 ;
      RECT  8980.0 21320.0 9942.5 21390.0 ;
      RECT  8945.0 22170.0 9015.0 22240.0 ;
      RECT  8945.0 22135.0 9015.0 22205.0 ;
      RECT  8980.0 22170.0 9942.5 22240.0 ;
      RECT  8945.0 24010.0 9015.0 24080.0 ;
      RECT  8945.0 24045.0 9015.0 24115.0 ;
      RECT  8980.0 24010.0 9942.5 24080.0 ;
      RECT  8945.0 24860.0 9015.0 24930.0 ;
      RECT  8945.0 24825.0 9015.0 24895.0 ;
      RECT  8980.0 24860.0 9942.5 24930.0 ;
      RECT  8945.0 26700.0 9015.0 26770.0 ;
      RECT  8945.0 26735.0 9015.0 26805.0 ;
      RECT  8980.0 26700.0 9942.5 26770.0 ;
      RECT  8945.0 27550.0 9015.0 27620.0 ;
      RECT  8945.0 27515.0 9015.0 27585.0 ;
      RECT  8980.0 27550.0 9942.5 27620.0 ;
      RECT  8945.0 29390.0 9015.0 29460.0 ;
      RECT  8945.0 29425.0 9015.0 29495.0 ;
      RECT  8980.0 29390.0 9942.5 29460.0 ;
      RECT  8945.0 30240.0 9015.0 30310.0 ;
      RECT  8945.0 30205.0 9015.0 30275.0 ;
      RECT  8980.0 30240.0 9942.5 30310.0 ;
      RECT  8945.0 32080.0 9015.0 32150.0 ;
      RECT  8945.0 32115.0 9015.0 32185.0 ;
      RECT  8980.0 32080.0 9942.5 32150.0 ;
      RECT  8945.0 32930.0 9015.0 33000.0 ;
      RECT  8945.0 32895.0 9015.0 32965.0 ;
      RECT  8980.0 32930.0 9942.5 33000.0 ;
      RECT  8945.0 34770.0 9015.0 34840.0 ;
      RECT  8945.0 34805.0 9015.0 34875.0 ;
      RECT  8980.0 34770.0 9942.5 34840.0 ;
      RECT  8945.0 35620.0 9015.0 35690.0 ;
      RECT  8945.0 35585.0 9015.0 35655.0 ;
      RECT  8980.0 35620.0 9942.5 35690.0 ;
      RECT  8945.0 37460.0 9015.0 37530.0 ;
      RECT  8945.0 37495.0 9015.0 37565.0 ;
      RECT  8980.0 37460.0 9942.5 37530.0 ;
      RECT  8945.0 38310.0 9015.0 38380.0 ;
      RECT  8945.0 38275.0 9015.0 38345.0 ;
      RECT  8980.0 38310.0 9942.5 38380.0 ;
      RECT  8945.0 40150.0 9015.0 40220.0 ;
      RECT  8945.0 40185.0 9015.0 40255.0 ;
      RECT  8980.0 40150.0 9942.5 40220.0 ;
      RECT  9880.0 19695.0 9950.0 19765.0 ;
      RECT  10070.0 19695.0 10140.0 19765.0 ;
      RECT  9880.0 19730.0 9950.0 20092.5 ;
      RECT  9915.0 19695.0 10105.0 19765.0 ;
      RECT  10070.0 19387.5 10140.0 19730.0 ;
      RECT  9880.0 20092.5 9950.0 20227.5 ;
      RECT  10070.0 19252.5 10140.0 19387.5 ;
      RECT  10172.5 19695.0 10037.5 19765.0 ;
      RECT  8805.0 19650.0 8875.0 19785.0 ;
      RECT  8945.0 19377.5 9015.0 19512.5 ;
      RECT  9942.5 19480.0 9807.5 19550.0 ;
      RECT  9880.0 21175.0 9950.0 21105.0 ;
      RECT  10070.0 21175.0 10140.0 21105.0 ;
      RECT  9880.0 21140.0 9950.0 20777.5 ;
      RECT  9915.0 21175.0 10105.0 21105.0 ;
      RECT  10070.0 21482.5 10140.0 21140.0 ;
      RECT  9880.0 20777.5 9950.0 20642.5 ;
      RECT  10070.0 21617.5 10140.0 21482.5 ;
      RECT  10172.5 21175.0 10037.5 21105.0 ;
      RECT  8805.0 21085.0 8875.0 21220.0 ;
      RECT  8945.0 21357.5 9015.0 21492.5 ;
      RECT  9942.5 21320.0 9807.5 21390.0 ;
      RECT  9880.0 22385.0 9950.0 22455.0 ;
      RECT  10070.0 22385.0 10140.0 22455.0 ;
      RECT  9880.0 22420.0 9950.0 22782.5 ;
      RECT  9915.0 22385.0 10105.0 22455.0 ;
      RECT  10070.0 22077.5 10140.0 22420.0 ;
      RECT  9880.0 22782.5 9950.0 22917.5 ;
      RECT  10070.0 21942.5 10140.0 22077.5 ;
      RECT  10172.5 22385.0 10037.5 22455.0 ;
      RECT  8805.0 22340.0 8875.0 22475.0 ;
      RECT  8945.0 22067.5 9015.0 22202.5 ;
      RECT  9942.5 22170.0 9807.5 22240.0 ;
      RECT  9880.0 23865.0 9950.0 23795.0 ;
      RECT  10070.0 23865.0 10140.0 23795.0 ;
      RECT  9880.0 23830.0 9950.0 23467.5 ;
      RECT  9915.0 23865.0 10105.0 23795.0 ;
      RECT  10070.0 24172.5 10140.0 23830.0 ;
      RECT  9880.0 23467.5 9950.0 23332.5 ;
      RECT  10070.0 24307.5 10140.0 24172.5 ;
      RECT  10172.5 23865.0 10037.5 23795.0 ;
      RECT  8805.0 23775.0 8875.0 23910.0 ;
      RECT  8945.0 24047.5 9015.0 24182.5 ;
      RECT  9942.5 24010.0 9807.5 24080.0 ;
      RECT  9880.0 25075.0 9950.0 25145.0 ;
      RECT  10070.0 25075.0 10140.0 25145.0 ;
      RECT  9880.0 25110.0 9950.0 25472.5 ;
      RECT  9915.0 25075.0 10105.0 25145.0 ;
      RECT  10070.0 24767.5 10140.0 25110.0 ;
      RECT  9880.0 25472.5 9950.0 25607.5 ;
      RECT  10070.0 24632.5 10140.0 24767.5 ;
      RECT  10172.5 25075.0 10037.5 25145.0 ;
      RECT  8805.0 25030.0 8875.0 25165.0 ;
      RECT  8945.0 24757.5 9015.0 24892.5 ;
      RECT  9942.5 24860.0 9807.5 24930.0 ;
      RECT  9880.0 26555.0 9950.0 26485.0 ;
      RECT  10070.0 26555.0 10140.0 26485.0 ;
      RECT  9880.0 26520.0 9950.0 26157.5 ;
      RECT  9915.0 26555.0 10105.0 26485.0 ;
      RECT  10070.0 26862.5 10140.0 26520.0 ;
      RECT  9880.0 26157.5 9950.0 26022.5 ;
      RECT  10070.0 26997.5 10140.0 26862.5 ;
      RECT  10172.5 26555.0 10037.5 26485.0 ;
      RECT  8805.0 26465.0 8875.0 26600.0 ;
      RECT  8945.0 26737.5 9015.0 26872.5 ;
      RECT  9942.5 26700.0 9807.5 26770.0 ;
      RECT  9880.0 27765.0 9950.0 27835.0 ;
      RECT  10070.0 27765.0 10140.0 27835.0 ;
      RECT  9880.0 27800.0 9950.0 28162.5 ;
      RECT  9915.0 27765.0 10105.0 27835.0 ;
      RECT  10070.0 27457.5 10140.0 27800.0 ;
      RECT  9880.0 28162.5 9950.0 28297.5 ;
      RECT  10070.0 27322.5 10140.0 27457.5 ;
      RECT  10172.5 27765.0 10037.5 27835.0 ;
      RECT  8805.0 27720.0 8875.0 27855.0 ;
      RECT  8945.0 27447.5 9015.0 27582.5 ;
      RECT  9942.5 27550.0 9807.5 27620.0 ;
      RECT  9880.0 29245.0 9950.0 29175.0 ;
      RECT  10070.0 29245.0 10140.0 29175.0 ;
      RECT  9880.0 29210.0 9950.0 28847.5 ;
      RECT  9915.0 29245.0 10105.0 29175.0 ;
      RECT  10070.0 29552.5 10140.0 29210.0 ;
      RECT  9880.0 28847.5 9950.0 28712.5 ;
      RECT  10070.0 29687.5 10140.0 29552.5 ;
      RECT  10172.5 29245.0 10037.5 29175.0 ;
      RECT  8805.0 29155.0 8875.0 29290.0 ;
      RECT  8945.0 29427.5 9015.0 29562.5 ;
      RECT  9942.5 29390.0 9807.5 29460.0 ;
      RECT  9880.0 30455.0 9950.0 30525.0 ;
      RECT  10070.0 30455.0 10140.0 30525.0 ;
      RECT  9880.0 30490.0 9950.0 30852.5 ;
      RECT  9915.0 30455.0 10105.0 30525.0 ;
      RECT  10070.0 30147.5 10140.0 30490.0 ;
      RECT  9880.0 30852.5 9950.0 30987.5 ;
      RECT  10070.0 30012.5 10140.0 30147.5 ;
      RECT  10172.5 30455.0 10037.5 30525.0 ;
      RECT  8805.0 30410.0 8875.0 30545.0 ;
      RECT  8945.0 30137.5 9015.0 30272.5 ;
      RECT  9942.5 30240.0 9807.5 30310.0 ;
      RECT  9880.0 31935.0 9950.0 31865.0 ;
      RECT  10070.0 31935.0 10140.0 31865.0 ;
      RECT  9880.0 31900.0 9950.0 31537.5 ;
      RECT  9915.0 31935.0 10105.0 31865.0 ;
      RECT  10070.0 32242.5 10140.0 31900.0 ;
      RECT  9880.0 31537.5 9950.0 31402.5 ;
      RECT  10070.0 32377.5 10140.0 32242.5 ;
      RECT  10172.5 31935.0 10037.5 31865.0 ;
      RECT  8805.0 31845.0 8875.0 31980.0 ;
      RECT  8945.0 32117.5 9015.0 32252.5 ;
      RECT  9942.5 32080.0 9807.5 32150.0 ;
      RECT  9880.0 33145.0 9950.0 33215.0 ;
      RECT  10070.0 33145.0 10140.0 33215.0 ;
      RECT  9880.0 33180.0 9950.0 33542.5 ;
      RECT  9915.0 33145.0 10105.0 33215.0 ;
      RECT  10070.0 32837.5 10140.0 33180.0 ;
      RECT  9880.0 33542.5 9950.0 33677.5 ;
      RECT  10070.0 32702.5 10140.0 32837.5 ;
      RECT  10172.5 33145.0 10037.5 33215.0 ;
      RECT  8805.0 33100.0 8875.0 33235.0 ;
      RECT  8945.0 32827.5 9015.0 32962.5 ;
      RECT  9942.5 32930.0 9807.5 33000.0 ;
      RECT  9880.0 34625.0 9950.0 34555.0 ;
      RECT  10070.0 34625.0 10140.0 34555.0 ;
      RECT  9880.0 34590.0 9950.0 34227.5 ;
      RECT  9915.0 34625.0 10105.0 34555.0 ;
      RECT  10070.0 34932.5 10140.0 34590.0 ;
      RECT  9880.0 34227.5 9950.0 34092.5 ;
      RECT  10070.0 35067.5 10140.0 34932.5 ;
      RECT  10172.5 34625.0 10037.5 34555.0 ;
      RECT  8805.0 34535.0 8875.0 34670.0 ;
      RECT  8945.0 34807.5 9015.0 34942.5 ;
      RECT  9942.5 34770.0 9807.5 34840.0 ;
      RECT  9880.0 35835.0 9950.0 35905.0 ;
      RECT  10070.0 35835.0 10140.0 35905.0 ;
      RECT  9880.0 35870.0 9950.0 36232.5 ;
      RECT  9915.0 35835.0 10105.0 35905.0 ;
      RECT  10070.0 35527.5 10140.0 35870.0 ;
      RECT  9880.0 36232.5 9950.0 36367.5 ;
      RECT  10070.0 35392.5 10140.0 35527.5 ;
      RECT  10172.5 35835.0 10037.5 35905.0 ;
      RECT  8805.0 35790.0 8875.0 35925.0 ;
      RECT  8945.0 35517.5 9015.0 35652.5 ;
      RECT  9942.5 35620.0 9807.5 35690.0 ;
      RECT  9880.0 37315.0 9950.0 37245.0 ;
      RECT  10070.0 37315.0 10140.0 37245.0 ;
      RECT  9880.0 37280.0 9950.0 36917.5 ;
      RECT  9915.0 37315.0 10105.0 37245.0 ;
      RECT  10070.0 37622.5 10140.0 37280.0 ;
      RECT  9880.0 36917.5 9950.0 36782.5 ;
      RECT  10070.0 37757.5 10140.0 37622.5 ;
      RECT  10172.5 37315.0 10037.5 37245.0 ;
      RECT  8805.0 37225.0 8875.0 37360.0 ;
      RECT  8945.0 37497.5 9015.0 37632.5 ;
      RECT  9942.5 37460.0 9807.5 37530.0 ;
      RECT  9880.0 38525.0 9950.0 38595.0 ;
      RECT  10070.0 38525.0 10140.0 38595.0 ;
      RECT  9880.0 38560.0 9950.0 38922.5 ;
      RECT  9915.0 38525.0 10105.0 38595.0 ;
      RECT  10070.0 38217.5 10140.0 38560.0 ;
      RECT  9880.0 38922.5 9950.0 39057.5 ;
      RECT  10070.0 38082.5 10140.0 38217.5 ;
      RECT  10172.5 38525.0 10037.5 38595.0 ;
      RECT  8805.0 38480.0 8875.0 38615.0 ;
      RECT  8945.0 38207.5 9015.0 38342.5 ;
      RECT  9942.5 38310.0 9807.5 38380.0 ;
      RECT  9880.0 40005.0 9950.0 39935.0 ;
      RECT  10070.0 40005.0 10140.0 39935.0 ;
      RECT  9880.0 39970.0 9950.0 39607.5 ;
      RECT  9915.0 40005.0 10105.0 39935.0 ;
      RECT  10070.0 40312.5 10140.0 39970.0 ;
      RECT  9880.0 39607.5 9950.0 39472.5 ;
      RECT  10070.0 40447.5 10140.0 40312.5 ;
      RECT  10172.5 40005.0 10037.5 39935.0 ;
      RECT  8805.0 39915.0 8875.0 40050.0 ;
      RECT  8945.0 40187.5 9015.0 40322.5 ;
      RECT  9942.5 40150.0 9807.5 40220.0 ;
      RECT  8805.0 19090.0 8875.0 40610.0 ;
      RECT  4655.0 7920.0 11095.0 7215.0 ;
      RECT  4655.0 6510.0 11095.0 7215.0 ;
      RECT  4655.0 6510.0 11095.0 5805.0 ;
      RECT  4655.0 5100.0 11095.0 5805.0 ;
      RECT  4655.0 7602.5 4800.0 7532.5 ;
      RECT  4655.0 6897.5 4800.0 6827.5 ;
      RECT  4655.0 6192.5 4800.0 6122.5 ;
      RECT  4655.0 5487.5 4800.0 5417.5 ;
      RECT  10825.0 7602.5 11095.0 7532.5 ;
      RECT  10407.5 7757.5 11095.0 7687.5 ;
      RECT  10825.0 6897.5 11095.0 6827.5 ;
      RECT  10407.5 6742.5 11095.0 6672.5 ;
      RECT  10825.0 6192.5 11095.0 6122.5 ;
      RECT  10407.5 6347.5 11095.0 6277.5 ;
      RECT  10825.0 5487.5 11095.0 5417.5 ;
      RECT  10407.5 5332.5 11095.0 5262.5 ;
      RECT  4655.0 7955.0 11095.0 7885.0 ;
      RECT  4655.0 7250.0 11095.0 7180.0 ;
      RECT  4655.0 6545.0 11095.0 6475.0 ;
      RECT  4655.0 5840.0 11095.0 5770.0 ;
      RECT  4655.0 5135.0 11095.0 5065.0 ;
      RECT  14627.5 440.0 14697.5 575.0 ;
      RECT  15332.5 440.0 15402.5 575.0 ;
      RECT  14837.5 0.0 14907.5 135.0 ;
      RECT  15542.5 0.0 15612.5 135.0 ;
      RECT  12427.5 19125.0 12562.5 19055.0 ;
      RECT  12427.5 21815.0 12562.5 21745.0 ;
      RECT  12427.5 24505.0 12562.5 24435.0 ;
      RECT  12427.5 27195.0 12562.5 27125.0 ;
      RECT  12427.5 29885.0 12562.5 29815.0 ;
      RECT  12427.5 32575.0 12562.5 32505.0 ;
      RECT  12427.5 35265.0 12562.5 35195.0 ;
      RECT  12427.5 37955.0 12562.5 37885.0 ;
      RECT  12427.5 40645.0 12562.5 40575.0 ;
      RECT  11095.0 8500.0 10960.0 8570.0 ;
      RECT  11505.0 8500.0 11370.0 8570.0 ;
      RECT  10820.0 9845.0 10685.0 9915.0 ;
      RECT  11710.0 9845.0 11575.0 9915.0 ;
      RECT  11095.0 13880.0 10960.0 13950.0 ;
      RECT  11915.0 13880.0 11780.0 13950.0 ;
      RECT  10820.0 15225.0 10685.0 15295.0 ;
      RECT  12120.0 15225.0 11985.0 15295.0 ;
      RECT  11300.0 8295.0 11165.0 8365.0 ;
      RECT  11300.0 8295.0 11165.0 8365.0 ;
      RECT  12360.0 8365.0 12495.0 8295.0 ;
      RECT  11300.0 10985.0 11165.0 11055.0 ;
      RECT  11300.0 10985.0 11165.0 11055.0 ;
      RECT  12360.0 11055.0 12495.0 10985.0 ;
      RECT  11300.0 13675.0 11165.0 13745.0 ;
      RECT  11300.0 13675.0 11165.0 13745.0 ;
      RECT  12360.0 13745.0 12495.0 13675.0 ;
      RECT  11300.0 16365.0 11165.0 16435.0 ;
      RECT  11300.0 16365.0 11165.0 16435.0 ;
      RECT  12360.0 16435.0 12495.0 16365.0 ;
      RECT  11162.5 7532.5 11027.5 7602.5 ;
      RECT  11505.0 7532.5 11370.0 7602.5 ;
      RECT  11162.5 6827.5 11027.5 6897.5 ;
      RECT  11710.0 6827.5 11575.0 6897.5 ;
      RECT  11162.5 6122.5 11027.5 6192.5 ;
      RECT  11915.0 6122.5 11780.0 6192.5 ;
      RECT  11162.5 5417.5 11027.5 5487.5 ;
      RECT  12120.0 5417.5 11985.0 5487.5 ;
      RECT  11230.0 7885.0 11095.0 7955.0 ;
      RECT  12562.5 7885.0 12427.5 7955.0 ;
      RECT  11230.0 7180.0 11095.0 7250.0 ;
      RECT  12562.5 7180.0 12427.5 7250.0 ;
      RECT  11230.0 6475.0 11095.0 6545.0 ;
      RECT  12562.5 6475.0 12427.5 6545.0 ;
      RECT  11230.0 5770.0 11095.0 5840.0 ;
      RECT  12562.5 5770.0 12427.5 5840.0 ;
      RECT  11230.0 5065.0 11095.0 5135.0 ;
      RECT  12562.5 5065.0 12427.5 5135.0 ;
      RECT  13700.0 3792.5 13565.0 3862.5 ;
      RECT  13290.0 1607.5 13155.0 1677.5 ;
      RECT  13495.0 3155.0 13360.0 3225.0 ;
      RECT  13700.0 41585.0 13565.0 41655.0 ;
      RECT  13905.0 10295.0 13770.0 10365.0 ;
      RECT  14110.0 14320.0 13975.0 14390.0 ;
      RECT  13085.0 8090.0 12950.0 8160.0 ;
      RECT  8907.5 40780.0 8772.5 40850.0 ;
      RECT  13085.0 40780.0 12950.0 40850.0 ;
      RECT  12777.5 3025.0 12642.5 3095.0 ;
      RECT  12777.5 14450.0 12642.5 14520.0 ;
      RECT  12777.5 3952.5 12642.5 4022.5 ;
      RECT  12777.5 11227.5 12642.5 11297.5 ;
      RECT  14837.5 0.0 14907.5 140.0 ;
      RECT  15542.5 0.0 15612.5 140.0 ;
      RECT  14007.5 0.0 14077.5 42337.5 ;
      RECT  13802.5 0.0 13872.5 42337.5 ;
      RECT  13187.5 0.0 13257.5 42337.5 ;
      RECT  13392.5 0.0 13462.5 42337.5 ;
      RECT  13597.5 0.0 13667.5 42337.5 ;
      RECT  12982.5 0.0 13052.5 42337.5 ;
      RECT  12427.5 0.0 12777.5 42337.5 ;
      RECT  4035.0 26490.0 8.881784197e-13 26560.0 ;
      RECT  4035.0 26695.0 8.881784197e-13 26765.0 ;
      RECT  4035.0 26900.0 8.881784197e-13 26970.0 ;
      RECT  4035.0 27310.0 8.881784197e-13 27380.0 ;
      RECT  3422.5 22000.0 2690.0 22070.0 ;
      RECT  2520.0 19467.5 2450.0 26115.0 ;
      RECT  4035.0 26285.0 3830.0 26355.0 ;
      RECT  2895.0 27105.0 2690.0 27175.0 ;
      RECT  1550.0 26285.0 1345.0 26355.0 ;
      RECT  205.0 27105.0 8.881784197e-13 27175.0 ;
      RECT  165.0 19230.0 870.0 25670.0 ;
      RECT  1575.0 19230.0 870.0 25670.0 ;
      RECT  1575.0 19230.0 2280.0 25670.0 ;
      RECT  482.5 19230.0 552.5 19375.0 ;
      RECT  1187.5 19230.0 1257.5 19375.0 ;
      RECT  1892.5 19230.0 1962.5 19375.0 ;
      RECT  482.5 25400.0 552.5 25670.0 ;
      RECT  327.5 24982.5 397.5 25670.0 ;
      RECT  1187.5 25400.0 1257.5 25670.0 ;
      RECT  1342.5 24982.5 1412.5 25670.0 ;
      RECT  1892.5 25400.0 1962.5 25670.0 ;
      RECT  1737.5 24982.5 1807.5 25670.0 ;
      RECT  130.0 19230.0 200.0 25670.0 ;
      RECT  835.0 19230.0 905.0 25670.0 ;
      RECT  1540.0 19230.0 1610.0 25670.0 ;
      RECT  2245.0 19230.0 2315.0 25670.0 ;
      RECT  3737.5 28560.0 3032.5 28630.0 ;
      RECT  3382.5 28180.0 3312.5 28250.0 ;
      RECT  3382.5 28560.0 3312.5 28630.0 ;
      RECT  3347.5 28180.0 3032.5 28250.0 ;
      RECT  3382.5 28215.0 3312.5 28595.0 ;
      RECT  3737.5 28560.0 3347.5 28630.0 ;
      RECT  3032.5 28180.0 2897.5 28250.0 ;
      RECT  3032.5 28560.0 2897.5 28630.0 ;
      RECT  3872.5 28560.0 3737.5 28630.0 ;
      RECT  3415.0 28560.0 3280.0 28630.0 ;
      RECT  1895.0 28370.0 1965.0 28440.0 ;
      RECT  1930.0 28370.0 2280.0 28440.0 ;
      RECT  1895.0 28405.0 1965.0 28475.0 ;
      RECT  1495.0 28370.0 1565.0 28440.0 ;
      RECT  1495.0 28247.5 1565.0 28405.0 ;
      RECT  1530.0 28370.0 1930.0 28440.0 ;
      RECT  2280.0 28370.0 2415.0 28440.0 ;
      RECT  1495.0 28282.5 1565.0 28147.5 ;
      RECT  1895.0 28542.5 1965.0 28407.5 ;
      RECT  1950.0 29325.0 2020.0 29395.0 ;
      RECT  1950.0 29515.0 2020.0 29585.0 ;
      RECT  1985.0 29325.0 2347.5 29395.0 ;
      RECT  1950.0 29360.0 2020.0 29550.0 ;
      RECT  1642.5 29515.0 1985.0 29585.0 ;
      RECT  2347.5 29325.0 2482.5 29395.0 ;
      RECT  1507.5 29515.0 1642.5 29585.0 ;
      RECT  1950.0 29617.5 2020.0 29482.5 ;
      RECT  1047.5 29120.0 342.5 29190.0 ;
      RECT  692.5 28740.0 622.5 28810.0 ;
      RECT  692.5 29120.0 622.5 29190.0 ;
      RECT  657.5 28740.0 342.5 28810.0 ;
      RECT  692.5 28775.0 622.5 29155.0 ;
      RECT  1047.5 29120.0 657.5 29190.0 ;
      RECT  342.5 28740.0 207.5 28810.0 ;
      RECT  342.5 29120.0 207.5 29190.0 ;
      RECT  1182.5 29120.0 1047.5 29190.0 ;
      RECT  725.0 29120.0 590.0 29190.0 ;
      RECT  397.5 25737.5 327.5 25602.5 ;
      RECT  397.5 27412.5 327.5 27277.5 ;
      RECT  552.5 25737.5 482.5 25602.5 ;
      RECT  552.5 26592.5 482.5 26457.5 ;
      RECT  1412.5 25737.5 1342.5 25602.5 ;
      RECT  1412.5 26797.5 1342.5 26662.5 ;
      RECT  1807.5 25737.5 1737.5 25602.5 ;
      RECT  1807.5 27002.5 1737.5 26867.5 ;
      RECT  200.0 25737.5 130.0 25602.5 ;
      RECT  200.0 26387.5 130.0 26252.5 ;
      RECT  905.0 25737.5 835.0 25602.5 ;
      RECT  905.0 26387.5 835.0 26252.5 ;
      RECT  1610.0 25737.5 1540.0 25602.5 ;
      RECT  1610.0 26387.5 1540.0 26252.5 ;
      RECT  2315.0 25737.5 2245.0 25602.5 ;
      RECT  2315.0 26387.5 2245.0 26252.5 ;
      RECT  1380.0 31895.0 1310.0 36955.0 ;
      RECT  970.0 31895.0 900.0 36645.0 ;
      RECT  265.0 31895.0 195.0 36645.0 ;
      RECT  1207.5 32062.5 1137.5 32660.0 ;
      RECT  785.0 32062.5 715.0 32342.5 ;
      RECT  3372.5 34457.5 3442.5 34852.5 ;
      RECT  2655.0 34982.5 2725.0 35052.5 ;
      RECT  2655.0 35062.5 2725.0 35132.5 ;
      RECT  2690.0 34982.5 3407.5 35052.5 ;
      RECT  2655.0 35017.5 2725.0 35097.5 ;
      RECT  1972.5 35062.5 2690.0 35132.5 ;
      RECT  1937.5 34537.5 2007.5 34932.5 ;
      RECT  3340.0 34817.5 3475.0 34887.5 ;
      RECT  1905.0 35062.5 2040.0 35132.5 ;
      RECT  1905.0 34502.5 2040.0 34572.5 ;
      RECT  3340.0 34422.5 3475.0 34492.5 ;
      RECT  3340.0 34982.5 3475.0 35052.5 ;
      RECT  1905.0 34897.5 2040.0 34967.5 ;
      RECT  935.0 33800.0 225.0 32455.0 ;
      RECT  935.0 33800.0 230.0 35145.0 ;
      RECT  935.0 36490.0 230.0 35145.0 ;
      RECT  785.0 33700.0 715.0 36645.0 ;
      RECT  450.0 33700.0 380.0 36645.0 ;
      RECT  970.0 33700.0 900.0 36645.0 ;
      RECT  265.0 33700.0 195.0 36645.0 ;
      RECT  1347.5 33872.5 1277.5 34007.5 ;
      RECT  1347.5 36282.5 1277.5 36417.5 ;
      RECT  1345.0 34135.0 1275.0 34270.0 ;
      RECT  1380.0 31760.0 1310.0 31895.0 ;
      RECT  867.5 31860.0 1002.5 31930.0 ;
      RECT  162.5 31860.0 297.5 31930.0 ;
      RECT  1105.0 32625.0 1240.0 32695.0 ;
      RECT  1105.0 32027.5 1240.0 32097.5 ;
      RECT  682.5 32027.5 817.5 32097.5 ;
      RECT  3457.5 26182.5 3387.5 26047.5 ;
      RECT  3457.5 22102.5 3387.5 21967.5 ;
      RECT  2725.0 22102.5 2655.0 21967.5 ;
      RECT  2725.0 27617.5 2655.0 27482.5 ;
      RECT  2520.0 19535.0 2450.0 19400.0 ;
      RECT  1965.0 26182.5 1895.0 26047.5 ;
      RECT  1750.0 26592.5 1680.0 26457.5 ;
      RECT  2020.0 29130.0 1950.0 28995.0 ;
      RECT  2020.0 29130.0 1950.0 28995.0 ;
      RECT  2020.0 27617.5 1950.0 27482.5 ;
      RECT  1805.0 29387.5 1735.0 29252.5 ;
      RECT  1805.0 29387.5 1735.0 29252.5 ;
      RECT  1805.0 27412.5 1735.0 27277.5 ;
      RECT  3382.5 27617.5 3312.5 27482.5 ;
      RECT  3522.5 27412.5 3452.5 27277.5 ;
      RECT  3662.5 26797.5 3592.5 26662.5 ;
      RECT  692.5 27617.5 622.5 27482.5 ;
      RECT  832.5 26797.5 762.5 26662.5 ;
      RECT  972.5 27002.5 902.5 26867.5 ;
      RECT  1997.5 28810.0 1862.5 28880.0 ;
      RECT  2052.5 29955.0 1917.5 30025.0 ;
      RECT  785.0 31140.0 650.0 31210.0 ;
      RECT  2040.0 30180.0 1905.0 30250.0 ;
      RECT  4070.0 26387.5 4000.0 26252.5 ;
      RECT  2725.0 27207.5 2655.0 27072.5 ;
      RECT  1380.0 26387.5 1310.0 26252.5 ;
      RECT  35.0 27207.5 -35.0 27072.5 ;
      RECT  4035.0 30180.0 1972.5 30250.0 ;
      RECT  4035.0 31140.0 717.5 31210.0 ;
      RECT  4035.0 28810.0 1930.0 28880.0 ;
      RECT  4035.0 29955.0 1985.0 30025.0 ;
      RECT  4035.0 27515.0 8.881784197e-13 27585.0 ;
      RECT  4035.0 26080.0 0.0 26150.0 ;
      RECT  4035.0 27105.0 8.881784197e-13 27175.0 ;
      RECT  4035.0 26285.0 0.0 26355.0 ;
      RECT  14110.0 30180.0 13975.0 30250.0 ;
      RECT  4035.0 30180.0 3900.0 30250.0 ;
      RECT  13905.0 31140.0 13770.0 31210.0 ;
      RECT  4035.0 31140.0 3900.0 31210.0 ;
      RECT  13495.0 28810.0 13360.0 28880.0 ;
      RECT  4035.0 28810.0 3900.0 28880.0 ;
      RECT  13290.0 29955.0 13155.0 30025.0 ;
      RECT  4035.0 29955.0 3900.0 30025.0 ;
      RECT  13700.0 27515.0 13565.0 27585.0 ;
      RECT  4035.0 27515.0 3900.0 27585.0 ;
      RECT  13085.0 26080.0 12950.0 26150.0 ;
      RECT  4035.0 26080.0 3900.0 26150.0 ;
      RECT  4417.5 27105.0 4282.5 27175.0 ;
      RECT  12670.0 26285.0 12535.0 26355.0 ;
      RECT  4035.0 26285.0 3900.0 26355.0 ;
   LAYER  metal3 ;
      RECT  4035.0 30180.0 14042.5 30250.0 ;
      RECT  4035.0 31140.0 13837.5 31210.0 ;
      RECT  4035.0 28810.0 13427.5 28880.0 ;
      RECT  4035.0 29955.0 13222.5 30025.0 ;
      RECT  4035.0 27515.0 13632.5 27585.0 ;
      RECT  4035.0 26080.0 13017.5 26150.0 ;
      RECT  4035.0 26285.0 12602.5 26355.0 ;
      RECT  14627.5 18985.0 14697.5 19055.0 ;
      RECT  14627.5 475.0 14697.5 19020.0 ;
      RECT  14662.5 18985.0 14832.5 19055.0 ;
      RECT  15332.5 18985.0 15402.5 19055.0 ;
      RECT  15332.5 475.0 15402.5 19020.0 ;
      RECT  15367.5 18985.0 15537.5 19055.0 ;
      RECT  14837.5 0.0 14907.5 3590.0 ;
      RECT  15542.5 0.0 15612.5 3590.0 ;
      RECT  11232.5 8295.0 12427.5 8365.0 ;
      RECT  11232.5 10985.0 12427.5 11055.0 ;
      RECT  11232.5 13675.0 12427.5 13745.0 ;
      RECT  11232.5 16365.0 12427.5 16435.0 ;
      RECT  14832.5 18950.0 14902.5 19090.0 ;
      RECT  15537.5 18950.0 15607.5 19090.0 ;
      RECT  14837.5 3590.0 14907.5 3730.0 ;
      RECT  15542.5 3590.0 15612.5 3730.0 ;
      RECT  4655.0 7602.5 4795.0 7532.5 ;
      RECT  4655.0 6897.5 4795.0 6827.5 ;
      RECT  4655.0 6192.5 4795.0 6122.5 ;
      RECT  4655.0 5487.5 4795.0 5417.5 ;
      RECT  14627.5 440.0 14697.5 575.0 ;
      RECT  15332.5 440.0 15402.5 575.0 ;
      RECT  14837.5 0.0 14907.5 135.0 ;
      RECT  15542.5 0.0 15612.5 135.0 ;
      RECT  11300.0 8295.0 11165.0 8365.0 ;
      RECT  12360.0 8365.0 12495.0 8295.0 ;
      RECT  11300.0 10985.0 11165.0 11055.0 ;
      RECT  12360.0 11055.0 12495.0 10985.0 ;
      RECT  11300.0 13675.0 11165.0 13745.0 ;
      RECT  12360.0 13745.0 12495.0 13675.0 ;
      RECT  11300.0 16365.0 11165.0 16435.0 ;
      RECT  12360.0 16435.0 12495.0 16365.0 ;
      RECT  4175.0 7532.5 4655.0 7602.5 ;
      RECT  4175.0 6827.5 4655.0 6897.5 ;
      RECT  4175.0 6122.5 4655.0 6192.5 ;
      RECT  4175.0 5417.5 4655.0 5487.5 ;
      RECT  397.5 25670.0 327.5 27345.0 ;
      RECT  552.5 25670.0 482.5 26525.0 ;
      RECT  1412.5 25670.0 1342.5 26730.0 ;
      RECT  1807.5 25670.0 1737.5 26935.0 ;
      RECT  200.0 25670.0 130.0 26320.0 ;
      RECT  905.0 25670.0 835.0 26320.0 ;
      RECT  1610.0 25670.0 1540.0 26320.0 ;
      RECT  2315.0 25670.0 2245.0 26320.0 ;
      RECT  2725.0 22035.0 2655.0 27550.0 ;
      RECT  2020.0 27550.0 1950.0 29062.5 ;
      RECT  1805.0 27345.0 1735.0 29320.0 ;
      RECT  482.5 19230.0 552.5 19370.0 ;
      RECT  1187.5 19230.0 1257.5 19370.0 ;
      RECT  1892.5 19230.0 1962.5 19370.0 ;
      RECT  397.5 25737.5 327.5 25602.5 ;
      RECT  397.5 27412.5 327.5 27277.5 ;
      RECT  552.5 25737.5 482.5 25602.5 ;
      RECT  552.5 26592.5 482.5 26457.5 ;
      RECT  1412.5 25737.5 1342.5 25602.5 ;
      RECT  1412.5 26797.5 1342.5 26662.5 ;
      RECT  1807.5 25737.5 1737.5 25602.5 ;
      RECT  1807.5 27002.5 1737.5 26867.5 ;
      RECT  200.0 25737.5 130.0 25602.5 ;
      RECT  200.0 26387.5 130.0 26252.5 ;
      RECT  905.0 25737.5 835.0 25602.5 ;
      RECT  905.0 26387.5 835.0 26252.5 ;
      RECT  1610.0 25737.5 1540.0 25602.5 ;
      RECT  1610.0 26387.5 1540.0 26252.5 ;
      RECT  2315.0 25737.5 2245.0 25602.5 ;
      RECT  2315.0 26387.5 2245.0 26252.5 ;
      RECT  2725.0 22102.5 2655.0 21967.5 ;
      RECT  2725.0 27617.5 2655.0 27482.5 ;
      RECT  2020.0 29130.0 1950.0 28995.0 ;
      RECT  2020.0 27617.5 1950.0 27482.5 ;
      RECT  1805.0 29387.5 1735.0 29252.5 ;
      RECT  1805.0 27412.5 1735.0 27277.5 ;
      RECT  1257.5 19230.0 1187.5 19370.0 ;
      RECT  1962.5 19230.0 1892.5 19370.0 ;
      RECT  552.5 19230.0 482.5 19370.0 ;
      RECT  14110.0 30180.0 13975.0 30250.0 ;
      RECT  4035.0 30180.0 3900.0 30250.0 ;
      RECT  13905.0 31140.0 13770.0 31210.0 ;
      RECT  4035.0 31140.0 3900.0 31210.0 ;
      RECT  13495.0 28810.0 13360.0 28880.0 ;
      RECT  4035.0 28810.0 3900.0 28880.0 ;
      RECT  13290.0 29955.0 13155.0 30025.0 ;
      RECT  4035.0 29955.0 3900.0 30025.0 ;
      RECT  13700.0 27515.0 13565.0 27585.0 ;
      RECT  4035.0 27515.0 3900.0 27585.0 ;
      RECT  13085.0 26080.0 12950.0 26150.0 ;
      RECT  4035.0 26080.0 3900.0 26150.0 ;
      RECT  12670.0 26285.0 12535.0 26355.0 ;
      RECT  4035.0 26285.0 3900.0 26355.0 ;
   END
   END    sram_2_16_1_freepdk45
END    LIBRARY
