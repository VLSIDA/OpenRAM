MACRO sram_2_16_1_scn3me_subm
    CLASS RING ;
    ORIGIN 53.7 0.0 ;
    FOREIGN  sram 0.0 0.0 ;
    SIZE 201.0 BY 444.3 ;
    SYMMETRY X Y R90 ;
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  143.4 0.0 147.9 444.3 ;
        RECT  143.4 0.0 147.9 444.3 ;
        RECT  0.0 0.0 4.5 444.3 ;
        RECT  0.0 0.0 4.5 444.3 ;
        END
    END vdd
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal2 ;
        RECT  92.85 0.0 97.35 444.3 ;
        RECT  92.85 0.0 97.35 444.3 ;
        END
    END gnd
    PIN DATA[0]
        DIRECTION INOUT ;
        PORT
        LAYER metal2 ;
        RECT  124.8 0.0 125.7 1.8 ;
        RECT  124.8 0.0 125.7 1.8 ;
        END
    END DATA[0]
    PIN DATA[1]
        DIRECTION INOUT ;
        PORT
        LAYER metal2 ;
        RECT  135.0 0.0 135.9 1.8 ;
        RECT  135.0 0.0 135.9 1.8 ;
        END
    END DATA[1]
    PIN ADDR[0]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 75.0 7.2 76.5 ;
        RECT  0.0 75.0 7.2 76.5 ;
        END
    END ADDR[0]
    PIN ADDR[1]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 64.8 7.2 66.3 ;
        RECT  0.0 64.8 7.2 66.3 ;
        END
    END ADDR[1]
    PIN ADDR[2]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 54.6 7.2 56.1 ;
        RECT  0.0 54.6 7.2 56.1 ;
        END
    END ADDR[2]
    PIN ADDR[3]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 44.4 7.2 45.9 ;
        RECT  0.0 44.4 7.2 45.9 ;
        END
    END ADDR[3]
    PIN CSb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        END
    END CSb
    PIN OEb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        END
    END OEb
    PIN WEb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        END
    END WEb
    PIN clk
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -9.9 202.2 -9.0 203.1 ;
        RECT  -9.9 202.2 -9.0 203.1 ;
        RECT  -9.9 202.2 -9.0 204.3 ;
        END
    END clk
    OBS
        LAYER  metal1 ;
        RECT  1.8 316.95 2.7 319.65 ;
        RECT  -9.9 202.2 -9.0 203.1 ;
        RECT  143.4 0.0 147.9 444.3 ;
        RECT  0.0 0.0 4.5 444.3 ;
        RECT  44.7 205.2 45.6 206.1 ;
        RECT  44.7 207.3 45.6 208.2 ;
        RECT  40.5 205.2 45.15 206.1 ;
        RECT  44.7 205.65 45.6 207.75 ;
        RECT  45.15 207.3 49.8 208.2 ;
        RECT  83.85 205.2 84.75 206.1 ;
        RECT  83.85 201.45 84.75 202.35 ;
        RECT  82.2 205.2 84.3 206.1 ;
        RECT  83.85 201.9 84.75 205.65 ;
        RECT  84.3 201.45 119.7 202.35 ;
        RECT  44.7 220.5 45.6 221.4 ;
        RECT  44.7 218.4 45.6 219.3 ;
        RECT  40.5 220.5 45.15 221.4 ;
        RECT  44.7 218.85 45.6 220.95 ;
        RECT  45.15 218.4 49.8 219.3 ;
        RECT  83.85 220.5 84.75 221.4 ;
        RECT  83.85 224.25 84.75 225.15 ;
        RECT  82.2 220.5 84.3 221.4 ;
        RECT  83.85 220.95 84.75 224.7 ;
        RECT  84.3 224.25 119.7 225.15 ;
        RECT  44.7 233.4 45.6 234.3 ;
        RECT  44.7 235.5 45.6 236.4 ;
        RECT  40.5 233.4 45.15 234.3 ;
        RECT  44.7 233.85 45.6 235.95 ;
        RECT  45.15 235.5 49.8 236.4 ;
        RECT  83.85 233.4 84.75 234.3 ;
        RECT  83.85 229.65 84.75 230.55 ;
        RECT  82.2 233.4 84.3 234.3 ;
        RECT  83.85 230.1 84.75 233.85 ;
        RECT  84.3 229.65 119.7 230.55 ;
        RECT  44.7 248.7 45.6 249.6 ;
        RECT  44.7 246.6 45.6 247.5 ;
        RECT  40.5 248.7 45.15 249.6 ;
        RECT  44.7 247.05 45.6 249.15 ;
        RECT  45.15 246.6 49.8 247.5 ;
        RECT  83.85 248.7 84.75 249.6 ;
        RECT  83.85 252.45 84.75 253.35 ;
        RECT  82.2 248.7 84.3 249.6 ;
        RECT  83.85 249.15 84.75 252.9 ;
        RECT  84.3 252.45 119.7 253.35 ;
        RECT  44.7 261.6 45.6 262.5 ;
        RECT  44.7 263.7 45.6 264.6 ;
        RECT  40.5 261.6 45.15 262.5 ;
        RECT  44.7 262.05 45.6 264.15 ;
        RECT  45.15 263.7 49.8 264.6 ;
        RECT  83.85 261.6 84.75 262.5 ;
        RECT  83.85 257.85 84.75 258.75 ;
        RECT  82.2 261.6 84.3 262.5 ;
        RECT  83.85 258.3 84.75 262.05 ;
        RECT  84.3 257.85 119.7 258.75 ;
        RECT  44.7 276.9 45.6 277.8 ;
        RECT  44.7 274.8 45.6 275.7 ;
        RECT  40.5 276.9 45.15 277.8 ;
        RECT  44.7 275.25 45.6 277.35 ;
        RECT  45.15 274.8 49.8 275.7 ;
        RECT  83.85 276.9 84.75 277.8 ;
        RECT  83.85 280.65 84.75 281.55 ;
        RECT  82.2 276.9 84.3 277.8 ;
        RECT  83.85 277.35 84.75 281.1 ;
        RECT  84.3 280.65 119.7 281.55 ;
        RECT  44.7 289.8 45.6 290.7 ;
        RECT  44.7 291.9 45.6 292.8 ;
        RECT  40.5 289.8 45.15 290.7 ;
        RECT  44.7 290.25 45.6 292.35 ;
        RECT  45.15 291.9 49.8 292.8 ;
        RECT  83.85 289.8 84.75 290.7 ;
        RECT  83.85 286.05 84.75 286.95 ;
        RECT  82.2 289.8 84.3 290.7 ;
        RECT  83.85 286.5 84.75 290.25 ;
        RECT  84.3 286.05 119.7 286.95 ;
        RECT  44.7 305.1 45.6 306.0 ;
        RECT  44.7 303.0 45.6 303.9 ;
        RECT  40.5 305.1 45.15 306.0 ;
        RECT  44.7 303.45 45.6 305.55 ;
        RECT  45.15 303.0 49.8 303.9 ;
        RECT  83.85 305.1 84.75 306.0 ;
        RECT  83.85 308.85 84.75 309.75 ;
        RECT  82.2 305.1 84.3 306.0 ;
        RECT  83.85 305.55 84.75 309.3 ;
        RECT  84.3 308.85 119.7 309.75 ;
        RECT  44.7 318.0 45.6 318.9 ;
        RECT  44.7 320.1 45.6 321.0 ;
        RECT  40.5 318.0 45.15 318.9 ;
        RECT  44.7 318.45 45.6 320.55 ;
        RECT  45.15 320.1 49.8 321.0 ;
        RECT  83.85 318.0 84.75 318.9 ;
        RECT  83.85 314.25 84.75 315.15 ;
        RECT  82.2 318.0 84.3 318.9 ;
        RECT  83.85 314.7 84.75 318.45 ;
        RECT  84.3 314.25 119.7 315.15 ;
        RECT  44.7 333.3 45.6 334.2 ;
        RECT  44.7 331.2 45.6 332.1 ;
        RECT  40.5 333.3 45.15 334.2 ;
        RECT  44.7 331.65 45.6 333.75 ;
        RECT  45.15 331.2 49.8 332.1 ;
        RECT  83.85 333.3 84.75 334.2 ;
        RECT  83.85 337.05 84.75 337.95 ;
        RECT  82.2 333.3 84.3 334.2 ;
        RECT  83.85 333.75 84.75 337.5 ;
        RECT  84.3 337.05 119.7 337.95 ;
        RECT  44.7 346.2 45.6 347.1 ;
        RECT  44.7 348.3 45.6 349.2 ;
        RECT  40.5 346.2 45.15 347.1 ;
        RECT  44.7 346.65 45.6 348.75 ;
        RECT  45.15 348.3 49.8 349.2 ;
        RECT  83.85 346.2 84.75 347.1 ;
        RECT  83.85 342.45 84.75 343.35 ;
        RECT  82.2 346.2 84.3 347.1 ;
        RECT  83.85 342.9 84.75 346.65 ;
        RECT  84.3 342.45 119.7 343.35 ;
        RECT  44.7 361.5 45.6 362.4 ;
        RECT  44.7 359.4 45.6 360.3 ;
        RECT  40.5 361.5 45.15 362.4 ;
        RECT  44.7 359.85 45.6 361.95 ;
        RECT  45.15 359.4 49.8 360.3 ;
        RECT  83.85 361.5 84.75 362.4 ;
        RECT  83.85 365.25 84.75 366.15 ;
        RECT  82.2 361.5 84.3 362.4 ;
        RECT  83.85 361.95 84.75 365.7 ;
        RECT  84.3 365.25 119.7 366.15 ;
        RECT  44.7 374.4 45.6 375.3 ;
        RECT  44.7 376.5 45.6 377.4 ;
        RECT  40.5 374.4 45.15 375.3 ;
        RECT  44.7 374.85 45.6 376.95 ;
        RECT  45.15 376.5 49.8 377.4 ;
        RECT  83.85 374.4 84.75 375.3 ;
        RECT  83.85 370.65 84.75 371.55 ;
        RECT  82.2 374.4 84.3 375.3 ;
        RECT  83.85 371.1 84.75 374.85 ;
        RECT  84.3 370.65 119.7 371.55 ;
        RECT  44.7 389.7 45.6 390.6 ;
        RECT  44.7 387.6 45.6 388.5 ;
        RECT  40.5 389.7 45.15 390.6 ;
        RECT  44.7 388.05 45.6 390.15 ;
        RECT  45.15 387.6 49.8 388.5 ;
        RECT  83.85 389.7 84.75 390.6 ;
        RECT  83.85 393.45 84.75 394.35 ;
        RECT  82.2 389.7 84.3 390.6 ;
        RECT  83.85 390.15 84.75 393.9 ;
        RECT  84.3 393.45 119.7 394.35 ;
        RECT  44.7 402.6 45.6 403.5 ;
        RECT  44.7 404.7 45.6 405.6 ;
        RECT  40.5 402.6 45.15 403.5 ;
        RECT  44.7 403.05 45.6 405.15 ;
        RECT  45.15 404.7 49.8 405.6 ;
        RECT  83.85 402.6 84.75 403.5 ;
        RECT  83.85 398.85 84.75 399.75 ;
        RECT  82.2 402.6 84.3 403.5 ;
        RECT  83.85 399.3 84.75 403.05 ;
        RECT  84.3 398.85 119.7 399.75 ;
        RECT  44.7 417.9 45.6 418.8 ;
        RECT  44.7 415.8 45.6 416.7 ;
        RECT  40.5 417.9 45.15 418.8 ;
        RECT  44.7 416.25 45.6 418.35 ;
        RECT  45.15 415.8 49.8 416.7 ;
        RECT  83.85 417.9 84.75 418.8 ;
        RECT  83.85 421.65 84.75 422.55 ;
        RECT  82.2 417.9 84.3 418.8 ;
        RECT  83.85 418.35 84.75 422.1 ;
        RECT  84.3 421.65 119.7 422.55 ;
        RECT  51.0 198.75 120.3 199.65 ;
        RECT  51.0 226.95 120.3 227.85 ;
        RECT  51.0 255.15 120.3 256.05 ;
        RECT  51.0 283.35 120.3 284.25 ;
        RECT  51.0 311.55 120.3 312.45 ;
        RECT  51.0 339.75 120.3 340.65 ;
        RECT  51.0 367.95 120.3 368.85 ;
        RECT  51.0 396.15 120.3 397.05 ;
        RECT  51.0 424.35 120.3 425.25 ;
        RECT  0.0 212.85 147.9 213.75 ;
        RECT  0.0 241.05 147.9 241.95 ;
        RECT  0.0 269.25 147.9 270.15 ;
        RECT  0.0 297.45 147.9 298.35 ;
        RECT  0.0 325.65 147.9 326.55 ;
        RECT  0.0 353.85 147.9 354.75 ;
        RECT  0.0 382.05 147.9 382.95 ;
        RECT  0.0 410.25 147.9 411.15 ;
        RECT  75.3 88.65 80.25 89.55 ;
        RECT  72.3 102.75 82.95 103.65 ;
        RECT  75.3 145.05 85.65 145.95 ;
        RECT  72.3 159.15 88.35 160.05 ;
        RECT  75.3 85.95 76.8 86.85 ;
        RECT  75.3 114.15 76.8 115.05 ;
        RECT  75.3 142.35 76.8 143.25 ;
        RECT  75.3 170.55 76.8 171.45 ;
        RECT  0.0 100.05 75.3 100.95 ;
        RECT  0.0 128.25 75.3 129.15 ;
        RECT  0.0 156.45 75.3 157.35 ;
        RECT  0.0 184.65 75.3 185.55 ;
        RECT  66.3 75.45 80.25 76.35 ;
        RECT  66.3 65.25 82.95 66.15 ;
        RECT  66.3 55.05 85.65 55.95 ;
        RECT  66.3 44.85 88.35 45.75 ;
        RECT  66.3 70.35 94.05 71.25 ;
        RECT  66.3 49.95 94.05 50.85 ;
        RECT  62.7 37.65 63.6 38.55 ;
        RECT  62.7 38.1 63.6 40.2 ;
        RECT  0.0 37.65 63.15 38.55 ;
        RECT  108.6 32.4 120.3 33.3 ;
        RECT  103.2 27.9 120.3 28.8 ;
        RECT  105.9 25.5 120.3 26.4 ;
        RECT  108.6 431.4 120.3 432.3 ;
        RECT  111.3 96.9 120.3 97.8 ;
        RECT  114.0 195.0 120.3 195.9 ;
        RECT  8.7 82.65 9.6 83.55 ;
        RECT  8.7 81.0 9.6 83.1 ;
        RECT  9.15 82.65 100.95 83.55 ;
        RECT  47.85 426.45 100.95 427.35 ;
        RECT  120.3 443.4 143.4 444.3 ;
        RECT  120.3 167.7 143.4 168.6 ;
        RECT  120.3 99.0 143.4 99.9 ;
        RECT  120.3 86.4 143.4 87.3 ;
        RECT  120.3 9.6 143.4 10.5 ;
        RECT  97.35 23.4 120.3 24.3 ;
        RECT  97.35 192.9 120.3 193.8 ;
        RECT  97.35 94.8 120.3 95.7 ;
        RECT  143.4 0.0 147.9 444.3 ;
        RECT  0.0 0.0 4.5 444.3 ;
        RECT  119.7 257.7 141.3 258.9 ;
        RECT  119.7 201.3 141.3 202.5 ;
        RECT  119.7 229.5 141.3 230.7 ;
        RECT  119.7 421.5 141.3 422.7 ;
        RECT  119.7 314.1 141.3 315.3 ;
        RECT  119.7 285.9 141.3 287.1 ;
        RECT  119.7 393.3 141.3 394.5 ;
        RECT  119.7 365.1 141.3 366.3 ;
        RECT  119.7 252.3 141.3 253.5 ;
        RECT  119.7 280.5 141.3 281.7 ;
        RECT  119.7 224.1 141.3 225.3 ;
        RECT  119.7 398.7 141.3 399.9 ;
        RECT  119.7 342.3 141.3 343.5 ;
        RECT  119.7 336.9 141.3 338.1 ;
        RECT  119.7 212.7 141.3 213.6 ;
        RECT  119.7 240.9 141.3 241.8 ;
        RECT  119.7 269.1 141.3 270.0 ;
        RECT  119.7 297.3 141.3 298.2 ;
        RECT  119.7 325.5 141.3 326.4 ;
        RECT  119.7 353.7 141.3 354.6 ;
        RECT  119.7 381.9 141.3 382.8 ;
        RECT  119.7 410.1 141.3 411.0 ;
        RECT  119.7 370.5 141.3 371.7 ;
        RECT  119.7 308.7 141.3 309.9 ;
        RECT  126.0 199.2 128.7 200.4 ;
        RECT  121.8 199.2 124.5 200.4 ;
        RECT  119.7 201.3 131.1 202.5 ;
        RECT  125.4 202.5 126.6 202.8 ;
        RECT  129.9 204.0 131.1 209.7 ;
        RECT  127.5 204.0 128.7 205.2 ;
        RECT  123.3 204.0 124.5 205.2 ;
        RECT  127.2 205.2 128.4 205.8 ;
        RECT  126.6 205.8 128.4 207.0 ;
        RECT  127.2 207.0 128.4 210.6 ;
        RECT  123.6 205.2 124.8 208.5 ;
        RECT  123.6 208.5 126.0 209.7 ;
        RECT  120.9 204.0 122.1 209.7 ;
        RECT  123.6 209.7 124.8 210.6 ;
        RECT  129.9 210.6 131.1 212.7 ;
        RECT  126.9 210.6 128.1 211.8 ;
        RECT  123.9 210.6 125.1 211.8 ;
        RECT  120.9 210.6 122.1 212.7 ;
        RECT  119.7 212.7 131.1 213.9 ;
        RECT  119.7 201.3 131.1 202.5 ;
        RECT  119.7 212.7 131.1 213.9 ;
        RECT  126.0 226.2 128.7 227.4 ;
        RECT  121.8 226.2 124.5 227.4 ;
        RECT  119.7 224.1 131.1 225.3 ;
        RECT  125.4 223.8 126.6 224.1 ;
        RECT  129.9 216.9 131.1 222.6 ;
        RECT  127.5 221.4 128.7 222.6 ;
        RECT  123.3 221.4 124.5 222.6 ;
        RECT  127.2 220.8 128.4 221.4 ;
        RECT  126.6 219.6 128.4 220.8 ;
        RECT  127.2 216.0 128.4 219.6 ;
        RECT  123.6 218.1 124.8 221.4 ;
        RECT  123.6 216.9 126.0 218.1 ;
        RECT  120.9 216.9 122.1 222.6 ;
        RECT  123.6 216.0 124.8 216.9 ;
        RECT  129.9 213.9 131.1 216.0 ;
        RECT  126.9 214.8 128.1 216.0 ;
        RECT  123.9 214.8 125.1 216.0 ;
        RECT  120.9 213.9 122.1 216.0 ;
        RECT  119.7 212.7 131.1 213.9 ;
        RECT  119.7 224.1 131.1 225.3 ;
        RECT  119.7 212.7 131.1 213.9 ;
        RECT  126.0 227.4 128.7 228.6 ;
        RECT  121.8 227.4 124.5 228.6 ;
        RECT  119.7 229.5 131.1 230.7 ;
        RECT  125.4 230.7 126.6 231.0 ;
        RECT  129.9 232.2 131.1 237.9 ;
        RECT  127.5 232.2 128.7 233.4 ;
        RECT  123.3 232.2 124.5 233.4 ;
        RECT  127.2 233.4 128.4 234.0 ;
        RECT  126.6 234.0 128.4 235.2 ;
        RECT  127.2 235.2 128.4 238.8 ;
        RECT  123.6 233.4 124.8 236.7 ;
        RECT  123.6 236.7 126.0 237.9 ;
        RECT  120.9 232.2 122.1 237.9 ;
        RECT  123.6 237.9 124.8 238.8 ;
        RECT  129.9 238.8 131.1 240.9 ;
        RECT  126.9 238.8 128.1 240.0 ;
        RECT  123.9 238.8 125.1 240.0 ;
        RECT  120.9 238.8 122.1 240.9 ;
        RECT  119.7 240.9 131.1 242.1 ;
        RECT  119.7 229.5 131.1 230.7 ;
        RECT  119.7 240.9 131.1 242.1 ;
        RECT  126.0 254.4 128.7 255.6 ;
        RECT  121.8 254.4 124.5 255.6 ;
        RECT  119.7 252.3 131.1 253.5 ;
        RECT  125.4 252.0 126.6 252.3 ;
        RECT  129.9 245.1 131.1 250.8 ;
        RECT  127.5 249.6 128.7 250.8 ;
        RECT  123.3 249.6 124.5 250.8 ;
        RECT  127.2 249.0 128.4 249.6 ;
        RECT  126.6 247.8 128.4 249.0 ;
        RECT  127.2 244.2 128.4 247.8 ;
        RECT  123.6 246.3 124.8 249.6 ;
        RECT  123.6 245.1 126.0 246.3 ;
        RECT  120.9 245.1 122.1 250.8 ;
        RECT  123.6 244.2 124.8 245.1 ;
        RECT  129.9 242.1 131.1 244.2 ;
        RECT  126.9 243.0 128.1 244.2 ;
        RECT  123.9 243.0 125.1 244.2 ;
        RECT  120.9 242.1 122.1 244.2 ;
        RECT  119.7 240.9 131.1 242.1 ;
        RECT  119.7 252.3 131.1 253.5 ;
        RECT  119.7 240.9 131.1 242.1 ;
        RECT  126.0 255.6 128.7 256.8 ;
        RECT  121.8 255.6 124.5 256.8 ;
        RECT  119.7 257.7 131.1 258.9 ;
        RECT  125.4 258.9 126.6 259.2 ;
        RECT  129.9 260.4 131.1 266.1 ;
        RECT  127.5 260.4 128.7 261.6 ;
        RECT  123.3 260.4 124.5 261.6 ;
        RECT  127.2 261.6 128.4 262.2 ;
        RECT  126.6 262.2 128.4 263.4 ;
        RECT  127.2 263.4 128.4 267.0 ;
        RECT  123.6 261.6 124.8 264.9 ;
        RECT  123.6 264.9 126.0 266.1 ;
        RECT  120.9 260.4 122.1 266.1 ;
        RECT  123.6 266.1 124.8 267.0 ;
        RECT  129.9 267.0 131.1 269.1 ;
        RECT  126.9 267.0 128.1 268.2 ;
        RECT  123.9 267.0 125.1 268.2 ;
        RECT  120.9 267.0 122.1 269.1 ;
        RECT  119.7 269.1 131.1 270.3 ;
        RECT  119.7 257.7 131.1 258.9 ;
        RECT  119.7 269.1 131.1 270.3 ;
        RECT  126.0 282.6 128.7 283.8 ;
        RECT  121.8 282.6 124.5 283.8 ;
        RECT  119.7 280.5 131.1 281.7 ;
        RECT  125.4 280.2 126.6 280.5 ;
        RECT  129.9 273.3 131.1 279.0 ;
        RECT  127.5 277.8 128.7 279.0 ;
        RECT  123.3 277.8 124.5 279.0 ;
        RECT  127.2 277.2 128.4 277.8 ;
        RECT  126.6 276.0 128.4 277.2 ;
        RECT  127.2 272.4 128.4 276.0 ;
        RECT  123.6 274.5 124.8 277.8 ;
        RECT  123.6 273.3 126.0 274.5 ;
        RECT  120.9 273.3 122.1 279.0 ;
        RECT  123.6 272.4 124.8 273.3 ;
        RECT  129.9 270.3 131.1 272.4 ;
        RECT  126.9 271.2 128.1 272.4 ;
        RECT  123.9 271.2 125.1 272.4 ;
        RECT  120.9 270.3 122.1 272.4 ;
        RECT  119.7 269.1 131.1 270.3 ;
        RECT  119.7 280.5 131.1 281.7 ;
        RECT  119.7 269.1 131.1 270.3 ;
        RECT  126.0 283.8 128.7 285.0 ;
        RECT  121.8 283.8 124.5 285.0 ;
        RECT  119.7 285.9 131.1 287.1 ;
        RECT  125.4 287.1 126.6 287.4 ;
        RECT  129.9 288.6 131.1 294.3 ;
        RECT  127.5 288.6 128.7 289.8 ;
        RECT  123.3 288.6 124.5 289.8 ;
        RECT  127.2 289.8 128.4 290.4 ;
        RECT  126.6 290.4 128.4 291.6 ;
        RECT  127.2 291.6 128.4 295.2 ;
        RECT  123.6 289.8 124.8 293.1 ;
        RECT  123.6 293.1 126.0 294.3 ;
        RECT  120.9 288.6 122.1 294.3 ;
        RECT  123.6 294.3 124.8 295.2 ;
        RECT  129.9 295.2 131.1 297.3 ;
        RECT  126.9 295.2 128.1 296.4 ;
        RECT  123.9 295.2 125.1 296.4 ;
        RECT  120.9 295.2 122.1 297.3 ;
        RECT  119.7 297.3 131.1 298.5 ;
        RECT  119.7 285.9 131.1 287.1 ;
        RECT  119.7 297.3 131.1 298.5 ;
        RECT  126.0 310.8 128.7 312.0 ;
        RECT  121.8 310.8 124.5 312.0 ;
        RECT  119.7 308.7 131.1 309.9 ;
        RECT  125.4 308.4 126.6 308.7 ;
        RECT  129.9 301.5 131.1 307.2 ;
        RECT  127.5 306.0 128.7 307.2 ;
        RECT  123.3 306.0 124.5 307.2 ;
        RECT  127.2 305.4 128.4 306.0 ;
        RECT  126.6 304.2 128.4 305.4 ;
        RECT  127.2 300.6 128.4 304.2 ;
        RECT  123.6 302.7 124.8 306.0 ;
        RECT  123.6 301.5 126.0 302.7 ;
        RECT  120.9 301.5 122.1 307.2 ;
        RECT  123.6 300.6 124.8 301.5 ;
        RECT  129.9 298.5 131.1 300.6 ;
        RECT  126.9 299.4 128.1 300.6 ;
        RECT  123.9 299.4 125.1 300.6 ;
        RECT  120.9 298.5 122.1 300.6 ;
        RECT  119.7 297.3 131.1 298.5 ;
        RECT  119.7 308.7 131.1 309.9 ;
        RECT  119.7 297.3 131.1 298.5 ;
        RECT  126.0 312.0 128.7 313.2 ;
        RECT  121.8 312.0 124.5 313.2 ;
        RECT  119.7 314.1 131.1 315.3 ;
        RECT  125.4 315.3 126.6 315.6 ;
        RECT  129.9 316.8 131.1 322.5 ;
        RECT  127.5 316.8 128.7 318.0 ;
        RECT  123.3 316.8 124.5 318.0 ;
        RECT  127.2 318.0 128.4 318.6 ;
        RECT  126.6 318.6 128.4 319.8 ;
        RECT  127.2 319.8 128.4 323.4 ;
        RECT  123.6 318.0 124.8 321.3 ;
        RECT  123.6 321.3 126.0 322.5 ;
        RECT  120.9 316.8 122.1 322.5 ;
        RECT  123.6 322.5 124.8 323.4 ;
        RECT  129.9 323.4 131.1 325.5 ;
        RECT  126.9 323.4 128.1 324.6 ;
        RECT  123.9 323.4 125.1 324.6 ;
        RECT  120.9 323.4 122.1 325.5 ;
        RECT  119.7 325.5 131.1 326.7 ;
        RECT  119.7 314.1 131.1 315.3 ;
        RECT  119.7 325.5 131.1 326.7 ;
        RECT  126.0 339.0 128.7 340.2 ;
        RECT  121.8 339.0 124.5 340.2 ;
        RECT  119.7 336.9 131.1 338.1 ;
        RECT  125.4 336.6 126.6 336.9 ;
        RECT  129.9 329.7 131.1 335.4 ;
        RECT  127.5 334.2 128.7 335.4 ;
        RECT  123.3 334.2 124.5 335.4 ;
        RECT  127.2 333.6 128.4 334.2 ;
        RECT  126.6 332.4 128.4 333.6 ;
        RECT  127.2 328.8 128.4 332.4 ;
        RECT  123.6 330.9 124.8 334.2 ;
        RECT  123.6 329.7 126.0 330.9 ;
        RECT  120.9 329.7 122.1 335.4 ;
        RECT  123.6 328.8 124.8 329.7 ;
        RECT  129.9 326.7 131.1 328.8 ;
        RECT  126.9 327.6 128.1 328.8 ;
        RECT  123.9 327.6 125.1 328.8 ;
        RECT  120.9 326.7 122.1 328.8 ;
        RECT  119.7 325.5 131.1 326.7 ;
        RECT  119.7 336.9 131.1 338.1 ;
        RECT  119.7 325.5 131.1 326.7 ;
        RECT  126.0 340.2 128.7 341.4 ;
        RECT  121.8 340.2 124.5 341.4 ;
        RECT  119.7 342.3 131.1 343.5 ;
        RECT  125.4 343.5 126.6 343.8 ;
        RECT  129.9 345.0 131.1 350.7 ;
        RECT  127.5 345.0 128.7 346.2 ;
        RECT  123.3 345.0 124.5 346.2 ;
        RECT  127.2 346.2 128.4 346.8 ;
        RECT  126.6 346.8 128.4 348.0 ;
        RECT  127.2 348.0 128.4 351.6 ;
        RECT  123.6 346.2 124.8 349.5 ;
        RECT  123.6 349.5 126.0 350.7 ;
        RECT  120.9 345.0 122.1 350.7 ;
        RECT  123.6 350.7 124.8 351.6 ;
        RECT  129.9 351.6 131.1 353.7 ;
        RECT  126.9 351.6 128.1 352.8 ;
        RECT  123.9 351.6 125.1 352.8 ;
        RECT  120.9 351.6 122.1 353.7 ;
        RECT  119.7 353.7 131.1 354.9 ;
        RECT  119.7 342.3 131.1 343.5 ;
        RECT  119.7 353.7 131.1 354.9 ;
        RECT  126.0 367.2 128.7 368.4 ;
        RECT  121.8 367.2 124.5 368.4 ;
        RECT  119.7 365.1 131.1 366.3 ;
        RECT  125.4 364.8 126.6 365.1 ;
        RECT  129.9 357.9 131.1 363.6 ;
        RECT  127.5 362.4 128.7 363.6 ;
        RECT  123.3 362.4 124.5 363.6 ;
        RECT  127.2 361.8 128.4 362.4 ;
        RECT  126.6 360.6 128.4 361.8 ;
        RECT  127.2 357.0 128.4 360.6 ;
        RECT  123.6 359.1 124.8 362.4 ;
        RECT  123.6 357.9 126.0 359.1 ;
        RECT  120.9 357.9 122.1 363.6 ;
        RECT  123.6 357.0 124.8 357.9 ;
        RECT  129.9 354.9 131.1 357.0 ;
        RECT  126.9 355.8 128.1 357.0 ;
        RECT  123.9 355.8 125.1 357.0 ;
        RECT  120.9 354.9 122.1 357.0 ;
        RECT  119.7 353.7 131.1 354.9 ;
        RECT  119.7 365.1 131.1 366.3 ;
        RECT  119.7 353.7 131.1 354.9 ;
        RECT  126.0 368.4 128.7 369.6 ;
        RECT  121.8 368.4 124.5 369.6 ;
        RECT  119.7 370.5 131.1 371.7 ;
        RECT  125.4 371.7 126.6 372.0 ;
        RECT  129.9 373.2 131.1 378.9 ;
        RECT  127.5 373.2 128.7 374.4 ;
        RECT  123.3 373.2 124.5 374.4 ;
        RECT  127.2 374.4 128.4 375.0 ;
        RECT  126.6 375.0 128.4 376.2 ;
        RECT  127.2 376.2 128.4 379.8 ;
        RECT  123.6 374.4 124.8 377.7 ;
        RECT  123.6 377.7 126.0 378.9 ;
        RECT  120.9 373.2 122.1 378.9 ;
        RECT  123.6 378.9 124.8 379.8 ;
        RECT  129.9 379.8 131.1 381.9 ;
        RECT  126.9 379.8 128.1 381.0 ;
        RECT  123.9 379.8 125.1 381.0 ;
        RECT  120.9 379.8 122.1 381.9 ;
        RECT  119.7 381.9 131.1 383.1 ;
        RECT  119.7 370.5 131.1 371.7 ;
        RECT  119.7 381.9 131.1 383.1 ;
        RECT  126.0 395.4 128.7 396.6 ;
        RECT  121.8 395.4 124.5 396.6 ;
        RECT  119.7 393.3 131.1 394.5 ;
        RECT  125.4 393.0 126.6 393.3 ;
        RECT  129.9 386.1 131.1 391.8 ;
        RECT  127.5 390.6 128.7 391.8 ;
        RECT  123.3 390.6 124.5 391.8 ;
        RECT  127.2 390.0 128.4 390.6 ;
        RECT  126.6 388.8 128.4 390.0 ;
        RECT  127.2 385.2 128.4 388.8 ;
        RECT  123.6 387.3 124.8 390.6 ;
        RECT  123.6 386.1 126.0 387.3 ;
        RECT  120.9 386.1 122.1 391.8 ;
        RECT  123.6 385.2 124.8 386.1 ;
        RECT  129.9 383.1 131.1 385.2 ;
        RECT  126.9 384.0 128.1 385.2 ;
        RECT  123.9 384.0 125.1 385.2 ;
        RECT  120.9 383.1 122.1 385.2 ;
        RECT  119.7 381.9 131.1 383.1 ;
        RECT  119.7 393.3 131.1 394.5 ;
        RECT  119.7 381.9 131.1 383.1 ;
        RECT  126.0 396.6 128.7 397.8 ;
        RECT  121.8 396.6 124.5 397.8 ;
        RECT  119.7 398.7 131.1 399.9 ;
        RECT  125.4 399.9 126.6 400.2 ;
        RECT  129.9 401.4 131.1 407.1 ;
        RECT  127.5 401.4 128.7 402.6 ;
        RECT  123.3 401.4 124.5 402.6 ;
        RECT  127.2 402.6 128.4 403.2 ;
        RECT  126.6 403.2 128.4 404.4 ;
        RECT  127.2 404.4 128.4 408.0 ;
        RECT  123.6 402.6 124.8 405.9 ;
        RECT  123.6 405.9 126.0 407.1 ;
        RECT  120.9 401.4 122.1 407.1 ;
        RECT  123.6 407.1 124.8 408.0 ;
        RECT  129.9 408.0 131.1 410.1 ;
        RECT  126.9 408.0 128.1 409.2 ;
        RECT  123.9 408.0 125.1 409.2 ;
        RECT  120.9 408.0 122.1 410.1 ;
        RECT  119.7 410.1 131.1 411.3 ;
        RECT  119.7 398.7 131.1 399.9 ;
        RECT  119.7 410.1 131.1 411.3 ;
        RECT  126.0 423.6 128.7 424.8 ;
        RECT  121.8 423.6 124.5 424.8 ;
        RECT  119.7 421.5 131.1 422.7 ;
        RECT  125.4 421.2 126.6 421.5 ;
        RECT  129.9 414.3 131.1 420.0 ;
        RECT  127.5 418.8 128.7 420.0 ;
        RECT  123.3 418.8 124.5 420.0 ;
        RECT  127.2 418.2 128.4 418.8 ;
        RECT  126.6 417.0 128.4 418.2 ;
        RECT  127.2 413.4 128.4 417.0 ;
        RECT  123.6 415.5 124.8 418.8 ;
        RECT  123.6 414.3 126.0 415.5 ;
        RECT  120.9 414.3 122.1 420.0 ;
        RECT  123.6 413.4 124.8 414.3 ;
        RECT  129.9 411.3 131.1 413.4 ;
        RECT  126.9 412.2 128.1 413.4 ;
        RECT  123.9 412.2 125.1 413.4 ;
        RECT  120.9 411.3 122.1 413.4 ;
        RECT  119.7 410.1 131.1 411.3 ;
        RECT  119.7 421.5 131.1 422.7 ;
        RECT  119.7 410.1 131.1 411.3 ;
        RECT  136.2 199.2 138.9 200.4 ;
        RECT  132.0 199.2 134.7 200.4 ;
        RECT  129.9 201.3 141.3 202.5 ;
        RECT  135.6 202.5 136.8 202.8 ;
        RECT  140.1 204.0 141.3 209.7 ;
        RECT  137.7 204.0 138.9 205.2 ;
        RECT  133.5 204.0 134.7 205.2 ;
        RECT  137.4 205.2 138.6 205.8 ;
        RECT  136.8 205.8 138.6 207.0 ;
        RECT  137.4 207.0 138.6 210.6 ;
        RECT  133.8 205.2 135.0 208.5 ;
        RECT  133.8 208.5 136.2 209.7 ;
        RECT  131.1 204.0 132.3 209.7 ;
        RECT  133.8 209.7 135.0 210.6 ;
        RECT  140.1 210.6 141.3 212.7 ;
        RECT  137.1 210.6 138.3 211.8 ;
        RECT  134.1 210.6 135.3 211.8 ;
        RECT  131.1 210.6 132.3 212.7 ;
        RECT  129.9 212.7 141.3 213.9 ;
        RECT  129.9 201.3 141.3 202.5 ;
        RECT  129.9 212.7 141.3 213.9 ;
        RECT  136.2 226.2 138.9 227.4 ;
        RECT  132.0 226.2 134.7 227.4 ;
        RECT  129.9 224.1 141.3 225.3 ;
        RECT  135.6 223.8 136.8 224.1 ;
        RECT  140.1 216.9 141.3 222.6 ;
        RECT  137.7 221.4 138.9 222.6 ;
        RECT  133.5 221.4 134.7 222.6 ;
        RECT  137.4 220.8 138.6 221.4 ;
        RECT  136.8 219.6 138.6 220.8 ;
        RECT  137.4 216.0 138.6 219.6 ;
        RECT  133.8 218.1 135.0 221.4 ;
        RECT  133.8 216.9 136.2 218.1 ;
        RECT  131.1 216.9 132.3 222.6 ;
        RECT  133.8 216.0 135.0 216.9 ;
        RECT  140.1 213.9 141.3 216.0 ;
        RECT  137.1 214.8 138.3 216.0 ;
        RECT  134.1 214.8 135.3 216.0 ;
        RECT  131.1 213.9 132.3 216.0 ;
        RECT  129.9 212.7 141.3 213.9 ;
        RECT  129.9 224.1 141.3 225.3 ;
        RECT  129.9 212.7 141.3 213.9 ;
        RECT  136.2 227.4 138.9 228.6 ;
        RECT  132.0 227.4 134.7 228.6 ;
        RECT  129.9 229.5 141.3 230.7 ;
        RECT  135.6 230.7 136.8 231.0 ;
        RECT  140.1 232.2 141.3 237.9 ;
        RECT  137.7 232.2 138.9 233.4 ;
        RECT  133.5 232.2 134.7 233.4 ;
        RECT  137.4 233.4 138.6 234.0 ;
        RECT  136.8 234.0 138.6 235.2 ;
        RECT  137.4 235.2 138.6 238.8 ;
        RECT  133.8 233.4 135.0 236.7 ;
        RECT  133.8 236.7 136.2 237.9 ;
        RECT  131.1 232.2 132.3 237.9 ;
        RECT  133.8 237.9 135.0 238.8 ;
        RECT  140.1 238.8 141.3 240.9 ;
        RECT  137.1 238.8 138.3 240.0 ;
        RECT  134.1 238.8 135.3 240.0 ;
        RECT  131.1 238.8 132.3 240.9 ;
        RECT  129.9 240.9 141.3 242.1 ;
        RECT  129.9 229.5 141.3 230.7 ;
        RECT  129.9 240.9 141.3 242.1 ;
        RECT  136.2 254.4 138.9 255.6 ;
        RECT  132.0 254.4 134.7 255.6 ;
        RECT  129.9 252.3 141.3 253.5 ;
        RECT  135.6 252.0 136.8 252.3 ;
        RECT  140.1 245.1 141.3 250.8 ;
        RECT  137.7 249.6 138.9 250.8 ;
        RECT  133.5 249.6 134.7 250.8 ;
        RECT  137.4 249.0 138.6 249.6 ;
        RECT  136.8 247.8 138.6 249.0 ;
        RECT  137.4 244.2 138.6 247.8 ;
        RECT  133.8 246.3 135.0 249.6 ;
        RECT  133.8 245.1 136.2 246.3 ;
        RECT  131.1 245.1 132.3 250.8 ;
        RECT  133.8 244.2 135.0 245.1 ;
        RECT  140.1 242.1 141.3 244.2 ;
        RECT  137.1 243.0 138.3 244.2 ;
        RECT  134.1 243.0 135.3 244.2 ;
        RECT  131.1 242.1 132.3 244.2 ;
        RECT  129.9 240.9 141.3 242.1 ;
        RECT  129.9 252.3 141.3 253.5 ;
        RECT  129.9 240.9 141.3 242.1 ;
        RECT  136.2 255.6 138.9 256.8 ;
        RECT  132.0 255.6 134.7 256.8 ;
        RECT  129.9 257.7 141.3 258.9 ;
        RECT  135.6 258.9 136.8 259.2 ;
        RECT  140.1 260.4 141.3 266.1 ;
        RECT  137.7 260.4 138.9 261.6 ;
        RECT  133.5 260.4 134.7 261.6 ;
        RECT  137.4 261.6 138.6 262.2 ;
        RECT  136.8 262.2 138.6 263.4 ;
        RECT  137.4 263.4 138.6 267.0 ;
        RECT  133.8 261.6 135.0 264.9 ;
        RECT  133.8 264.9 136.2 266.1 ;
        RECT  131.1 260.4 132.3 266.1 ;
        RECT  133.8 266.1 135.0 267.0 ;
        RECT  140.1 267.0 141.3 269.1 ;
        RECT  137.1 267.0 138.3 268.2 ;
        RECT  134.1 267.0 135.3 268.2 ;
        RECT  131.1 267.0 132.3 269.1 ;
        RECT  129.9 269.1 141.3 270.3 ;
        RECT  129.9 257.7 141.3 258.9 ;
        RECT  129.9 269.1 141.3 270.3 ;
        RECT  136.2 282.6 138.9 283.8 ;
        RECT  132.0 282.6 134.7 283.8 ;
        RECT  129.9 280.5 141.3 281.7 ;
        RECT  135.6 280.2 136.8 280.5 ;
        RECT  140.1 273.3 141.3 279.0 ;
        RECT  137.7 277.8 138.9 279.0 ;
        RECT  133.5 277.8 134.7 279.0 ;
        RECT  137.4 277.2 138.6 277.8 ;
        RECT  136.8 276.0 138.6 277.2 ;
        RECT  137.4 272.4 138.6 276.0 ;
        RECT  133.8 274.5 135.0 277.8 ;
        RECT  133.8 273.3 136.2 274.5 ;
        RECT  131.1 273.3 132.3 279.0 ;
        RECT  133.8 272.4 135.0 273.3 ;
        RECT  140.1 270.3 141.3 272.4 ;
        RECT  137.1 271.2 138.3 272.4 ;
        RECT  134.1 271.2 135.3 272.4 ;
        RECT  131.1 270.3 132.3 272.4 ;
        RECT  129.9 269.1 141.3 270.3 ;
        RECT  129.9 280.5 141.3 281.7 ;
        RECT  129.9 269.1 141.3 270.3 ;
        RECT  136.2 283.8 138.9 285.0 ;
        RECT  132.0 283.8 134.7 285.0 ;
        RECT  129.9 285.9 141.3 287.1 ;
        RECT  135.6 287.1 136.8 287.4 ;
        RECT  140.1 288.6 141.3 294.3 ;
        RECT  137.7 288.6 138.9 289.8 ;
        RECT  133.5 288.6 134.7 289.8 ;
        RECT  137.4 289.8 138.6 290.4 ;
        RECT  136.8 290.4 138.6 291.6 ;
        RECT  137.4 291.6 138.6 295.2 ;
        RECT  133.8 289.8 135.0 293.1 ;
        RECT  133.8 293.1 136.2 294.3 ;
        RECT  131.1 288.6 132.3 294.3 ;
        RECT  133.8 294.3 135.0 295.2 ;
        RECT  140.1 295.2 141.3 297.3 ;
        RECT  137.1 295.2 138.3 296.4 ;
        RECT  134.1 295.2 135.3 296.4 ;
        RECT  131.1 295.2 132.3 297.3 ;
        RECT  129.9 297.3 141.3 298.5 ;
        RECT  129.9 285.9 141.3 287.1 ;
        RECT  129.9 297.3 141.3 298.5 ;
        RECT  136.2 310.8 138.9 312.0 ;
        RECT  132.0 310.8 134.7 312.0 ;
        RECT  129.9 308.7 141.3 309.9 ;
        RECT  135.6 308.4 136.8 308.7 ;
        RECT  140.1 301.5 141.3 307.2 ;
        RECT  137.7 306.0 138.9 307.2 ;
        RECT  133.5 306.0 134.7 307.2 ;
        RECT  137.4 305.4 138.6 306.0 ;
        RECT  136.8 304.2 138.6 305.4 ;
        RECT  137.4 300.6 138.6 304.2 ;
        RECT  133.8 302.7 135.0 306.0 ;
        RECT  133.8 301.5 136.2 302.7 ;
        RECT  131.1 301.5 132.3 307.2 ;
        RECT  133.8 300.6 135.0 301.5 ;
        RECT  140.1 298.5 141.3 300.6 ;
        RECT  137.1 299.4 138.3 300.6 ;
        RECT  134.1 299.4 135.3 300.6 ;
        RECT  131.1 298.5 132.3 300.6 ;
        RECT  129.9 297.3 141.3 298.5 ;
        RECT  129.9 308.7 141.3 309.9 ;
        RECT  129.9 297.3 141.3 298.5 ;
        RECT  136.2 312.0 138.9 313.2 ;
        RECT  132.0 312.0 134.7 313.2 ;
        RECT  129.9 314.1 141.3 315.3 ;
        RECT  135.6 315.3 136.8 315.6 ;
        RECT  140.1 316.8 141.3 322.5 ;
        RECT  137.7 316.8 138.9 318.0 ;
        RECT  133.5 316.8 134.7 318.0 ;
        RECT  137.4 318.0 138.6 318.6 ;
        RECT  136.8 318.6 138.6 319.8 ;
        RECT  137.4 319.8 138.6 323.4 ;
        RECT  133.8 318.0 135.0 321.3 ;
        RECT  133.8 321.3 136.2 322.5 ;
        RECT  131.1 316.8 132.3 322.5 ;
        RECT  133.8 322.5 135.0 323.4 ;
        RECT  140.1 323.4 141.3 325.5 ;
        RECT  137.1 323.4 138.3 324.6 ;
        RECT  134.1 323.4 135.3 324.6 ;
        RECT  131.1 323.4 132.3 325.5 ;
        RECT  129.9 325.5 141.3 326.7 ;
        RECT  129.9 314.1 141.3 315.3 ;
        RECT  129.9 325.5 141.3 326.7 ;
        RECT  136.2 339.0 138.9 340.2 ;
        RECT  132.0 339.0 134.7 340.2 ;
        RECT  129.9 336.9 141.3 338.1 ;
        RECT  135.6 336.6 136.8 336.9 ;
        RECT  140.1 329.7 141.3 335.4 ;
        RECT  137.7 334.2 138.9 335.4 ;
        RECT  133.5 334.2 134.7 335.4 ;
        RECT  137.4 333.6 138.6 334.2 ;
        RECT  136.8 332.4 138.6 333.6 ;
        RECT  137.4 328.8 138.6 332.4 ;
        RECT  133.8 330.9 135.0 334.2 ;
        RECT  133.8 329.7 136.2 330.9 ;
        RECT  131.1 329.7 132.3 335.4 ;
        RECT  133.8 328.8 135.0 329.7 ;
        RECT  140.1 326.7 141.3 328.8 ;
        RECT  137.1 327.6 138.3 328.8 ;
        RECT  134.1 327.6 135.3 328.8 ;
        RECT  131.1 326.7 132.3 328.8 ;
        RECT  129.9 325.5 141.3 326.7 ;
        RECT  129.9 336.9 141.3 338.1 ;
        RECT  129.9 325.5 141.3 326.7 ;
        RECT  136.2 340.2 138.9 341.4 ;
        RECT  132.0 340.2 134.7 341.4 ;
        RECT  129.9 342.3 141.3 343.5 ;
        RECT  135.6 343.5 136.8 343.8 ;
        RECT  140.1 345.0 141.3 350.7 ;
        RECT  137.7 345.0 138.9 346.2 ;
        RECT  133.5 345.0 134.7 346.2 ;
        RECT  137.4 346.2 138.6 346.8 ;
        RECT  136.8 346.8 138.6 348.0 ;
        RECT  137.4 348.0 138.6 351.6 ;
        RECT  133.8 346.2 135.0 349.5 ;
        RECT  133.8 349.5 136.2 350.7 ;
        RECT  131.1 345.0 132.3 350.7 ;
        RECT  133.8 350.7 135.0 351.6 ;
        RECT  140.1 351.6 141.3 353.7 ;
        RECT  137.1 351.6 138.3 352.8 ;
        RECT  134.1 351.6 135.3 352.8 ;
        RECT  131.1 351.6 132.3 353.7 ;
        RECT  129.9 353.7 141.3 354.9 ;
        RECT  129.9 342.3 141.3 343.5 ;
        RECT  129.9 353.7 141.3 354.9 ;
        RECT  136.2 367.2 138.9 368.4 ;
        RECT  132.0 367.2 134.7 368.4 ;
        RECT  129.9 365.1 141.3 366.3 ;
        RECT  135.6 364.8 136.8 365.1 ;
        RECT  140.1 357.9 141.3 363.6 ;
        RECT  137.7 362.4 138.9 363.6 ;
        RECT  133.5 362.4 134.7 363.6 ;
        RECT  137.4 361.8 138.6 362.4 ;
        RECT  136.8 360.6 138.6 361.8 ;
        RECT  137.4 357.0 138.6 360.6 ;
        RECT  133.8 359.1 135.0 362.4 ;
        RECT  133.8 357.9 136.2 359.1 ;
        RECT  131.1 357.9 132.3 363.6 ;
        RECT  133.8 357.0 135.0 357.9 ;
        RECT  140.1 354.9 141.3 357.0 ;
        RECT  137.1 355.8 138.3 357.0 ;
        RECT  134.1 355.8 135.3 357.0 ;
        RECT  131.1 354.9 132.3 357.0 ;
        RECT  129.9 353.7 141.3 354.9 ;
        RECT  129.9 365.1 141.3 366.3 ;
        RECT  129.9 353.7 141.3 354.9 ;
        RECT  136.2 368.4 138.9 369.6 ;
        RECT  132.0 368.4 134.7 369.6 ;
        RECT  129.9 370.5 141.3 371.7 ;
        RECT  135.6 371.7 136.8 372.0 ;
        RECT  140.1 373.2 141.3 378.9 ;
        RECT  137.7 373.2 138.9 374.4 ;
        RECT  133.5 373.2 134.7 374.4 ;
        RECT  137.4 374.4 138.6 375.0 ;
        RECT  136.8 375.0 138.6 376.2 ;
        RECT  137.4 376.2 138.6 379.8 ;
        RECT  133.8 374.4 135.0 377.7 ;
        RECT  133.8 377.7 136.2 378.9 ;
        RECT  131.1 373.2 132.3 378.9 ;
        RECT  133.8 378.9 135.0 379.8 ;
        RECT  140.1 379.8 141.3 381.9 ;
        RECT  137.1 379.8 138.3 381.0 ;
        RECT  134.1 379.8 135.3 381.0 ;
        RECT  131.1 379.8 132.3 381.9 ;
        RECT  129.9 381.9 141.3 383.1 ;
        RECT  129.9 370.5 141.3 371.7 ;
        RECT  129.9 381.9 141.3 383.1 ;
        RECT  136.2 395.4 138.9 396.6 ;
        RECT  132.0 395.4 134.7 396.6 ;
        RECT  129.9 393.3 141.3 394.5 ;
        RECT  135.6 393.0 136.8 393.3 ;
        RECT  140.1 386.1 141.3 391.8 ;
        RECT  137.7 390.6 138.9 391.8 ;
        RECT  133.5 390.6 134.7 391.8 ;
        RECT  137.4 390.0 138.6 390.6 ;
        RECT  136.8 388.8 138.6 390.0 ;
        RECT  137.4 385.2 138.6 388.8 ;
        RECT  133.8 387.3 135.0 390.6 ;
        RECT  133.8 386.1 136.2 387.3 ;
        RECT  131.1 386.1 132.3 391.8 ;
        RECT  133.8 385.2 135.0 386.1 ;
        RECT  140.1 383.1 141.3 385.2 ;
        RECT  137.1 384.0 138.3 385.2 ;
        RECT  134.1 384.0 135.3 385.2 ;
        RECT  131.1 383.1 132.3 385.2 ;
        RECT  129.9 381.9 141.3 383.1 ;
        RECT  129.9 393.3 141.3 394.5 ;
        RECT  129.9 381.9 141.3 383.1 ;
        RECT  136.2 396.6 138.9 397.8 ;
        RECT  132.0 396.6 134.7 397.8 ;
        RECT  129.9 398.7 141.3 399.9 ;
        RECT  135.6 399.9 136.8 400.2 ;
        RECT  140.1 401.4 141.3 407.1 ;
        RECT  137.7 401.4 138.9 402.6 ;
        RECT  133.5 401.4 134.7 402.6 ;
        RECT  137.4 402.6 138.6 403.2 ;
        RECT  136.8 403.2 138.6 404.4 ;
        RECT  137.4 404.4 138.6 408.0 ;
        RECT  133.8 402.6 135.0 405.9 ;
        RECT  133.8 405.9 136.2 407.1 ;
        RECT  131.1 401.4 132.3 407.1 ;
        RECT  133.8 407.1 135.0 408.0 ;
        RECT  140.1 408.0 141.3 410.1 ;
        RECT  137.1 408.0 138.3 409.2 ;
        RECT  134.1 408.0 135.3 409.2 ;
        RECT  131.1 408.0 132.3 410.1 ;
        RECT  129.9 410.1 141.3 411.3 ;
        RECT  129.9 398.7 141.3 399.9 ;
        RECT  129.9 410.1 141.3 411.3 ;
        RECT  136.2 423.6 138.9 424.8 ;
        RECT  132.0 423.6 134.7 424.8 ;
        RECT  129.9 421.5 141.3 422.7 ;
        RECT  135.6 421.2 136.8 421.5 ;
        RECT  140.1 414.3 141.3 420.0 ;
        RECT  137.7 418.8 138.9 420.0 ;
        RECT  133.5 418.8 134.7 420.0 ;
        RECT  137.4 418.2 138.6 418.8 ;
        RECT  136.8 417.0 138.6 418.2 ;
        RECT  137.4 413.4 138.6 417.0 ;
        RECT  133.8 415.5 135.0 418.8 ;
        RECT  133.8 414.3 136.2 415.5 ;
        RECT  131.1 414.3 132.3 420.0 ;
        RECT  133.8 413.4 135.0 414.3 ;
        RECT  140.1 411.3 141.3 413.4 ;
        RECT  137.1 412.2 138.3 413.4 ;
        RECT  134.1 412.2 135.3 413.4 ;
        RECT  131.1 411.3 132.3 413.4 ;
        RECT  129.9 410.1 141.3 411.3 ;
        RECT  129.9 421.5 141.3 422.7 ;
        RECT  129.9 410.1 141.3 411.3 ;
        RECT  120.3 431.4 140.7 432.3 ;
        RECT  120.3 443.4 140.7 444.3 ;
        RECT  125.7 435.9 126.6 444.3 ;
        RECT  120.3 443.4 130.5 444.3 ;
        RECT  120.3 431.4 130.5 432.3 ;
        RECT  123.3 427.5 124.5 428.7 ;
        RECT  125.7 427.5 126.9 428.7 ;
        RECT  123.3 427.5 124.5 428.7 ;
        RECT  125.7 427.5 126.9 428.7 ;
        RECT  123.3 435.9 124.5 437.1 ;
        RECT  125.7 435.9 126.9 437.1 ;
        RECT  123.3 435.9 124.5 437.1 ;
        RECT  125.7 435.9 126.9 437.1 ;
        RECT  125.7 435.9 126.9 437.1 ;
        RECT  128.1 435.9 129.3 437.1 ;
        RECT  125.7 435.9 126.9 437.1 ;
        RECT  128.1 435.9 129.3 437.1 ;
        RECT  124.2 431.4 125.4 432.6 ;
        RECT  125.7 441.3 126.9 442.5 ;
        RECT  123.3 435.9 124.5 437.1 ;
        RECT  128.1 435.9 129.3 437.1 ;
        RECT  123.3 427.5 124.5 428.7 ;
        RECT  125.7 427.5 126.9 428.7 ;
        RECT  135.9 435.9 136.8 444.3 ;
        RECT  130.5 443.4 140.7 444.3 ;
        RECT  130.5 431.4 140.7 432.3 ;
        RECT  133.5 427.5 134.7 428.7 ;
        RECT  135.9 427.5 137.1 428.7 ;
        RECT  133.5 427.5 134.7 428.7 ;
        RECT  135.9 427.5 137.1 428.7 ;
        RECT  133.5 435.9 134.7 437.1 ;
        RECT  135.9 435.9 137.1 437.1 ;
        RECT  133.5 435.9 134.7 437.1 ;
        RECT  135.9 435.9 137.1 437.1 ;
        RECT  135.9 435.9 137.1 437.1 ;
        RECT  138.3 435.9 139.5 437.1 ;
        RECT  135.9 435.9 137.1 437.1 ;
        RECT  138.3 435.9 139.5 437.1 ;
        RECT  134.4 431.4 135.6 432.6 ;
        RECT  135.9 441.3 137.1 442.5 ;
        RECT  133.5 435.9 134.7 437.1 ;
        RECT  138.3 435.9 139.5 437.1 ;
        RECT  133.5 427.5 134.7 428.7 ;
        RECT  135.9 427.5 137.1 428.7 ;
        RECT  120.3 195.0 140.7 195.9 ;
        RECT  120.3 167.7 140.7 168.6 ;
        RECT  120.3 192.9 140.7 193.8 ;
        RECT  119.7 195.0 131.1 196.2 ;
        RECT  119.7 192.9 131.1 194.1 ;
        RECT  125.1 189.3 126.3 192.0 ;
        RECT  127.5 189.3 128.7 192.9 ;
        RECT  129.9 191.7 131.1 192.9 ;
        RECT  125.1 185.4 126.0 189.3 ;
        RECT  122.4 171.0 123.6 185.4 ;
        RECT  124.8 182.7 126.0 185.4 ;
        RECT  127.2 181.8 128.4 185.4 ;
        RECT  127.2 180.6 129.3 181.8 ;
        RECT  124.8 173.7 126.0 179.1 ;
        RECT  127.2 173.7 128.4 180.6 ;
        RECT  124.8 172.8 125.7 173.7 ;
        RECT  124.8 171.9 126.6 172.8 ;
        RECT  122.4 169.8 124.2 171.0 ;
        RECT  125.7 170.1 126.6 171.9 ;
        RECT  125.7 168.9 126.9 170.1 ;
        RECT  119.7 167.7 131.1 168.9 ;
        RECT  123.0 166.5 124.2 166.8 ;
        RECT  122.1 165.6 124.2 166.5 ;
        RECT  129.0 165.6 130.5 166.8 ;
        RECT  122.1 163.5 123.0 165.6 ;
        RECT  124.2 163.5 125.4 164.7 ;
        RECT  122.1 157.2 123.3 163.5 ;
        RECT  121.2 156.3 123.3 157.2 ;
        RECT  124.5 156.3 125.7 163.5 ;
        RECT  126.9 156.3 128.1 164.7 ;
        RECT  129.6 163.5 130.5 165.6 ;
        RECT  129.3 156.3 130.5 163.5 ;
        RECT  121.2 153.6 122.4 156.3 ;
        RECT  119.7 195.0 131.1 196.2 ;
        RECT  119.7 167.7 131.1 168.9 ;
        RECT  119.7 192.9 131.1 194.1 ;
        RECT  129.9 195.0 141.3 196.2 ;
        RECT  129.9 192.9 141.3 194.1 ;
        RECT  135.3 189.3 136.5 192.0 ;
        RECT  137.7 189.3 138.9 192.9 ;
        RECT  140.1 191.7 141.3 192.9 ;
        RECT  135.3 185.4 136.2 189.3 ;
        RECT  132.6 171.0 133.8 185.4 ;
        RECT  135.0 182.7 136.2 185.4 ;
        RECT  137.4 181.8 138.6 185.4 ;
        RECT  137.4 180.6 139.5 181.8 ;
        RECT  135.0 173.7 136.2 179.1 ;
        RECT  137.4 173.7 138.6 180.6 ;
        RECT  135.0 172.8 135.9 173.7 ;
        RECT  135.0 171.9 136.8 172.8 ;
        RECT  132.6 169.8 134.4 171.0 ;
        RECT  135.9 170.1 136.8 171.9 ;
        RECT  135.9 168.9 137.1 170.1 ;
        RECT  129.9 167.7 141.3 168.9 ;
        RECT  133.2 166.5 134.4 166.8 ;
        RECT  132.3 165.6 134.4 166.5 ;
        RECT  139.2 165.6 140.7 166.8 ;
        RECT  132.3 163.5 133.2 165.6 ;
        RECT  134.4 163.5 135.6 164.7 ;
        RECT  132.3 157.2 133.5 163.5 ;
        RECT  131.4 156.3 133.5 157.2 ;
        RECT  134.7 156.3 135.9 163.5 ;
        RECT  137.1 156.3 138.3 164.7 ;
        RECT  139.8 163.5 140.7 165.6 ;
        RECT  139.5 156.3 140.7 163.5 ;
        RECT  131.4 153.6 132.6 156.3 ;
        RECT  129.9 195.0 141.3 196.2 ;
        RECT  129.9 167.7 141.3 168.9 ;
        RECT  129.9 192.9 141.3 194.1 ;
        RECT  120.3 96.9 140.7 97.8 ;
        RECT  120.3 99.0 140.7 99.9 ;
        RECT  120.3 94.8 140.7 95.7 ;
        RECT  121.8 147.0 123.0 148.2 ;
        RECT  121.8 146.4 122.7 147.0 ;
        RECT  121.5 142.8 122.7 146.4 ;
        RECT  123.9 142.8 125.1 146.4 ;
        RECT  126.3 142.8 127.5 147.6 ;
        RECT  128.7 144.0 130.2 145.2 ;
        RECT  124.2 140.4 125.1 142.8 ;
        RECT  121.5 127.2 122.7 139.8 ;
        RECT  124.2 139.2 128.4 140.4 ;
        RECT  123.6 136.8 128.4 138.0 ;
        RECT  123.9 132.9 125.1 136.8 ;
        RECT  126.3 132.3 127.5 134.1 ;
        RECT  129.3 132.3 130.2 144.0 ;
        RECT  126.3 131.1 130.2 132.3 ;
        RECT  123.9 126.3 125.1 129.3 ;
        RECT  126.3 127.2 127.5 131.1 ;
        RECT  120.3 125.1 131.1 126.3 ;
        RECT  121.8 120.9 123.0 123.9 ;
        RECT  124.2 121.8 125.4 125.1 ;
        RECT  126.6 120.9 127.8 123.9 ;
        RECT  121.8 120.0 127.8 120.9 ;
        RECT  121.8 114.3 123.0 120.0 ;
        RECT  126.6 119.7 127.8 120.0 ;
        RECT  126.6 118.5 128.4 119.7 ;
        RECT  124.2 114.3 125.4 116.4 ;
        RECT  126.6 115.5 127.8 116.4 ;
        RECT  126.6 114.3 130.5 115.5 ;
        RECT  127.2 112.2 129.6 113.4 ;
        RECT  121.2 111.0 122.4 112.2 ;
        RECT  121.5 108.9 122.4 111.0 ;
        RECT  121.2 105.0 122.4 108.9 ;
        RECT  123.6 106.8 124.8 108.9 ;
        RECT  126.0 106.8 127.2 110.1 ;
        RECT  121.2 104.1 124.8 105.0 ;
        RECT  121.2 100.2 122.4 103.2 ;
        RECT  123.6 101.1 124.8 104.1 ;
        RECT  126.0 100.2 127.2 103.2 ;
        RECT  128.4 101.1 129.6 112.2 ;
        RECT  120.3 99.0 131.1 100.2 ;
        RECT  120.3 96.9 131.1 98.1 ;
        RECT  120.3 94.8 131.1 96.0 ;
        RECT  123.9 92.7 126.3 93.9 ;
        RECT  120.3 96.9 131.1 98.1 ;
        RECT  120.3 99.0 131.1 100.2 ;
        RECT  120.3 94.8 131.1 96.0 ;
        RECT  132.0 147.0 133.2 148.2 ;
        RECT  132.0 146.4 132.9 147.0 ;
        RECT  131.7 142.8 132.9 146.4 ;
        RECT  134.1 142.8 135.3 146.4 ;
        RECT  136.5 142.8 137.7 147.6 ;
        RECT  138.9 144.0 140.4 145.2 ;
        RECT  134.4 140.4 135.3 142.8 ;
        RECT  131.7 127.2 132.9 139.8 ;
        RECT  134.4 139.2 138.6 140.4 ;
        RECT  133.8 136.8 138.6 138.0 ;
        RECT  134.1 132.9 135.3 136.8 ;
        RECT  136.5 132.3 137.7 134.1 ;
        RECT  139.5 132.3 140.4 144.0 ;
        RECT  136.5 131.1 140.4 132.3 ;
        RECT  134.1 126.3 135.3 129.3 ;
        RECT  136.5 127.2 137.7 131.1 ;
        RECT  130.5 125.1 141.3 126.3 ;
        RECT  132.0 120.9 133.2 123.9 ;
        RECT  134.4 121.8 135.6 125.1 ;
        RECT  136.8 120.9 138.0 123.9 ;
        RECT  132.0 120.0 138.0 120.9 ;
        RECT  132.0 114.3 133.2 120.0 ;
        RECT  136.8 119.7 138.0 120.0 ;
        RECT  136.8 118.5 138.6 119.7 ;
        RECT  134.4 114.3 135.6 116.4 ;
        RECT  136.8 115.5 138.0 116.4 ;
        RECT  136.8 114.3 140.7 115.5 ;
        RECT  137.4 112.2 139.8 113.4 ;
        RECT  131.4 111.0 132.6 112.2 ;
        RECT  131.7 108.9 132.6 111.0 ;
        RECT  131.4 105.0 132.6 108.9 ;
        RECT  133.8 106.8 135.0 108.9 ;
        RECT  136.2 106.8 137.4 110.1 ;
        RECT  131.4 104.1 135.0 105.0 ;
        RECT  131.4 100.2 132.6 103.2 ;
        RECT  133.8 101.1 135.0 104.1 ;
        RECT  136.2 100.2 137.4 103.2 ;
        RECT  138.6 101.1 139.8 112.2 ;
        RECT  130.5 99.0 141.3 100.2 ;
        RECT  130.5 96.9 141.3 98.1 ;
        RECT  130.5 94.8 141.3 96.0 ;
        RECT  134.1 92.7 136.5 93.9 ;
        RECT  130.5 96.9 141.3 98.1 ;
        RECT  130.5 99.0 141.3 100.2 ;
        RECT  130.5 94.8 141.3 96.0 ;
        RECT  120.3 32.4 140.7 33.3 ;
        RECT  120.3 86.4 140.7 87.3 ;
        RECT  119.7 86.4 131.1 87.3 ;
        RECT  119.7 83.1 120.9 86.4 ;
        RECT  122.1 84.6 128.7 85.5 ;
        RECT  122.1 84.3 125.1 84.6 ;
        RECT  127.5 84.3 128.7 84.6 ;
        RECT  119.7 81.9 123.9 83.1 ;
        RECT  127.5 81.9 131.1 83.1 ;
        RECT  119.7 78.3 120.9 81.9 ;
        RECT  125.1 81.0 126.3 81.9 ;
        RECT  125.1 80.7 127.5 81.0 ;
        RECT  122.1 79.8 128.7 80.7 ;
        RECT  122.1 79.5 123.9 79.8 ;
        RECT  127.5 79.5 128.7 79.8 ;
        RECT  119.7 77.1 123.9 78.3 ;
        RECT  119.7 63.3 120.9 77.1 ;
        RECT  125.4 76.5 126.6 78.9 ;
        RECT  130.2 78.3 131.1 81.9 ;
        RECT  127.5 77.1 131.1 78.3 ;
        RECT  129.9 75.9 131.1 77.1 ;
        RECT  122.1 73.5 123.3 74.7 ;
        RECT  124.2 74.4 126.6 75.6 ;
        RECT  122.1 72.6 128.7 73.5 ;
        RECT  122.1 72.3 123.9 72.6 ;
        RECT  127.5 72.3 128.7 72.6 ;
        RECT  122.1 70.2 128.7 71.1 ;
        RECT  122.1 69.9 123.9 70.2 ;
        RECT  126.3 69.9 128.7 70.2 ;
        RECT  122.1 67.8 128.7 68.7 ;
        RECT  122.1 67.5 123.9 67.8 ;
        RECT  126.3 67.5 128.7 67.8 ;
        RECT  125.1 65.7 126.3 66.6 ;
        RECT  122.1 64.8 128.7 65.7 ;
        RECT  122.1 64.5 125.1 64.8 ;
        RECT  127.5 64.5 128.7 64.8 ;
        RECT  119.7 62.1 123.9 63.3 ;
        RECT  119.7 57.6 120.9 62.1 ;
        RECT  124.8 61.2 126.0 63.6 ;
        RECT  130.2 63.3 131.1 75.9 ;
        RECT  127.5 62.1 131.1 63.3 ;
        RECT  122.1 60.0 123.3 61.2 ;
        RECT  122.1 59.1 128.7 60.0 ;
        RECT  122.1 58.8 123.9 59.1 ;
        RECT  127.5 58.8 128.7 59.1 ;
        RECT  130.2 57.6 131.1 62.1 ;
        RECT  119.7 56.4 123.9 57.6 ;
        RECT  119.7 52.8 120.9 56.4 ;
        RECT  125.4 55.5 126.6 56.7 ;
        RECT  127.5 56.4 131.1 57.6 ;
        RECT  122.1 55.2 127.5 55.5 ;
        RECT  122.1 54.6 128.7 55.2 ;
        RECT  122.1 54.0 123.9 54.6 ;
        RECT  126.3 54.3 128.7 54.6 ;
        RECT  127.5 54.0 128.7 54.3 ;
        RECT  119.7 51.6 123.9 52.8 ;
        RECT  119.7 36.6 120.9 51.6 ;
        RECT  125.4 51.0 126.6 53.4 ;
        RECT  130.2 52.8 131.1 56.4 ;
        RECT  127.5 51.6 131.1 52.8 ;
        RECT  129.9 50.4 131.1 51.6 ;
        RECT  122.1 47.1 123.3 48.3 ;
        RECT  124.2 48.0 126.6 49.2 ;
        RECT  122.1 46.2 128.7 47.1 ;
        RECT  122.1 45.9 123.9 46.2 ;
        RECT  127.5 45.9 128.7 46.2 ;
        RECT  122.1 43.8 128.7 44.7 ;
        RECT  122.1 43.5 123.9 43.8 ;
        RECT  126.3 43.5 128.7 43.8 ;
        RECT  122.1 41.4 128.7 42.3 ;
        RECT  122.1 41.1 123.9 41.4 ;
        RECT  126.3 41.1 128.7 41.4 ;
        RECT  125.1 39.3 126.3 40.2 ;
        RECT  122.1 38.4 128.7 39.3 ;
        RECT  122.1 38.1 125.1 38.4 ;
        RECT  127.5 38.1 128.7 38.4 ;
        RECT  130.2 36.9 131.1 50.4 ;
        RECT  122.1 36.6 123.9 36.9 ;
        RECT  119.7 35.7 123.9 36.6 ;
        RECT  127.5 36.0 131.1 36.9 ;
        RECT  127.5 35.7 128.7 36.0 ;
        RECT  122.7 34.2 123.9 35.7 ;
        RECT  124.8 33.3 126.0 34.2 ;
        RECT  119.7 32.4 131.1 33.3 ;
        RECT  119.7 32.4 131.1 33.3 ;
        RECT  119.7 86.4 131.1 87.3 ;
        RECT  129.9 86.4 141.3 87.3 ;
        RECT  140.1 83.1 141.3 86.4 ;
        RECT  132.3 84.6 138.9 85.5 ;
        RECT  135.9 84.3 138.9 84.6 ;
        RECT  132.3 84.3 133.5 84.6 ;
        RECT  137.1 81.9 141.3 83.1 ;
        RECT  129.9 81.9 133.5 83.1 ;
        RECT  140.1 78.3 141.3 81.9 ;
        RECT  134.7 81.0 135.9 81.9 ;
        RECT  133.5 80.7 135.9 81.0 ;
        RECT  132.3 79.8 138.9 80.7 ;
        RECT  137.1 79.5 138.9 79.8 ;
        RECT  132.3 79.5 133.5 79.8 ;
        RECT  137.1 77.1 141.3 78.3 ;
        RECT  140.1 63.3 141.3 77.1 ;
        RECT  134.4 76.5 135.6 78.9 ;
        RECT  129.9 78.3 130.8 81.9 ;
        RECT  129.9 77.1 133.5 78.3 ;
        RECT  129.9 75.9 131.1 77.1 ;
        RECT  137.7 73.5 138.9 74.7 ;
        RECT  134.4 74.4 136.8 75.6 ;
        RECT  132.3 72.6 138.9 73.5 ;
        RECT  137.1 72.3 138.9 72.6 ;
        RECT  132.3 72.3 133.5 72.6 ;
        RECT  132.3 70.2 138.9 71.1 ;
        RECT  137.1 69.9 138.9 70.2 ;
        RECT  132.3 69.9 134.7 70.2 ;
        RECT  132.3 67.8 138.9 68.7 ;
        RECT  137.1 67.5 138.9 67.8 ;
        RECT  132.3 67.5 134.7 67.8 ;
        RECT  134.7 65.7 135.9 66.6 ;
        RECT  132.3 64.8 138.9 65.7 ;
        RECT  135.9 64.5 138.9 64.8 ;
        RECT  132.3 64.5 133.5 64.8 ;
        RECT  137.1 62.1 141.3 63.3 ;
        RECT  140.1 57.6 141.3 62.1 ;
        RECT  135.0 61.2 136.2 63.6 ;
        RECT  129.9 63.3 130.8 75.9 ;
        RECT  129.9 62.1 133.5 63.3 ;
        RECT  137.7 60.0 138.9 61.2 ;
        RECT  132.3 59.1 138.9 60.0 ;
        RECT  137.1 58.8 138.9 59.1 ;
        RECT  132.3 58.8 133.5 59.1 ;
        RECT  129.9 57.6 130.8 62.1 ;
        RECT  137.1 56.4 141.3 57.6 ;
        RECT  140.1 52.8 141.3 56.4 ;
        RECT  134.4 55.5 135.6 56.7 ;
        RECT  129.9 56.4 133.5 57.6 ;
        RECT  133.5 55.2 138.9 55.5 ;
        RECT  132.3 54.6 138.9 55.2 ;
        RECT  137.1 54.0 138.9 54.6 ;
        RECT  132.3 54.3 134.7 54.6 ;
        RECT  132.3 54.0 133.5 54.3 ;
        RECT  137.1 51.6 141.3 52.8 ;
        RECT  140.1 36.6 141.3 51.6 ;
        RECT  134.4 51.0 135.6 53.4 ;
        RECT  129.9 52.8 130.8 56.4 ;
        RECT  129.9 51.6 133.5 52.8 ;
        RECT  129.9 50.4 131.1 51.6 ;
        RECT  137.7 47.1 138.9 48.3 ;
        RECT  134.4 48.0 136.8 49.2 ;
        RECT  132.3 46.2 138.9 47.1 ;
        RECT  137.1 45.9 138.9 46.2 ;
        RECT  132.3 45.9 133.5 46.2 ;
        RECT  132.3 43.8 138.9 44.7 ;
        RECT  137.1 43.5 138.9 43.8 ;
        RECT  132.3 43.5 134.7 43.8 ;
        RECT  132.3 41.4 138.9 42.3 ;
        RECT  137.1 41.1 138.9 41.4 ;
        RECT  132.3 41.1 134.7 41.4 ;
        RECT  134.7 39.3 135.9 40.2 ;
        RECT  132.3 38.4 138.9 39.3 ;
        RECT  135.9 38.1 138.9 38.4 ;
        RECT  132.3 38.1 133.5 38.4 ;
        RECT  129.9 36.9 130.8 50.4 ;
        RECT  137.1 36.6 138.9 36.9 ;
        RECT  137.1 35.7 141.3 36.6 ;
        RECT  129.9 36.0 133.5 36.9 ;
        RECT  132.3 35.7 133.5 36.0 ;
        RECT  137.1 34.2 138.3 35.7 ;
        RECT  135.0 33.3 136.2 34.2 ;
        RECT  129.9 32.4 141.3 33.3 ;
        RECT  129.9 32.4 141.3 33.3 ;
        RECT  129.9 86.4 141.3 87.3 ;
        RECT  120.3 25.5 140.7 26.4 ;
        RECT  120.3 9.6 140.7 10.5 ;
        RECT  120.3 23.4 140.7 24.3 ;
        RECT  120.3 27.9 140.7 28.8 ;
        RECT  120.3 49.5 131.1 50.7 ;
        RECT  121.2 45.9 122.7 48.3 ;
        RECT  123.9 45.9 125.1 49.5 ;
        RECT  126.3 45.9 127.5 48.3 ;
        RECT  128.7 45.9 129.9 48.3 ;
        RECT  121.2 42.6 122.1 45.9 ;
        RECT  123.0 43.8 124.2 45.0 ;
        RECT  121.2 41.4 126.3 42.6 ;
        RECT  129.0 41.4 129.9 45.9 ;
        RECT  121.2 39.3 122.1 41.4 ;
        RECT  127.8 40.2 129.9 41.4 ;
        RECT  129.0 39.3 129.9 40.2 ;
        RECT  121.2 38.1 122.7 39.3 ;
        RECT  123.9 36.9 125.1 39.3 ;
        RECT  126.3 38.1 127.5 39.3 ;
        RECT  128.7 38.1 129.9 39.3 ;
        RECT  120.3 35.7 131.1 36.9 ;
        RECT  120.3 33.6 131.1 34.8 ;
        RECT  120.3 31.2 131.1 32.4 ;
        RECT  120.3 33.6 131.1 34.8 ;
        RECT  120.3 49.5 131.1 50.7 ;
        RECT  120.3 35.7 131.1 36.9 ;
        RECT  120.3 35.7 131.1 36.9 ;
        RECT  120.3 31.2 131.1 32.4 ;
        RECT  130.5 49.5 141.3 50.7 ;
        RECT  131.4 45.9 132.9 48.3 ;
        RECT  134.1 45.9 135.3 49.5 ;
        RECT  136.5 45.9 137.7 48.3 ;
        RECT  138.9 45.9 140.1 48.3 ;
        RECT  131.4 42.6 132.3 45.9 ;
        RECT  133.2 43.8 134.4 45.0 ;
        RECT  131.4 41.4 136.5 42.6 ;
        RECT  139.2 41.4 140.1 45.9 ;
        RECT  131.4 39.3 132.3 41.4 ;
        RECT  138.0 40.2 140.1 41.4 ;
        RECT  139.2 39.3 140.1 40.2 ;
        RECT  131.4 38.1 132.9 39.3 ;
        RECT  134.1 36.9 135.3 39.3 ;
        RECT  136.5 38.1 137.7 39.3 ;
        RECT  138.9 38.1 140.1 39.3 ;
        RECT  130.5 35.7 141.3 36.9 ;
        RECT  130.5 33.6 141.3 34.8 ;
        RECT  130.5 31.2 141.3 32.4 ;
        RECT  130.5 33.6 141.3 34.8 ;
        RECT  130.5 49.5 141.3 50.7 ;
        RECT  130.5 35.7 141.3 36.9 ;
        RECT  130.5 35.7 141.3 36.9 ;
        RECT  130.5 31.2 141.3 32.4 ;
        RECT  35.1 205.2 36.0 206.1 ;
        RECT  35.1 220.5 36.0 221.4 ;
        RECT  35.1 233.4 36.0 234.3 ;
        RECT  35.1 248.7 36.0 249.6 ;
        RECT  35.1 261.6 36.0 262.5 ;
        RECT  35.1 276.9 36.0 277.8 ;
        RECT  35.1 289.8 36.0 290.7 ;
        RECT  35.1 305.1 36.0 306.0 ;
        RECT  35.1 318.0 36.0 318.9 ;
        RECT  35.1 333.3 36.0 334.2 ;
        RECT  35.1 346.2 36.0 347.1 ;
        RECT  35.1 361.5 36.0 362.4 ;
        RECT  35.1 374.4 36.0 375.3 ;
        RECT  35.1 389.7 36.0 390.6 ;
        RECT  35.1 402.6 36.0 403.5 ;
        RECT  35.1 417.9 36.0 418.8 ;
        RECT  6.3 92.4 23.1 93.3 ;
        RECT  8.4 107.7 23.1 108.6 ;
        RECT  10.5 120.6 23.1 121.5 ;
        RECT  12.6 135.9 23.1 136.8 ;
        RECT  14.7 148.8 23.1 149.7 ;
        RECT  16.8 164.1 23.1 165.0 ;
        RECT  18.9 177.0 23.1 177.9 ;
        RECT  21.0 192.3 23.1 193.2 ;
        RECT  6.3 207.3 23.1 208.2 ;
        RECT  14.7 204.6 23.1 205.5 ;
        RECT  6.3 218.4 23.1 219.3 ;
        RECT  16.8 221.1 23.1 222.0 ;
        RECT  6.3 235.5 23.1 236.4 ;
        RECT  18.9 232.8 23.1 233.7 ;
        RECT  6.3 246.6 23.1 247.5 ;
        RECT  21.0 249.3 23.1 250.2 ;
        RECT  8.4 263.7 23.1 264.6 ;
        RECT  14.7 261.0 23.1 261.9 ;
        RECT  8.4 274.8 23.1 275.7 ;
        RECT  16.8 277.5 23.1 278.4 ;
        RECT  8.4 291.9 23.1 292.8 ;
        RECT  18.9 289.2 23.1 290.1 ;
        RECT  8.4 303.0 23.1 303.9 ;
        RECT  21.0 305.7 23.1 306.6 ;
        RECT  10.5 320.1 23.1 321.0 ;
        RECT  14.7 317.4 23.1 318.3 ;
        RECT  10.5 331.2 23.1 332.1 ;
        RECT  16.8 333.9 23.1 334.8 ;
        RECT  10.5 348.3 23.1 349.2 ;
        RECT  18.9 345.6 23.1 346.5 ;
        RECT  10.5 359.4 23.1 360.3 ;
        RECT  21.0 362.1 23.1 363.0 ;
        RECT  12.6 376.5 23.1 377.4 ;
        RECT  14.7 373.8 23.1 374.7 ;
        RECT  12.6 387.6 23.1 388.5 ;
        RECT  16.8 390.3 23.1 391.2 ;
        RECT  12.6 404.7 23.1 405.6 ;
        RECT  18.9 402.0 23.1 402.9 ;
        RECT  12.6 415.8 23.1 416.7 ;
        RECT  21.0 418.5 23.1 419.4 ;
        RECT  40.5 306.0 44.7 306.9 ;
        RECT  40.5 277.8 44.7 278.7 ;
        RECT  40.5 346.2 44.7 347.1 ;
        RECT  40.5 221.4 44.7 222.3 ;
        RECT  40.5 249.6 44.7 250.5 ;
        RECT  40.5 374.4 44.7 375.3 ;
        RECT  40.5 318.0 44.7 318.9 ;
        RECT  40.5 402.6 44.7 403.5 ;
        RECT  40.5 289.8 44.7 290.7 ;
        RECT  40.5 205.2 44.7 206.1 ;
        RECT  40.5 261.6 44.7 262.5 ;
        RECT  40.5 233.4 44.7 234.3 ;
        RECT  40.5 390.6 44.7 391.5 ;
        RECT  40.5 334.2 44.7 335.1 ;
        RECT  40.5 418.8 44.7 419.7 ;
        RECT  40.5 362.4 44.7 363.3 ;
        RECT  6.3 100.05 75.3 100.95 ;
        RECT  6.3 128.25 75.3 129.15 ;
        RECT  6.3 156.45 75.3 157.35 ;
        RECT  6.3 184.65 75.3 185.55 ;
        RECT  6.3 212.85 75.3 213.75 ;
        RECT  6.3 241.05 75.3 241.95 ;
        RECT  6.3 269.25 75.3 270.15 ;
        RECT  6.3 297.45 75.3 298.35 ;
        RECT  6.3 325.65 75.3 326.55 ;
        RECT  6.3 353.85 75.3 354.75 ;
        RECT  6.3 382.05 75.3 382.95 ;
        RECT  6.3 410.25 75.3 411.15 ;
        RECT  6.3 85.95 75.3 86.85 ;
        RECT  6.3 114.15 75.3 115.05 ;
        RECT  6.3 142.35 75.3 143.25 ;
        RECT  6.3 170.55 75.3 171.45 ;
        RECT  6.3 198.75 75.3 199.65 ;
        RECT  6.3 226.95 75.3 227.85 ;
        RECT  6.3 255.15 75.3 256.05 ;
        RECT  6.3 283.35 75.3 284.25 ;
        RECT  6.3 311.55 75.3 312.45 ;
        RECT  6.3 339.75 75.3 340.65 ;
        RECT  6.3 367.95 75.3 368.85 ;
        RECT  6.3 396.15 75.3 397.05 ;
        RECT  6.3 424.35 75.3 425.25 ;
        RECT  31.8 92.4 32.7 93.3 ;
        RECT  31.8 107.7 32.7 108.6 ;
        RECT  31.8 120.6 32.7 121.5 ;
        RECT  31.8 135.9 32.7 136.8 ;
        RECT  55.8 97.8 59.7 98.7 ;
        RECT  58.8 92.4 59.7 97.8 ;
        RECT  69.3 92.4 75.3 93.3 ;
        RECT  52.8 111.9 59.7 112.8 ;
        RECT  58.8 107.7 59.7 111.9 ;
        RECT  69.3 107.7 72.3 108.6 ;
        RECT  49.8 116.4 75.3 117.3 ;
        RECT  46.8 130.5 72.3 131.4 ;
        RECT  44.7 94.5 56.7 95.4 ;
        RECT  44.7 91.8 53.7 92.7 ;
        RECT  44.7 105.6 50.7 106.5 ;
        RECT  44.7 108.3 53.7 109.2 ;
        RECT  44.7 122.7 56.7 123.6 ;
        RECT  44.7 120.0 47.7 120.9 ;
        RECT  44.7 133.8 50.7 134.7 ;
        RECT  44.7 136.5 47.7 137.4 ;
        RECT  23.1 135.9 27.3 136.8 ;
        RECT  23.1 120.6 27.3 121.5 ;
        RECT  23.1 92.4 27.3 93.3 ;
        RECT  23.1 107.7 27.3 108.6 ;
        RECT  22.2 100.05 75.3 100.95 ;
        RECT  22.2 128.25 75.3 129.15 ;
        RECT  22.2 85.95 75.3 86.85 ;
        RECT  22.2 114.15 75.3 115.05 ;
        RECT  22.2 142.35 75.3 143.25 ;
        RECT  61.5 72.75 62.7 75.15 ;
        RECT  61.5 84.15 62.7 85.95 ;
        RECT  66.3 85.05 67.5 85.95 ;
        RECT  66.3 72.75 67.5 73.95 ;
        RECT  63.9 75.0 65.1 83.85 ;
        RECT  67.2 79.5 69.3 80.4 ;
        RECT  59.7 79.5 63.9 80.4 ;
        RECT  59.7 71.85 69.3 72.75 ;
        RECT  59.7 85.95 69.3 86.85 ;
        RECT  66.3 83.85 67.5 85.05 ;
        RECT  63.9 83.85 65.1 85.05 ;
        RECT  66.3 82.65 67.5 83.85 ;
        RECT  63.9 82.65 65.1 83.85 ;
        RECT  66.3 73.95 67.5 75.15 ;
        RECT  63.9 73.95 65.1 75.15 ;
        RECT  66.3 73.95 67.5 75.15 ;
        RECT  63.9 73.95 65.1 75.15 ;
        RECT  61.5 73.95 62.7 75.15 ;
        RECT  61.5 83.85 62.7 85.05 ;
        RECT  66.0 79.35 67.2 80.55 ;
        RECT  61.5 125.85 62.7 128.25 ;
        RECT  61.5 115.05 62.7 116.85 ;
        RECT  66.3 115.05 67.5 115.95 ;
        RECT  66.3 127.05 67.5 128.25 ;
        RECT  63.9 117.15 65.1 126.0 ;
        RECT  67.2 120.6 69.3 121.5 ;
        RECT  59.7 120.6 63.9 121.5 ;
        RECT  59.7 128.25 69.3 129.15 ;
        RECT  59.7 114.15 69.3 115.05 ;
        RECT  66.3 120.75 67.5 121.95 ;
        RECT  63.9 120.75 65.1 121.95 ;
        RECT  66.3 119.55 67.5 120.75 ;
        RECT  63.9 119.55 65.1 120.75 ;
        RECT  66.3 119.85 67.5 121.05 ;
        RECT  63.9 119.85 65.1 121.05 ;
        RECT  66.3 119.85 67.5 121.05 ;
        RECT  63.9 119.85 65.1 121.05 ;
        RECT  61.5 124.65 62.7 125.85 ;
        RECT  61.5 114.75 62.7 115.95 ;
        RECT  66.0 119.25 67.2 120.45 ;
        RECT  24.9 72.75 26.1 75.15 ;
        RECT  24.9 84.15 26.1 85.95 ;
        RECT  29.7 85.05 30.9 85.95 ;
        RECT  29.7 72.75 30.9 73.95 ;
        RECT  27.3 75.0 28.5 83.85 ;
        RECT  30.6 79.5 32.7 80.4 ;
        RECT  23.1 79.5 27.3 80.4 ;
        RECT  23.1 71.85 32.7 72.75 ;
        RECT  23.1 85.95 32.7 86.85 ;
        RECT  29.7 83.85 30.9 85.05 ;
        RECT  27.3 83.85 28.5 85.05 ;
        RECT  29.7 82.65 30.9 83.85 ;
        RECT  27.3 82.65 28.5 83.85 ;
        RECT  29.7 73.95 30.9 75.15 ;
        RECT  27.3 73.95 28.5 75.15 ;
        RECT  29.7 73.95 30.9 75.15 ;
        RECT  27.3 73.95 28.5 75.15 ;
        RECT  24.9 73.95 26.1 75.15 ;
        RECT  24.9 83.85 26.1 85.05 ;
        RECT  29.4 79.35 30.6 80.55 ;
        RECT  24.9 125.85 26.1 128.25 ;
        RECT  24.9 115.05 26.1 116.85 ;
        RECT  29.7 115.05 30.9 115.95 ;
        RECT  29.7 127.05 30.9 128.25 ;
        RECT  27.3 117.15 28.5 126.0 ;
        RECT  30.6 120.6 32.7 121.5 ;
        RECT  23.1 120.6 27.3 121.5 ;
        RECT  23.1 128.25 32.7 129.15 ;
        RECT  23.1 114.15 32.7 115.05 ;
        RECT  29.7 120.75 30.9 121.95 ;
        RECT  27.3 120.75 28.5 121.95 ;
        RECT  29.7 119.55 30.9 120.75 ;
        RECT  27.3 119.55 28.5 120.75 ;
        RECT  29.7 119.85 30.9 121.05 ;
        RECT  27.3 119.85 28.5 121.05 ;
        RECT  29.7 119.85 30.9 121.05 ;
        RECT  27.3 119.85 28.5 121.05 ;
        RECT  24.9 124.65 26.1 125.85 ;
        RECT  24.9 114.75 26.1 115.95 ;
        RECT  29.4 119.25 30.6 120.45 ;
        RECT  24.9 100.95 26.1 103.35 ;
        RECT  24.9 112.35 26.1 114.15 ;
        RECT  29.7 113.25 30.9 114.15 ;
        RECT  29.7 100.95 30.9 102.15 ;
        RECT  27.3 103.2 28.5 112.05 ;
        RECT  30.6 107.7 32.7 108.6 ;
        RECT  23.1 107.7 27.3 108.6 ;
        RECT  23.1 100.05 32.7 100.95 ;
        RECT  23.1 114.15 32.7 115.05 ;
        RECT  29.7 112.05 30.9 113.25 ;
        RECT  27.3 112.05 28.5 113.25 ;
        RECT  29.7 110.85 30.9 112.05 ;
        RECT  27.3 110.85 28.5 112.05 ;
        RECT  29.7 102.15 30.9 103.35 ;
        RECT  27.3 102.15 28.5 103.35 ;
        RECT  29.7 102.15 30.9 103.35 ;
        RECT  27.3 102.15 28.5 103.35 ;
        RECT  24.9 102.15 26.1 103.35 ;
        RECT  24.9 112.05 26.1 113.25 ;
        RECT  29.4 107.55 30.6 108.75 ;
        RECT  24.9 154.05 26.1 156.45 ;
        RECT  24.9 143.25 26.1 145.05 ;
        RECT  29.7 143.25 30.9 144.15 ;
        RECT  29.7 155.25 30.9 156.45 ;
        RECT  27.3 145.35 28.5 154.2 ;
        RECT  30.6 148.8 32.7 149.7 ;
        RECT  23.1 148.8 27.3 149.7 ;
        RECT  23.1 156.45 32.7 157.35 ;
        RECT  23.1 142.35 32.7 143.25 ;
        RECT  29.7 148.95 30.9 150.15 ;
        RECT  27.3 148.95 28.5 150.15 ;
        RECT  29.7 147.75 30.9 148.95 ;
        RECT  27.3 147.75 28.5 148.95 ;
        RECT  29.7 148.05 30.9 149.25 ;
        RECT  27.3 148.05 28.5 149.25 ;
        RECT  29.7 148.05 30.9 149.25 ;
        RECT  27.3 148.05 28.5 149.25 ;
        RECT  24.9 152.85 26.1 154.05 ;
        RECT  24.9 142.95 26.1 144.15 ;
        RECT  29.4 147.45 30.6 148.65 ;
        RECT  34.8 72.3 35.7 75.15 ;
        RECT  34.8 84.0 35.7 86.4 ;
        RECT  41.85 72.3 42.75 75.15 ;
        RECT  37.05 72.3 37.95 75.15 ;
        RECT  41.85 83.55 42.75 86.4 ;
        RECT  36.6 77.4 37.5 78.3 ;
        RECT  39.6 77.4 40.5 78.3 ;
        RECT  36.6 77.85 37.5 84.75 ;
        RECT  37.05 77.4 40.05 78.3 ;
        RECT  39.6 75.15 40.5 77.85 ;
        RECT  42.6 77.4 44.7 78.3 ;
        RECT  32.7 79.5 37.05 80.4 ;
        RECT  39.6 80.1 44.7 81.0 ;
        RECT  32.7 71.85 44.7 72.75 ;
        RECT  32.7 85.95 44.7 86.85 ;
        RECT  41.7 83.55 42.9 84.75 ;
        RECT  39.3 83.55 40.5 84.75 ;
        RECT  41.7 82.35 42.9 83.55 ;
        RECT  39.3 82.35 40.5 83.55 ;
        RECT  39.3 83.55 40.5 84.75 ;
        RECT  36.9 83.55 38.1 84.75 ;
        RECT  39.3 82.35 40.5 83.55 ;
        RECT  36.9 82.35 38.1 83.55 ;
        RECT  41.7 73.95 42.9 75.15 ;
        RECT  39.3 73.95 40.5 75.15 ;
        RECT  41.7 73.95 42.9 75.15 ;
        RECT  39.3 73.95 40.5 75.15 ;
        RECT  39.3 73.95 40.5 75.15 ;
        RECT  36.9 73.95 38.1 75.15 ;
        RECT  39.3 73.95 40.5 75.15 ;
        RECT  36.9 73.95 38.1 75.15 ;
        RECT  34.5 73.95 35.7 75.15 ;
        RECT  34.5 83.55 35.7 84.75 ;
        RECT  41.4 77.4 42.6 78.6 ;
        RECT  38.4 80.1 39.6 81.3 ;
        RECT  34.8 125.85 35.7 128.7 ;
        RECT  34.8 114.6 35.7 117.0 ;
        RECT  41.85 125.85 42.75 128.7 ;
        RECT  37.05 125.85 37.95 128.7 ;
        RECT  41.85 114.6 42.75 117.45 ;
        RECT  36.6 122.7 37.5 123.6 ;
        RECT  39.6 122.7 40.5 123.6 ;
        RECT  36.6 116.25 37.5 123.15 ;
        RECT  37.05 122.7 40.05 123.6 ;
        RECT  39.6 123.15 40.5 125.85 ;
        RECT  42.6 122.7 44.7 123.6 ;
        RECT  32.7 120.6 37.05 121.5 ;
        RECT  39.6 120.0 44.7 120.9 ;
        RECT  32.7 128.25 44.7 129.15 ;
        RECT  32.7 114.15 44.7 115.05 ;
        RECT  41.7 122.25 42.9 123.45 ;
        RECT  39.3 122.25 40.5 123.45 ;
        RECT  41.7 121.05 42.9 122.25 ;
        RECT  39.3 121.05 40.5 122.25 ;
        RECT  39.3 122.25 40.5 123.45 ;
        RECT  36.9 122.25 38.1 123.45 ;
        RECT  39.3 121.05 40.5 122.25 ;
        RECT  36.9 121.05 38.1 122.25 ;
        RECT  41.7 119.85 42.9 121.05 ;
        RECT  39.3 119.85 40.5 121.05 ;
        RECT  41.7 119.85 42.9 121.05 ;
        RECT  39.3 119.85 40.5 121.05 ;
        RECT  39.3 119.85 40.5 121.05 ;
        RECT  36.9 119.85 38.1 121.05 ;
        RECT  39.3 119.85 40.5 121.05 ;
        RECT  36.9 119.85 38.1 121.05 ;
        RECT  34.5 124.65 35.7 125.85 ;
        RECT  34.5 115.05 35.7 116.25 ;
        RECT  41.4 121.2 42.6 122.4 ;
        RECT  38.4 118.5 39.6 119.7 ;
        RECT  34.8 100.5 35.7 103.35 ;
        RECT  34.8 112.2 35.7 114.6 ;
        RECT  41.85 100.5 42.75 103.35 ;
        RECT  37.05 100.5 37.95 103.35 ;
        RECT  41.85 111.75 42.75 114.6 ;
        RECT  36.6 105.6 37.5 106.5 ;
        RECT  39.6 105.6 40.5 106.5 ;
        RECT  36.6 106.05 37.5 112.95 ;
        RECT  37.05 105.6 40.05 106.5 ;
        RECT  39.6 103.35 40.5 106.05 ;
        RECT  42.6 105.6 44.7 106.5 ;
        RECT  32.7 107.7 37.05 108.6 ;
        RECT  39.6 108.3 44.7 109.2 ;
        RECT  32.7 100.05 44.7 100.95 ;
        RECT  32.7 114.15 44.7 115.05 ;
        RECT  41.7 111.75 42.9 112.95 ;
        RECT  39.3 111.75 40.5 112.95 ;
        RECT  41.7 110.55 42.9 111.75 ;
        RECT  39.3 110.55 40.5 111.75 ;
        RECT  39.3 111.75 40.5 112.95 ;
        RECT  36.9 111.75 38.1 112.95 ;
        RECT  39.3 110.55 40.5 111.75 ;
        RECT  36.9 110.55 38.1 111.75 ;
        RECT  41.7 102.15 42.9 103.35 ;
        RECT  39.3 102.15 40.5 103.35 ;
        RECT  41.7 102.15 42.9 103.35 ;
        RECT  39.3 102.15 40.5 103.35 ;
        RECT  39.3 102.15 40.5 103.35 ;
        RECT  36.9 102.15 38.1 103.35 ;
        RECT  39.3 102.15 40.5 103.35 ;
        RECT  36.9 102.15 38.1 103.35 ;
        RECT  34.5 102.15 35.7 103.35 ;
        RECT  34.5 111.75 35.7 112.95 ;
        RECT  41.4 105.6 42.6 106.8 ;
        RECT  38.4 108.3 39.6 109.5 ;
        RECT  34.8 154.05 35.7 156.9 ;
        RECT  34.8 142.8 35.7 145.2 ;
        RECT  41.85 154.05 42.75 156.9 ;
        RECT  37.05 154.05 37.95 156.9 ;
        RECT  41.85 142.8 42.75 145.65 ;
        RECT  36.6 150.9 37.5 151.8 ;
        RECT  39.6 150.9 40.5 151.8 ;
        RECT  36.6 144.45 37.5 151.35 ;
        RECT  37.05 150.9 40.05 151.8 ;
        RECT  39.6 151.35 40.5 154.05 ;
        RECT  42.6 150.9 44.7 151.8 ;
        RECT  32.7 148.8 37.05 149.7 ;
        RECT  39.6 148.2 44.7 149.1 ;
        RECT  32.7 156.45 44.7 157.35 ;
        RECT  32.7 142.35 44.7 143.25 ;
        RECT  41.7 150.45 42.9 151.65 ;
        RECT  39.3 150.45 40.5 151.65 ;
        RECT  41.7 149.25 42.9 150.45 ;
        RECT  39.3 149.25 40.5 150.45 ;
        RECT  39.3 150.45 40.5 151.65 ;
        RECT  36.9 150.45 38.1 151.65 ;
        RECT  39.3 149.25 40.5 150.45 ;
        RECT  36.9 149.25 38.1 150.45 ;
        RECT  41.7 148.05 42.9 149.25 ;
        RECT  39.3 148.05 40.5 149.25 ;
        RECT  41.7 148.05 42.9 149.25 ;
        RECT  39.3 148.05 40.5 149.25 ;
        RECT  39.3 148.05 40.5 149.25 ;
        RECT  36.9 148.05 38.1 149.25 ;
        RECT  39.3 148.05 40.5 149.25 ;
        RECT  36.9 148.05 38.1 149.25 ;
        RECT  34.5 152.85 35.7 154.05 ;
        RECT  34.5 143.25 35.7 144.45 ;
        RECT  41.4 149.4 42.6 150.6 ;
        RECT  38.4 146.7 39.6 147.9 ;
        RECT  55.8 96.45 57.0 97.65 ;
        RECT  74.4 91.05 75.6 92.25 ;
        RECT  52.8 110.55 54.0 111.75 ;
        RECT  71.4 106.35 72.6 107.55 ;
        RECT  74.4 115.05 75.6 116.25 ;
        RECT  49.8 115.05 51.0 116.25 ;
        RECT  71.4 129.15 72.6 130.35 ;
        RECT  46.8 129.15 48.0 130.35 ;
        RECT  55.8 93.15 57.0 94.35 ;
        RECT  52.8 90.45 54.0 91.65 ;
        RECT  49.8 104.25 51.0 105.45 ;
        RECT  52.8 106.95 54.0 108.15 ;
        RECT  55.8 121.35 57.0 122.55 ;
        RECT  46.8 118.65 48.0 119.85 ;
        RECT  49.8 132.45 51.0 133.65 ;
        RECT  46.8 135.15 48.0 136.35 ;
        RECT  31.8 148.8 32.7 149.7 ;
        RECT  31.8 164.1 32.7 165.0 ;
        RECT  31.8 177.0 32.7 177.9 ;
        RECT  31.8 192.3 32.7 193.2 ;
        RECT  55.8 154.2 59.7 155.1 ;
        RECT  58.8 148.8 59.7 154.2 ;
        RECT  69.3 148.8 75.3 149.7 ;
        RECT  52.8 168.3 59.7 169.2 ;
        RECT  58.8 164.1 59.7 168.3 ;
        RECT  69.3 164.1 72.3 165.0 ;
        RECT  49.8 172.8 75.3 173.7 ;
        RECT  46.8 186.9 72.3 187.8 ;
        RECT  44.7 150.9 56.7 151.8 ;
        RECT  44.7 148.2 53.7 149.1 ;
        RECT  44.7 162.0 50.7 162.9 ;
        RECT  44.7 164.7 53.7 165.6 ;
        RECT  44.7 179.1 56.7 180.0 ;
        RECT  44.7 176.4 47.7 177.3 ;
        RECT  44.7 190.2 50.7 191.1 ;
        RECT  44.7 192.9 47.7 193.8 ;
        RECT  23.1 192.3 27.3 193.2 ;
        RECT  23.1 177.0 27.3 177.9 ;
        RECT  23.1 148.8 27.3 149.7 ;
        RECT  23.1 164.1 27.3 165.0 ;
        RECT  22.2 156.45 75.3 157.35 ;
        RECT  22.2 184.65 75.3 185.55 ;
        RECT  22.2 142.35 75.3 143.25 ;
        RECT  22.2 170.55 75.3 171.45 ;
        RECT  22.2 198.75 75.3 199.65 ;
        RECT  61.5 129.15 62.7 131.55 ;
        RECT  61.5 140.55 62.7 142.35 ;
        RECT  66.3 141.45 67.5 142.35 ;
        RECT  66.3 129.15 67.5 130.35 ;
        RECT  63.9 131.4 65.1 140.25 ;
        RECT  67.2 135.9 69.3 136.8 ;
        RECT  59.7 135.9 63.9 136.8 ;
        RECT  59.7 128.25 69.3 129.15 ;
        RECT  59.7 142.35 69.3 143.25 ;
        RECT  66.3 140.25 67.5 141.45 ;
        RECT  63.9 140.25 65.1 141.45 ;
        RECT  66.3 139.05 67.5 140.25 ;
        RECT  63.9 139.05 65.1 140.25 ;
        RECT  66.3 130.35 67.5 131.55 ;
        RECT  63.9 130.35 65.1 131.55 ;
        RECT  66.3 130.35 67.5 131.55 ;
        RECT  63.9 130.35 65.1 131.55 ;
        RECT  61.5 130.35 62.7 131.55 ;
        RECT  61.5 140.25 62.7 141.45 ;
        RECT  66.0 135.75 67.2 136.95 ;
        RECT  61.5 182.25 62.7 184.65 ;
        RECT  61.5 171.45 62.7 173.25 ;
        RECT  66.3 171.45 67.5 172.35 ;
        RECT  66.3 183.45 67.5 184.65 ;
        RECT  63.9 173.55 65.1 182.4 ;
        RECT  67.2 177.0 69.3 177.9 ;
        RECT  59.7 177.0 63.9 177.9 ;
        RECT  59.7 184.65 69.3 185.55 ;
        RECT  59.7 170.55 69.3 171.45 ;
        RECT  66.3 177.15 67.5 178.35 ;
        RECT  63.9 177.15 65.1 178.35 ;
        RECT  66.3 175.95 67.5 177.15 ;
        RECT  63.9 175.95 65.1 177.15 ;
        RECT  66.3 176.25 67.5 177.45 ;
        RECT  63.9 176.25 65.1 177.45 ;
        RECT  66.3 176.25 67.5 177.45 ;
        RECT  63.9 176.25 65.1 177.45 ;
        RECT  61.5 181.05 62.7 182.25 ;
        RECT  61.5 171.15 62.7 172.35 ;
        RECT  66.0 175.65 67.2 176.85 ;
        RECT  24.9 129.15 26.1 131.55 ;
        RECT  24.9 140.55 26.1 142.35 ;
        RECT  29.7 141.45 30.9 142.35 ;
        RECT  29.7 129.15 30.9 130.35 ;
        RECT  27.3 131.4 28.5 140.25 ;
        RECT  30.6 135.9 32.7 136.8 ;
        RECT  23.1 135.9 27.3 136.8 ;
        RECT  23.1 128.25 32.7 129.15 ;
        RECT  23.1 142.35 32.7 143.25 ;
        RECT  29.7 140.25 30.9 141.45 ;
        RECT  27.3 140.25 28.5 141.45 ;
        RECT  29.7 139.05 30.9 140.25 ;
        RECT  27.3 139.05 28.5 140.25 ;
        RECT  29.7 130.35 30.9 131.55 ;
        RECT  27.3 130.35 28.5 131.55 ;
        RECT  29.7 130.35 30.9 131.55 ;
        RECT  27.3 130.35 28.5 131.55 ;
        RECT  24.9 130.35 26.1 131.55 ;
        RECT  24.9 140.25 26.1 141.45 ;
        RECT  29.4 135.75 30.6 136.95 ;
        RECT  24.9 182.25 26.1 184.65 ;
        RECT  24.9 171.45 26.1 173.25 ;
        RECT  29.7 171.45 30.9 172.35 ;
        RECT  29.7 183.45 30.9 184.65 ;
        RECT  27.3 173.55 28.5 182.4 ;
        RECT  30.6 177.0 32.7 177.9 ;
        RECT  23.1 177.0 27.3 177.9 ;
        RECT  23.1 184.65 32.7 185.55 ;
        RECT  23.1 170.55 32.7 171.45 ;
        RECT  29.7 177.15 30.9 178.35 ;
        RECT  27.3 177.15 28.5 178.35 ;
        RECT  29.7 175.95 30.9 177.15 ;
        RECT  27.3 175.95 28.5 177.15 ;
        RECT  29.7 176.25 30.9 177.45 ;
        RECT  27.3 176.25 28.5 177.45 ;
        RECT  29.7 176.25 30.9 177.45 ;
        RECT  27.3 176.25 28.5 177.45 ;
        RECT  24.9 181.05 26.1 182.25 ;
        RECT  24.9 171.15 26.1 172.35 ;
        RECT  29.4 175.65 30.6 176.85 ;
        RECT  24.9 157.35 26.1 159.75 ;
        RECT  24.9 168.75 26.1 170.55 ;
        RECT  29.7 169.65 30.9 170.55 ;
        RECT  29.7 157.35 30.9 158.55 ;
        RECT  27.3 159.6 28.5 168.45 ;
        RECT  30.6 164.1 32.7 165.0 ;
        RECT  23.1 164.1 27.3 165.0 ;
        RECT  23.1 156.45 32.7 157.35 ;
        RECT  23.1 170.55 32.7 171.45 ;
        RECT  29.7 168.45 30.9 169.65 ;
        RECT  27.3 168.45 28.5 169.65 ;
        RECT  29.7 167.25 30.9 168.45 ;
        RECT  27.3 167.25 28.5 168.45 ;
        RECT  29.7 158.55 30.9 159.75 ;
        RECT  27.3 158.55 28.5 159.75 ;
        RECT  29.7 158.55 30.9 159.75 ;
        RECT  27.3 158.55 28.5 159.75 ;
        RECT  24.9 158.55 26.1 159.75 ;
        RECT  24.9 168.45 26.1 169.65 ;
        RECT  29.4 163.95 30.6 165.15 ;
        RECT  24.9 210.45 26.1 212.85 ;
        RECT  24.9 199.65 26.1 201.45 ;
        RECT  29.7 199.65 30.9 200.55 ;
        RECT  29.7 211.65 30.9 212.85 ;
        RECT  27.3 201.75 28.5 210.6 ;
        RECT  30.6 205.2 32.7 206.1 ;
        RECT  23.1 205.2 27.3 206.1 ;
        RECT  23.1 212.85 32.7 213.75 ;
        RECT  23.1 198.75 32.7 199.65 ;
        RECT  29.7 205.35 30.9 206.55 ;
        RECT  27.3 205.35 28.5 206.55 ;
        RECT  29.7 204.15 30.9 205.35 ;
        RECT  27.3 204.15 28.5 205.35 ;
        RECT  29.7 204.45 30.9 205.65 ;
        RECT  27.3 204.45 28.5 205.65 ;
        RECT  29.7 204.45 30.9 205.65 ;
        RECT  27.3 204.45 28.5 205.65 ;
        RECT  24.9 209.25 26.1 210.45 ;
        RECT  24.9 199.35 26.1 200.55 ;
        RECT  29.4 203.85 30.6 205.05 ;
        RECT  34.8 128.7 35.7 131.55 ;
        RECT  34.8 140.4 35.7 142.8 ;
        RECT  41.85 128.7 42.75 131.55 ;
        RECT  37.05 128.7 37.95 131.55 ;
        RECT  41.85 139.95 42.75 142.8 ;
        RECT  36.6 133.8 37.5 134.7 ;
        RECT  39.6 133.8 40.5 134.7 ;
        RECT  36.6 134.25 37.5 141.15 ;
        RECT  37.05 133.8 40.05 134.7 ;
        RECT  39.6 131.55 40.5 134.25 ;
        RECT  42.6 133.8 44.7 134.7 ;
        RECT  32.7 135.9 37.05 136.8 ;
        RECT  39.6 136.5 44.7 137.4 ;
        RECT  32.7 128.25 44.7 129.15 ;
        RECT  32.7 142.35 44.7 143.25 ;
        RECT  41.7 139.95 42.9 141.15 ;
        RECT  39.3 139.95 40.5 141.15 ;
        RECT  41.7 138.75 42.9 139.95 ;
        RECT  39.3 138.75 40.5 139.95 ;
        RECT  39.3 139.95 40.5 141.15 ;
        RECT  36.9 139.95 38.1 141.15 ;
        RECT  39.3 138.75 40.5 139.95 ;
        RECT  36.9 138.75 38.1 139.95 ;
        RECT  41.7 130.35 42.9 131.55 ;
        RECT  39.3 130.35 40.5 131.55 ;
        RECT  41.7 130.35 42.9 131.55 ;
        RECT  39.3 130.35 40.5 131.55 ;
        RECT  39.3 130.35 40.5 131.55 ;
        RECT  36.9 130.35 38.1 131.55 ;
        RECT  39.3 130.35 40.5 131.55 ;
        RECT  36.9 130.35 38.1 131.55 ;
        RECT  34.5 130.35 35.7 131.55 ;
        RECT  34.5 139.95 35.7 141.15 ;
        RECT  41.4 133.8 42.6 135.0 ;
        RECT  38.4 136.5 39.6 137.7 ;
        RECT  34.8 182.25 35.7 185.1 ;
        RECT  34.8 171.0 35.7 173.4 ;
        RECT  41.85 182.25 42.75 185.1 ;
        RECT  37.05 182.25 37.95 185.1 ;
        RECT  41.85 171.0 42.75 173.85 ;
        RECT  36.6 179.1 37.5 180.0 ;
        RECT  39.6 179.1 40.5 180.0 ;
        RECT  36.6 172.65 37.5 179.55 ;
        RECT  37.05 179.1 40.05 180.0 ;
        RECT  39.6 179.55 40.5 182.25 ;
        RECT  42.6 179.1 44.7 180.0 ;
        RECT  32.7 177.0 37.05 177.9 ;
        RECT  39.6 176.4 44.7 177.3 ;
        RECT  32.7 184.65 44.7 185.55 ;
        RECT  32.7 170.55 44.7 171.45 ;
        RECT  41.7 178.65 42.9 179.85 ;
        RECT  39.3 178.65 40.5 179.85 ;
        RECT  41.7 177.45 42.9 178.65 ;
        RECT  39.3 177.45 40.5 178.65 ;
        RECT  39.3 178.65 40.5 179.85 ;
        RECT  36.9 178.65 38.1 179.85 ;
        RECT  39.3 177.45 40.5 178.65 ;
        RECT  36.9 177.45 38.1 178.65 ;
        RECT  41.7 176.25 42.9 177.45 ;
        RECT  39.3 176.25 40.5 177.45 ;
        RECT  41.7 176.25 42.9 177.45 ;
        RECT  39.3 176.25 40.5 177.45 ;
        RECT  39.3 176.25 40.5 177.45 ;
        RECT  36.9 176.25 38.1 177.45 ;
        RECT  39.3 176.25 40.5 177.45 ;
        RECT  36.9 176.25 38.1 177.45 ;
        RECT  34.5 181.05 35.7 182.25 ;
        RECT  34.5 171.45 35.7 172.65 ;
        RECT  41.4 177.6 42.6 178.8 ;
        RECT  38.4 174.9 39.6 176.1 ;
        RECT  34.8 156.9 35.7 159.75 ;
        RECT  34.8 168.6 35.7 171.0 ;
        RECT  41.85 156.9 42.75 159.75 ;
        RECT  37.05 156.9 37.95 159.75 ;
        RECT  41.85 168.15 42.75 171.0 ;
        RECT  36.6 162.0 37.5 162.9 ;
        RECT  39.6 162.0 40.5 162.9 ;
        RECT  36.6 162.45 37.5 169.35 ;
        RECT  37.05 162.0 40.05 162.9 ;
        RECT  39.6 159.75 40.5 162.45 ;
        RECT  42.6 162.0 44.7 162.9 ;
        RECT  32.7 164.1 37.05 165.0 ;
        RECT  39.6 164.7 44.7 165.6 ;
        RECT  32.7 156.45 44.7 157.35 ;
        RECT  32.7 170.55 44.7 171.45 ;
        RECT  41.7 168.15 42.9 169.35 ;
        RECT  39.3 168.15 40.5 169.35 ;
        RECT  41.7 166.95 42.9 168.15 ;
        RECT  39.3 166.95 40.5 168.15 ;
        RECT  39.3 168.15 40.5 169.35 ;
        RECT  36.9 168.15 38.1 169.35 ;
        RECT  39.3 166.95 40.5 168.15 ;
        RECT  36.9 166.95 38.1 168.15 ;
        RECT  41.7 158.55 42.9 159.75 ;
        RECT  39.3 158.55 40.5 159.75 ;
        RECT  41.7 158.55 42.9 159.75 ;
        RECT  39.3 158.55 40.5 159.75 ;
        RECT  39.3 158.55 40.5 159.75 ;
        RECT  36.9 158.55 38.1 159.75 ;
        RECT  39.3 158.55 40.5 159.75 ;
        RECT  36.9 158.55 38.1 159.75 ;
        RECT  34.5 158.55 35.7 159.75 ;
        RECT  34.5 168.15 35.7 169.35 ;
        RECT  41.4 162.0 42.6 163.2 ;
        RECT  38.4 164.7 39.6 165.9 ;
        RECT  34.8 210.45 35.7 213.3 ;
        RECT  34.8 199.2 35.7 201.6 ;
        RECT  41.85 210.45 42.75 213.3 ;
        RECT  37.05 210.45 37.95 213.3 ;
        RECT  41.85 199.2 42.75 202.05 ;
        RECT  36.6 207.3 37.5 208.2 ;
        RECT  39.6 207.3 40.5 208.2 ;
        RECT  36.6 200.85 37.5 207.75 ;
        RECT  37.05 207.3 40.05 208.2 ;
        RECT  39.6 207.75 40.5 210.45 ;
        RECT  42.6 207.3 44.7 208.2 ;
        RECT  32.7 205.2 37.05 206.1 ;
        RECT  39.6 204.6 44.7 205.5 ;
        RECT  32.7 212.85 44.7 213.75 ;
        RECT  32.7 198.75 44.7 199.65 ;
        RECT  41.7 206.85 42.9 208.05 ;
        RECT  39.3 206.85 40.5 208.05 ;
        RECT  41.7 205.65 42.9 206.85 ;
        RECT  39.3 205.65 40.5 206.85 ;
        RECT  39.3 206.85 40.5 208.05 ;
        RECT  36.9 206.85 38.1 208.05 ;
        RECT  39.3 205.65 40.5 206.85 ;
        RECT  36.9 205.65 38.1 206.85 ;
        RECT  41.7 204.45 42.9 205.65 ;
        RECT  39.3 204.45 40.5 205.65 ;
        RECT  41.7 204.45 42.9 205.65 ;
        RECT  39.3 204.45 40.5 205.65 ;
        RECT  39.3 204.45 40.5 205.65 ;
        RECT  36.9 204.45 38.1 205.65 ;
        RECT  39.3 204.45 40.5 205.65 ;
        RECT  36.9 204.45 38.1 205.65 ;
        RECT  34.5 209.25 35.7 210.45 ;
        RECT  34.5 199.65 35.7 200.85 ;
        RECT  41.4 205.8 42.6 207.0 ;
        RECT  38.4 203.1 39.6 204.3 ;
        RECT  55.8 152.85 57.0 154.05 ;
        RECT  74.4 147.45 75.6 148.65 ;
        RECT  52.8 166.95 54.0 168.15 ;
        RECT  71.4 162.75 72.6 163.95 ;
        RECT  74.4 171.45 75.6 172.65 ;
        RECT  49.8 171.45 51.0 172.65 ;
        RECT  71.4 185.55 72.6 186.75 ;
        RECT  46.8 185.55 48.0 186.75 ;
        RECT  55.8 149.55 57.0 150.75 ;
        RECT  52.8 146.85 54.0 148.05 ;
        RECT  49.8 160.65 51.0 161.85 ;
        RECT  52.8 163.35 54.0 164.55 ;
        RECT  55.8 177.75 57.0 178.95 ;
        RECT  46.8 175.05 48.0 176.25 ;
        RECT  49.8 188.85 51.0 190.05 ;
        RECT  46.8 191.55 48.0 192.75 ;
        RECT  32.1 210.45 33.0 213.3 ;
        RECT  32.1 199.2 33.0 201.6 ;
        RECT  25.05 210.45 25.95 213.3 ;
        RECT  29.85 210.45 30.75 213.3 ;
        RECT  25.05 199.2 25.95 202.05 ;
        RECT  30.3 207.3 31.2 208.2 ;
        RECT  27.3 207.3 28.2 208.2 ;
        RECT  30.3 200.85 31.2 207.75 ;
        RECT  27.75 207.3 30.75 208.2 ;
        RECT  27.3 207.75 28.2 210.45 ;
        RECT  23.1 207.3 25.2 208.2 ;
        RECT  30.75 205.2 35.1 206.1 ;
        RECT  23.1 204.6 28.2 205.5 ;
        RECT  23.1 212.85 35.1 213.75 ;
        RECT  23.1 198.75 35.1 199.65 ;
        RECT  24.9 200.85 26.1 202.05 ;
        RECT  27.3 200.85 28.5 202.05 ;
        RECT  24.9 202.05 26.1 203.25 ;
        RECT  27.3 202.05 28.5 203.25 ;
        RECT  27.3 200.85 28.5 202.05 ;
        RECT  29.7 200.85 30.9 202.05 ;
        RECT  27.3 202.05 28.5 203.25 ;
        RECT  29.7 202.05 30.9 203.25 ;
        RECT  24.9 210.45 26.1 211.65 ;
        RECT  27.3 210.45 28.5 211.65 ;
        RECT  24.9 210.45 26.1 211.65 ;
        RECT  27.3 210.45 28.5 211.65 ;
        RECT  27.3 210.45 28.5 211.65 ;
        RECT  29.7 210.45 30.9 211.65 ;
        RECT  27.3 210.45 28.5 211.65 ;
        RECT  29.7 210.45 30.9 211.65 ;
        RECT  32.1 210.45 33.3 211.65 ;
        RECT  32.1 200.85 33.3 202.05 ;
        RECT  25.2 207.0 26.4 208.2 ;
        RECT  28.2 204.3 29.4 205.5 ;
        RECT  32.1 213.3 33.0 216.15 ;
        RECT  32.1 225.0 33.0 227.4 ;
        RECT  25.05 213.3 25.95 216.15 ;
        RECT  29.85 213.3 30.75 216.15 ;
        RECT  25.05 224.55 25.95 227.4 ;
        RECT  30.3 218.4 31.2 219.3 ;
        RECT  27.3 218.4 28.2 219.3 ;
        RECT  30.3 218.85 31.2 225.75 ;
        RECT  27.75 218.4 30.75 219.3 ;
        RECT  27.3 216.15 28.2 218.85 ;
        RECT  23.1 218.4 25.2 219.3 ;
        RECT  30.75 220.5 35.1 221.4 ;
        RECT  23.1 221.1 28.2 222.0 ;
        RECT  23.1 212.85 35.1 213.75 ;
        RECT  23.1 226.95 35.1 227.85 ;
        RECT  24.9 218.55 26.1 219.75 ;
        RECT  27.3 218.55 28.5 219.75 ;
        RECT  24.9 219.75 26.1 220.95 ;
        RECT  27.3 219.75 28.5 220.95 ;
        RECT  27.3 218.55 28.5 219.75 ;
        RECT  29.7 218.55 30.9 219.75 ;
        RECT  27.3 219.75 28.5 220.95 ;
        RECT  29.7 219.75 30.9 220.95 ;
        RECT  24.9 220.95 26.1 222.15 ;
        RECT  27.3 220.95 28.5 222.15 ;
        RECT  24.9 220.95 26.1 222.15 ;
        RECT  27.3 220.95 28.5 222.15 ;
        RECT  27.3 220.95 28.5 222.15 ;
        RECT  29.7 220.95 30.9 222.15 ;
        RECT  27.3 220.95 28.5 222.15 ;
        RECT  29.7 220.95 30.9 222.15 ;
        RECT  32.1 216.15 33.3 217.35 ;
        RECT  32.1 225.75 33.3 226.95 ;
        RECT  25.2 219.6 26.4 220.8 ;
        RECT  28.2 222.3 29.4 223.5 ;
        RECT  32.1 238.65 33.0 241.5 ;
        RECT  32.1 227.4 33.0 229.8 ;
        RECT  25.05 238.65 25.95 241.5 ;
        RECT  29.85 238.65 30.75 241.5 ;
        RECT  25.05 227.4 25.95 230.25 ;
        RECT  30.3 235.5 31.2 236.4 ;
        RECT  27.3 235.5 28.2 236.4 ;
        RECT  30.3 229.05 31.2 235.95 ;
        RECT  27.75 235.5 30.75 236.4 ;
        RECT  27.3 235.95 28.2 238.65 ;
        RECT  23.1 235.5 25.2 236.4 ;
        RECT  30.75 233.4 35.1 234.3 ;
        RECT  23.1 232.8 28.2 233.7 ;
        RECT  23.1 241.05 35.1 241.95 ;
        RECT  23.1 226.95 35.1 227.85 ;
        RECT  24.9 229.05 26.1 230.25 ;
        RECT  27.3 229.05 28.5 230.25 ;
        RECT  24.9 230.25 26.1 231.45 ;
        RECT  27.3 230.25 28.5 231.45 ;
        RECT  27.3 229.05 28.5 230.25 ;
        RECT  29.7 229.05 30.9 230.25 ;
        RECT  27.3 230.25 28.5 231.45 ;
        RECT  29.7 230.25 30.9 231.45 ;
        RECT  24.9 238.65 26.1 239.85 ;
        RECT  27.3 238.65 28.5 239.85 ;
        RECT  24.9 238.65 26.1 239.85 ;
        RECT  27.3 238.65 28.5 239.85 ;
        RECT  27.3 238.65 28.5 239.85 ;
        RECT  29.7 238.65 30.9 239.85 ;
        RECT  27.3 238.65 28.5 239.85 ;
        RECT  29.7 238.65 30.9 239.85 ;
        RECT  32.1 238.65 33.3 239.85 ;
        RECT  32.1 229.05 33.3 230.25 ;
        RECT  25.2 235.2 26.4 236.4 ;
        RECT  28.2 232.5 29.4 233.7 ;
        RECT  32.1 241.5 33.0 244.35 ;
        RECT  32.1 253.2 33.0 255.6 ;
        RECT  25.05 241.5 25.95 244.35 ;
        RECT  29.85 241.5 30.75 244.35 ;
        RECT  25.05 252.75 25.95 255.6 ;
        RECT  30.3 246.6 31.2 247.5 ;
        RECT  27.3 246.6 28.2 247.5 ;
        RECT  30.3 247.05 31.2 253.95 ;
        RECT  27.75 246.6 30.75 247.5 ;
        RECT  27.3 244.35 28.2 247.05 ;
        RECT  23.1 246.6 25.2 247.5 ;
        RECT  30.75 248.7 35.1 249.6 ;
        RECT  23.1 249.3 28.2 250.2 ;
        RECT  23.1 241.05 35.1 241.95 ;
        RECT  23.1 255.15 35.1 256.05 ;
        RECT  24.9 246.75 26.1 247.95 ;
        RECT  27.3 246.75 28.5 247.95 ;
        RECT  24.9 247.95 26.1 249.15 ;
        RECT  27.3 247.95 28.5 249.15 ;
        RECT  27.3 246.75 28.5 247.95 ;
        RECT  29.7 246.75 30.9 247.95 ;
        RECT  27.3 247.95 28.5 249.15 ;
        RECT  29.7 247.95 30.9 249.15 ;
        RECT  24.9 249.15 26.1 250.35 ;
        RECT  27.3 249.15 28.5 250.35 ;
        RECT  24.9 249.15 26.1 250.35 ;
        RECT  27.3 249.15 28.5 250.35 ;
        RECT  27.3 249.15 28.5 250.35 ;
        RECT  29.7 249.15 30.9 250.35 ;
        RECT  27.3 249.15 28.5 250.35 ;
        RECT  29.7 249.15 30.9 250.35 ;
        RECT  32.1 244.35 33.3 245.55 ;
        RECT  32.1 253.95 33.3 255.15 ;
        RECT  25.2 247.8 26.4 249.0 ;
        RECT  28.2 250.5 29.4 251.7 ;
        RECT  32.1 266.85 33.0 269.7 ;
        RECT  32.1 255.6 33.0 258.0 ;
        RECT  25.05 266.85 25.95 269.7 ;
        RECT  29.85 266.85 30.75 269.7 ;
        RECT  25.05 255.6 25.95 258.45 ;
        RECT  30.3 263.7 31.2 264.6 ;
        RECT  27.3 263.7 28.2 264.6 ;
        RECT  30.3 257.25 31.2 264.15 ;
        RECT  27.75 263.7 30.75 264.6 ;
        RECT  27.3 264.15 28.2 266.85 ;
        RECT  23.1 263.7 25.2 264.6 ;
        RECT  30.75 261.6 35.1 262.5 ;
        RECT  23.1 261.0 28.2 261.9 ;
        RECT  23.1 269.25 35.1 270.15 ;
        RECT  23.1 255.15 35.1 256.05 ;
        RECT  24.9 257.25 26.1 258.45 ;
        RECT  27.3 257.25 28.5 258.45 ;
        RECT  24.9 258.45 26.1 259.65 ;
        RECT  27.3 258.45 28.5 259.65 ;
        RECT  27.3 257.25 28.5 258.45 ;
        RECT  29.7 257.25 30.9 258.45 ;
        RECT  27.3 258.45 28.5 259.65 ;
        RECT  29.7 258.45 30.9 259.65 ;
        RECT  24.9 266.85 26.1 268.05 ;
        RECT  27.3 266.85 28.5 268.05 ;
        RECT  24.9 266.85 26.1 268.05 ;
        RECT  27.3 266.85 28.5 268.05 ;
        RECT  27.3 266.85 28.5 268.05 ;
        RECT  29.7 266.85 30.9 268.05 ;
        RECT  27.3 266.85 28.5 268.05 ;
        RECT  29.7 266.85 30.9 268.05 ;
        RECT  32.1 266.85 33.3 268.05 ;
        RECT  32.1 257.25 33.3 258.45 ;
        RECT  25.2 263.4 26.4 264.6 ;
        RECT  28.2 260.7 29.4 261.9 ;
        RECT  32.1 269.7 33.0 272.55 ;
        RECT  32.1 281.4 33.0 283.8 ;
        RECT  25.05 269.7 25.95 272.55 ;
        RECT  29.85 269.7 30.75 272.55 ;
        RECT  25.05 280.95 25.95 283.8 ;
        RECT  30.3 274.8 31.2 275.7 ;
        RECT  27.3 274.8 28.2 275.7 ;
        RECT  30.3 275.25 31.2 282.15 ;
        RECT  27.75 274.8 30.75 275.7 ;
        RECT  27.3 272.55 28.2 275.25 ;
        RECT  23.1 274.8 25.2 275.7 ;
        RECT  30.75 276.9 35.1 277.8 ;
        RECT  23.1 277.5 28.2 278.4 ;
        RECT  23.1 269.25 35.1 270.15 ;
        RECT  23.1 283.35 35.1 284.25 ;
        RECT  24.9 274.95 26.1 276.15 ;
        RECT  27.3 274.95 28.5 276.15 ;
        RECT  24.9 276.15 26.1 277.35 ;
        RECT  27.3 276.15 28.5 277.35 ;
        RECT  27.3 274.95 28.5 276.15 ;
        RECT  29.7 274.95 30.9 276.15 ;
        RECT  27.3 276.15 28.5 277.35 ;
        RECT  29.7 276.15 30.9 277.35 ;
        RECT  24.9 277.35 26.1 278.55 ;
        RECT  27.3 277.35 28.5 278.55 ;
        RECT  24.9 277.35 26.1 278.55 ;
        RECT  27.3 277.35 28.5 278.55 ;
        RECT  27.3 277.35 28.5 278.55 ;
        RECT  29.7 277.35 30.9 278.55 ;
        RECT  27.3 277.35 28.5 278.55 ;
        RECT  29.7 277.35 30.9 278.55 ;
        RECT  32.1 272.55 33.3 273.75 ;
        RECT  32.1 282.15 33.3 283.35 ;
        RECT  25.2 276.0 26.4 277.2 ;
        RECT  28.2 278.7 29.4 279.9 ;
        RECT  32.1 295.05 33.0 297.9 ;
        RECT  32.1 283.8 33.0 286.2 ;
        RECT  25.05 295.05 25.95 297.9 ;
        RECT  29.85 295.05 30.75 297.9 ;
        RECT  25.05 283.8 25.95 286.65 ;
        RECT  30.3 291.9 31.2 292.8 ;
        RECT  27.3 291.9 28.2 292.8 ;
        RECT  30.3 285.45 31.2 292.35 ;
        RECT  27.75 291.9 30.75 292.8 ;
        RECT  27.3 292.35 28.2 295.05 ;
        RECT  23.1 291.9 25.2 292.8 ;
        RECT  30.75 289.8 35.1 290.7 ;
        RECT  23.1 289.2 28.2 290.1 ;
        RECT  23.1 297.45 35.1 298.35 ;
        RECT  23.1 283.35 35.1 284.25 ;
        RECT  24.9 285.45 26.1 286.65 ;
        RECT  27.3 285.45 28.5 286.65 ;
        RECT  24.9 286.65 26.1 287.85 ;
        RECT  27.3 286.65 28.5 287.85 ;
        RECT  27.3 285.45 28.5 286.65 ;
        RECT  29.7 285.45 30.9 286.65 ;
        RECT  27.3 286.65 28.5 287.85 ;
        RECT  29.7 286.65 30.9 287.85 ;
        RECT  24.9 295.05 26.1 296.25 ;
        RECT  27.3 295.05 28.5 296.25 ;
        RECT  24.9 295.05 26.1 296.25 ;
        RECT  27.3 295.05 28.5 296.25 ;
        RECT  27.3 295.05 28.5 296.25 ;
        RECT  29.7 295.05 30.9 296.25 ;
        RECT  27.3 295.05 28.5 296.25 ;
        RECT  29.7 295.05 30.9 296.25 ;
        RECT  32.1 295.05 33.3 296.25 ;
        RECT  32.1 285.45 33.3 286.65 ;
        RECT  25.2 291.6 26.4 292.8 ;
        RECT  28.2 288.9 29.4 290.1 ;
        RECT  32.1 297.9 33.0 300.75 ;
        RECT  32.1 309.6 33.0 312.0 ;
        RECT  25.05 297.9 25.95 300.75 ;
        RECT  29.85 297.9 30.75 300.75 ;
        RECT  25.05 309.15 25.95 312.0 ;
        RECT  30.3 303.0 31.2 303.9 ;
        RECT  27.3 303.0 28.2 303.9 ;
        RECT  30.3 303.45 31.2 310.35 ;
        RECT  27.75 303.0 30.75 303.9 ;
        RECT  27.3 300.75 28.2 303.45 ;
        RECT  23.1 303.0 25.2 303.9 ;
        RECT  30.75 305.1 35.1 306.0 ;
        RECT  23.1 305.7 28.2 306.6 ;
        RECT  23.1 297.45 35.1 298.35 ;
        RECT  23.1 311.55 35.1 312.45 ;
        RECT  24.9 303.15 26.1 304.35 ;
        RECT  27.3 303.15 28.5 304.35 ;
        RECT  24.9 304.35 26.1 305.55 ;
        RECT  27.3 304.35 28.5 305.55 ;
        RECT  27.3 303.15 28.5 304.35 ;
        RECT  29.7 303.15 30.9 304.35 ;
        RECT  27.3 304.35 28.5 305.55 ;
        RECT  29.7 304.35 30.9 305.55 ;
        RECT  24.9 305.55 26.1 306.75 ;
        RECT  27.3 305.55 28.5 306.75 ;
        RECT  24.9 305.55 26.1 306.75 ;
        RECT  27.3 305.55 28.5 306.75 ;
        RECT  27.3 305.55 28.5 306.75 ;
        RECT  29.7 305.55 30.9 306.75 ;
        RECT  27.3 305.55 28.5 306.75 ;
        RECT  29.7 305.55 30.9 306.75 ;
        RECT  32.1 300.75 33.3 301.95 ;
        RECT  32.1 310.35 33.3 311.55 ;
        RECT  25.2 304.2 26.4 305.4 ;
        RECT  28.2 306.9 29.4 308.1 ;
        RECT  32.1 323.25 33.0 326.1 ;
        RECT  32.1 312.0 33.0 314.4 ;
        RECT  25.05 323.25 25.95 326.1 ;
        RECT  29.85 323.25 30.75 326.1 ;
        RECT  25.05 312.0 25.95 314.85 ;
        RECT  30.3 320.1 31.2 321.0 ;
        RECT  27.3 320.1 28.2 321.0 ;
        RECT  30.3 313.65 31.2 320.55 ;
        RECT  27.75 320.1 30.75 321.0 ;
        RECT  27.3 320.55 28.2 323.25 ;
        RECT  23.1 320.1 25.2 321.0 ;
        RECT  30.75 318.0 35.1 318.9 ;
        RECT  23.1 317.4 28.2 318.3 ;
        RECT  23.1 325.65 35.1 326.55 ;
        RECT  23.1 311.55 35.1 312.45 ;
        RECT  24.9 313.65 26.1 314.85 ;
        RECT  27.3 313.65 28.5 314.85 ;
        RECT  24.9 314.85 26.1 316.05 ;
        RECT  27.3 314.85 28.5 316.05 ;
        RECT  27.3 313.65 28.5 314.85 ;
        RECT  29.7 313.65 30.9 314.85 ;
        RECT  27.3 314.85 28.5 316.05 ;
        RECT  29.7 314.85 30.9 316.05 ;
        RECT  24.9 323.25 26.1 324.45 ;
        RECT  27.3 323.25 28.5 324.45 ;
        RECT  24.9 323.25 26.1 324.45 ;
        RECT  27.3 323.25 28.5 324.45 ;
        RECT  27.3 323.25 28.5 324.45 ;
        RECT  29.7 323.25 30.9 324.45 ;
        RECT  27.3 323.25 28.5 324.45 ;
        RECT  29.7 323.25 30.9 324.45 ;
        RECT  32.1 323.25 33.3 324.45 ;
        RECT  32.1 313.65 33.3 314.85 ;
        RECT  25.2 319.8 26.4 321.0 ;
        RECT  28.2 317.1 29.4 318.3 ;
        RECT  32.1 326.1 33.0 328.95 ;
        RECT  32.1 337.8 33.0 340.2 ;
        RECT  25.05 326.1 25.95 328.95 ;
        RECT  29.85 326.1 30.75 328.95 ;
        RECT  25.05 337.35 25.95 340.2 ;
        RECT  30.3 331.2 31.2 332.1 ;
        RECT  27.3 331.2 28.2 332.1 ;
        RECT  30.3 331.65 31.2 338.55 ;
        RECT  27.75 331.2 30.75 332.1 ;
        RECT  27.3 328.95 28.2 331.65 ;
        RECT  23.1 331.2 25.2 332.1 ;
        RECT  30.75 333.3 35.1 334.2 ;
        RECT  23.1 333.9 28.2 334.8 ;
        RECT  23.1 325.65 35.1 326.55 ;
        RECT  23.1 339.75 35.1 340.65 ;
        RECT  24.9 331.35 26.1 332.55 ;
        RECT  27.3 331.35 28.5 332.55 ;
        RECT  24.9 332.55 26.1 333.75 ;
        RECT  27.3 332.55 28.5 333.75 ;
        RECT  27.3 331.35 28.5 332.55 ;
        RECT  29.7 331.35 30.9 332.55 ;
        RECT  27.3 332.55 28.5 333.75 ;
        RECT  29.7 332.55 30.9 333.75 ;
        RECT  24.9 333.75 26.1 334.95 ;
        RECT  27.3 333.75 28.5 334.95 ;
        RECT  24.9 333.75 26.1 334.95 ;
        RECT  27.3 333.75 28.5 334.95 ;
        RECT  27.3 333.75 28.5 334.95 ;
        RECT  29.7 333.75 30.9 334.95 ;
        RECT  27.3 333.75 28.5 334.95 ;
        RECT  29.7 333.75 30.9 334.95 ;
        RECT  32.1 328.95 33.3 330.15 ;
        RECT  32.1 338.55 33.3 339.75 ;
        RECT  25.2 332.4 26.4 333.6 ;
        RECT  28.2 335.1 29.4 336.3 ;
        RECT  32.1 351.45 33.0 354.3 ;
        RECT  32.1 340.2 33.0 342.6 ;
        RECT  25.05 351.45 25.95 354.3 ;
        RECT  29.85 351.45 30.75 354.3 ;
        RECT  25.05 340.2 25.95 343.05 ;
        RECT  30.3 348.3 31.2 349.2 ;
        RECT  27.3 348.3 28.2 349.2 ;
        RECT  30.3 341.85 31.2 348.75 ;
        RECT  27.75 348.3 30.75 349.2 ;
        RECT  27.3 348.75 28.2 351.45 ;
        RECT  23.1 348.3 25.2 349.2 ;
        RECT  30.75 346.2 35.1 347.1 ;
        RECT  23.1 345.6 28.2 346.5 ;
        RECT  23.1 353.85 35.1 354.75 ;
        RECT  23.1 339.75 35.1 340.65 ;
        RECT  24.9 341.85 26.1 343.05 ;
        RECT  27.3 341.85 28.5 343.05 ;
        RECT  24.9 343.05 26.1 344.25 ;
        RECT  27.3 343.05 28.5 344.25 ;
        RECT  27.3 341.85 28.5 343.05 ;
        RECT  29.7 341.85 30.9 343.05 ;
        RECT  27.3 343.05 28.5 344.25 ;
        RECT  29.7 343.05 30.9 344.25 ;
        RECT  24.9 351.45 26.1 352.65 ;
        RECT  27.3 351.45 28.5 352.65 ;
        RECT  24.9 351.45 26.1 352.65 ;
        RECT  27.3 351.45 28.5 352.65 ;
        RECT  27.3 351.45 28.5 352.65 ;
        RECT  29.7 351.45 30.9 352.65 ;
        RECT  27.3 351.45 28.5 352.65 ;
        RECT  29.7 351.45 30.9 352.65 ;
        RECT  32.1 351.45 33.3 352.65 ;
        RECT  32.1 341.85 33.3 343.05 ;
        RECT  25.2 348.0 26.4 349.2 ;
        RECT  28.2 345.3 29.4 346.5 ;
        RECT  32.1 354.3 33.0 357.15 ;
        RECT  32.1 366.0 33.0 368.4 ;
        RECT  25.05 354.3 25.95 357.15 ;
        RECT  29.85 354.3 30.75 357.15 ;
        RECT  25.05 365.55 25.95 368.4 ;
        RECT  30.3 359.4 31.2 360.3 ;
        RECT  27.3 359.4 28.2 360.3 ;
        RECT  30.3 359.85 31.2 366.75 ;
        RECT  27.75 359.4 30.75 360.3 ;
        RECT  27.3 357.15 28.2 359.85 ;
        RECT  23.1 359.4 25.2 360.3 ;
        RECT  30.75 361.5 35.1 362.4 ;
        RECT  23.1 362.1 28.2 363.0 ;
        RECT  23.1 353.85 35.1 354.75 ;
        RECT  23.1 367.95 35.1 368.85 ;
        RECT  24.9 359.55 26.1 360.75 ;
        RECT  27.3 359.55 28.5 360.75 ;
        RECT  24.9 360.75 26.1 361.95 ;
        RECT  27.3 360.75 28.5 361.95 ;
        RECT  27.3 359.55 28.5 360.75 ;
        RECT  29.7 359.55 30.9 360.75 ;
        RECT  27.3 360.75 28.5 361.95 ;
        RECT  29.7 360.75 30.9 361.95 ;
        RECT  24.9 361.95 26.1 363.15 ;
        RECT  27.3 361.95 28.5 363.15 ;
        RECT  24.9 361.95 26.1 363.15 ;
        RECT  27.3 361.95 28.5 363.15 ;
        RECT  27.3 361.95 28.5 363.15 ;
        RECT  29.7 361.95 30.9 363.15 ;
        RECT  27.3 361.95 28.5 363.15 ;
        RECT  29.7 361.95 30.9 363.15 ;
        RECT  32.1 357.15 33.3 358.35 ;
        RECT  32.1 366.75 33.3 367.95 ;
        RECT  25.2 360.6 26.4 361.8 ;
        RECT  28.2 363.3 29.4 364.5 ;
        RECT  32.1 379.65 33.0 382.5 ;
        RECT  32.1 368.4 33.0 370.8 ;
        RECT  25.05 379.65 25.95 382.5 ;
        RECT  29.85 379.65 30.75 382.5 ;
        RECT  25.05 368.4 25.95 371.25 ;
        RECT  30.3 376.5 31.2 377.4 ;
        RECT  27.3 376.5 28.2 377.4 ;
        RECT  30.3 370.05 31.2 376.95 ;
        RECT  27.75 376.5 30.75 377.4 ;
        RECT  27.3 376.95 28.2 379.65 ;
        RECT  23.1 376.5 25.2 377.4 ;
        RECT  30.75 374.4 35.1 375.3 ;
        RECT  23.1 373.8 28.2 374.7 ;
        RECT  23.1 382.05 35.1 382.95 ;
        RECT  23.1 367.95 35.1 368.85 ;
        RECT  24.9 370.05 26.1 371.25 ;
        RECT  27.3 370.05 28.5 371.25 ;
        RECT  24.9 371.25 26.1 372.45 ;
        RECT  27.3 371.25 28.5 372.45 ;
        RECT  27.3 370.05 28.5 371.25 ;
        RECT  29.7 370.05 30.9 371.25 ;
        RECT  27.3 371.25 28.5 372.45 ;
        RECT  29.7 371.25 30.9 372.45 ;
        RECT  24.9 379.65 26.1 380.85 ;
        RECT  27.3 379.65 28.5 380.85 ;
        RECT  24.9 379.65 26.1 380.85 ;
        RECT  27.3 379.65 28.5 380.85 ;
        RECT  27.3 379.65 28.5 380.85 ;
        RECT  29.7 379.65 30.9 380.85 ;
        RECT  27.3 379.65 28.5 380.85 ;
        RECT  29.7 379.65 30.9 380.85 ;
        RECT  32.1 379.65 33.3 380.85 ;
        RECT  32.1 370.05 33.3 371.25 ;
        RECT  25.2 376.2 26.4 377.4 ;
        RECT  28.2 373.5 29.4 374.7 ;
        RECT  32.1 382.5 33.0 385.35 ;
        RECT  32.1 394.2 33.0 396.6 ;
        RECT  25.05 382.5 25.95 385.35 ;
        RECT  29.85 382.5 30.75 385.35 ;
        RECT  25.05 393.75 25.95 396.6 ;
        RECT  30.3 387.6 31.2 388.5 ;
        RECT  27.3 387.6 28.2 388.5 ;
        RECT  30.3 388.05 31.2 394.95 ;
        RECT  27.75 387.6 30.75 388.5 ;
        RECT  27.3 385.35 28.2 388.05 ;
        RECT  23.1 387.6 25.2 388.5 ;
        RECT  30.75 389.7 35.1 390.6 ;
        RECT  23.1 390.3 28.2 391.2 ;
        RECT  23.1 382.05 35.1 382.95 ;
        RECT  23.1 396.15 35.1 397.05 ;
        RECT  24.9 387.75 26.1 388.95 ;
        RECT  27.3 387.75 28.5 388.95 ;
        RECT  24.9 388.95 26.1 390.15 ;
        RECT  27.3 388.95 28.5 390.15 ;
        RECT  27.3 387.75 28.5 388.95 ;
        RECT  29.7 387.75 30.9 388.95 ;
        RECT  27.3 388.95 28.5 390.15 ;
        RECT  29.7 388.95 30.9 390.15 ;
        RECT  24.9 390.15 26.1 391.35 ;
        RECT  27.3 390.15 28.5 391.35 ;
        RECT  24.9 390.15 26.1 391.35 ;
        RECT  27.3 390.15 28.5 391.35 ;
        RECT  27.3 390.15 28.5 391.35 ;
        RECT  29.7 390.15 30.9 391.35 ;
        RECT  27.3 390.15 28.5 391.35 ;
        RECT  29.7 390.15 30.9 391.35 ;
        RECT  32.1 385.35 33.3 386.55 ;
        RECT  32.1 394.95 33.3 396.15 ;
        RECT  25.2 388.8 26.4 390.0 ;
        RECT  28.2 391.5 29.4 392.7 ;
        RECT  32.1 407.85 33.0 410.7 ;
        RECT  32.1 396.6 33.0 399.0 ;
        RECT  25.05 407.85 25.95 410.7 ;
        RECT  29.85 407.85 30.75 410.7 ;
        RECT  25.05 396.6 25.95 399.45 ;
        RECT  30.3 404.7 31.2 405.6 ;
        RECT  27.3 404.7 28.2 405.6 ;
        RECT  30.3 398.25 31.2 405.15 ;
        RECT  27.75 404.7 30.75 405.6 ;
        RECT  27.3 405.15 28.2 407.85 ;
        RECT  23.1 404.7 25.2 405.6 ;
        RECT  30.75 402.6 35.1 403.5 ;
        RECT  23.1 402.0 28.2 402.9 ;
        RECT  23.1 410.25 35.1 411.15 ;
        RECT  23.1 396.15 35.1 397.05 ;
        RECT  24.9 398.25 26.1 399.45 ;
        RECT  27.3 398.25 28.5 399.45 ;
        RECT  24.9 399.45 26.1 400.65 ;
        RECT  27.3 399.45 28.5 400.65 ;
        RECT  27.3 398.25 28.5 399.45 ;
        RECT  29.7 398.25 30.9 399.45 ;
        RECT  27.3 399.45 28.5 400.65 ;
        RECT  29.7 399.45 30.9 400.65 ;
        RECT  24.9 407.85 26.1 409.05 ;
        RECT  27.3 407.85 28.5 409.05 ;
        RECT  24.9 407.85 26.1 409.05 ;
        RECT  27.3 407.85 28.5 409.05 ;
        RECT  27.3 407.85 28.5 409.05 ;
        RECT  29.7 407.85 30.9 409.05 ;
        RECT  27.3 407.85 28.5 409.05 ;
        RECT  29.7 407.85 30.9 409.05 ;
        RECT  32.1 407.85 33.3 409.05 ;
        RECT  32.1 398.25 33.3 399.45 ;
        RECT  25.2 404.4 26.4 405.6 ;
        RECT  28.2 401.7 29.4 402.9 ;
        RECT  32.1 410.7 33.0 413.55 ;
        RECT  32.1 422.4 33.0 424.8 ;
        RECT  25.05 410.7 25.95 413.55 ;
        RECT  29.85 410.7 30.75 413.55 ;
        RECT  25.05 421.95 25.95 424.8 ;
        RECT  30.3 415.8 31.2 416.7 ;
        RECT  27.3 415.8 28.2 416.7 ;
        RECT  30.3 416.25 31.2 423.15 ;
        RECT  27.75 415.8 30.75 416.7 ;
        RECT  27.3 413.55 28.2 416.25 ;
        RECT  23.1 415.8 25.2 416.7 ;
        RECT  30.75 417.9 35.1 418.8 ;
        RECT  23.1 418.5 28.2 419.4 ;
        RECT  23.1 410.25 35.1 411.15 ;
        RECT  23.1 424.35 35.1 425.25 ;
        RECT  24.9 415.95 26.1 417.15 ;
        RECT  27.3 415.95 28.5 417.15 ;
        RECT  24.9 417.15 26.1 418.35 ;
        RECT  27.3 417.15 28.5 418.35 ;
        RECT  27.3 415.95 28.5 417.15 ;
        RECT  29.7 415.95 30.9 417.15 ;
        RECT  27.3 417.15 28.5 418.35 ;
        RECT  29.7 417.15 30.9 418.35 ;
        RECT  24.9 418.35 26.1 419.55 ;
        RECT  27.3 418.35 28.5 419.55 ;
        RECT  24.9 418.35 26.1 419.55 ;
        RECT  27.3 418.35 28.5 419.55 ;
        RECT  27.3 418.35 28.5 419.55 ;
        RECT  29.7 418.35 30.9 419.55 ;
        RECT  27.3 418.35 28.5 419.55 ;
        RECT  29.7 418.35 30.9 419.55 ;
        RECT  32.1 413.55 33.3 414.75 ;
        RECT  32.1 423.15 33.3 424.35 ;
        RECT  25.2 417.0 26.4 418.2 ;
        RECT  28.2 419.7 29.4 420.9 ;
        RECT  41.7 210.45 42.9 212.85 ;
        RECT  41.7 199.65 42.9 201.45 ;
        RECT  36.9 199.65 38.1 200.55 ;
        RECT  36.9 211.65 38.1 212.85 ;
        RECT  39.3 201.75 40.5 210.6 ;
        RECT  35.1 205.2 37.2 206.1 ;
        RECT  40.5 205.2 44.7 206.1 ;
        RECT  35.1 212.85 44.7 213.75 ;
        RECT  35.1 198.75 44.7 199.65 ;
        RECT  36.9 200.55 38.1 201.75 ;
        RECT  39.3 200.55 40.5 201.75 ;
        RECT  36.9 201.75 38.1 202.95 ;
        RECT  39.3 201.75 40.5 202.95 ;
        RECT  36.9 210.45 38.1 211.65 ;
        RECT  39.3 210.45 40.5 211.65 ;
        RECT  36.9 210.45 38.1 211.65 ;
        RECT  39.3 210.45 40.5 211.65 ;
        RECT  41.7 210.45 42.9 211.65 ;
        RECT  41.7 200.55 42.9 201.75 ;
        RECT  37.2 205.05 38.4 206.25 ;
        RECT  41.7 213.75 42.9 216.15 ;
        RECT  41.7 225.15 42.9 226.95 ;
        RECT  36.9 226.05 38.1 226.95 ;
        RECT  36.9 213.75 38.1 214.95 ;
        RECT  39.3 216.0 40.5 224.85 ;
        RECT  35.1 220.5 37.2 221.4 ;
        RECT  40.5 220.5 44.7 221.4 ;
        RECT  35.1 212.85 44.7 213.75 ;
        RECT  35.1 226.95 44.7 227.85 ;
        RECT  36.9 220.05 38.1 221.25 ;
        RECT  39.3 220.05 40.5 221.25 ;
        RECT  36.9 221.25 38.1 222.45 ;
        RECT  39.3 221.25 40.5 222.45 ;
        RECT  36.9 220.95 38.1 222.15 ;
        RECT  39.3 220.95 40.5 222.15 ;
        RECT  36.9 220.95 38.1 222.15 ;
        RECT  39.3 220.95 40.5 222.15 ;
        RECT  41.7 216.15 42.9 217.35 ;
        RECT  41.7 226.05 42.9 227.25 ;
        RECT  37.2 221.55 38.4 222.75 ;
        RECT  41.7 238.65 42.9 241.05 ;
        RECT  41.7 227.85 42.9 229.65 ;
        RECT  36.9 227.85 38.1 228.75 ;
        RECT  36.9 239.85 38.1 241.05 ;
        RECT  39.3 229.95 40.5 238.8 ;
        RECT  35.1 233.4 37.2 234.3 ;
        RECT  40.5 233.4 44.7 234.3 ;
        RECT  35.1 241.05 44.7 241.95 ;
        RECT  35.1 226.95 44.7 227.85 ;
        RECT  36.9 228.75 38.1 229.95 ;
        RECT  39.3 228.75 40.5 229.95 ;
        RECT  36.9 229.95 38.1 231.15 ;
        RECT  39.3 229.95 40.5 231.15 ;
        RECT  36.9 238.65 38.1 239.85 ;
        RECT  39.3 238.65 40.5 239.85 ;
        RECT  36.9 238.65 38.1 239.85 ;
        RECT  39.3 238.65 40.5 239.85 ;
        RECT  41.7 238.65 42.9 239.85 ;
        RECT  41.7 228.75 42.9 229.95 ;
        RECT  37.2 233.25 38.4 234.45 ;
        RECT  41.7 241.95 42.9 244.35 ;
        RECT  41.7 253.35 42.9 255.15 ;
        RECT  36.9 254.25 38.1 255.15 ;
        RECT  36.9 241.95 38.1 243.15 ;
        RECT  39.3 244.2 40.5 253.05 ;
        RECT  35.1 248.7 37.2 249.6 ;
        RECT  40.5 248.7 44.7 249.6 ;
        RECT  35.1 241.05 44.7 241.95 ;
        RECT  35.1 255.15 44.7 256.05 ;
        RECT  36.9 248.25 38.1 249.45 ;
        RECT  39.3 248.25 40.5 249.45 ;
        RECT  36.9 249.45 38.1 250.65 ;
        RECT  39.3 249.45 40.5 250.65 ;
        RECT  36.9 249.15 38.1 250.35 ;
        RECT  39.3 249.15 40.5 250.35 ;
        RECT  36.9 249.15 38.1 250.35 ;
        RECT  39.3 249.15 40.5 250.35 ;
        RECT  41.7 244.35 42.9 245.55 ;
        RECT  41.7 254.25 42.9 255.45 ;
        RECT  37.2 249.75 38.4 250.95 ;
        RECT  41.7 266.85 42.9 269.25 ;
        RECT  41.7 256.05 42.9 257.85 ;
        RECT  36.9 256.05 38.1 256.95 ;
        RECT  36.9 268.05 38.1 269.25 ;
        RECT  39.3 258.15 40.5 267.0 ;
        RECT  35.1 261.6 37.2 262.5 ;
        RECT  40.5 261.6 44.7 262.5 ;
        RECT  35.1 269.25 44.7 270.15 ;
        RECT  35.1 255.15 44.7 256.05 ;
        RECT  36.9 256.95 38.1 258.15 ;
        RECT  39.3 256.95 40.5 258.15 ;
        RECT  36.9 258.15 38.1 259.35 ;
        RECT  39.3 258.15 40.5 259.35 ;
        RECT  36.9 266.85 38.1 268.05 ;
        RECT  39.3 266.85 40.5 268.05 ;
        RECT  36.9 266.85 38.1 268.05 ;
        RECT  39.3 266.85 40.5 268.05 ;
        RECT  41.7 266.85 42.9 268.05 ;
        RECT  41.7 256.95 42.9 258.15 ;
        RECT  37.2 261.45 38.4 262.65 ;
        RECT  41.7 270.15 42.9 272.55 ;
        RECT  41.7 281.55 42.9 283.35 ;
        RECT  36.9 282.45 38.1 283.35 ;
        RECT  36.9 270.15 38.1 271.35 ;
        RECT  39.3 272.4 40.5 281.25 ;
        RECT  35.1 276.9 37.2 277.8 ;
        RECT  40.5 276.9 44.7 277.8 ;
        RECT  35.1 269.25 44.7 270.15 ;
        RECT  35.1 283.35 44.7 284.25 ;
        RECT  36.9 276.45 38.1 277.65 ;
        RECT  39.3 276.45 40.5 277.65 ;
        RECT  36.9 277.65 38.1 278.85 ;
        RECT  39.3 277.65 40.5 278.85 ;
        RECT  36.9 277.35 38.1 278.55 ;
        RECT  39.3 277.35 40.5 278.55 ;
        RECT  36.9 277.35 38.1 278.55 ;
        RECT  39.3 277.35 40.5 278.55 ;
        RECT  41.7 272.55 42.9 273.75 ;
        RECT  41.7 282.45 42.9 283.65 ;
        RECT  37.2 277.95 38.4 279.15 ;
        RECT  41.7 295.05 42.9 297.45 ;
        RECT  41.7 284.25 42.9 286.05 ;
        RECT  36.9 284.25 38.1 285.15 ;
        RECT  36.9 296.25 38.1 297.45 ;
        RECT  39.3 286.35 40.5 295.2 ;
        RECT  35.1 289.8 37.2 290.7 ;
        RECT  40.5 289.8 44.7 290.7 ;
        RECT  35.1 297.45 44.7 298.35 ;
        RECT  35.1 283.35 44.7 284.25 ;
        RECT  36.9 285.15 38.1 286.35 ;
        RECT  39.3 285.15 40.5 286.35 ;
        RECT  36.9 286.35 38.1 287.55 ;
        RECT  39.3 286.35 40.5 287.55 ;
        RECT  36.9 295.05 38.1 296.25 ;
        RECT  39.3 295.05 40.5 296.25 ;
        RECT  36.9 295.05 38.1 296.25 ;
        RECT  39.3 295.05 40.5 296.25 ;
        RECT  41.7 295.05 42.9 296.25 ;
        RECT  41.7 285.15 42.9 286.35 ;
        RECT  37.2 289.65 38.4 290.85 ;
        RECT  41.7 298.35 42.9 300.75 ;
        RECT  41.7 309.75 42.9 311.55 ;
        RECT  36.9 310.65 38.1 311.55 ;
        RECT  36.9 298.35 38.1 299.55 ;
        RECT  39.3 300.6 40.5 309.45 ;
        RECT  35.1 305.1 37.2 306.0 ;
        RECT  40.5 305.1 44.7 306.0 ;
        RECT  35.1 297.45 44.7 298.35 ;
        RECT  35.1 311.55 44.7 312.45 ;
        RECT  36.9 304.65 38.1 305.85 ;
        RECT  39.3 304.65 40.5 305.85 ;
        RECT  36.9 305.85 38.1 307.05 ;
        RECT  39.3 305.85 40.5 307.05 ;
        RECT  36.9 305.55 38.1 306.75 ;
        RECT  39.3 305.55 40.5 306.75 ;
        RECT  36.9 305.55 38.1 306.75 ;
        RECT  39.3 305.55 40.5 306.75 ;
        RECT  41.7 300.75 42.9 301.95 ;
        RECT  41.7 310.65 42.9 311.85 ;
        RECT  37.2 306.15 38.4 307.35 ;
        RECT  41.7 323.25 42.9 325.65 ;
        RECT  41.7 312.45 42.9 314.25 ;
        RECT  36.9 312.45 38.1 313.35 ;
        RECT  36.9 324.45 38.1 325.65 ;
        RECT  39.3 314.55 40.5 323.4 ;
        RECT  35.1 318.0 37.2 318.9 ;
        RECT  40.5 318.0 44.7 318.9 ;
        RECT  35.1 325.65 44.7 326.55 ;
        RECT  35.1 311.55 44.7 312.45 ;
        RECT  36.9 313.35 38.1 314.55 ;
        RECT  39.3 313.35 40.5 314.55 ;
        RECT  36.9 314.55 38.1 315.75 ;
        RECT  39.3 314.55 40.5 315.75 ;
        RECT  36.9 323.25 38.1 324.45 ;
        RECT  39.3 323.25 40.5 324.45 ;
        RECT  36.9 323.25 38.1 324.45 ;
        RECT  39.3 323.25 40.5 324.45 ;
        RECT  41.7 323.25 42.9 324.45 ;
        RECT  41.7 313.35 42.9 314.55 ;
        RECT  37.2 317.85 38.4 319.05 ;
        RECT  41.7 326.55 42.9 328.95 ;
        RECT  41.7 337.95 42.9 339.75 ;
        RECT  36.9 338.85 38.1 339.75 ;
        RECT  36.9 326.55 38.1 327.75 ;
        RECT  39.3 328.8 40.5 337.65 ;
        RECT  35.1 333.3 37.2 334.2 ;
        RECT  40.5 333.3 44.7 334.2 ;
        RECT  35.1 325.65 44.7 326.55 ;
        RECT  35.1 339.75 44.7 340.65 ;
        RECT  36.9 332.85 38.1 334.05 ;
        RECT  39.3 332.85 40.5 334.05 ;
        RECT  36.9 334.05 38.1 335.25 ;
        RECT  39.3 334.05 40.5 335.25 ;
        RECT  36.9 333.75 38.1 334.95 ;
        RECT  39.3 333.75 40.5 334.95 ;
        RECT  36.9 333.75 38.1 334.95 ;
        RECT  39.3 333.75 40.5 334.95 ;
        RECT  41.7 328.95 42.9 330.15 ;
        RECT  41.7 338.85 42.9 340.05 ;
        RECT  37.2 334.35 38.4 335.55 ;
        RECT  41.7 351.45 42.9 353.85 ;
        RECT  41.7 340.65 42.9 342.45 ;
        RECT  36.9 340.65 38.1 341.55 ;
        RECT  36.9 352.65 38.1 353.85 ;
        RECT  39.3 342.75 40.5 351.6 ;
        RECT  35.1 346.2 37.2 347.1 ;
        RECT  40.5 346.2 44.7 347.1 ;
        RECT  35.1 353.85 44.7 354.75 ;
        RECT  35.1 339.75 44.7 340.65 ;
        RECT  36.9 341.55 38.1 342.75 ;
        RECT  39.3 341.55 40.5 342.75 ;
        RECT  36.9 342.75 38.1 343.95 ;
        RECT  39.3 342.75 40.5 343.95 ;
        RECT  36.9 351.45 38.1 352.65 ;
        RECT  39.3 351.45 40.5 352.65 ;
        RECT  36.9 351.45 38.1 352.65 ;
        RECT  39.3 351.45 40.5 352.65 ;
        RECT  41.7 351.45 42.9 352.65 ;
        RECT  41.7 341.55 42.9 342.75 ;
        RECT  37.2 346.05 38.4 347.25 ;
        RECT  41.7 354.75 42.9 357.15 ;
        RECT  41.7 366.15 42.9 367.95 ;
        RECT  36.9 367.05 38.1 367.95 ;
        RECT  36.9 354.75 38.1 355.95 ;
        RECT  39.3 357.0 40.5 365.85 ;
        RECT  35.1 361.5 37.2 362.4 ;
        RECT  40.5 361.5 44.7 362.4 ;
        RECT  35.1 353.85 44.7 354.75 ;
        RECT  35.1 367.95 44.7 368.85 ;
        RECT  36.9 361.05 38.1 362.25 ;
        RECT  39.3 361.05 40.5 362.25 ;
        RECT  36.9 362.25 38.1 363.45 ;
        RECT  39.3 362.25 40.5 363.45 ;
        RECT  36.9 361.95 38.1 363.15 ;
        RECT  39.3 361.95 40.5 363.15 ;
        RECT  36.9 361.95 38.1 363.15 ;
        RECT  39.3 361.95 40.5 363.15 ;
        RECT  41.7 357.15 42.9 358.35 ;
        RECT  41.7 367.05 42.9 368.25 ;
        RECT  37.2 362.55 38.4 363.75 ;
        RECT  41.7 379.65 42.9 382.05 ;
        RECT  41.7 368.85 42.9 370.65 ;
        RECT  36.9 368.85 38.1 369.75 ;
        RECT  36.9 380.85 38.1 382.05 ;
        RECT  39.3 370.95 40.5 379.8 ;
        RECT  35.1 374.4 37.2 375.3 ;
        RECT  40.5 374.4 44.7 375.3 ;
        RECT  35.1 382.05 44.7 382.95 ;
        RECT  35.1 367.95 44.7 368.85 ;
        RECT  36.9 369.75 38.1 370.95 ;
        RECT  39.3 369.75 40.5 370.95 ;
        RECT  36.9 370.95 38.1 372.15 ;
        RECT  39.3 370.95 40.5 372.15 ;
        RECT  36.9 379.65 38.1 380.85 ;
        RECT  39.3 379.65 40.5 380.85 ;
        RECT  36.9 379.65 38.1 380.85 ;
        RECT  39.3 379.65 40.5 380.85 ;
        RECT  41.7 379.65 42.9 380.85 ;
        RECT  41.7 369.75 42.9 370.95 ;
        RECT  37.2 374.25 38.4 375.45 ;
        RECT  41.7 382.95 42.9 385.35 ;
        RECT  41.7 394.35 42.9 396.15 ;
        RECT  36.9 395.25 38.1 396.15 ;
        RECT  36.9 382.95 38.1 384.15 ;
        RECT  39.3 385.2 40.5 394.05 ;
        RECT  35.1 389.7 37.2 390.6 ;
        RECT  40.5 389.7 44.7 390.6 ;
        RECT  35.1 382.05 44.7 382.95 ;
        RECT  35.1 396.15 44.7 397.05 ;
        RECT  36.9 389.25 38.1 390.45 ;
        RECT  39.3 389.25 40.5 390.45 ;
        RECT  36.9 390.45 38.1 391.65 ;
        RECT  39.3 390.45 40.5 391.65 ;
        RECT  36.9 390.15 38.1 391.35 ;
        RECT  39.3 390.15 40.5 391.35 ;
        RECT  36.9 390.15 38.1 391.35 ;
        RECT  39.3 390.15 40.5 391.35 ;
        RECT  41.7 385.35 42.9 386.55 ;
        RECT  41.7 395.25 42.9 396.45 ;
        RECT  37.2 390.75 38.4 391.95 ;
        RECT  41.7 407.85 42.9 410.25 ;
        RECT  41.7 397.05 42.9 398.85 ;
        RECT  36.9 397.05 38.1 397.95 ;
        RECT  36.9 409.05 38.1 410.25 ;
        RECT  39.3 399.15 40.5 408.0 ;
        RECT  35.1 402.6 37.2 403.5 ;
        RECT  40.5 402.6 44.7 403.5 ;
        RECT  35.1 410.25 44.7 411.15 ;
        RECT  35.1 396.15 44.7 397.05 ;
        RECT  36.9 397.95 38.1 399.15 ;
        RECT  39.3 397.95 40.5 399.15 ;
        RECT  36.9 399.15 38.1 400.35 ;
        RECT  39.3 399.15 40.5 400.35 ;
        RECT  36.9 407.85 38.1 409.05 ;
        RECT  39.3 407.85 40.5 409.05 ;
        RECT  36.9 407.85 38.1 409.05 ;
        RECT  39.3 407.85 40.5 409.05 ;
        RECT  41.7 407.85 42.9 409.05 ;
        RECT  41.7 397.95 42.9 399.15 ;
        RECT  37.2 402.45 38.4 403.65 ;
        RECT  41.7 411.15 42.9 413.55 ;
        RECT  41.7 422.55 42.9 424.35 ;
        RECT  36.9 423.45 38.1 424.35 ;
        RECT  36.9 411.15 38.1 412.35 ;
        RECT  39.3 413.4 40.5 422.25 ;
        RECT  35.1 417.9 37.2 418.8 ;
        RECT  40.5 417.9 44.7 418.8 ;
        RECT  35.1 410.25 44.7 411.15 ;
        RECT  35.1 424.35 44.7 425.25 ;
        RECT  36.9 417.45 38.1 418.65 ;
        RECT  39.3 417.45 40.5 418.65 ;
        RECT  36.9 418.65 38.1 419.85 ;
        RECT  39.3 418.65 40.5 419.85 ;
        RECT  36.9 418.35 38.1 419.55 ;
        RECT  39.3 418.35 40.5 419.55 ;
        RECT  36.9 418.35 38.1 419.55 ;
        RECT  39.3 418.35 40.5 419.55 ;
        RECT  41.7 413.55 42.9 414.75 ;
        RECT  41.7 423.45 42.9 424.65 ;
        RECT  37.2 418.95 38.4 420.15 ;
        RECT  6.3 92.4 7.5 93.6 ;
        RECT  8.4 107.7 9.6 108.9 ;
        RECT  10.5 120.6 11.7 121.8 ;
        RECT  12.6 135.9 13.8 137.1 ;
        RECT  14.7 148.8 15.9 150.0 ;
        RECT  16.8 164.1 18.0 165.3 ;
        RECT  18.9 177.0 20.1 178.2 ;
        RECT  21.0 192.3 22.2 193.5 ;
        RECT  6.3 207.3 7.5 208.5 ;
        RECT  14.7 204.6 15.9 205.8 ;
        RECT  6.3 218.4 7.5 219.6 ;
        RECT  16.8 221.1 18.0 222.3 ;
        RECT  6.3 235.5 7.5 236.7 ;
        RECT  18.9 232.8 20.1 234.0 ;
        RECT  6.3 246.6 7.5 247.8 ;
        RECT  21.0 249.3 22.2 250.5 ;
        RECT  8.4 263.7 9.6 264.9 ;
        RECT  14.7 261.0 15.9 262.2 ;
        RECT  8.4 274.8 9.6 276.0 ;
        RECT  16.8 277.5 18.0 278.7 ;
        RECT  8.4 291.9 9.6 293.1 ;
        RECT  18.9 289.2 20.1 290.4 ;
        RECT  8.4 303.0 9.6 304.2 ;
        RECT  21.0 305.7 22.2 306.9 ;
        RECT  10.5 320.1 11.7 321.3 ;
        RECT  14.7 317.4 15.9 318.6 ;
        RECT  10.5 331.2 11.7 332.4 ;
        RECT  16.8 333.9 18.0 335.1 ;
        RECT  10.5 348.3 11.7 349.5 ;
        RECT  18.9 345.6 20.1 346.8 ;
        RECT  10.5 359.4 11.7 360.6 ;
        RECT  21.0 362.1 22.2 363.3 ;
        RECT  12.6 376.5 13.8 377.7 ;
        RECT  14.7 373.8 15.9 375.0 ;
        RECT  12.6 387.6 13.8 388.8 ;
        RECT  16.8 390.3 18.0 391.5 ;
        RECT  12.6 404.7 13.8 405.9 ;
        RECT  18.9 402.0 20.1 403.2 ;
        RECT  12.6 415.8 13.8 417.0 ;
        RECT  21.0 418.5 22.2 419.7 ;
        RECT  47.85 205.2 51.0 206.1 ;
        RECT  60.15 205.2 61.05 206.1 ;
        RECT  60.15 204.6 61.05 205.5 ;
        RECT  56.4 205.2 60.6 206.1 ;
        RECT  60.15 205.05 61.05 205.65 ;
        RECT  60.6 204.6 65.7 205.5 ;
        RECT  68.25 205.2 72.6 206.1 ;
        RECT  72.6 205.2 74.7 206.1 ;
        RECT  47.85 220.5 51.0 221.4 ;
        RECT  60.15 220.5 61.05 221.4 ;
        RECT  60.15 221.1 61.05 222.0 ;
        RECT  56.4 220.5 60.6 221.4 ;
        RECT  60.15 220.95 61.05 221.55 ;
        RECT  60.6 221.1 65.7 222.0 ;
        RECT  68.25 220.5 72.6 221.4 ;
        RECT  72.6 220.5 74.7 221.4 ;
        RECT  47.85 233.4 51.0 234.3 ;
        RECT  60.15 233.4 61.05 234.3 ;
        RECT  60.15 232.8 61.05 233.7 ;
        RECT  56.4 233.4 60.6 234.3 ;
        RECT  60.15 233.25 61.05 233.85 ;
        RECT  60.6 232.8 65.7 233.7 ;
        RECT  68.25 233.4 72.6 234.3 ;
        RECT  72.6 233.4 74.7 234.3 ;
        RECT  47.85 248.7 51.0 249.6 ;
        RECT  60.15 248.7 61.05 249.6 ;
        RECT  60.15 249.3 61.05 250.2 ;
        RECT  56.4 248.7 60.6 249.6 ;
        RECT  60.15 249.15 61.05 249.75 ;
        RECT  60.6 249.3 65.7 250.2 ;
        RECT  68.25 248.7 72.6 249.6 ;
        RECT  72.6 248.7 74.7 249.6 ;
        RECT  47.85 261.6 51.0 262.5 ;
        RECT  60.15 261.6 61.05 262.5 ;
        RECT  60.15 261.0 61.05 261.9 ;
        RECT  56.4 261.6 60.6 262.5 ;
        RECT  60.15 261.45 61.05 262.05 ;
        RECT  60.6 261.0 65.7 261.9 ;
        RECT  68.25 261.6 72.6 262.5 ;
        RECT  72.6 261.6 74.7 262.5 ;
        RECT  47.85 276.9 51.0 277.8 ;
        RECT  60.15 276.9 61.05 277.8 ;
        RECT  60.15 277.5 61.05 278.4 ;
        RECT  56.4 276.9 60.6 277.8 ;
        RECT  60.15 277.35 61.05 277.95 ;
        RECT  60.6 277.5 65.7 278.4 ;
        RECT  68.25 276.9 72.6 277.8 ;
        RECT  72.6 276.9 74.7 277.8 ;
        RECT  47.85 289.8 51.0 290.7 ;
        RECT  60.15 289.8 61.05 290.7 ;
        RECT  60.15 289.2 61.05 290.1 ;
        RECT  56.4 289.8 60.6 290.7 ;
        RECT  60.15 289.65 61.05 290.25 ;
        RECT  60.6 289.2 65.7 290.1 ;
        RECT  68.25 289.8 72.6 290.7 ;
        RECT  72.6 289.8 74.7 290.7 ;
        RECT  47.85 305.1 51.0 306.0 ;
        RECT  60.15 305.1 61.05 306.0 ;
        RECT  60.15 305.7 61.05 306.6 ;
        RECT  56.4 305.1 60.6 306.0 ;
        RECT  60.15 305.55 61.05 306.15 ;
        RECT  60.6 305.7 65.7 306.6 ;
        RECT  68.25 305.1 72.6 306.0 ;
        RECT  72.6 305.1 74.7 306.0 ;
        RECT  47.85 318.0 51.0 318.9 ;
        RECT  60.15 318.0 61.05 318.9 ;
        RECT  60.15 317.4 61.05 318.3 ;
        RECT  56.4 318.0 60.6 318.9 ;
        RECT  60.15 317.85 61.05 318.45 ;
        RECT  60.6 317.4 65.7 318.3 ;
        RECT  68.25 318.0 72.6 318.9 ;
        RECT  72.6 318.0 74.7 318.9 ;
        RECT  47.85 333.3 51.0 334.2 ;
        RECT  60.15 333.3 61.05 334.2 ;
        RECT  60.15 333.9 61.05 334.8 ;
        RECT  56.4 333.3 60.6 334.2 ;
        RECT  60.15 333.75 61.05 334.35 ;
        RECT  60.6 333.9 65.7 334.8 ;
        RECT  68.25 333.3 72.6 334.2 ;
        RECT  72.6 333.3 74.7 334.2 ;
        RECT  47.85 346.2 51.0 347.1 ;
        RECT  60.15 346.2 61.05 347.1 ;
        RECT  60.15 345.6 61.05 346.5 ;
        RECT  56.4 346.2 60.6 347.1 ;
        RECT  60.15 346.05 61.05 346.65 ;
        RECT  60.6 345.6 65.7 346.5 ;
        RECT  68.25 346.2 72.6 347.1 ;
        RECT  72.6 346.2 74.7 347.1 ;
        RECT  47.85 361.5 51.0 362.4 ;
        RECT  60.15 361.5 61.05 362.4 ;
        RECT  60.15 362.1 61.05 363.0 ;
        RECT  56.4 361.5 60.6 362.4 ;
        RECT  60.15 361.95 61.05 362.55 ;
        RECT  60.6 362.1 65.7 363.0 ;
        RECT  68.25 361.5 72.6 362.4 ;
        RECT  72.6 361.5 74.7 362.4 ;
        RECT  47.85 374.4 51.0 375.3 ;
        RECT  60.15 374.4 61.05 375.3 ;
        RECT  60.15 373.8 61.05 374.7 ;
        RECT  56.4 374.4 60.6 375.3 ;
        RECT  60.15 374.25 61.05 374.85 ;
        RECT  60.6 373.8 65.7 374.7 ;
        RECT  68.25 374.4 72.6 375.3 ;
        RECT  72.6 374.4 74.7 375.3 ;
        RECT  47.85 389.7 51.0 390.6 ;
        RECT  60.15 389.7 61.05 390.6 ;
        RECT  60.15 390.3 61.05 391.2 ;
        RECT  56.4 389.7 60.6 390.6 ;
        RECT  60.15 390.15 61.05 390.75 ;
        RECT  60.6 390.3 65.7 391.2 ;
        RECT  68.25 389.7 72.6 390.6 ;
        RECT  72.6 389.7 74.7 390.6 ;
        RECT  47.85 402.6 51.0 403.5 ;
        RECT  60.15 402.6 61.05 403.5 ;
        RECT  60.15 402.0 61.05 402.9 ;
        RECT  56.4 402.6 60.6 403.5 ;
        RECT  60.15 402.45 61.05 403.05 ;
        RECT  60.6 402.0 65.7 402.9 ;
        RECT  68.25 402.6 72.6 403.5 ;
        RECT  72.6 402.6 74.7 403.5 ;
        RECT  47.85 417.9 51.0 418.8 ;
        RECT  60.15 417.9 61.05 418.8 ;
        RECT  60.15 418.5 61.05 419.4 ;
        RECT  56.4 417.9 60.6 418.8 ;
        RECT  60.15 418.35 61.05 418.95 ;
        RECT  60.6 418.5 65.7 419.4 ;
        RECT  68.25 417.9 72.6 418.8 ;
        RECT  72.6 417.9 74.7 418.8 ;
        RECT  81.3 261.6 82.2 262.5 ;
        RECT  44.7 246.6 49.8 247.5 ;
        RECT  81.3 205.2 82.2 206.1 ;
        RECT  44.7 303.0 49.8 303.9 ;
        RECT  81.3 233.4 82.2 234.3 ;
        RECT  44.7 218.4 49.8 219.3 ;
        RECT  44.7 274.8 49.8 275.7 ;
        RECT  44.7 320.1 49.8 321.0 ;
        RECT  81.3 417.9 82.2 418.8 ;
        RECT  44.7 348.3 49.8 349.2 ;
        RECT  81.3 318.0 82.2 318.9 ;
        RECT  44.7 404.7 49.8 405.6 ;
        RECT  44.7 376.5 49.8 377.4 ;
        RECT  81.3 289.8 82.2 290.7 ;
        RECT  81.3 389.7 82.2 390.6 ;
        RECT  81.3 361.5 82.2 362.4 ;
        RECT  81.3 248.7 82.2 249.6 ;
        RECT  44.7 235.5 49.8 236.4 ;
        RECT  81.3 276.9 82.2 277.8 ;
        RECT  81.3 220.5 82.2 221.4 ;
        RECT  44.7 207.3 49.8 208.2 ;
        RECT  44.7 263.7 49.8 264.6 ;
        RECT  44.7 291.9 49.8 292.8 ;
        RECT  44.7 331.2 49.8 332.1 ;
        RECT  44.7 359.4 49.8 360.3 ;
        RECT  81.3 402.6 82.2 403.5 ;
        RECT  44.7 415.8 49.8 416.7 ;
        RECT  81.3 346.2 82.2 347.1 ;
        RECT  81.3 333.3 82.2 334.2 ;
        RECT  44.7 212.85 51.0 213.75 ;
        RECT  44.7 241.05 51.0 241.95 ;
        RECT  44.7 269.25 51.0 270.15 ;
        RECT  44.7 297.45 51.0 298.35 ;
        RECT  44.7 325.65 51.0 326.55 ;
        RECT  44.7 353.85 51.0 354.75 ;
        RECT  44.7 382.05 51.0 382.95 ;
        RECT  44.7 410.25 51.0 411.15 ;
        RECT  44.7 198.75 51.0 199.65 ;
        RECT  44.7 226.95 51.0 227.85 ;
        RECT  44.7 255.15 51.0 256.05 ;
        RECT  44.7 283.35 51.0 284.25 ;
        RECT  44.7 311.55 51.0 312.45 ;
        RECT  44.7 339.75 51.0 340.65 ;
        RECT  44.7 367.95 51.0 368.85 ;
        RECT  44.7 396.15 51.0 397.05 ;
        RECT  44.7 424.35 51.0 425.25 ;
        RECT  44.7 387.6 49.8 388.5 ;
        RECT  81.3 374.4 82.2 375.3 ;
        RECT  81.3 305.1 82.2 306.0 ;
        RECT  57.6 210.45 58.8 212.85 ;
        RECT  57.6 199.65 58.8 201.45 ;
        RECT  52.8 199.65 54.0 200.55 ;
        RECT  52.8 211.65 54.0 212.85 ;
        RECT  55.2 201.75 56.4 210.6 ;
        RECT  51.0 205.2 53.1 206.1 ;
        RECT  56.4 205.2 60.6 206.1 ;
        RECT  51.0 212.85 60.6 213.75 ;
        RECT  51.0 198.75 60.6 199.65 ;
        RECT  52.8 200.55 54.0 201.75 ;
        RECT  55.2 200.55 56.4 201.75 ;
        RECT  52.8 201.75 54.0 202.95 ;
        RECT  55.2 201.75 56.4 202.95 ;
        RECT  52.8 210.45 54.0 211.65 ;
        RECT  55.2 210.45 56.4 211.65 ;
        RECT  52.8 210.45 54.0 211.65 ;
        RECT  55.2 210.45 56.4 211.65 ;
        RECT  57.6 210.45 58.8 211.65 ;
        RECT  57.6 200.55 58.8 201.75 ;
        RECT  53.1 205.05 54.3 206.25 ;
        RECT  69.6 210.45 70.5 213.3 ;
        RECT  69.6 199.2 70.5 201.6 ;
        RECT  62.55 210.45 63.45 213.3 ;
        RECT  67.35 210.45 68.25 213.3 ;
        RECT  62.55 199.2 63.45 202.05 ;
        RECT  67.8 207.3 68.7 208.2 ;
        RECT  64.8 207.3 65.7 208.2 ;
        RECT  67.8 200.85 68.7 207.75 ;
        RECT  65.25 207.3 68.25 208.2 ;
        RECT  64.8 207.75 65.7 210.45 ;
        RECT  60.6 207.3 62.7 208.2 ;
        RECT  68.25 205.2 72.6 206.1 ;
        RECT  60.6 204.6 65.7 205.5 ;
        RECT  60.6 212.85 72.6 213.75 ;
        RECT  60.6 198.75 72.6 199.65 ;
        RECT  62.4 200.85 63.6 202.05 ;
        RECT  64.8 200.85 66.0 202.05 ;
        RECT  62.4 202.05 63.6 203.25 ;
        RECT  64.8 202.05 66.0 203.25 ;
        RECT  64.8 200.85 66.0 202.05 ;
        RECT  67.2 200.85 68.4 202.05 ;
        RECT  64.8 202.05 66.0 203.25 ;
        RECT  67.2 202.05 68.4 203.25 ;
        RECT  62.4 210.45 63.6 211.65 ;
        RECT  64.8 210.45 66.0 211.65 ;
        RECT  62.4 210.45 63.6 211.65 ;
        RECT  64.8 210.45 66.0 211.65 ;
        RECT  64.8 210.45 66.0 211.65 ;
        RECT  67.2 210.45 68.4 211.65 ;
        RECT  64.8 210.45 66.0 211.65 ;
        RECT  67.2 210.45 68.4 211.65 ;
        RECT  69.6 210.45 70.8 211.65 ;
        RECT  69.6 200.85 70.8 202.05 ;
        RECT  62.7 207.0 63.9 208.2 ;
        RECT  65.7 204.3 66.9 205.5 ;
        RECT  79.2 210.45 80.4 212.85 ;
        RECT  79.2 199.65 80.4 201.45 ;
        RECT  74.4 199.65 75.6 200.55 ;
        RECT  74.4 211.65 75.6 212.85 ;
        RECT  76.8 201.75 78.0 210.6 ;
        RECT  72.6 205.2 74.7 206.1 ;
        RECT  78.0 205.2 82.2 206.1 ;
        RECT  72.6 212.85 82.2 213.75 ;
        RECT  72.6 198.75 82.2 199.65 ;
        RECT  74.4 200.55 75.6 201.75 ;
        RECT  76.8 200.55 78.0 201.75 ;
        RECT  74.4 201.75 75.6 202.95 ;
        RECT  76.8 201.75 78.0 202.95 ;
        RECT  74.4 210.45 75.6 211.65 ;
        RECT  76.8 210.45 78.0 211.65 ;
        RECT  74.4 210.45 75.6 211.65 ;
        RECT  76.8 210.45 78.0 211.65 ;
        RECT  79.2 210.45 80.4 211.65 ;
        RECT  79.2 200.55 80.4 201.75 ;
        RECT  74.7 205.05 75.9 206.25 ;
        RECT  47.25 205.05 48.45 206.25 ;
        RECT  49.2 207.15 50.4 208.35 ;
        RECT  60.6 207.15 61.8 208.35 ;
        RECT  57.6 213.75 58.8 216.15 ;
        RECT  57.6 225.15 58.8 226.95 ;
        RECT  52.8 226.05 54.0 226.95 ;
        RECT  52.8 213.75 54.0 214.95 ;
        RECT  55.2 216.0 56.4 224.85 ;
        RECT  51.0 220.5 53.1 221.4 ;
        RECT  56.4 220.5 60.6 221.4 ;
        RECT  51.0 212.85 60.6 213.75 ;
        RECT  51.0 226.95 60.6 227.85 ;
        RECT  52.8 220.05 54.0 221.25 ;
        RECT  55.2 220.05 56.4 221.25 ;
        RECT  52.8 221.25 54.0 222.45 ;
        RECT  55.2 221.25 56.4 222.45 ;
        RECT  52.8 220.95 54.0 222.15 ;
        RECT  55.2 220.95 56.4 222.15 ;
        RECT  52.8 220.95 54.0 222.15 ;
        RECT  55.2 220.95 56.4 222.15 ;
        RECT  57.6 216.15 58.8 217.35 ;
        RECT  57.6 226.05 58.8 227.25 ;
        RECT  53.1 221.55 54.3 222.75 ;
        RECT  69.6 213.3 70.5 216.15 ;
        RECT  69.6 225.0 70.5 227.4 ;
        RECT  62.55 213.3 63.45 216.15 ;
        RECT  67.35 213.3 68.25 216.15 ;
        RECT  62.55 224.55 63.45 227.4 ;
        RECT  67.8 218.4 68.7 219.3 ;
        RECT  64.8 218.4 65.7 219.3 ;
        RECT  67.8 218.85 68.7 225.75 ;
        RECT  65.25 218.4 68.25 219.3 ;
        RECT  64.8 216.15 65.7 218.85 ;
        RECT  60.6 218.4 62.7 219.3 ;
        RECT  68.25 220.5 72.6 221.4 ;
        RECT  60.6 221.1 65.7 222.0 ;
        RECT  60.6 212.85 72.6 213.75 ;
        RECT  60.6 226.95 72.6 227.85 ;
        RECT  62.4 218.55 63.6 219.75 ;
        RECT  64.8 218.55 66.0 219.75 ;
        RECT  62.4 219.75 63.6 220.95 ;
        RECT  64.8 219.75 66.0 220.95 ;
        RECT  64.8 218.55 66.0 219.75 ;
        RECT  67.2 218.55 68.4 219.75 ;
        RECT  64.8 219.75 66.0 220.95 ;
        RECT  67.2 219.75 68.4 220.95 ;
        RECT  62.4 220.95 63.6 222.15 ;
        RECT  64.8 220.95 66.0 222.15 ;
        RECT  62.4 220.95 63.6 222.15 ;
        RECT  64.8 220.95 66.0 222.15 ;
        RECT  64.8 220.95 66.0 222.15 ;
        RECT  67.2 220.95 68.4 222.15 ;
        RECT  64.8 220.95 66.0 222.15 ;
        RECT  67.2 220.95 68.4 222.15 ;
        RECT  69.6 216.15 70.8 217.35 ;
        RECT  69.6 225.75 70.8 226.95 ;
        RECT  62.7 219.6 63.9 220.8 ;
        RECT  65.7 222.3 66.9 223.5 ;
        RECT  79.2 213.75 80.4 216.15 ;
        RECT  79.2 225.15 80.4 226.95 ;
        RECT  74.4 226.05 75.6 226.95 ;
        RECT  74.4 213.75 75.6 214.95 ;
        RECT  76.8 216.0 78.0 224.85 ;
        RECT  72.6 220.5 74.7 221.4 ;
        RECT  78.0 220.5 82.2 221.4 ;
        RECT  72.6 212.85 82.2 213.75 ;
        RECT  72.6 226.95 82.2 227.85 ;
        RECT  74.4 220.05 75.6 221.25 ;
        RECT  76.8 220.05 78.0 221.25 ;
        RECT  74.4 221.25 75.6 222.45 ;
        RECT  76.8 221.25 78.0 222.45 ;
        RECT  74.4 220.95 75.6 222.15 ;
        RECT  76.8 220.95 78.0 222.15 ;
        RECT  74.4 220.95 75.6 222.15 ;
        RECT  76.8 220.95 78.0 222.15 ;
        RECT  79.2 216.15 80.4 217.35 ;
        RECT  79.2 226.05 80.4 227.25 ;
        RECT  74.7 221.55 75.9 222.75 ;
        RECT  47.25 220.35 48.45 221.55 ;
        RECT  49.2 218.25 50.4 219.45 ;
        RECT  60.6 218.25 61.8 219.45 ;
        RECT  57.6 238.65 58.8 241.05 ;
        RECT  57.6 227.85 58.8 229.65 ;
        RECT  52.8 227.85 54.0 228.75 ;
        RECT  52.8 239.85 54.0 241.05 ;
        RECT  55.2 229.95 56.4 238.8 ;
        RECT  51.0 233.4 53.1 234.3 ;
        RECT  56.4 233.4 60.6 234.3 ;
        RECT  51.0 241.05 60.6 241.95 ;
        RECT  51.0 226.95 60.6 227.85 ;
        RECT  52.8 228.75 54.0 229.95 ;
        RECT  55.2 228.75 56.4 229.95 ;
        RECT  52.8 229.95 54.0 231.15 ;
        RECT  55.2 229.95 56.4 231.15 ;
        RECT  52.8 238.65 54.0 239.85 ;
        RECT  55.2 238.65 56.4 239.85 ;
        RECT  52.8 238.65 54.0 239.85 ;
        RECT  55.2 238.65 56.4 239.85 ;
        RECT  57.6 238.65 58.8 239.85 ;
        RECT  57.6 228.75 58.8 229.95 ;
        RECT  53.1 233.25 54.3 234.45 ;
        RECT  69.6 238.65 70.5 241.5 ;
        RECT  69.6 227.4 70.5 229.8 ;
        RECT  62.55 238.65 63.45 241.5 ;
        RECT  67.35 238.65 68.25 241.5 ;
        RECT  62.55 227.4 63.45 230.25 ;
        RECT  67.8 235.5 68.7 236.4 ;
        RECT  64.8 235.5 65.7 236.4 ;
        RECT  67.8 229.05 68.7 235.95 ;
        RECT  65.25 235.5 68.25 236.4 ;
        RECT  64.8 235.95 65.7 238.65 ;
        RECT  60.6 235.5 62.7 236.4 ;
        RECT  68.25 233.4 72.6 234.3 ;
        RECT  60.6 232.8 65.7 233.7 ;
        RECT  60.6 241.05 72.6 241.95 ;
        RECT  60.6 226.95 72.6 227.85 ;
        RECT  62.4 229.05 63.6 230.25 ;
        RECT  64.8 229.05 66.0 230.25 ;
        RECT  62.4 230.25 63.6 231.45 ;
        RECT  64.8 230.25 66.0 231.45 ;
        RECT  64.8 229.05 66.0 230.25 ;
        RECT  67.2 229.05 68.4 230.25 ;
        RECT  64.8 230.25 66.0 231.45 ;
        RECT  67.2 230.25 68.4 231.45 ;
        RECT  62.4 238.65 63.6 239.85 ;
        RECT  64.8 238.65 66.0 239.85 ;
        RECT  62.4 238.65 63.6 239.85 ;
        RECT  64.8 238.65 66.0 239.85 ;
        RECT  64.8 238.65 66.0 239.85 ;
        RECT  67.2 238.65 68.4 239.85 ;
        RECT  64.8 238.65 66.0 239.85 ;
        RECT  67.2 238.65 68.4 239.85 ;
        RECT  69.6 238.65 70.8 239.85 ;
        RECT  69.6 229.05 70.8 230.25 ;
        RECT  62.7 235.2 63.9 236.4 ;
        RECT  65.7 232.5 66.9 233.7 ;
        RECT  79.2 238.65 80.4 241.05 ;
        RECT  79.2 227.85 80.4 229.65 ;
        RECT  74.4 227.85 75.6 228.75 ;
        RECT  74.4 239.85 75.6 241.05 ;
        RECT  76.8 229.95 78.0 238.8 ;
        RECT  72.6 233.4 74.7 234.3 ;
        RECT  78.0 233.4 82.2 234.3 ;
        RECT  72.6 241.05 82.2 241.95 ;
        RECT  72.6 226.95 82.2 227.85 ;
        RECT  74.4 228.75 75.6 229.95 ;
        RECT  76.8 228.75 78.0 229.95 ;
        RECT  74.4 229.95 75.6 231.15 ;
        RECT  76.8 229.95 78.0 231.15 ;
        RECT  74.4 238.65 75.6 239.85 ;
        RECT  76.8 238.65 78.0 239.85 ;
        RECT  74.4 238.65 75.6 239.85 ;
        RECT  76.8 238.65 78.0 239.85 ;
        RECT  79.2 238.65 80.4 239.85 ;
        RECT  79.2 228.75 80.4 229.95 ;
        RECT  74.7 233.25 75.9 234.45 ;
        RECT  47.25 233.25 48.45 234.45 ;
        RECT  49.2 235.35 50.4 236.55 ;
        RECT  60.6 235.35 61.8 236.55 ;
        RECT  57.6 241.95 58.8 244.35 ;
        RECT  57.6 253.35 58.8 255.15 ;
        RECT  52.8 254.25 54.0 255.15 ;
        RECT  52.8 241.95 54.0 243.15 ;
        RECT  55.2 244.2 56.4 253.05 ;
        RECT  51.0 248.7 53.1 249.6 ;
        RECT  56.4 248.7 60.6 249.6 ;
        RECT  51.0 241.05 60.6 241.95 ;
        RECT  51.0 255.15 60.6 256.05 ;
        RECT  52.8 248.25 54.0 249.45 ;
        RECT  55.2 248.25 56.4 249.45 ;
        RECT  52.8 249.45 54.0 250.65 ;
        RECT  55.2 249.45 56.4 250.65 ;
        RECT  52.8 249.15 54.0 250.35 ;
        RECT  55.2 249.15 56.4 250.35 ;
        RECT  52.8 249.15 54.0 250.35 ;
        RECT  55.2 249.15 56.4 250.35 ;
        RECT  57.6 244.35 58.8 245.55 ;
        RECT  57.6 254.25 58.8 255.45 ;
        RECT  53.1 249.75 54.3 250.95 ;
        RECT  69.6 241.5 70.5 244.35 ;
        RECT  69.6 253.2 70.5 255.6 ;
        RECT  62.55 241.5 63.45 244.35 ;
        RECT  67.35 241.5 68.25 244.35 ;
        RECT  62.55 252.75 63.45 255.6 ;
        RECT  67.8 246.6 68.7 247.5 ;
        RECT  64.8 246.6 65.7 247.5 ;
        RECT  67.8 247.05 68.7 253.95 ;
        RECT  65.25 246.6 68.25 247.5 ;
        RECT  64.8 244.35 65.7 247.05 ;
        RECT  60.6 246.6 62.7 247.5 ;
        RECT  68.25 248.7 72.6 249.6 ;
        RECT  60.6 249.3 65.7 250.2 ;
        RECT  60.6 241.05 72.6 241.95 ;
        RECT  60.6 255.15 72.6 256.05 ;
        RECT  62.4 246.75 63.6 247.95 ;
        RECT  64.8 246.75 66.0 247.95 ;
        RECT  62.4 247.95 63.6 249.15 ;
        RECT  64.8 247.95 66.0 249.15 ;
        RECT  64.8 246.75 66.0 247.95 ;
        RECT  67.2 246.75 68.4 247.95 ;
        RECT  64.8 247.95 66.0 249.15 ;
        RECT  67.2 247.95 68.4 249.15 ;
        RECT  62.4 249.15 63.6 250.35 ;
        RECT  64.8 249.15 66.0 250.35 ;
        RECT  62.4 249.15 63.6 250.35 ;
        RECT  64.8 249.15 66.0 250.35 ;
        RECT  64.8 249.15 66.0 250.35 ;
        RECT  67.2 249.15 68.4 250.35 ;
        RECT  64.8 249.15 66.0 250.35 ;
        RECT  67.2 249.15 68.4 250.35 ;
        RECT  69.6 244.35 70.8 245.55 ;
        RECT  69.6 253.95 70.8 255.15 ;
        RECT  62.7 247.8 63.9 249.0 ;
        RECT  65.7 250.5 66.9 251.7 ;
        RECT  79.2 241.95 80.4 244.35 ;
        RECT  79.2 253.35 80.4 255.15 ;
        RECT  74.4 254.25 75.6 255.15 ;
        RECT  74.4 241.95 75.6 243.15 ;
        RECT  76.8 244.2 78.0 253.05 ;
        RECT  72.6 248.7 74.7 249.6 ;
        RECT  78.0 248.7 82.2 249.6 ;
        RECT  72.6 241.05 82.2 241.95 ;
        RECT  72.6 255.15 82.2 256.05 ;
        RECT  74.4 248.25 75.6 249.45 ;
        RECT  76.8 248.25 78.0 249.45 ;
        RECT  74.4 249.45 75.6 250.65 ;
        RECT  76.8 249.45 78.0 250.65 ;
        RECT  74.4 249.15 75.6 250.35 ;
        RECT  76.8 249.15 78.0 250.35 ;
        RECT  74.4 249.15 75.6 250.35 ;
        RECT  76.8 249.15 78.0 250.35 ;
        RECT  79.2 244.35 80.4 245.55 ;
        RECT  79.2 254.25 80.4 255.45 ;
        RECT  74.7 249.75 75.9 250.95 ;
        RECT  47.25 248.55 48.45 249.75 ;
        RECT  49.2 246.45 50.4 247.65 ;
        RECT  60.6 246.45 61.8 247.65 ;
        RECT  57.6 266.85 58.8 269.25 ;
        RECT  57.6 256.05 58.8 257.85 ;
        RECT  52.8 256.05 54.0 256.95 ;
        RECT  52.8 268.05 54.0 269.25 ;
        RECT  55.2 258.15 56.4 267.0 ;
        RECT  51.0 261.6 53.1 262.5 ;
        RECT  56.4 261.6 60.6 262.5 ;
        RECT  51.0 269.25 60.6 270.15 ;
        RECT  51.0 255.15 60.6 256.05 ;
        RECT  52.8 256.95 54.0 258.15 ;
        RECT  55.2 256.95 56.4 258.15 ;
        RECT  52.8 258.15 54.0 259.35 ;
        RECT  55.2 258.15 56.4 259.35 ;
        RECT  52.8 266.85 54.0 268.05 ;
        RECT  55.2 266.85 56.4 268.05 ;
        RECT  52.8 266.85 54.0 268.05 ;
        RECT  55.2 266.85 56.4 268.05 ;
        RECT  57.6 266.85 58.8 268.05 ;
        RECT  57.6 256.95 58.8 258.15 ;
        RECT  53.1 261.45 54.3 262.65 ;
        RECT  69.6 266.85 70.5 269.7 ;
        RECT  69.6 255.6 70.5 258.0 ;
        RECT  62.55 266.85 63.45 269.7 ;
        RECT  67.35 266.85 68.25 269.7 ;
        RECT  62.55 255.6 63.45 258.45 ;
        RECT  67.8 263.7 68.7 264.6 ;
        RECT  64.8 263.7 65.7 264.6 ;
        RECT  67.8 257.25 68.7 264.15 ;
        RECT  65.25 263.7 68.25 264.6 ;
        RECT  64.8 264.15 65.7 266.85 ;
        RECT  60.6 263.7 62.7 264.6 ;
        RECT  68.25 261.6 72.6 262.5 ;
        RECT  60.6 261.0 65.7 261.9 ;
        RECT  60.6 269.25 72.6 270.15 ;
        RECT  60.6 255.15 72.6 256.05 ;
        RECT  62.4 257.25 63.6 258.45 ;
        RECT  64.8 257.25 66.0 258.45 ;
        RECT  62.4 258.45 63.6 259.65 ;
        RECT  64.8 258.45 66.0 259.65 ;
        RECT  64.8 257.25 66.0 258.45 ;
        RECT  67.2 257.25 68.4 258.45 ;
        RECT  64.8 258.45 66.0 259.65 ;
        RECT  67.2 258.45 68.4 259.65 ;
        RECT  62.4 266.85 63.6 268.05 ;
        RECT  64.8 266.85 66.0 268.05 ;
        RECT  62.4 266.85 63.6 268.05 ;
        RECT  64.8 266.85 66.0 268.05 ;
        RECT  64.8 266.85 66.0 268.05 ;
        RECT  67.2 266.85 68.4 268.05 ;
        RECT  64.8 266.85 66.0 268.05 ;
        RECT  67.2 266.85 68.4 268.05 ;
        RECT  69.6 266.85 70.8 268.05 ;
        RECT  69.6 257.25 70.8 258.45 ;
        RECT  62.7 263.4 63.9 264.6 ;
        RECT  65.7 260.7 66.9 261.9 ;
        RECT  79.2 266.85 80.4 269.25 ;
        RECT  79.2 256.05 80.4 257.85 ;
        RECT  74.4 256.05 75.6 256.95 ;
        RECT  74.4 268.05 75.6 269.25 ;
        RECT  76.8 258.15 78.0 267.0 ;
        RECT  72.6 261.6 74.7 262.5 ;
        RECT  78.0 261.6 82.2 262.5 ;
        RECT  72.6 269.25 82.2 270.15 ;
        RECT  72.6 255.15 82.2 256.05 ;
        RECT  74.4 256.95 75.6 258.15 ;
        RECT  76.8 256.95 78.0 258.15 ;
        RECT  74.4 258.15 75.6 259.35 ;
        RECT  76.8 258.15 78.0 259.35 ;
        RECT  74.4 266.85 75.6 268.05 ;
        RECT  76.8 266.85 78.0 268.05 ;
        RECT  74.4 266.85 75.6 268.05 ;
        RECT  76.8 266.85 78.0 268.05 ;
        RECT  79.2 266.85 80.4 268.05 ;
        RECT  79.2 256.95 80.4 258.15 ;
        RECT  74.7 261.45 75.9 262.65 ;
        RECT  47.25 261.45 48.45 262.65 ;
        RECT  49.2 263.55 50.4 264.75 ;
        RECT  60.6 263.55 61.8 264.75 ;
        RECT  57.6 270.15 58.8 272.55 ;
        RECT  57.6 281.55 58.8 283.35 ;
        RECT  52.8 282.45 54.0 283.35 ;
        RECT  52.8 270.15 54.0 271.35 ;
        RECT  55.2 272.4 56.4 281.25 ;
        RECT  51.0 276.9 53.1 277.8 ;
        RECT  56.4 276.9 60.6 277.8 ;
        RECT  51.0 269.25 60.6 270.15 ;
        RECT  51.0 283.35 60.6 284.25 ;
        RECT  52.8 276.45 54.0 277.65 ;
        RECT  55.2 276.45 56.4 277.65 ;
        RECT  52.8 277.65 54.0 278.85 ;
        RECT  55.2 277.65 56.4 278.85 ;
        RECT  52.8 277.35 54.0 278.55 ;
        RECT  55.2 277.35 56.4 278.55 ;
        RECT  52.8 277.35 54.0 278.55 ;
        RECT  55.2 277.35 56.4 278.55 ;
        RECT  57.6 272.55 58.8 273.75 ;
        RECT  57.6 282.45 58.8 283.65 ;
        RECT  53.1 277.95 54.3 279.15 ;
        RECT  69.6 269.7 70.5 272.55 ;
        RECT  69.6 281.4 70.5 283.8 ;
        RECT  62.55 269.7 63.45 272.55 ;
        RECT  67.35 269.7 68.25 272.55 ;
        RECT  62.55 280.95 63.45 283.8 ;
        RECT  67.8 274.8 68.7 275.7 ;
        RECT  64.8 274.8 65.7 275.7 ;
        RECT  67.8 275.25 68.7 282.15 ;
        RECT  65.25 274.8 68.25 275.7 ;
        RECT  64.8 272.55 65.7 275.25 ;
        RECT  60.6 274.8 62.7 275.7 ;
        RECT  68.25 276.9 72.6 277.8 ;
        RECT  60.6 277.5 65.7 278.4 ;
        RECT  60.6 269.25 72.6 270.15 ;
        RECT  60.6 283.35 72.6 284.25 ;
        RECT  62.4 274.95 63.6 276.15 ;
        RECT  64.8 274.95 66.0 276.15 ;
        RECT  62.4 276.15 63.6 277.35 ;
        RECT  64.8 276.15 66.0 277.35 ;
        RECT  64.8 274.95 66.0 276.15 ;
        RECT  67.2 274.95 68.4 276.15 ;
        RECT  64.8 276.15 66.0 277.35 ;
        RECT  67.2 276.15 68.4 277.35 ;
        RECT  62.4 277.35 63.6 278.55 ;
        RECT  64.8 277.35 66.0 278.55 ;
        RECT  62.4 277.35 63.6 278.55 ;
        RECT  64.8 277.35 66.0 278.55 ;
        RECT  64.8 277.35 66.0 278.55 ;
        RECT  67.2 277.35 68.4 278.55 ;
        RECT  64.8 277.35 66.0 278.55 ;
        RECT  67.2 277.35 68.4 278.55 ;
        RECT  69.6 272.55 70.8 273.75 ;
        RECT  69.6 282.15 70.8 283.35 ;
        RECT  62.7 276.0 63.9 277.2 ;
        RECT  65.7 278.7 66.9 279.9 ;
        RECT  79.2 270.15 80.4 272.55 ;
        RECT  79.2 281.55 80.4 283.35 ;
        RECT  74.4 282.45 75.6 283.35 ;
        RECT  74.4 270.15 75.6 271.35 ;
        RECT  76.8 272.4 78.0 281.25 ;
        RECT  72.6 276.9 74.7 277.8 ;
        RECT  78.0 276.9 82.2 277.8 ;
        RECT  72.6 269.25 82.2 270.15 ;
        RECT  72.6 283.35 82.2 284.25 ;
        RECT  74.4 276.45 75.6 277.65 ;
        RECT  76.8 276.45 78.0 277.65 ;
        RECT  74.4 277.65 75.6 278.85 ;
        RECT  76.8 277.65 78.0 278.85 ;
        RECT  74.4 277.35 75.6 278.55 ;
        RECT  76.8 277.35 78.0 278.55 ;
        RECT  74.4 277.35 75.6 278.55 ;
        RECT  76.8 277.35 78.0 278.55 ;
        RECT  79.2 272.55 80.4 273.75 ;
        RECT  79.2 282.45 80.4 283.65 ;
        RECT  74.7 277.95 75.9 279.15 ;
        RECT  47.25 276.75 48.45 277.95 ;
        RECT  49.2 274.65 50.4 275.85 ;
        RECT  60.6 274.65 61.8 275.85 ;
        RECT  57.6 295.05 58.8 297.45 ;
        RECT  57.6 284.25 58.8 286.05 ;
        RECT  52.8 284.25 54.0 285.15 ;
        RECT  52.8 296.25 54.0 297.45 ;
        RECT  55.2 286.35 56.4 295.2 ;
        RECT  51.0 289.8 53.1 290.7 ;
        RECT  56.4 289.8 60.6 290.7 ;
        RECT  51.0 297.45 60.6 298.35 ;
        RECT  51.0 283.35 60.6 284.25 ;
        RECT  52.8 285.15 54.0 286.35 ;
        RECT  55.2 285.15 56.4 286.35 ;
        RECT  52.8 286.35 54.0 287.55 ;
        RECT  55.2 286.35 56.4 287.55 ;
        RECT  52.8 295.05 54.0 296.25 ;
        RECT  55.2 295.05 56.4 296.25 ;
        RECT  52.8 295.05 54.0 296.25 ;
        RECT  55.2 295.05 56.4 296.25 ;
        RECT  57.6 295.05 58.8 296.25 ;
        RECT  57.6 285.15 58.8 286.35 ;
        RECT  53.1 289.65 54.3 290.85 ;
        RECT  69.6 295.05 70.5 297.9 ;
        RECT  69.6 283.8 70.5 286.2 ;
        RECT  62.55 295.05 63.45 297.9 ;
        RECT  67.35 295.05 68.25 297.9 ;
        RECT  62.55 283.8 63.45 286.65 ;
        RECT  67.8 291.9 68.7 292.8 ;
        RECT  64.8 291.9 65.7 292.8 ;
        RECT  67.8 285.45 68.7 292.35 ;
        RECT  65.25 291.9 68.25 292.8 ;
        RECT  64.8 292.35 65.7 295.05 ;
        RECT  60.6 291.9 62.7 292.8 ;
        RECT  68.25 289.8 72.6 290.7 ;
        RECT  60.6 289.2 65.7 290.1 ;
        RECT  60.6 297.45 72.6 298.35 ;
        RECT  60.6 283.35 72.6 284.25 ;
        RECT  62.4 285.45 63.6 286.65 ;
        RECT  64.8 285.45 66.0 286.65 ;
        RECT  62.4 286.65 63.6 287.85 ;
        RECT  64.8 286.65 66.0 287.85 ;
        RECT  64.8 285.45 66.0 286.65 ;
        RECT  67.2 285.45 68.4 286.65 ;
        RECT  64.8 286.65 66.0 287.85 ;
        RECT  67.2 286.65 68.4 287.85 ;
        RECT  62.4 295.05 63.6 296.25 ;
        RECT  64.8 295.05 66.0 296.25 ;
        RECT  62.4 295.05 63.6 296.25 ;
        RECT  64.8 295.05 66.0 296.25 ;
        RECT  64.8 295.05 66.0 296.25 ;
        RECT  67.2 295.05 68.4 296.25 ;
        RECT  64.8 295.05 66.0 296.25 ;
        RECT  67.2 295.05 68.4 296.25 ;
        RECT  69.6 295.05 70.8 296.25 ;
        RECT  69.6 285.45 70.8 286.65 ;
        RECT  62.7 291.6 63.9 292.8 ;
        RECT  65.7 288.9 66.9 290.1 ;
        RECT  79.2 295.05 80.4 297.45 ;
        RECT  79.2 284.25 80.4 286.05 ;
        RECT  74.4 284.25 75.6 285.15 ;
        RECT  74.4 296.25 75.6 297.45 ;
        RECT  76.8 286.35 78.0 295.2 ;
        RECT  72.6 289.8 74.7 290.7 ;
        RECT  78.0 289.8 82.2 290.7 ;
        RECT  72.6 297.45 82.2 298.35 ;
        RECT  72.6 283.35 82.2 284.25 ;
        RECT  74.4 285.15 75.6 286.35 ;
        RECT  76.8 285.15 78.0 286.35 ;
        RECT  74.4 286.35 75.6 287.55 ;
        RECT  76.8 286.35 78.0 287.55 ;
        RECT  74.4 295.05 75.6 296.25 ;
        RECT  76.8 295.05 78.0 296.25 ;
        RECT  74.4 295.05 75.6 296.25 ;
        RECT  76.8 295.05 78.0 296.25 ;
        RECT  79.2 295.05 80.4 296.25 ;
        RECT  79.2 285.15 80.4 286.35 ;
        RECT  74.7 289.65 75.9 290.85 ;
        RECT  47.25 289.65 48.45 290.85 ;
        RECT  49.2 291.75 50.4 292.95 ;
        RECT  60.6 291.75 61.8 292.95 ;
        RECT  57.6 298.35 58.8 300.75 ;
        RECT  57.6 309.75 58.8 311.55 ;
        RECT  52.8 310.65 54.0 311.55 ;
        RECT  52.8 298.35 54.0 299.55 ;
        RECT  55.2 300.6 56.4 309.45 ;
        RECT  51.0 305.1 53.1 306.0 ;
        RECT  56.4 305.1 60.6 306.0 ;
        RECT  51.0 297.45 60.6 298.35 ;
        RECT  51.0 311.55 60.6 312.45 ;
        RECT  52.8 304.65 54.0 305.85 ;
        RECT  55.2 304.65 56.4 305.85 ;
        RECT  52.8 305.85 54.0 307.05 ;
        RECT  55.2 305.85 56.4 307.05 ;
        RECT  52.8 305.55 54.0 306.75 ;
        RECT  55.2 305.55 56.4 306.75 ;
        RECT  52.8 305.55 54.0 306.75 ;
        RECT  55.2 305.55 56.4 306.75 ;
        RECT  57.6 300.75 58.8 301.95 ;
        RECT  57.6 310.65 58.8 311.85 ;
        RECT  53.1 306.15 54.3 307.35 ;
        RECT  69.6 297.9 70.5 300.75 ;
        RECT  69.6 309.6 70.5 312.0 ;
        RECT  62.55 297.9 63.45 300.75 ;
        RECT  67.35 297.9 68.25 300.75 ;
        RECT  62.55 309.15 63.45 312.0 ;
        RECT  67.8 303.0 68.7 303.9 ;
        RECT  64.8 303.0 65.7 303.9 ;
        RECT  67.8 303.45 68.7 310.35 ;
        RECT  65.25 303.0 68.25 303.9 ;
        RECT  64.8 300.75 65.7 303.45 ;
        RECT  60.6 303.0 62.7 303.9 ;
        RECT  68.25 305.1 72.6 306.0 ;
        RECT  60.6 305.7 65.7 306.6 ;
        RECT  60.6 297.45 72.6 298.35 ;
        RECT  60.6 311.55 72.6 312.45 ;
        RECT  62.4 303.15 63.6 304.35 ;
        RECT  64.8 303.15 66.0 304.35 ;
        RECT  62.4 304.35 63.6 305.55 ;
        RECT  64.8 304.35 66.0 305.55 ;
        RECT  64.8 303.15 66.0 304.35 ;
        RECT  67.2 303.15 68.4 304.35 ;
        RECT  64.8 304.35 66.0 305.55 ;
        RECT  67.2 304.35 68.4 305.55 ;
        RECT  62.4 305.55 63.6 306.75 ;
        RECT  64.8 305.55 66.0 306.75 ;
        RECT  62.4 305.55 63.6 306.75 ;
        RECT  64.8 305.55 66.0 306.75 ;
        RECT  64.8 305.55 66.0 306.75 ;
        RECT  67.2 305.55 68.4 306.75 ;
        RECT  64.8 305.55 66.0 306.75 ;
        RECT  67.2 305.55 68.4 306.75 ;
        RECT  69.6 300.75 70.8 301.95 ;
        RECT  69.6 310.35 70.8 311.55 ;
        RECT  62.7 304.2 63.9 305.4 ;
        RECT  65.7 306.9 66.9 308.1 ;
        RECT  79.2 298.35 80.4 300.75 ;
        RECT  79.2 309.75 80.4 311.55 ;
        RECT  74.4 310.65 75.6 311.55 ;
        RECT  74.4 298.35 75.6 299.55 ;
        RECT  76.8 300.6 78.0 309.45 ;
        RECT  72.6 305.1 74.7 306.0 ;
        RECT  78.0 305.1 82.2 306.0 ;
        RECT  72.6 297.45 82.2 298.35 ;
        RECT  72.6 311.55 82.2 312.45 ;
        RECT  74.4 304.65 75.6 305.85 ;
        RECT  76.8 304.65 78.0 305.85 ;
        RECT  74.4 305.85 75.6 307.05 ;
        RECT  76.8 305.85 78.0 307.05 ;
        RECT  74.4 305.55 75.6 306.75 ;
        RECT  76.8 305.55 78.0 306.75 ;
        RECT  74.4 305.55 75.6 306.75 ;
        RECT  76.8 305.55 78.0 306.75 ;
        RECT  79.2 300.75 80.4 301.95 ;
        RECT  79.2 310.65 80.4 311.85 ;
        RECT  74.7 306.15 75.9 307.35 ;
        RECT  47.25 304.95 48.45 306.15 ;
        RECT  49.2 302.85 50.4 304.05 ;
        RECT  60.6 302.85 61.8 304.05 ;
        RECT  57.6 323.25 58.8 325.65 ;
        RECT  57.6 312.45 58.8 314.25 ;
        RECT  52.8 312.45 54.0 313.35 ;
        RECT  52.8 324.45 54.0 325.65 ;
        RECT  55.2 314.55 56.4 323.4 ;
        RECT  51.0 318.0 53.1 318.9 ;
        RECT  56.4 318.0 60.6 318.9 ;
        RECT  51.0 325.65 60.6 326.55 ;
        RECT  51.0 311.55 60.6 312.45 ;
        RECT  52.8 313.35 54.0 314.55 ;
        RECT  55.2 313.35 56.4 314.55 ;
        RECT  52.8 314.55 54.0 315.75 ;
        RECT  55.2 314.55 56.4 315.75 ;
        RECT  52.8 323.25 54.0 324.45 ;
        RECT  55.2 323.25 56.4 324.45 ;
        RECT  52.8 323.25 54.0 324.45 ;
        RECT  55.2 323.25 56.4 324.45 ;
        RECT  57.6 323.25 58.8 324.45 ;
        RECT  57.6 313.35 58.8 314.55 ;
        RECT  53.1 317.85 54.3 319.05 ;
        RECT  69.6 323.25 70.5 326.1 ;
        RECT  69.6 312.0 70.5 314.4 ;
        RECT  62.55 323.25 63.45 326.1 ;
        RECT  67.35 323.25 68.25 326.1 ;
        RECT  62.55 312.0 63.45 314.85 ;
        RECT  67.8 320.1 68.7 321.0 ;
        RECT  64.8 320.1 65.7 321.0 ;
        RECT  67.8 313.65 68.7 320.55 ;
        RECT  65.25 320.1 68.25 321.0 ;
        RECT  64.8 320.55 65.7 323.25 ;
        RECT  60.6 320.1 62.7 321.0 ;
        RECT  68.25 318.0 72.6 318.9 ;
        RECT  60.6 317.4 65.7 318.3 ;
        RECT  60.6 325.65 72.6 326.55 ;
        RECT  60.6 311.55 72.6 312.45 ;
        RECT  62.4 313.65 63.6 314.85 ;
        RECT  64.8 313.65 66.0 314.85 ;
        RECT  62.4 314.85 63.6 316.05 ;
        RECT  64.8 314.85 66.0 316.05 ;
        RECT  64.8 313.65 66.0 314.85 ;
        RECT  67.2 313.65 68.4 314.85 ;
        RECT  64.8 314.85 66.0 316.05 ;
        RECT  67.2 314.85 68.4 316.05 ;
        RECT  62.4 323.25 63.6 324.45 ;
        RECT  64.8 323.25 66.0 324.45 ;
        RECT  62.4 323.25 63.6 324.45 ;
        RECT  64.8 323.25 66.0 324.45 ;
        RECT  64.8 323.25 66.0 324.45 ;
        RECT  67.2 323.25 68.4 324.45 ;
        RECT  64.8 323.25 66.0 324.45 ;
        RECT  67.2 323.25 68.4 324.45 ;
        RECT  69.6 323.25 70.8 324.45 ;
        RECT  69.6 313.65 70.8 314.85 ;
        RECT  62.7 319.8 63.9 321.0 ;
        RECT  65.7 317.1 66.9 318.3 ;
        RECT  79.2 323.25 80.4 325.65 ;
        RECT  79.2 312.45 80.4 314.25 ;
        RECT  74.4 312.45 75.6 313.35 ;
        RECT  74.4 324.45 75.6 325.65 ;
        RECT  76.8 314.55 78.0 323.4 ;
        RECT  72.6 318.0 74.7 318.9 ;
        RECT  78.0 318.0 82.2 318.9 ;
        RECT  72.6 325.65 82.2 326.55 ;
        RECT  72.6 311.55 82.2 312.45 ;
        RECT  74.4 313.35 75.6 314.55 ;
        RECT  76.8 313.35 78.0 314.55 ;
        RECT  74.4 314.55 75.6 315.75 ;
        RECT  76.8 314.55 78.0 315.75 ;
        RECT  74.4 323.25 75.6 324.45 ;
        RECT  76.8 323.25 78.0 324.45 ;
        RECT  74.4 323.25 75.6 324.45 ;
        RECT  76.8 323.25 78.0 324.45 ;
        RECT  79.2 323.25 80.4 324.45 ;
        RECT  79.2 313.35 80.4 314.55 ;
        RECT  74.7 317.85 75.9 319.05 ;
        RECT  47.25 317.85 48.45 319.05 ;
        RECT  49.2 319.95 50.4 321.15 ;
        RECT  60.6 319.95 61.8 321.15 ;
        RECT  57.6 326.55 58.8 328.95 ;
        RECT  57.6 337.95 58.8 339.75 ;
        RECT  52.8 338.85 54.0 339.75 ;
        RECT  52.8 326.55 54.0 327.75 ;
        RECT  55.2 328.8 56.4 337.65 ;
        RECT  51.0 333.3 53.1 334.2 ;
        RECT  56.4 333.3 60.6 334.2 ;
        RECT  51.0 325.65 60.6 326.55 ;
        RECT  51.0 339.75 60.6 340.65 ;
        RECT  52.8 332.85 54.0 334.05 ;
        RECT  55.2 332.85 56.4 334.05 ;
        RECT  52.8 334.05 54.0 335.25 ;
        RECT  55.2 334.05 56.4 335.25 ;
        RECT  52.8 333.75 54.0 334.95 ;
        RECT  55.2 333.75 56.4 334.95 ;
        RECT  52.8 333.75 54.0 334.95 ;
        RECT  55.2 333.75 56.4 334.95 ;
        RECT  57.6 328.95 58.8 330.15 ;
        RECT  57.6 338.85 58.8 340.05 ;
        RECT  53.1 334.35 54.3 335.55 ;
        RECT  69.6 326.1 70.5 328.95 ;
        RECT  69.6 337.8 70.5 340.2 ;
        RECT  62.55 326.1 63.45 328.95 ;
        RECT  67.35 326.1 68.25 328.95 ;
        RECT  62.55 337.35 63.45 340.2 ;
        RECT  67.8 331.2 68.7 332.1 ;
        RECT  64.8 331.2 65.7 332.1 ;
        RECT  67.8 331.65 68.7 338.55 ;
        RECT  65.25 331.2 68.25 332.1 ;
        RECT  64.8 328.95 65.7 331.65 ;
        RECT  60.6 331.2 62.7 332.1 ;
        RECT  68.25 333.3 72.6 334.2 ;
        RECT  60.6 333.9 65.7 334.8 ;
        RECT  60.6 325.65 72.6 326.55 ;
        RECT  60.6 339.75 72.6 340.65 ;
        RECT  62.4 331.35 63.6 332.55 ;
        RECT  64.8 331.35 66.0 332.55 ;
        RECT  62.4 332.55 63.6 333.75 ;
        RECT  64.8 332.55 66.0 333.75 ;
        RECT  64.8 331.35 66.0 332.55 ;
        RECT  67.2 331.35 68.4 332.55 ;
        RECT  64.8 332.55 66.0 333.75 ;
        RECT  67.2 332.55 68.4 333.75 ;
        RECT  62.4 333.75 63.6 334.95 ;
        RECT  64.8 333.75 66.0 334.95 ;
        RECT  62.4 333.75 63.6 334.95 ;
        RECT  64.8 333.75 66.0 334.95 ;
        RECT  64.8 333.75 66.0 334.95 ;
        RECT  67.2 333.75 68.4 334.95 ;
        RECT  64.8 333.75 66.0 334.95 ;
        RECT  67.2 333.75 68.4 334.95 ;
        RECT  69.6 328.95 70.8 330.15 ;
        RECT  69.6 338.55 70.8 339.75 ;
        RECT  62.7 332.4 63.9 333.6 ;
        RECT  65.7 335.1 66.9 336.3 ;
        RECT  79.2 326.55 80.4 328.95 ;
        RECT  79.2 337.95 80.4 339.75 ;
        RECT  74.4 338.85 75.6 339.75 ;
        RECT  74.4 326.55 75.6 327.75 ;
        RECT  76.8 328.8 78.0 337.65 ;
        RECT  72.6 333.3 74.7 334.2 ;
        RECT  78.0 333.3 82.2 334.2 ;
        RECT  72.6 325.65 82.2 326.55 ;
        RECT  72.6 339.75 82.2 340.65 ;
        RECT  74.4 332.85 75.6 334.05 ;
        RECT  76.8 332.85 78.0 334.05 ;
        RECT  74.4 334.05 75.6 335.25 ;
        RECT  76.8 334.05 78.0 335.25 ;
        RECT  74.4 333.75 75.6 334.95 ;
        RECT  76.8 333.75 78.0 334.95 ;
        RECT  74.4 333.75 75.6 334.95 ;
        RECT  76.8 333.75 78.0 334.95 ;
        RECT  79.2 328.95 80.4 330.15 ;
        RECT  79.2 338.85 80.4 340.05 ;
        RECT  74.7 334.35 75.9 335.55 ;
        RECT  47.25 333.15 48.45 334.35 ;
        RECT  49.2 331.05 50.4 332.25 ;
        RECT  60.6 331.05 61.8 332.25 ;
        RECT  57.6 351.45 58.8 353.85 ;
        RECT  57.6 340.65 58.8 342.45 ;
        RECT  52.8 340.65 54.0 341.55 ;
        RECT  52.8 352.65 54.0 353.85 ;
        RECT  55.2 342.75 56.4 351.6 ;
        RECT  51.0 346.2 53.1 347.1 ;
        RECT  56.4 346.2 60.6 347.1 ;
        RECT  51.0 353.85 60.6 354.75 ;
        RECT  51.0 339.75 60.6 340.65 ;
        RECT  52.8 341.55 54.0 342.75 ;
        RECT  55.2 341.55 56.4 342.75 ;
        RECT  52.8 342.75 54.0 343.95 ;
        RECT  55.2 342.75 56.4 343.95 ;
        RECT  52.8 351.45 54.0 352.65 ;
        RECT  55.2 351.45 56.4 352.65 ;
        RECT  52.8 351.45 54.0 352.65 ;
        RECT  55.2 351.45 56.4 352.65 ;
        RECT  57.6 351.45 58.8 352.65 ;
        RECT  57.6 341.55 58.8 342.75 ;
        RECT  53.1 346.05 54.3 347.25 ;
        RECT  69.6 351.45 70.5 354.3 ;
        RECT  69.6 340.2 70.5 342.6 ;
        RECT  62.55 351.45 63.45 354.3 ;
        RECT  67.35 351.45 68.25 354.3 ;
        RECT  62.55 340.2 63.45 343.05 ;
        RECT  67.8 348.3 68.7 349.2 ;
        RECT  64.8 348.3 65.7 349.2 ;
        RECT  67.8 341.85 68.7 348.75 ;
        RECT  65.25 348.3 68.25 349.2 ;
        RECT  64.8 348.75 65.7 351.45 ;
        RECT  60.6 348.3 62.7 349.2 ;
        RECT  68.25 346.2 72.6 347.1 ;
        RECT  60.6 345.6 65.7 346.5 ;
        RECT  60.6 353.85 72.6 354.75 ;
        RECT  60.6 339.75 72.6 340.65 ;
        RECT  62.4 341.85 63.6 343.05 ;
        RECT  64.8 341.85 66.0 343.05 ;
        RECT  62.4 343.05 63.6 344.25 ;
        RECT  64.8 343.05 66.0 344.25 ;
        RECT  64.8 341.85 66.0 343.05 ;
        RECT  67.2 341.85 68.4 343.05 ;
        RECT  64.8 343.05 66.0 344.25 ;
        RECT  67.2 343.05 68.4 344.25 ;
        RECT  62.4 351.45 63.6 352.65 ;
        RECT  64.8 351.45 66.0 352.65 ;
        RECT  62.4 351.45 63.6 352.65 ;
        RECT  64.8 351.45 66.0 352.65 ;
        RECT  64.8 351.45 66.0 352.65 ;
        RECT  67.2 351.45 68.4 352.65 ;
        RECT  64.8 351.45 66.0 352.65 ;
        RECT  67.2 351.45 68.4 352.65 ;
        RECT  69.6 351.45 70.8 352.65 ;
        RECT  69.6 341.85 70.8 343.05 ;
        RECT  62.7 348.0 63.9 349.2 ;
        RECT  65.7 345.3 66.9 346.5 ;
        RECT  79.2 351.45 80.4 353.85 ;
        RECT  79.2 340.65 80.4 342.45 ;
        RECT  74.4 340.65 75.6 341.55 ;
        RECT  74.4 352.65 75.6 353.85 ;
        RECT  76.8 342.75 78.0 351.6 ;
        RECT  72.6 346.2 74.7 347.1 ;
        RECT  78.0 346.2 82.2 347.1 ;
        RECT  72.6 353.85 82.2 354.75 ;
        RECT  72.6 339.75 82.2 340.65 ;
        RECT  74.4 341.55 75.6 342.75 ;
        RECT  76.8 341.55 78.0 342.75 ;
        RECT  74.4 342.75 75.6 343.95 ;
        RECT  76.8 342.75 78.0 343.95 ;
        RECT  74.4 351.45 75.6 352.65 ;
        RECT  76.8 351.45 78.0 352.65 ;
        RECT  74.4 351.45 75.6 352.65 ;
        RECT  76.8 351.45 78.0 352.65 ;
        RECT  79.2 351.45 80.4 352.65 ;
        RECT  79.2 341.55 80.4 342.75 ;
        RECT  74.7 346.05 75.9 347.25 ;
        RECT  47.25 346.05 48.45 347.25 ;
        RECT  49.2 348.15 50.4 349.35 ;
        RECT  60.6 348.15 61.8 349.35 ;
        RECT  57.6 354.75 58.8 357.15 ;
        RECT  57.6 366.15 58.8 367.95 ;
        RECT  52.8 367.05 54.0 367.95 ;
        RECT  52.8 354.75 54.0 355.95 ;
        RECT  55.2 357.0 56.4 365.85 ;
        RECT  51.0 361.5 53.1 362.4 ;
        RECT  56.4 361.5 60.6 362.4 ;
        RECT  51.0 353.85 60.6 354.75 ;
        RECT  51.0 367.95 60.6 368.85 ;
        RECT  52.8 361.05 54.0 362.25 ;
        RECT  55.2 361.05 56.4 362.25 ;
        RECT  52.8 362.25 54.0 363.45 ;
        RECT  55.2 362.25 56.4 363.45 ;
        RECT  52.8 361.95 54.0 363.15 ;
        RECT  55.2 361.95 56.4 363.15 ;
        RECT  52.8 361.95 54.0 363.15 ;
        RECT  55.2 361.95 56.4 363.15 ;
        RECT  57.6 357.15 58.8 358.35 ;
        RECT  57.6 367.05 58.8 368.25 ;
        RECT  53.1 362.55 54.3 363.75 ;
        RECT  69.6 354.3 70.5 357.15 ;
        RECT  69.6 366.0 70.5 368.4 ;
        RECT  62.55 354.3 63.45 357.15 ;
        RECT  67.35 354.3 68.25 357.15 ;
        RECT  62.55 365.55 63.45 368.4 ;
        RECT  67.8 359.4 68.7 360.3 ;
        RECT  64.8 359.4 65.7 360.3 ;
        RECT  67.8 359.85 68.7 366.75 ;
        RECT  65.25 359.4 68.25 360.3 ;
        RECT  64.8 357.15 65.7 359.85 ;
        RECT  60.6 359.4 62.7 360.3 ;
        RECT  68.25 361.5 72.6 362.4 ;
        RECT  60.6 362.1 65.7 363.0 ;
        RECT  60.6 353.85 72.6 354.75 ;
        RECT  60.6 367.95 72.6 368.85 ;
        RECT  62.4 359.55 63.6 360.75 ;
        RECT  64.8 359.55 66.0 360.75 ;
        RECT  62.4 360.75 63.6 361.95 ;
        RECT  64.8 360.75 66.0 361.95 ;
        RECT  64.8 359.55 66.0 360.75 ;
        RECT  67.2 359.55 68.4 360.75 ;
        RECT  64.8 360.75 66.0 361.95 ;
        RECT  67.2 360.75 68.4 361.95 ;
        RECT  62.4 361.95 63.6 363.15 ;
        RECT  64.8 361.95 66.0 363.15 ;
        RECT  62.4 361.95 63.6 363.15 ;
        RECT  64.8 361.95 66.0 363.15 ;
        RECT  64.8 361.95 66.0 363.15 ;
        RECT  67.2 361.95 68.4 363.15 ;
        RECT  64.8 361.95 66.0 363.15 ;
        RECT  67.2 361.95 68.4 363.15 ;
        RECT  69.6 357.15 70.8 358.35 ;
        RECT  69.6 366.75 70.8 367.95 ;
        RECT  62.7 360.6 63.9 361.8 ;
        RECT  65.7 363.3 66.9 364.5 ;
        RECT  79.2 354.75 80.4 357.15 ;
        RECT  79.2 366.15 80.4 367.95 ;
        RECT  74.4 367.05 75.6 367.95 ;
        RECT  74.4 354.75 75.6 355.95 ;
        RECT  76.8 357.0 78.0 365.85 ;
        RECT  72.6 361.5 74.7 362.4 ;
        RECT  78.0 361.5 82.2 362.4 ;
        RECT  72.6 353.85 82.2 354.75 ;
        RECT  72.6 367.95 82.2 368.85 ;
        RECT  74.4 361.05 75.6 362.25 ;
        RECT  76.8 361.05 78.0 362.25 ;
        RECT  74.4 362.25 75.6 363.45 ;
        RECT  76.8 362.25 78.0 363.45 ;
        RECT  74.4 361.95 75.6 363.15 ;
        RECT  76.8 361.95 78.0 363.15 ;
        RECT  74.4 361.95 75.6 363.15 ;
        RECT  76.8 361.95 78.0 363.15 ;
        RECT  79.2 357.15 80.4 358.35 ;
        RECT  79.2 367.05 80.4 368.25 ;
        RECT  74.7 362.55 75.9 363.75 ;
        RECT  47.25 361.35 48.45 362.55 ;
        RECT  49.2 359.25 50.4 360.45 ;
        RECT  60.6 359.25 61.8 360.45 ;
        RECT  57.6 379.65 58.8 382.05 ;
        RECT  57.6 368.85 58.8 370.65 ;
        RECT  52.8 368.85 54.0 369.75 ;
        RECT  52.8 380.85 54.0 382.05 ;
        RECT  55.2 370.95 56.4 379.8 ;
        RECT  51.0 374.4 53.1 375.3 ;
        RECT  56.4 374.4 60.6 375.3 ;
        RECT  51.0 382.05 60.6 382.95 ;
        RECT  51.0 367.95 60.6 368.85 ;
        RECT  52.8 369.75 54.0 370.95 ;
        RECT  55.2 369.75 56.4 370.95 ;
        RECT  52.8 370.95 54.0 372.15 ;
        RECT  55.2 370.95 56.4 372.15 ;
        RECT  52.8 379.65 54.0 380.85 ;
        RECT  55.2 379.65 56.4 380.85 ;
        RECT  52.8 379.65 54.0 380.85 ;
        RECT  55.2 379.65 56.4 380.85 ;
        RECT  57.6 379.65 58.8 380.85 ;
        RECT  57.6 369.75 58.8 370.95 ;
        RECT  53.1 374.25 54.3 375.45 ;
        RECT  69.6 379.65 70.5 382.5 ;
        RECT  69.6 368.4 70.5 370.8 ;
        RECT  62.55 379.65 63.45 382.5 ;
        RECT  67.35 379.65 68.25 382.5 ;
        RECT  62.55 368.4 63.45 371.25 ;
        RECT  67.8 376.5 68.7 377.4 ;
        RECT  64.8 376.5 65.7 377.4 ;
        RECT  67.8 370.05 68.7 376.95 ;
        RECT  65.25 376.5 68.25 377.4 ;
        RECT  64.8 376.95 65.7 379.65 ;
        RECT  60.6 376.5 62.7 377.4 ;
        RECT  68.25 374.4 72.6 375.3 ;
        RECT  60.6 373.8 65.7 374.7 ;
        RECT  60.6 382.05 72.6 382.95 ;
        RECT  60.6 367.95 72.6 368.85 ;
        RECT  62.4 370.05 63.6 371.25 ;
        RECT  64.8 370.05 66.0 371.25 ;
        RECT  62.4 371.25 63.6 372.45 ;
        RECT  64.8 371.25 66.0 372.45 ;
        RECT  64.8 370.05 66.0 371.25 ;
        RECT  67.2 370.05 68.4 371.25 ;
        RECT  64.8 371.25 66.0 372.45 ;
        RECT  67.2 371.25 68.4 372.45 ;
        RECT  62.4 379.65 63.6 380.85 ;
        RECT  64.8 379.65 66.0 380.85 ;
        RECT  62.4 379.65 63.6 380.85 ;
        RECT  64.8 379.65 66.0 380.85 ;
        RECT  64.8 379.65 66.0 380.85 ;
        RECT  67.2 379.65 68.4 380.85 ;
        RECT  64.8 379.65 66.0 380.85 ;
        RECT  67.2 379.65 68.4 380.85 ;
        RECT  69.6 379.65 70.8 380.85 ;
        RECT  69.6 370.05 70.8 371.25 ;
        RECT  62.7 376.2 63.9 377.4 ;
        RECT  65.7 373.5 66.9 374.7 ;
        RECT  79.2 379.65 80.4 382.05 ;
        RECT  79.2 368.85 80.4 370.65 ;
        RECT  74.4 368.85 75.6 369.75 ;
        RECT  74.4 380.85 75.6 382.05 ;
        RECT  76.8 370.95 78.0 379.8 ;
        RECT  72.6 374.4 74.7 375.3 ;
        RECT  78.0 374.4 82.2 375.3 ;
        RECT  72.6 382.05 82.2 382.95 ;
        RECT  72.6 367.95 82.2 368.85 ;
        RECT  74.4 369.75 75.6 370.95 ;
        RECT  76.8 369.75 78.0 370.95 ;
        RECT  74.4 370.95 75.6 372.15 ;
        RECT  76.8 370.95 78.0 372.15 ;
        RECT  74.4 379.65 75.6 380.85 ;
        RECT  76.8 379.65 78.0 380.85 ;
        RECT  74.4 379.65 75.6 380.85 ;
        RECT  76.8 379.65 78.0 380.85 ;
        RECT  79.2 379.65 80.4 380.85 ;
        RECT  79.2 369.75 80.4 370.95 ;
        RECT  74.7 374.25 75.9 375.45 ;
        RECT  47.25 374.25 48.45 375.45 ;
        RECT  49.2 376.35 50.4 377.55 ;
        RECT  60.6 376.35 61.8 377.55 ;
        RECT  57.6 382.95 58.8 385.35 ;
        RECT  57.6 394.35 58.8 396.15 ;
        RECT  52.8 395.25 54.0 396.15 ;
        RECT  52.8 382.95 54.0 384.15 ;
        RECT  55.2 385.2 56.4 394.05 ;
        RECT  51.0 389.7 53.1 390.6 ;
        RECT  56.4 389.7 60.6 390.6 ;
        RECT  51.0 382.05 60.6 382.95 ;
        RECT  51.0 396.15 60.6 397.05 ;
        RECT  52.8 389.25 54.0 390.45 ;
        RECT  55.2 389.25 56.4 390.45 ;
        RECT  52.8 390.45 54.0 391.65 ;
        RECT  55.2 390.45 56.4 391.65 ;
        RECT  52.8 390.15 54.0 391.35 ;
        RECT  55.2 390.15 56.4 391.35 ;
        RECT  52.8 390.15 54.0 391.35 ;
        RECT  55.2 390.15 56.4 391.35 ;
        RECT  57.6 385.35 58.8 386.55 ;
        RECT  57.6 395.25 58.8 396.45 ;
        RECT  53.1 390.75 54.3 391.95 ;
        RECT  69.6 382.5 70.5 385.35 ;
        RECT  69.6 394.2 70.5 396.6 ;
        RECT  62.55 382.5 63.45 385.35 ;
        RECT  67.35 382.5 68.25 385.35 ;
        RECT  62.55 393.75 63.45 396.6 ;
        RECT  67.8 387.6 68.7 388.5 ;
        RECT  64.8 387.6 65.7 388.5 ;
        RECT  67.8 388.05 68.7 394.95 ;
        RECT  65.25 387.6 68.25 388.5 ;
        RECT  64.8 385.35 65.7 388.05 ;
        RECT  60.6 387.6 62.7 388.5 ;
        RECT  68.25 389.7 72.6 390.6 ;
        RECT  60.6 390.3 65.7 391.2 ;
        RECT  60.6 382.05 72.6 382.95 ;
        RECT  60.6 396.15 72.6 397.05 ;
        RECT  62.4 387.75 63.6 388.95 ;
        RECT  64.8 387.75 66.0 388.95 ;
        RECT  62.4 388.95 63.6 390.15 ;
        RECT  64.8 388.95 66.0 390.15 ;
        RECT  64.8 387.75 66.0 388.95 ;
        RECT  67.2 387.75 68.4 388.95 ;
        RECT  64.8 388.95 66.0 390.15 ;
        RECT  67.2 388.95 68.4 390.15 ;
        RECT  62.4 390.15 63.6 391.35 ;
        RECT  64.8 390.15 66.0 391.35 ;
        RECT  62.4 390.15 63.6 391.35 ;
        RECT  64.8 390.15 66.0 391.35 ;
        RECT  64.8 390.15 66.0 391.35 ;
        RECT  67.2 390.15 68.4 391.35 ;
        RECT  64.8 390.15 66.0 391.35 ;
        RECT  67.2 390.15 68.4 391.35 ;
        RECT  69.6 385.35 70.8 386.55 ;
        RECT  69.6 394.95 70.8 396.15 ;
        RECT  62.7 388.8 63.9 390.0 ;
        RECT  65.7 391.5 66.9 392.7 ;
        RECT  79.2 382.95 80.4 385.35 ;
        RECT  79.2 394.35 80.4 396.15 ;
        RECT  74.4 395.25 75.6 396.15 ;
        RECT  74.4 382.95 75.6 384.15 ;
        RECT  76.8 385.2 78.0 394.05 ;
        RECT  72.6 389.7 74.7 390.6 ;
        RECT  78.0 389.7 82.2 390.6 ;
        RECT  72.6 382.05 82.2 382.95 ;
        RECT  72.6 396.15 82.2 397.05 ;
        RECT  74.4 389.25 75.6 390.45 ;
        RECT  76.8 389.25 78.0 390.45 ;
        RECT  74.4 390.45 75.6 391.65 ;
        RECT  76.8 390.45 78.0 391.65 ;
        RECT  74.4 390.15 75.6 391.35 ;
        RECT  76.8 390.15 78.0 391.35 ;
        RECT  74.4 390.15 75.6 391.35 ;
        RECT  76.8 390.15 78.0 391.35 ;
        RECT  79.2 385.35 80.4 386.55 ;
        RECT  79.2 395.25 80.4 396.45 ;
        RECT  74.7 390.75 75.9 391.95 ;
        RECT  47.25 389.55 48.45 390.75 ;
        RECT  49.2 387.45 50.4 388.65 ;
        RECT  60.6 387.45 61.8 388.65 ;
        RECT  57.6 407.85 58.8 410.25 ;
        RECT  57.6 397.05 58.8 398.85 ;
        RECT  52.8 397.05 54.0 397.95 ;
        RECT  52.8 409.05 54.0 410.25 ;
        RECT  55.2 399.15 56.4 408.0 ;
        RECT  51.0 402.6 53.1 403.5 ;
        RECT  56.4 402.6 60.6 403.5 ;
        RECT  51.0 410.25 60.6 411.15 ;
        RECT  51.0 396.15 60.6 397.05 ;
        RECT  52.8 397.95 54.0 399.15 ;
        RECT  55.2 397.95 56.4 399.15 ;
        RECT  52.8 399.15 54.0 400.35 ;
        RECT  55.2 399.15 56.4 400.35 ;
        RECT  52.8 407.85 54.0 409.05 ;
        RECT  55.2 407.85 56.4 409.05 ;
        RECT  52.8 407.85 54.0 409.05 ;
        RECT  55.2 407.85 56.4 409.05 ;
        RECT  57.6 407.85 58.8 409.05 ;
        RECT  57.6 397.95 58.8 399.15 ;
        RECT  53.1 402.45 54.3 403.65 ;
        RECT  69.6 407.85 70.5 410.7 ;
        RECT  69.6 396.6 70.5 399.0 ;
        RECT  62.55 407.85 63.45 410.7 ;
        RECT  67.35 407.85 68.25 410.7 ;
        RECT  62.55 396.6 63.45 399.45 ;
        RECT  67.8 404.7 68.7 405.6 ;
        RECT  64.8 404.7 65.7 405.6 ;
        RECT  67.8 398.25 68.7 405.15 ;
        RECT  65.25 404.7 68.25 405.6 ;
        RECT  64.8 405.15 65.7 407.85 ;
        RECT  60.6 404.7 62.7 405.6 ;
        RECT  68.25 402.6 72.6 403.5 ;
        RECT  60.6 402.0 65.7 402.9 ;
        RECT  60.6 410.25 72.6 411.15 ;
        RECT  60.6 396.15 72.6 397.05 ;
        RECT  62.4 398.25 63.6 399.45 ;
        RECT  64.8 398.25 66.0 399.45 ;
        RECT  62.4 399.45 63.6 400.65 ;
        RECT  64.8 399.45 66.0 400.65 ;
        RECT  64.8 398.25 66.0 399.45 ;
        RECT  67.2 398.25 68.4 399.45 ;
        RECT  64.8 399.45 66.0 400.65 ;
        RECT  67.2 399.45 68.4 400.65 ;
        RECT  62.4 407.85 63.6 409.05 ;
        RECT  64.8 407.85 66.0 409.05 ;
        RECT  62.4 407.85 63.6 409.05 ;
        RECT  64.8 407.85 66.0 409.05 ;
        RECT  64.8 407.85 66.0 409.05 ;
        RECT  67.2 407.85 68.4 409.05 ;
        RECT  64.8 407.85 66.0 409.05 ;
        RECT  67.2 407.85 68.4 409.05 ;
        RECT  69.6 407.85 70.8 409.05 ;
        RECT  69.6 398.25 70.8 399.45 ;
        RECT  62.7 404.4 63.9 405.6 ;
        RECT  65.7 401.7 66.9 402.9 ;
        RECT  79.2 407.85 80.4 410.25 ;
        RECT  79.2 397.05 80.4 398.85 ;
        RECT  74.4 397.05 75.6 397.95 ;
        RECT  74.4 409.05 75.6 410.25 ;
        RECT  76.8 399.15 78.0 408.0 ;
        RECT  72.6 402.6 74.7 403.5 ;
        RECT  78.0 402.6 82.2 403.5 ;
        RECT  72.6 410.25 82.2 411.15 ;
        RECT  72.6 396.15 82.2 397.05 ;
        RECT  74.4 397.95 75.6 399.15 ;
        RECT  76.8 397.95 78.0 399.15 ;
        RECT  74.4 399.15 75.6 400.35 ;
        RECT  76.8 399.15 78.0 400.35 ;
        RECT  74.4 407.85 75.6 409.05 ;
        RECT  76.8 407.85 78.0 409.05 ;
        RECT  74.4 407.85 75.6 409.05 ;
        RECT  76.8 407.85 78.0 409.05 ;
        RECT  79.2 407.85 80.4 409.05 ;
        RECT  79.2 397.95 80.4 399.15 ;
        RECT  74.7 402.45 75.9 403.65 ;
        RECT  47.25 402.45 48.45 403.65 ;
        RECT  49.2 404.55 50.4 405.75 ;
        RECT  60.6 404.55 61.8 405.75 ;
        RECT  57.6 411.15 58.8 413.55 ;
        RECT  57.6 422.55 58.8 424.35 ;
        RECT  52.8 423.45 54.0 424.35 ;
        RECT  52.8 411.15 54.0 412.35 ;
        RECT  55.2 413.4 56.4 422.25 ;
        RECT  51.0 417.9 53.1 418.8 ;
        RECT  56.4 417.9 60.6 418.8 ;
        RECT  51.0 410.25 60.6 411.15 ;
        RECT  51.0 424.35 60.6 425.25 ;
        RECT  52.8 417.45 54.0 418.65 ;
        RECT  55.2 417.45 56.4 418.65 ;
        RECT  52.8 418.65 54.0 419.85 ;
        RECT  55.2 418.65 56.4 419.85 ;
        RECT  52.8 418.35 54.0 419.55 ;
        RECT  55.2 418.35 56.4 419.55 ;
        RECT  52.8 418.35 54.0 419.55 ;
        RECT  55.2 418.35 56.4 419.55 ;
        RECT  57.6 413.55 58.8 414.75 ;
        RECT  57.6 423.45 58.8 424.65 ;
        RECT  53.1 418.95 54.3 420.15 ;
        RECT  69.6 410.7 70.5 413.55 ;
        RECT  69.6 422.4 70.5 424.8 ;
        RECT  62.55 410.7 63.45 413.55 ;
        RECT  67.35 410.7 68.25 413.55 ;
        RECT  62.55 421.95 63.45 424.8 ;
        RECT  67.8 415.8 68.7 416.7 ;
        RECT  64.8 415.8 65.7 416.7 ;
        RECT  67.8 416.25 68.7 423.15 ;
        RECT  65.25 415.8 68.25 416.7 ;
        RECT  64.8 413.55 65.7 416.25 ;
        RECT  60.6 415.8 62.7 416.7 ;
        RECT  68.25 417.9 72.6 418.8 ;
        RECT  60.6 418.5 65.7 419.4 ;
        RECT  60.6 410.25 72.6 411.15 ;
        RECT  60.6 424.35 72.6 425.25 ;
        RECT  62.4 415.95 63.6 417.15 ;
        RECT  64.8 415.95 66.0 417.15 ;
        RECT  62.4 417.15 63.6 418.35 ;
        RECT  64.8 417.15 66.0 418.35 ;
        RECT  64.8 415.95 66.0 417.15 ;
        RECT  67.2 415.95 68.4 417.15 ;
        RECT  64.8 417.15 66.0 418.35 ;
        RECT  67.2 417.15 68.4 418.35 ;
        RECT  62.4 418.35 63.6 419.55 ;
        RECT  64.8 418.35 66.0 419.55 ;
        RECT  62.4 418.35 63.6 419.55 ;
        RECT  64.8 418.35 66.0 419.55 ;
        RECT  64.8 418.35 66.0 419.55 ;
        RECT  67.2 418.35 68.4 419.55 ;
        RECT  64.8 418.35 66.0 419.55 ;
        RECT  67.2 418.35 68.4 419.55 ;
        RECT  69.6 413.55 70.8 414.75 ;
        RECT  69.6 423.15 70.8 424.35 ;
        RECT  62.7 417.0 63.9 418.2 ;
        RECT  65.7 419.7 66.9 420.9 ;
        RECT  79.2 411.15 80.4 413.55 ;
        RECT  79.2 422.55 80.4 424.35 ;
        RECT  74.4 423.45 75.6 424.35 ;
        RECT  74.4 411.15 75.6 412.35 ;
        RECT  76.8 413.4 78.0 422.25 ;
        RECT  72.6 417.9 74.7 418.8 ;
        RECT  78.0 417.9 82.2 418.8 ;
        RECT  72.6 410.25 82.2 411.15 ;
        RECT  72.6 424.35 82.2 425.25 ;
        RECT  74.4 417.45 75.6 418.65 ;
        RECT  76.8 417.45 78.0 418.65 ;
        RECT  74.4 418.65 75.6 419.85 ;
        RECT  76.8 418.65 78.0 419.85 ;
        RECT  74.4 418.35 75.6 419.55 ;
        RECT  76.8 418.35 78.0 419.55 ;
        RECT  74.4 418.35 75.6 419.55 ;
        RECT  76.8 418.35 78.0 419.55 ;
        RECT  79.2 413.55 80.4 414.75 ;
        RECT  79.2 423.45 80.4 424.65 ;
        RECT  74.7 418.95 75.9 420.15 ;
        RECT  47.25 417.75 48.45 418.95 ;
        RECT  49.2 415.65 50.4 416.85 ;
        RECT  60.6 415.65 61.8 416.85 ;
        RECT  8.7 40.2 9.6 81.0 ;
        RECT  62.7 40.2 63.6 81.0 ;
        RECT  62.7 70.2 63.6 81.6 ;
        RECT  59.4 80.4 62.7 81.6 ;
        RECT  60.9 72.6 61.8 79.2 ;
        RECT  60.6 76.2 60.9 79.2 ;
        RECT  60.6 72.6 60.9 73.8 ;
        RECT  58.2 77.4 59.4 81.6 ;
        RECT  58.2 70.2 59.4 73.8 ;
        RECT  54.6 80.4 58.2 81.6 ;
        RECT  57.3 75.0 58.2 76.2 ;
        RECT  57.0 73.8 57.3 76.2 ;
        RECT  56.1 72.6 57.0 79.2 ;
        RECT  55.8 77.4 56.1 79.2 ;
        RECT  55.8 72.6 56.1 73.8 ;
        RECT  53.4 77.4 54.6 81.6 ;
        RECT  39.6 80.4 53.4 81.6 ;
        RECT  52.8 74.7 55.2 75.9 ;
        RECT  54.6 70.2 58.2 71.1 ;
        RECT  53.4 70.2 54.6 73.8 ;
        RECT  52.2 70.2 53.4 71.4 ;
        RECT  49.8 78.0 51.0 79.2 ;
        RECT  50.7 74.7 51.9 77.1 ;
        RECT  48.9 72.6 49.8 79.2 ;
        RECT  48.6 77.4 48.9 79.2 ;
        RECT  48.6 72.6 48.9 73.8 ;
        RECT  46.5 72.6 47.4 79.2 ;
        RECT  46.2 77.4 46.5 79.2 ;
        RECT  46.2 72.6 46.5 75.0 ;
        RECT  44.1 72.6 45.0 79.2 ;
        RECT  43.8 77.4 44.1 79.2 ;
        RECT  43.8 72.6 44.1 75.0 ;
        RECT  42.0 75.0 42.9 76.2 ;
        RECT  41.1 72.6 42.0 79.2 ;
        RECT  40.8 76.2 41.1 79.2 ;
        RECT  40.8 72.6 41.1 73.8 ;
        RECT  38.4 77.4 39.6 81.6 ;
        RECT  33.9 80.4 38.4 81.6 ;
        RECT  37.5 75.3 39.9 76.5 ;
        RECT  39.6 70.2 52.2 71.1 ;
        RECT  38.4 70.2 39.6 73.8 ;
        RECT  36.3 78.0 37.5 79.2 ;
        RECT  35.4 72.6 36.3 79.2 ;
        RECT  35.1 77.4 35.4 79.2 ;
        RECT  35.1 72.6 35.4 73.8 ;
        RECT  33.9 70.2 38.4 71.1 ;
        RECT  32.7 77.4 33.9 81.6 ;
        RECT  29.1 80.4 32.7 81.6 ;
        RECT  31.8 74.7 33.0 75.9 ;
        RECT  32.7 70.2 33.9 73.8 ;
        RECT  31.5 73.8 31.8 79.2 ;
        RECT  30.9 72.6 31.5 79.2 ;
        RECT  30.3 77.4 30.9 79.2 ;
        RECT  30.6 72.6 30.9 75.0 ;
        RECT  30.3 72.6 30.6 73.8 ;
        RECT  27.9 77.4 29.1 81.6 ;
        RECT  12.9 80.4 27.9 81.6 ;
        RECT  27.3 74.7 29.7 75.9 ;
        RECT  29.1 70.2 32.7 71.1 ;
        RECT  27.9 70.2 29.1 73.8 ;
        RECT  26.7 70.2 27.9 71.4 ;
        RECT  23.4 78.0 24.6 79.2 ;
        RECT  24.3 74.7 25.5 77.1 ;
        RECT  22.5 72.6 23.4 79.2 ;
        RECT  22.2 77.4 22.5 79.2 ;
        RECT  22.2 72.6 22.5 73.8 ;
        RECT  20.1 72.6 21.0 79.2 ;
        RECT  19.8 77.4 20.1 79.2 ;
        RECT  19.8 72.6 20.1 75.0 ;
        RECT  17.7 72.6 18.6 79.2 ;
        RECT  17.4 77.4 17.7 79.2 ;
        RECT  17.4 72.6 17.7 75.0 ;
        RECT  15.6 75.0 16.5 76.2 ;
        RECT  14.7 72.6 15.6 79.2 ;
        RECT  14.4 76.2 14.7 79.2 ;
        RECT  14.4 72.6 14.7 73.8 ;
        RECT  13.2 70.2 26.7 71.1 ;
        RECT  12.9 77.4 13.2 79.2 ;
        RECT  12.0 77.4 12.9 81.6 ;
        RECT  12.3 70.2 13.2 73.8 ;
        RECT  12.0 72.6 12.3 73.8 ;
        RECT  10.5 77.4 12.0 78.6 ;
        RECT  9.6 75.3 10.5 76.5 ;
        RECT  8.7 70.2 9.6 81.6 ;
        RECT  8.7 70.2 9.6 81.6 ;
        RECT  62.7 70.2 63.6 81.6 ;
        RECT  62.7 60.0 63.6 71.4 ;
        RECT  59.4 60.0 62.7 61.2 ;
        RECT  60.9 62.4 61.8 69.0 ;
        RECT  60.6 62.4 60.9 65.4 ;
        RECT  60.6 67.8 60.9 69.0 ;
        RECT  58.2 60.0 59.4 64.2 ;
        RECT  58.2 67.8 59.4 71.4 ;
        RECT  54.6 60.0 58.2 61.2 ;
        RECT  57.3 65.4 58.2 66.6 ;
        RECT  57.0 65.4 57.3 67.8 ;
        RECT  56.1 62.4 57.0 69.0 ;
        RECT  55.8 62.4 56.1 64.2 ;
        RECT  55.8 67.8 56.1 69.0 ;
        RECT  53.4 60.0 54.6 64.2 ;
        RECT  39.6 60.0 53.4 61.2 ;
        RECT  52.8 65.7 55.2 66.9 ;
        RECT  54.6 70.5 58.2 71.4 ;
        RECT  53.4 67.8 54.6 71.4 ;
        RECT  52.2 70.2 53.4 71.4 ;
        RECT  49.8 62.4 51.0 63.6 ;
        RECT  50.7 64.5 51.9 66.9 ;
        RECT  48.9 62.4 49.8 69.0 ;
        RECT  48.6 62.4 48.9 64.2 ;
        RECT  48.6 67.8 48.9 69.0 ;
        RECT  46.5 62.4 47.4 69.0 ;
        RECT  46.2 62.4 46.5 64.2 ;
        RECT  46.2 66.6 46.5 69.0 ;
        RECT  44.1 62.4 45.0 69.0 ;
        RECT  43.8 62.4 44.1 64.2 ;
        RECT  43.8 66.6 44.1 69.0 ;
        RECT  42.0 65.4 42.9 66.6 ;
        RECT  41.1 62.4 42.0 69.0 ;
        RECT  40.8 62.4 41.1 65.4 ;
        RECT  40.8 67.8 41.1 69.0 ;
        RECT  38.4 60.0 39.6 64.2 ;
        RECT  33.9 60.0 38.4 61.2 ;
        RECT  37.5 65.1 39.9 66.3 ;
        RECT  39.6 70.5 52.2 71.4 ;
        RECT  38.4 67.8 39.6 71.4 ;
        RECT  36.3 62.4 37.5 63.6 ;
        RECT  35.4 62.4 36.3 69.0 ;
        RECT  35.1 62.4 35.4 64.2 ;
        RECT  35.1 67.8 35.4 69.0 ;
        RECT  33.9 70.5 38.4 71.4 ;
        RECT  32.7 60.0 33.9 64.2 ;
        RECT  29.1 60.0 32.7 61.2 ;
        RECT  31.8 65.7 33.0 66.9 ;
        RECT  32.7 67.8 33.9 71.4 ;
        RECT  31.5 62.4 31.8 67.8 ;
        RECT  30.9 62.4 31.5 69.0 ;
        RECT  30.3 62.4 30.9 64.2 ;
        RECT  30.6 66.6 30.9 69.0 ;
        RECT  30.3 67.8 30.6 69.0 ;
        RECT  27.9 60.0 29.1 64.2 ;
        RECT  12.9 60.0 27.9 61.2 ;
        RECT  27.3 65.7 29.7 66.9 ;
        RECT  29.1 70.5 32.7 71.4 ;
        RECT  27.9 67.8 29.1 71.4 ;
        RECT  26.7 70.2 27.9 71.4 ;
        RECT  23.4 62.4 24.6 63.6 ;
        RECT  24.3 64.5 25.5 66.9 ;
        RECT  22.5 62.4 23.4 69.0 ;
        RECT  22.2 62.4 22.5 64.2 ;
        RECT  22.2 67.8 22.5 69.0 ;
        RECT  20.1 62.4 21.0 69.0 ;
        RECT  19.8 62.4 20.1 64.2 ;
        RECT  19.8 66.6 20.1 69.0 ;
        RECT  17.7 62.4 18.6 69.0 ;
        RECT  17.4 62.4 17.7 64.2 ;
        RECT  17.4 66.6 17.7 69.0 ;
        RECT  15.6 65.4 16.5 66.6 ;
        RECT  14.7 62.4 15.6 69.0 ;
        RECT  14.4 62.4 14.7 65.4 ;
        RECT  14.4 67.8 14.7 69.0 ;
        RECT  13.2 70.5 26.7 71.4 ;
        RECT  12.9 62.4 13.2 64.2 ;
        RECT  12.0 60.0 12.9 64.2 ;
        RECT  12.3 67.8 13.2 71.4 ;
        RECT  12.0 67.8 12.3 69.0 ;
        RECT  10.5 63.0 12.0 64.2 ;
        RECT  9.6 65.1 10.5 66.3 ;
        RECT  8.7 60.0 9.6 71.4 ;
        RECT  8.7 60.0 9.6 71.4 ;
        RECT  62.7 60.0 63.6 71.4 ;
        RECT  62.7 49.8 63.6 61.2 ;
        RECT  59.4 60.0 62.7 61.2 ;
        RECT  60.9 52.2 61.8 58.8 ;
        RECT  60.6 55.8 60.9 58.8 ;
        RECT  60.6 52.2 60.9 53.4 ;
        RECT  58.2 57.0 59.4 61.2 ;
        RECT  58.2 49.8 59.4 53.4 ;
        RECT  54.6 60.0 58.2 61.2 ;
        RECT  57.3 54.6 58.2 55.8 ;
        RECT  57.0 53.4 57.3 55.8 ;
        RECT  56.1 52.2 57.0 58.8 ;
        RECT  55.8 57.0 56.1 58.8 ;
        RECT  55.8 52.2 56.1 53.4 ;
        RECT  53.4 57.0 54.6 61.2 ;
        RECT  39.6 60.0 53.4 61.2 ;
        RECT  52.8 54.3 55.2 55.5 ;
        RECT  54.6 49.8 58.2 50.7 ;
        RECT  53.4 49.8 54.6 53.4 ;
        RECT  52.2 49.8 53.4 51.0 ;
        RECT  49.8 57.6 51.0 58.8 ;
        RECT  50.7 54.3 51.9 56.7 ;
        RECT  48.9 52.2 49.8 58.8 ;
        RECT  48.6 57.0 48.9 58.8 ;
        RECT  48.6 52.2 48.9 53.4 ;
        RECT  46.5 52.2 47.4 58.8 ;
        RECT  46.2 57.0 46.5 58.8 ;
        RECT  46.2 52.2 46.5 54.6 ;
        RECT  44.1 52.2 45.0 58.8 ;
        RECT  43.8 57.0 44.1 58.8 ;
        RECT  43.8 52.2 44.1 54.6 ;
        RECT  42.0 54.6 42.9 55.8 ;
        RECT  41.1 52.2 42.0 58.8 ;
        RECT  40.8 55.8 41.1 58.8 ;
        RECT  40.8 52.2 41.1 53.4 ;
        RECT  38.4 57.0 39.6 61.2 ;
        RECT  33.9 60.0 38.4 61.2 ;
        RECT  37.5 54.9 39.9 56.1 ;
        RECT  39.6 49.8 52.2 50.7 ;
        RECT  38.4 49.8 39.6 53.4 ;
        RECT  36.3 57.6 37.5 58.8 ;
        RECT  35.4 52.2 36.3 58.8 ;
        RECT  35.1 57.0 35.4 58.8 ;
        RECT  35.1 52.2 35.4 53.4 ;
        RECT  33.9 49.8 38.4 50.7 ;
        RECT  32.7 57.0 33.9 61.2 ;
        RECT  29.1 60.0 32.7 61.2 ;
        RECT  31.8 54.3 33.0 55.5 ;
        RECT  32.7 49.8 33.9 53.4 ;
        RECT  31.5 53.4 31.8 58.8 ;
        RECT  30.9 52.2 31.5 58.8 ;
        RECT  30.3 57.0 30.9 58.8 ;
        RECT  30.6 52.2 30.9 54.6 ;
        RECT  30.3 52.2 30.6 53.4 ;
        RECT  27.9 57.0 29.1 61.2 ;
        RECT  12.9 60.0 27.9 61.2 ;
        RECT  27.3 54.3 29.7 55.5 ;
        RECT  29.1 49.8 32.7 50.7 ;
        RECT  27.9 49.8 29.1 53.4 ;
        RECT  26.7 49.8 27.9 51.0 ;
        RECT  23.4 57.6 24.6 58.8 ;
        RECT  24.3 54.3 25.5 56.7 ;
        RECT  22.5 52.2 23.4 58.8 ;
        RECT  22.2 57.0 22.5 58.8 ;
        RECT  22.2 52.2 22.5 53.4 ;
        RECT  20.1 52.2 21.0 58.8 ;
        RECT  19.8 57.0 20.1 58.8 ;
        RECT  19.8 52.2 20.1 54.6 ;
        RECT  17.7 52.2 18.6 58.8 ;
        RECT  17.4 57.0 17.7 58.8 ;
        RECT  17.4 52.2 17.7 54.6 ;
        RECT  15.6 54.6 16.5 55.8 ;
        RECT  14.7 52.2 15.6 58.8 ;
        RECT  14.4 55.8 14.7 58.8 ;
        RECT  14.4 52.2 14.7 53.4 ;
        RECT  13.2 49.8 26.7 50.7 ;
        RECT  12.9 57.0 13.2 58.8 ;
        RECT  12.0 57.0 12.9 61.2 ;
        RECT  12.3 49.8 13.2 53.4 ;
        RECT  12.0 52.2 12.3 53.4 ;
        RECT  10.5 57.0 12.0 58.2 ;
        RECT  9.6 54.9 10.5 56.1 ;
        RECT  8.7 49.8 9.6 61.2 ;
        RECT  8.7 49.8 9.6 61.2 ;
        RECT  62.7 49.8 63.6 61.2 ;
        RECT  62.7 39.6 63.6 51.0 ;
        RECT  59.4 39.6 62.7 40.8 ;
        RECT  60.9 42.0 61.8 48.6 ;
        RECT  60.6 42.0 60.9 45.0 ;
        RECT  60.6 47.4 60.9 48.6 ;
        RECT  58.2 39.6 59.4 43.8 ;
        RECT  58.2 47.4 59.4 51.0 ;
        RECT  54.6 39.6 58.2 40.8 ;
        RECT  57.3 45.0 58.2 46.2 ;
        RECT  57.0 45.0 57.3 47.4 ;
        RECT  56.1 42.0 57.0 48.6 ;
        RECT  55.8 42.0 56.1 43.8 ;
        RECT  55.8 47.4 56.1 48.6 ;
        RECT  53.4 39.6 54.6 43.8 ;
        RECT  39.6 39.6 53.4 40.8 ;
        RECT  52.8 45.3 55.2 46.5 ;
        RECT  54.6 50.1 58.2 51.0 ;
        RECT  53.4 47.4 54.6 51.0 ;
        RECT  52.2 49.8 53.4 51.0 ;
        RECT  49.8 42.0 51.0 43.2 ;
        RECT  50.7 44.1 51.9 46.5 ;
        RECT  48.9 42.0 49.8 48.6 ;
        RECT  48.6 42.0 48.9 43.8 ;
        RECT  48.6 47.4 48.9 48.6 ;
        RECT  46.5 42.0 47.4 48.6 ;
        RECT  46.2 42.0 46.5 43.8 ;
        RECT  46.2 46.2 46.5 48.6 ;
        RECT  44.1 42.0 45.0 48.6 ;
        RECT  43.8 42.0 44.1 43.8 ;
        RECT  43.8 46.2 44.1 48.6 ;
        RECT  42.0 45.0 42.9 46.2 ;
        RECT  41.1 42.0 42.0 48.6 ;
        RECT  40.8 42.0 41.1 45.0 ;
        RECT  40.8 47.4 41.1 48.6 ;
        RECT  38.4 39.6 39.6 43.8 ;
        RECT  33.9 39.6 38.4 40.8 ;
        RECT  37.5 44.7 39.9 45.9 ;
        RECT  39.6 50.1 52.2 51.0 ;
        RECT  38.4 47.4 39.6 51.0 ;
        RECT  36.3 42.0 37.5 43.2 ;
        RECT  35.4 42.0 36.3 48.6 ;
        RECT  35.1 42.0 35.4 43.8 ;
        RECT  35.1 47.4 35.4 48.6 ;
        RECT  33.9 50.1 38.4 51.0 ;
        RECT  32.7 39.6 33.9 43.8 ;
        RECT  29.1 39.6 32.7 40.8 ;
        RECT  31.8 45.3 33.0 46.5 ;
        RECT  32.7 47.4 33.9 51.0 ;
        RECT  31.5 42.0 31.8 47.4 ;
        RECT  30.9 42.0 31.5 48.6 ;
        RECT  30.3 42.0 30.9 43.8 ;
        RECT  30.6 46.2 30.9 48.6 ;
        RECT  30.3 47.4 30.6 48.6 ;
        RECT  27.9 39.6 29.1 43.8 ;
        RECT  12.9 39.6 27.9 40.8 ;
        RECT  27.3 45.3 29.7 46.5 ;
        RECT  29.1 50.1 32.7 51.0 ;
        RECT  27.9 47.4 29.1 51.0 ;
        RECT  26.7 49.8 27.9 51.0 ;
        RECT  23.4 42.0 24.6 43.2 ;
        RECT  24.3 44.1 25.5 46.5 ;
        RECT  22.5 42.0 23.4 48.6 ;
        RECT  22.2 42.0 22.5 43.8 ;
        RECT  22.2 47.4 22.5 48.6 ;
        RECT  20.1 42.0 21.0 48.6 ;
        RECT  19.8 42.0 20.1 43.8 ;
        RECT  19.8 46.2 20.1 48.6 ;
        RECT  17.7 42.0 18.6 48.6 ;
        RECT  17.4 42.0 17.7 43.8 ;
        RECT  17.4 46.2 17.7 48.6 ;
        RECT  15.6 45.0 16.5 46.2 ;
        RECT  14.7 42.0 15.6 48.6 ;
        RECT  14.4 42.0 14.7 45.0 ;
        RECT  14.4 47.4 14.7 48.6 ;
        RECT  13.2 50.1 26.7 51.0 ;
        RECT  12.9 42.0 13.2 43.8 ;
        RECT  12.0 39.6 12.9 43.8 ;
        RECT  12.3 47.4 13.2 51.0 ;
        RECT  12.0 47.4 12.3 48.6 ;
        RECT  10.5 42.6 12.0 43.8 ;
        RECT  9.6 44.7 10.5 45.9 ;
        RECT  8.7 39.6 9.6 51.0 ;
        RECT  8.7 39.6 9.6 51.0 ;
        RECT  62.7 39.6 63.6 51.0 ;
        RECT  92.85 198.6 94.05 199.8 ;
        RECT  92.85 226.8 94.05 228.0 ;
        RECT  92.85 255.0 94.05 256.2 ;
        RECT  92.85 283.2 94.05 284.4 ;
        RECT  92.85 311.4 94.05 312.6 ;
        RECT  92.85 339.6 94.05 340.8 ;
        RECT  92.85 367.8 94.05 369.0 ;
        RECT  92.85 396.0 94.05 397.2 ;
        RECT  92.85 424.2 94.05 425.4 ;
        RECT  74.1 88.65 75.3 89.85 ;
        RECT  79.05 88.65 80.25 89.85 ;
        RECT  71.1 102.75 72.3 103.95 ;
        RECT  81.75 102.75 82.95 103.95 ;
        RECT  74.1 145.05 75.3 146.25 ;
        RECT  84.45 145.05 85.65 146.25 ;
        RECT  71.1 159.15 72.3 160.35 ;
        RECT  87.15 159.15 88.35 160.35 ;
        RECT  76.2 85.8 77.4 87.0 ;
        RECT  76.2 114.0 77.4 115.2 ;
        RECT  76.2 142.2 77.4 143.4 ;
        RECT  76.2 170.4 77.4 171.6 ;
        RECT  66.3 75.3 67.5 76.5 ;
        RECT  79.05 75.45 80.25 76.65 ;
        RECT  66.3 65.1 67.5 66.3 ;
        RECT  81.75 65.25 82.95 66.45 ;
        RECT  66.3 54.9 67.5 56.1 ;
        RECT  84.45 55.05 85.65 56.25 ;
        RECT  66.3 44.7 67.5 45.9 ;
        RECT  87.15 44.85 88.35 46.05 ;
        RECT  66.3 70.2 67.5 71.4 ;
        RECT  92.85 70.35 94.05 71.55 ;
        RECT  66.3 49.8 67.5 51.0 ;
        RECT  92.85 49.95 94.05 51.15 ;
        RECT  108.0 32.25 109.2 33.45 ;
        RECT  102.6 27.75 103.8 28.95 ;
        RECT  105.3 25.35 106.5 26.55 ;
        RECT  108.0 431.25 109.2 432.45 ;
        RECT  110.7 96.75 111.9 97.95 ;
        RECT  113.4 194.85 114.6 196.05 ;
        RECT  100.05 82.65 101.25 83.85 ;
        RECT  47.25 426.3 48.45 427.5 ;
        RECT  100.05 426.45 101.25 427.65 ;
        RECT  96.15 23.4 97.35 24.6 ;
        RECT  96.15 192.9 97.35 194.1 ;
        RECT  96.15 94.8 97.35 96.0 ;
        RECT  -22.5 258.6 -17.55 259.5 ;
        RECT  -9.9 207.6 -9.0 214.2 ;
        RECT  -9.9 224.4 -9.0 231.0 ;
        RECT  -9.9 303.0 -9.0 306.15 ;
        RECT  -22.5 204.6 -19.8 205.5 ;
        RECT  -27.3 306.15 -26.4 330.0 ;
        RECT  -25.2 311.55 -24.3 330.0 ;
        RECT  -12.75 325.05 -11.85 330.0 ;
        RECT  -10.65 322.35 -9.75 330.0 ;
        RECT  -8.55 314.25 -7.65 330.0 ;
        RECT  -10.65 345.15 -9.0 346.05 ;
        RECT  -9.9 355.2 -9.0 386.1 ;
        RECT  -40.95 325.05 -40.05 339.6 ;
        RECT  -38.85 316.95 -37.95 339.6 ;
        RECT  -36.75 314.25 -35.85 339.6 ;
        RECT  -38.85 354.75 -37.2 355.65 ;
        RECT  -25.2 385.65 -24.3 386.55 ;
        RECT  -25.2 385.65 -24.75 386.55 ;
        RECT  -25.2 383.4 -24.3 386.1 ;
        RECT  -3.45 202.2 -2.55 383.4 ;
        RECT  -3.45 308.85 -2.55 330.0 ;
        RECT  -17.55 202.2 -16.65 383.4 ;
        RECT  -17.55 319.65 -16.65 330.0 ;
        RECT  -31.65 330.0 -30.75 383.4 ;
        RECT  -31.65 308.85 -30.75 330.0 ;
        RECT  -45.75 330.0 -44.85 383.4 ;
        RECT  -45.75 319.65 -44.85 330.0 ;
        RECT  -3.45 383.4 -2.55 386.1 ;
        RECT  -17.55 383.4 -16.65 386.1 ;
        RECT  -31.65 383.4 -30.75 386.1 ;
        RECT  -45.75 382.95 -44.85 383.85 ;
        RECT  -49.8 382.95 -48.9 383.85 ;
        RECT  -45.75 381.3 -44.85 383.4 ;
        RECT  -49.35 382.95 -45.3 383.85 ;
        RECT  -49.8 383.4 -48.9 386.1 ;
        RECT  -9.9 202.2 -9.0 203.1 ;
        RECT  -17.55 202.2 -16.65 203.1 ;
        RECT  -3.45 202.2 -2.55 203.1 ;
        RECT  -53.1 204.6 -22.5 205.5 ;
        RECT  -53.1 258.6 -22.5 259.5 ;
        RECT  -53.7 258.6 -42.3 259.5 ;
        RECT  -53.7 255.3 -52.5 258.6 ;
        RECT  -51.3 256.8 -44.7 257.7 ;
        RECT  -51.3 256.5 -48.3 256.8 ;
        RECT  -45.9 256.5 -44.7 256.8 ;
        RECT  -53.7 254.1 -49.5 255.3 ;
        RECT  -45.9 254.1 -42.3 255.3 ;
        RECT  -53.7 250.5 -52.5 254.1 ;
        RECT  -48.3 253.2 -47.1 254.1 ;
        RECT  -48.3 252.9 -45.9 253.2 ;
        RECT  -51.3 252.0 -44.7 252.9 ;
        RECT  -51.3 251.7 -49.5 252.0 ;
        RECT  -45.9 251.7 -44.7 252.0 ;
        RECT  -53.7 249.3 -49.5 250.5 ;
        RECT  -53.7 235.5 -52.5 249.3 ;
        RECT  -48.0 248.7 -46.8 251.1 ;
        RECT  -43.2 250.5 -42.3 254.1 ;
        RECT  -45.9 249.3 -42.3 250.5 ;
        RECT  -43.5 248.1 -42.3 249.3 ;
        RECT  -51.3 245.7 -50.1 246.9 ;
        RECT  -49.2 246.6 -46.8 247.8 ;
        RECT  -51.3 244.8 -44.7 245.7 ;
        RECT  -51.3 244.5 -49.5 244.8 ;
        RECT  -45.9 244.5 -44.7 244.8 ;
        RECT  -51.3 242.4 -44.7 243.3 ;
        RECT  -51.3 242.1 -49.5 242.4 ;
        RECT  -47.1 242.1 -44.7 242.4 ;
        RECT  -51.3 240.0 -44.7 240.9 ;
        RECT  -51.3 239.7 -49.5 240.0 ;
        RECT  -47.1 239.7 -44.7 240.0 ;
        RECT  -48.3 237.9 -47.1 238.8 ;
        RECT  -51.3 237.0 -44.7 237.9 ;
        RECT  -51.3 236.7 -48.3 237.0 ;
        RECT  -45.9 236.7 -44.7 237.0 ;
        RECT  -53.7 234.3 -49.5 235.5 ;
        RECT  -53.7 229.8 -52.5 234.3 ;
        RECT  -48.6 233.4 -47.4 235.8 ;
        RECT  -43.2 235.5 -42.3 248.1 ;
        RECT  -45.9 234.3 -42.3 235.5 ;
        RECT  -51.3 232.2 -50.1 233.4 ;
        RECT  -51.3 231.3 -44.7 232.2 ;
        RECT  -51.3 231.0 -49.5 231.3 ;
        RECT  -45.9 231.0 -44.7 231.3 ;
        RECT  -43.2 229.8 -42.3 234.3 ;
        RECT  -53.7 228.6 -49.5 229.8 ;
        RECT  -53.7 225.0 -52.5 228.6 ;
        RECT  -48.0 227.7 -46.8 228.9 ;
        RECT  -45.9 228.6 -42.3 229.8 ;
        RECT  -51.3 227.4 -45.9 227.7 ;
        RECT  -51.3 226.8 -44.7 227.4 ;
        RECT  -51.3 226.2 -49.5 226.8 ;
        RECT  -47.1 226.5 -44.7 226.8 ;
        RECT  -45.9 226.2 -44.7 226.5 ;
        RECT  -53.7 223.8 -49.5 225.0 ;
        RECT  -53.7 208.8 -52.5 223.8 ;
        RECT  -48.0 223.2 -46.8 225.6 ;
        RECT  -43.2 225.0 -42.3 228.6 ;
        RECT  -45.9 223.8 -42.3 225.0 ;
        RECT  -43.5 222.6 -42.3 223.8 ;
        RECT  -51.3 219.3 -50.1 220.5 ;
        RECT  -49.2 220.2 -46.8 221.4 ;
        RECT  -51.3 218.4 -44.7 219.3 ;
        RECT  -51.3 218.1 -49.5 218.4 ;
        RECT  -45.9 218.1 -44.7 218.4 ;
        RECT  -51.3 216.0 -44.7 216.9 ;
        RECT  -51.3 215.7 -49.5 216.0 ;
        RECT  -47.1 215.7 -44.7 216.0 ;
        RECT  -51.3 213.6 -44.7 214.5 ;
        RECT  -51.3 213.3 -49.5 213.6 ;
        RECT  -47.1 213.3 -44.7 213.6 ;
        RECT  -48.3 211.5 -47.1 212.4 ;
        RECT  -51.3 210.6 -44.7 211.5 ;
        RECT  -51.3 210.3 -48.3 210.6 ;
        RECT  -45.9 210.3 -44.7 210.6 ;
        RECT  -43.2 209.1 -42.3 222.6 ;
        RECT  -51.3 208.8 -49.5 209.1 ;
        RECT  -53.7 207.9 -49.5 208.8 ;
        RECT  -45.9 208.2 -42.3 209.1 ;
        RECT  -45.9 207.9 -44.7 208.2 ;
        RECT  -50.7 206.4 -49.5 207.9 ;
        RECT  -48.6 205.5 -47.4 206.4 ;
        RECT  -53.7 204.6 -42.3 205.5 ;
        RECT  -53.7 204.6 -42.3 205.5 ;
        RECT  -53.7 258.6 -42.3 259.5 ;
        RECT  -43.5 258.6 -32.1 259.5 ;
        RECT  -33.3 255.3 -32.1 258.6 ;
        RECT  -41.1 256.8 -34.5 257.7 ;
        RECT  -37.5 256.5 -34.5 256.8 ;
        RECT  -41.1 256.5 -39.9 256.8 ;
        RECT  -36.3 254.1 -32.1 255.3 ;
        RECT  -43.5 254.1 -39.9 255.3 ;
        RECT  -33.3 250.5 -32.1 254.1 ;
        RECT  -38.7 253.2 -37.5 254.1 ;
        RECT  -39.9 252.9 -37.5 253.2 ;
        RECT  -41.1 252.0 -34.5 252.9 ;
        RECT  -36.3 251.7 -34.5 252.0 ;
        RECT  -41.1 251.7 -39.9 252.0 ;
        RECT  -36.3 249.3 -32.1 250.5 ;
        RECT  -33.3 235.5 -32.1 249.3 ;
        RECT  -39.0 248.7 -37.8 251.1 ;
        RECT  -43.5 250.5 -42.6 254.1 ;
        RECT  -43.5 249.3 -39.9 250.5 ;
        RECT  -43.5 248.1 -42.3 249.3 ;
        RECT  -35.7 245.7 -34.5 246.9 ;
        RECT  -39.0 246.6 -36.6 247.8 ;
        RECT  -41.1 244.8 -34.5 245.7 ;
        RECT  -36.3 244.5 -34.5 244.8 ;
        RECT  -41.1 244.5 -39.9 244.8 ;
        RECT  -41.1 242.4 -34.5 243.3 ;
        RECT  -36.3 242.1 -34.5 242.4 ;
        RECT  -41.1 242.1 -38.7 242.4 ;
        RECT  -41.1 240.0 -34.5 240.9 ;
        RECT  -36.3 239.7 -34.5 240.0 ;
        RECT  -41.1 239.7 -38.7 240.0 ;
        RECT  -38.7 237.9 -37.5 238.8 ;
        RECT  -41.1 237.0 -34.5 237.9 ;
        RECT  -37.5 236.7 -34.5 237.0 ;
        RECT  -41.1 236.7 -39.9 237.0 ;
        RECT  -36.3 234.3 -32.1 235.5 ;
        RECT  -33.3 229.8 -32.1 234.3 ;
        RECT  -38.4 233.4 -37.2 235.8 ;
        RECT  -43.5 235.5 -42.6 248.1 ;
        RECT  -43.5 234.3 -39.9 235.5 ;
        RECT  -35.7 232.2 -34.5 233.4 ;
        RECT  -41.1 231.3 -34.5 232.2 ;
        RECT  -36.3 231.0 -34.5 231.3 ;
        RECT  -41.1 231.0 -39.9 231.3 ;
        RECT  -43.5 229.8 -42.6 234.3 ;
        RECT  -36.3 228.6 -32.1 229.8 ;
        RECT  -33.3 225.0 -32.1 228.6 ;
        RECT  -39.0 227.7 -37.8 228.9 ;
        RECT  -43.5 228.6 -39.9 229.8 ;
        RECT  -39.9 227.4 -34.5 227.7 ;
        RECT  -41.1 226.8 -34.5 227.4 ;
        RECT  -36.3 226.2 -34.5 226.8 ;
        RECT  -41.1 226.5 -38.7 226.8 ;
        RECT  -41.1 226.2 -39.9 226.5 ;
        RECT  -36.3 223.8 -32.1 225.0 ;
        RECT  -33.3 208.8 -32.1 223.8 ;
        RECT  -39.0 223.2 -37.8 225.6 ;
        RECT  -43.5 225.0 -42.6 228.6 ;
        RECT  -43.5 223.8 -39.9 225.0 ;
        RECT  -43.5 222.6 -42.3 223.8 ;
        RECT  -35.7 219.3 -34.5 220.5 ;
        RECT  -39.0 220.2 -36.6 221.4 ;
        RECT  -41.1 218.4 -34.5 219.3 ;
        RECT  -36.3 218.1 -34.5 218.4 ;
        RECT  -41.1 218.1 -39.9 218.4 ;
        RECT  -41.1 216.0 -34.5 216.9 ;
        RECT  -36.3 215.7 -34.5 216.0 ;
        RECT  -41.1 215.7 -38.7 216.0 ;
        RECT  -41.1 213.6 -34.5 214.5 ;
        RECT  -36.3 213.3 -34.5 213.6 ;
        RECT  -41.1 213.3 -38.7 213.6 ;
        RECT  -38.7 211.5 -37.5 212.4 ;
        RECT  -41.1 210.6 -34.5 211.5 ;
        RECT  -37.5 210.3 -34.5 210.6 ;
        RECT  -41.1 210.3 -39.9 210.6 ;
        RECT  -43.5 209.1 -42.6 222.6 ;
        RECT  -36.3 208.8 -34.5 209.1 ;
        RECT  -36.3 207.9 -32.1 208.8 ;
        RECT  -43.5 208.2 -39.9 209.1 ;
        RECT  -41.1 207.9 -39.9 208.2 ;
        RECT  -36.3 206.4 -35.1 207.9 ;
        RECT  -38.4 205.5 -37.2 206.4 ;
        RECT  -43.5 204.6 -32.1 205.5 ;
        RECT  -43.5 204.6 -32.1 205.5 ;
        RECT  -43.5 258.6 -32.1 259.5 ;
        RECT  -33.3 258.6 -21.9 259.5 ;
        RECT  -33.3 255.3 -32.1 258.6 ;
        RECT  -30.9 256.8 -24.3 257.7 ;
        RECT  -30.9 256.5 -27.9 256.8 ;
        RECT  -25.5 256.5 -24.3 256.8 ;
        RECT  -33.3 254.1 -29.1 255.3 ;
        RECT  -25.5 254.1 -21.9 255.3 ;
        RECT  -33.3 250.5 -32.1 254.1 ;
        RECT  -27.9 253.2 -26.7 254.1 ;
        RECT  -27.9 252.9 -25.5 253.2 ;
        RECT  -30.9 252.0 -24.3 252.9 ;
        RECT  -30.9 251.7 -29.1 252.0 ;
        RECT  -25.5 251.7 -24.3 252.0 ;
        RECT  -33.3 249.3 -29.1 250.5 ;
        RECT  -33.3 235.5 -32.1 249.3 ;
        RECT  -27.6 248.7 -26.4 251.1 ;
        RECT  -22.8 250.5 -21.9 254.1 ;
        RECT  -25.5 249.3 -21.9 250.5 ;
        RECT  -23.1 248.1 -21.9 249.3 ;
        RECT  -30.9 245.7 -29.7 246.9 ;
        RECT  -28.8 246.6 -26.4 247.8 ;
        RECT  -30.9 244.8 -24.3 245.7 ;
        RECT  -30.9 244.5 -29.1 244.8 ;
        RECT  -25.5 244.5 -24.3 244.8 ;
        RECT  -30.9 242.4 -24.3 243.3 ;
        RECT  -30.9 242.1 -29.1 242.4 ;
        RECT  -26.7 242.1 -24.3 242.4 ;
        RECT  -30.9 240.0 -24.3 240.9 ;
        RECT  -30.9 239.7 -29.1 240.0 ;
        RECT  -26.7 239.7 -24.3 240.0 ;
        RECT  -27.9 237.9 -26.7 238.8 ;
        RECT  -30.9 237.0 -24.3 237.9 ;
        RECT  -30.9 236.7 -27.9 237.0 ;
        RECT  -25.5 236.7 -24.3 237.0 ;
        RECT  -33.3 234.3 -29.1 235.5 ;
        RECT  -33.3 229.8 -32.1 234.3 ;
        RECT  -28.2 233.4 -27.0 235.8 ;
        RECT  -22.8 235.5 -21.9 248.1 ;
        RECT  -25.5 234.3 -21.9 235.5 ;
        RECT  -30.9 232.2 -29.7 233.4 ;
        RECT  -30.9 231.3 -24.3 232.2 ;
        RECT  -30.9 231.0 -29.1 231.3 ;
        RECT  -25.5 231.0 -24.3 231.3 ;
        RECT  -22.8 229.8 -21.9 234.3 ;
        RECT  -33.3 228.6 -29.1 229.8 ;
        RECT  -33.3 225.0 -32.1 228.6 ;
        RECT  -27.6 227.7 -26.4 228.9 ;
        RECT  -25.5 228.6 -21.9 229.8 ;
        RECT  -30.9 227.4 -25.5 227.7 ;
        RECT  -30.9 226.8 -24.3 227.4 ;
        RECT  -30.9 226.2 -29.1 226.8 ;
        RECT  -26.7 226.5 -24.3 226.8 ;
        RECT  -25.5 226.2 -24.3 226.5 ;
        RECT  -33.3 223.8 -29.1 225.0 ;
        RECT  -33.3 208.8 -32.1 223.8 ;
        RECT  -27.6 223.2 -26.4 225.6 ;
        RECT  -22.8 225.0 -21.9 228.6 ;
        RECT  -25.5 223.8 -21.9 225.0 ;
        RECT  -23.1 222.6 -21.9 223.8 ;
        RECT  -30.9 219.3 -29.7 220.5 ;
        RECT  -28.8 220.2 -26.4 221.4 ;
        RECT  -30.9 218.4 -24.3 219.3 ;
        RECT  -30.9 218.1 -29.1 218.4 ;
        RECT  -25.5 218.1 -24.3 218.4 ;
        RECT  -30.9 216.0 -24.3 216.9 ;
        RECT  -30.9 215.7 -29.1 216.0 ;
        RECT  -26.7 215.7 -24.3 216.0 ;
        RECT  -30.9 213.6 -24.3 214.5 ;
        RECT  -30.9 213.3 -29.1 213.6 ;
        RECT  -26.7 213.3 -24.3 213.6 ;
        RECT  -27.9 211.5 -26.7 212.4 ;
        RECT  -30.9 210.6 -24.3 211.5 ;
        RECT  -30.9 210.3 -27.9 210.6 ;
        RECT  -25.5 210.3 -24.3 210.6 ;
        RECT  -22.8 209.1 -21.9 222.6 ;
        RECT  -30.9 208.8 -29.1 209.1 ;
        RECT  -33.3 207.9 -29.1 208.8 ;
        RECT  -25.5 208.2 -21.9 209.1 ;
        RECT  -25.5 207.9 -24.3 208.2 ;
        RECT  -30.3 206.4 -29.1 207.9 ;
        RECT  -28.2 205.5 -27.0 206.4 ;
        RECT  -33.3 204.6 -21.9 205.5 ;
        RECT  -33.3 204.6 -21.9 205.5 ;
        RECT  -33.3 258.6 -21.9 259.5 ;
        RECT  -16.65 211.2 -14.25 212.4 ;
        RECT  -5.25 211.2 -3.45 212.4 ;
        RECT  -14.4 206.4 -5.55 207.6 ;
        RECT  -9.9 202.2 -9.0 204.3 ;
        RECT  -9.9 207.6 -9.0 214.2 ;
        RECT  -17.55 202.2 -16.65 214.2 ;
        RECT  -3.45 202.2 -2.55 214.2 ;
        RECT  -5.55 204.0 -4.35 205.2 ;
        RECT  -5.55 206.4 -4.35 207.6 ;
        RECT  -5.55 208.8 -4.35 210.0 ;
        RECT  -3.45 204.0 -2.55 204.9 ;
        RECT  -3.45 208.8 -2.55 209.7 ;
        RECT  -5.55 204.0 -3.45 204.9 ;
        RECT  -3.45 204.0 -3.0 204.9 ;
        RECT  -3.45 204.45 -2.55 209.25 ;
        RECT  -5.55 208.8 -3.0 209.7 ;
        RECT  -3.45 204.0 -2.55 209.7 ;
        RECT  -6.75 204.0 -5.55 205.2 ;
        RECT  -6.75 206.4 -5.55 207.6 ;
        RECT  -6.75 208.8 -5.55 210.0 ;
        RECT  -15.45 204.0 -14.25 205.2 ;
        RECT  -15.45 206.4 -14.25 207.6 ;
        RECT  -15.45 208.8 -14.25 210.0 ;
        RECT  -17.25 204.0 -16.35 204.9 ;
        RECT  -17.25 208.8 -16.35 209.7 ;
        RECT  -16.35 204.0 -14.25 204.9 ;
        RECT  -16.8 204.0 -16.35 204.9 ;
        RECT  -17.25 204.45 -16.35 209.25 ;
        RECT  -16.8 208.8 -14.25 209.7 ;
        RECT  -17.25 204.0 -16.35 209.7 ;
        RECT  -15.45 204.0 -14.25 205.2 ;
        RECT  -15.45 206.4 -14.25 207.6 ;
        RECT  -15.45 208.8 -14.25 210.0 ;
        RECT  -15.45 211.2 -14.25 212.4 ;
        RECT  -5.55 211.2 -4.35 212.4 ;
        RECT  -10.05 204.3 -8.85 205.5 ;
        RECT  -16.65 228.0 -14.25 229.2 ;
        RECT  -5.25 228.0 -3.45 229.2 ;
        RECT  -14.4 218.4 -5.55 219.6 ;
        RECT  -14.4 223.2 -5.55 224.4 ;
        RECT  -9.9 214.2 -9.0 216.3 ;
        RECT  -9.9 224.4 -9.0 231.0 ;
        RECT  -17.55 214.2 -16.65 231.0 ;
        RECT  -3.45 214.2 -2.55 231.0 ;
        RECT  -5.55 216.0 -4.35 217.2 ;
        RECT  -5.55 218.4 -4.35 219.6 ;
        RECT  -5.55 220.8 -4.35 222.0 ;
        RECT  -5.55 223.2 -4.35 224.4 ;
        RECT  -5.55 225.6 -4.35 226.8 ;
        RECT  -3.45 216.0 -2.55 216.9 ;
        RECT  -3.45 220.8 -2.55 221.7 ;
        RECT  -3.45 220.8 -2.55 221.7 ;
        RECT  -3.45 225.6 -2.55 226.5 ;
        RECT  -5.55 216.0 -3.45 216.9 ;
        RECT  -3.45 216.0 -3.0 216.9 ;
        RECT  -3.45 216.45 -2.55 221.25 ;
        RECT  -5.55 220.8 -3.0 221.7 ;
        RECT  -5.55 220.8 -3.45 221.7 ;
        RECT  -3.45 220.8 -3.0 221.7 ;
        RECT  -3.45 221.25 -2.55 226.05 ;
        RECT  -5.55 225.6 -3.0 226.5 ;
        RECT  -7.35 218.4 -6.45 219.3 ;
        RECT  -7.35 223.2 -6.45 224.1 ;
        RECT  -6.45 218.4 -5.55 219.3 ;
        RECT  -6.9 218.4 -6.45 219.3 ;
        RECT  -7.35 218.85 -6.45 223.65 ;
        RECT  -6.9 223.2 -5.55 224.1 ;
        RECT  -3.45 216.0 -2.55 226.5 ;
        RECT  -7.35 218.4 -6.45 224.1 ;
        RECT  -6.75 216.0 -5.55 217.2 ;
        RECT  -6.75 218.4 -5.55 219.6 ;
        RECT  -6.75 220.8 -5.55 222.0 ;
        RECT  -6.75 223.2 -5.55 224.4 ;
        RECT  -6.75 225.6 -5.55 226.8 ;
        RECT  -15.45 216.0 -14.25 217.2 ;
        RECT  -15.45 218.4 -14.25 219.6 ;
        RECT  -15.45 220.8 -14.25 222.0 ;
        RECT  -15.45 223.2 -14.25 224.4 ;
        RECT  -15.45 225.6 -14.25 226.8 ;
        RECT  -17.25 216.0 -16.35 216.9 ;
        RECT  -17.25 220.8 -16.35 221.7 ;
        RECT  -17.25 220.8 -16.35 221.7 ;
        RECT  -17.25 225.6 -16.35 226.5 ;
        RECT  -16.35 216.0 -14.25 216.9 ;
        RECT  -16.8 216.0 -16.35 216.9 ;
        RECT  -17.25 216.45 -16.35 221.25 ;
        RECT  -16.8 220.8 -14.25 221.7 ;
        RECT  -16.35 220.8 -14.25 221.7 ;
        RECT  -16.8 220.8 -16.35 221.7 ;
        RECT  -17.25 221.25 -16.35 226.05 ;
        RECT  -16.8 225.6 -14.25 226.5 ;
        RECT  -13.35 218.4 -12.45 219.3 ;
        RECT  -13.35 223.2 -12.45 224.1 ;
        RECT  -14.25 218.4 -13.35 219.3 ;
        RECT  -13.35 218.4 -12.9 219.3 ;
        RECT  -13.35 218.85 -12.45 223.65 ;
        RECT  -14.25 223.2 -12.9 224.1 ;
        RECT  -17.25 216.0 -16.35 226.5 ;
        RECT  -13.35 218.4 -12.45 224.1 ;
        RECT  -15.45 216.0 -14.25 217.2 ;
        RECT  -15.45 218.4 -14.25 219.6 ;
        RECT  -15.45 220.8 -14.25 222.0 ;
        RECT  -15.45 223.2 -14.25 224.4 ;
        RECT  -15.45 225.6 -14.25 226.8 ;
        RECT  -15.45 228.0 -14.25 229.2 ;
        RECT  -5.55 228.0 -4.35 229.2 ;
        RECT  -10.05 216.3 -8.85 217.5 ;
        RECT  -16.65 254.4 -14.25 255.6 ;
        RECT  -5.25 254.4 -3.45 255.6 ;
        RECT  -14.4 235.2 -5.55 236.4 ;
        RECT  -14.4 240.0 -5.55 241.2 ;
        RECT  -14.4 244.8 -5.55 246.0 ;
        RECT  -14.4 249.6 -5.55 250.8 ;
        RECT  -9.9 231.0 -9.0 233.1 ;
        RECT  -9.9 250.8 -9.0 257.4 ;
        RECT  -17.55 231.0 -16.65 257.4 ;
        RECT  -3.45 231.0 -2.55 257.4 ;
        RECT  -5.55 232.8 -4.35 234.0 ;
        RECT  -5.55 235.2 -4.35 236.4 ;
        RECT  -5.55 237.6 -4.35 238.8 ;
        RECT  -5.55 240.0 -4.35 241.2 ;
        RECT  -5.55 242.4 -4.35 243.6 ;
        RECT  -5.55 244.8 -4.35 246.0 ;
        RECT  -5.55 247.2 -4.35 248.4 ;
        RECT  -5.55 249.6 -4.35 250.8 ;
        RECT  -5.55 252.0 -4.35 253.2 ;
        RECT  -3.45 232.8 -2.55 233.7 ;
        RECT  -3.45 237.6 -2.55 238.5 ;
        RECT  -3.45 237.6 -2.55 238.5 ;
        RECT  -3.45 242.4 -2.55 243.3 ;
        RECT  -3.45 242.4 -2.55 243.3 ;
        RECT  -3.45 247.2 -2.55 248.1 ;
        RECT  -3.45 247.2 -2.55 248.1 ;
        RECT  -3.45 252.0 -2.55 252.9 ;
        RECT  -5.55 232.8 -3.45 233.7 ;
        RECT  -3.45 232.8 -3.0 233.7 ;
        RECT  -3.45 233.25 -2.55 238.05 ;
        RECT  -5.55 237.6 -3.0 238.5 ;
        RECT  -5.55 237.6 -3.45 238.5 ;
        RECT  -3.45 237.6 -3.0 238.5 ;
        RECT  -3.45 238.05 -2.55 242.85 ;
        RECT  -5.55 242.4 -3.0 243.3 ;
        RECT  -5.55 242.4 -3.45 243.3 ;
        RECT  -3.45 242.4 -3.0 243.3 ;
        RECT  -3.45 242.85 -2.55 247.65 ;
        RECT  -5.55 247.2 -3.0 248.1 ;
        RECT  -5.55 247.2 -3.45 248.1 ;
        RECT  -3.45 247.2 -3.0 248.1 ;
        RECT  -3.45 247.65 -2.55 252.45 ;
        RECT  -5.55 252.0 -3.0 252.9 ;
        RECT  -7.35 235.2 -6.45 236.1 ;
        RECT  -7.35 240.0 -6.45 240.9 ;
        RECT  -7.35 240.0 -6.45 240.9 ;
        RECT  -7.35 244.8 -6.45 245.7 ;
        RECT  -7.35 244.8 -6.45 245.7 ;
        RECT  -7.35 249.6 -6.45 250.5 ;
        RECT  -6.45 235.2 -5.55 236.1 ;
        RECT  -6.9 235.2 -6.45 236.1 ;
        RECT  -7.35 235.65 -6.45 240.45 ;
        RECT  -6.9 240.0 -5.55 240.9 ;
        RECT  -6.45 240.0 -5.55 240.9 ;
        RECT  -6.9 240.0 -6.45 240.9 ;
        RECT  -7.35 240.45 -6.45 245.25 ;
        RECT  -6.9 244.8 -5.55 245.7 ;
        RECT  -6.45 244.8 -5.55 245.7 ;
        RECT  -6.9 244.8 -6.45 245.7 ;
        RECT  -7.35 245.25 -6.45 250.05 ;
        RECT  -6.9 249.6 -5.55 250.5 ;
        RECT  -3.45 232.8 -2.55 252.9 ;
        RECT  -7.35 235.2 -6.45 250.5 ;
        RECT  -6.75 232.8 -5.55 234.0 ;
        RECT  -6.75 235.2 -5.55 236.4 ;
        RECT  -6.75 237.6 -5.55 238.8 ;
        RECT  -6.75 240.0 -5.55 241.2 ;
        RECT  -6.75 242.4 -5.55 243.6 ;
        RECT  -6.75 244.8 -5.55 246.0 ;
        RECT  -6.75 247.2 -5.55 248.4 ;
        RECT  -6.75 249.6 -5.55 250.8 ;
        RECT  -6.75 252.0 -5.55 253.2 ;
        RECT  -15.45 232.8 -14.25 234.0 ;
        RECT  -15.45 235.2 -14.25 236.4 ;
        RECT  -15.45 237.6 -14.25 238.8 ;
        RECT  -15.45 240.0 -14.25 241.2 ;
        RECT  -15.45 242.4 -14.25 243.6 ;
        RECT  -15.45 244.8 -14.25 246.0 ;
        RECT  -15.45 247.2 -14.25 248.4 ;
        RECT  -15.45 249.6 -14.25 250.8 ;
        RECT  -15.45 252.0 -14.25 253.2 ;
        RECT  -17.25 232.8 -16.35 233.7 ;
        RECT  -17.25 237.6 -16.35 238.5 ;
        RECT  -17.25 237.6 -16.35 238.5 ;
        RECT  -17.25 242.4 -16.35 243.3 ;
        RECT  -17.25 242.4 -16.35 243.3 ;
        RECT  -17.25 247.2 -16.35 248.1 ;
        RECT  -17.25 247.2 -16.35 248.1 ;
        RECT  -17.25 252.0 -16.35 252.9 ;
        RECT  -16.35 232.8 -14.25 233.7 ;
        RECT  -16.8 232.8 -16.35 233.7 ;
        RECT  -17.25 233.25 -16.35 238.05 ;
        RECT  -16.8 237.6 -14.25 238.5 ;
        RECT  -16.35 237.6 -14.25 238.5 ;
        RECT  -16.8 237.6 -16.35 238.5 ;
        RECT  -17.25 238.05 -16.35 242.85 ;
        RECT  -16.8 242.4 -14.25 243.3 ;
        RECT  -16.35 242.4 -14.25 243.3 ;
        RECT  -16.8 242.4 -16.35 243.3 ;
        RECT  -17.25 242.85 -16.35 247.65 ;
        RECT  -16.8 247.2 -14.25 248.1 ;
        RECT  -16.35 247.2 -14.25 248.1 ;
        RECT  -16.8 247.2 -16.35 248.1 ;
        RECT  -17.25 247.65 -16.35 252.45 ;
        RECT  -16.8 252.0 -14.25 252.9 ;
        RECT  -13.35 235.2 -12.45 236.1 ;
        RECT  -13.35 240.0 -12.45 240.9 ;
        RECT  -13.35 240.0 -12.45 240.9 ;
        RECT  -13.35 244.8 -12.45 245.7 ;
        RECT  -13.35 244.8 -12.45 245.7 ;
        RECT  -13.35 249.6 -12.45 250.5 ;
        RECT  -14.25 235.2 -13.35 236.1 ;
        RECT  -13.35 235.2 -12.9 236.1 ;
        RECT  -13.35 235.65 -12.45 240.45 ;
        RECT  -14.25 240.0 -12.9 240.9 ;
        RECT  -14.25 240.0 -13.35 240.9 ;
        RECT  -13.35 240.0 -12.9 240.9 ;
        RECT  -13.35 240.45 -12.45 245.25 ;
        RECT  -14.25 244.8 -12.9 245.7 ;
        RECT  -14.25 244.8 -13.35 245.7 ;
        RECT  -13.35 244.8 -12.9 245.7 ;
        RECT  -13.35 245.25 -12.45 250.05 ;
        RECT  -14.25 249.6 -12.9 250.5 ;
        RECT  -17.25 232.8 -16.35 252.9 ;
        RECT  -13.35 235.2 -12.45 250.5 ;
        RECT  -15.45 232.8 -14.25 234.0 ;
        RECT  -15.45 235.2 -14.25 236.4 ;
        RECT  -15.45 237.6 -14.25 238.8 ;
        RECT  -15.45 240.0 -14.25 241.2 ;
        RECT  -15.45 242.4 -14.25 243.6 ;
        RECT  -15.45 244.8 -14.25 246.0 ;
        RECT  -15.45 247.2 -14.25 248.4 ;
        RECT  -15.45 249.6 -14.25 250.8 ;
        RECT  -15.45 252.0 -14.25 253.2 ;
        RECT  -15.45 254.4 -14.25 255.6 ;
        RECT  -5.55 254.4 -4.35 255.6 ;
        RECT  -10.05 233.1 -8.85 234.3 ;
        RECT  -16.65 300.0 -14.25 301.2 ;
        RECT  -5.25 300.0 -3.45 301.2 ;
        RECT  -14.4 261.6 -5.55 262.8 ;
        RECT  -14.4 266.4 -5.55 267.6 ;
        RECT  -14.4 271.2 -5.55 272.4 ;
        RECT  -14.4 276.0 -5.55 277.2 ;
        RECT  -14.4 280.8 -5.55 282.0 ;
        RECT  -14.4 285.6 -5.55 286.8 ;
        RECT  -14.4 290.4 -5.55 291.6 ;
        RECT  -14.4 295.2 -5.55 296.4 ;
        RECT  -9.9 257.4 -9.0 259.5 ;
        RECT  -9.9 296.4 -9.0 303.0 ;
        RECT  -17.55 257.4 -16.65 303.0 ;
        RECT  -3.45 257.4 -2.55 303.0 ;
        RECT  -5.55 259.2 -4.35 260.4 ;
        RECT  -5.55 261.6 -4.35 262.8 ;
        RECT  -5.55 264.0 -4.35 265.2 ;
        RECT  -5.55 266.4 -4.35 267.6 ;
        RECT  -5.55 268.8 -4.35 270.0 ;
        RECT  -5.55 271.2 -4.35 272.4 ;
        RECT  -5.55 273.6 -4.35 274.8 ;
        RECT  -5.55 276.0 -4.35 277.2 ;
        RECT  -5.55 278.4 -4.35 279.6 ;
        RECT  -5.55 280.8 -4.35 282.0 ;
        RECT  -5.55 283.2 -4.35 284.4 ;
        RECT  -5.55 285.6 -4.35 286.8 ;
        RECT  -5.55 288.0 -4.35 289.2 ;
        RECT  -5.55 290.4 -4.35 291.6 ;
        RECT  -5.55 292.8 -4.35 294.0 ;
        RECT  -5.55 295.2 -4.35 296.4 ;
        RECT  -5.55 297.6 -4.35 298.8 ;
        RECT  -3.45 259.2 -2.55 260.1 ;
        RECT  -3.45 264.0 -2.55 264.9 ;
        RECT  -3.45 264.0 -2.55 264.9 ;
        RECT  -3.45 268.8 -2.55 269.7 ;
        RECT  -3.45 268.8 -2.55 269.7 ;
        RECT  -3.45 273.6 -2.55 274.5 ;
        RECT  -3.45 273.6 -2.55 274.5 ;
        RECT  -3.45 278.4 -2.55 279.3 ;
        RECT  -3.45 278.4 -2.55 279.3 ;
        RECT  -3.45 283.2 -2.55 284.1 ;
        RECT  -3.45 283.2 -2.55 284.1 ;
        RECT  -3.45 288.0 -2.55 288.9 ;
        RECT  -3.45 288.0 -2.55 288.9 ;
        RECT  -3.45 292.8 -2.55 293.7 ;
        RECT  -3.45 292.8 -2.55 293.7 ;
        RECT  -3.45 297.6 -2.55 298.5 ;
        RECT  -5.55 259.2 -3.45 260.1 ;
        RECT  -3.45 259.2 -3.0 260.1 ;
        RECT  -3.45 259.65 -2.55 264.45 ;
        RECT  -5.55 264.0 -3.0 264.9 ;
        RECT  -5.55 264.0 -3.45 264.9 ;
        RECT  -3.45 264.0 -3.0 264.9 ;
        RECT  -3.45 264.45 -2.55 269.25 ;
        RECT  -5.55 268.8 -3.0 269.7 ;
        RECT  -5.55 268.8 -3.45 269.7 ;
        RECT  -3.45 268.8 -3.0 269.7 ;
        RECT  -3.45 269.25 -2.55 274.05 ;
        RECT  -5.55 273.6 -3.0 274.5 ;
        RECT  -5.55 273.6 -3.45 274.5 ;
        RECT  -3.45 273.6 -3.0 274.5 ;
        RECT  -3.45 274.05 -2.55 278.85 ;
        RECT  -5.55 278.4 -3.0 279.3 ;
        RECT  -5.55 278.4 -3.45 279.3 ;
        RECT  -3.45 278.4 -3.0 279.3 ;
        RECT  -3.45 278.85 -2.55 283.65 ;
        RECT  -5.55 283.2 -3.0 284.1 ;
        RECT  -5.55 283.2 -3.45 284.1 ;
        RECT  -3.45 283.2 -3.0 284.1 ;
        RECT  -3.45 283.65 -2.55 288.45 ;
        RECT  -5.55 288.0 -3.0 288.9 ;
        RECT  -5.55 288.0 -3.45 288.9 ;
        RECT  -3.45 288.0 -3.0 288.9 ;
        RECT  -3.45 288.45 -2.55 293.25 ;
        RECT  -5.55 292.8 -3.0 293.7 ;
        RECT  -5.55 292.8 -3.45 293.7 ;
        RECT  -3.45 292.8 -3.0 293.7 ;
        RECT  -3.45 293.25 -2.55 298.05 ;
        RECT  -5.55 297.6 -3.0 298.5 ;
        RECT  -7.35 261.6 -6.45 262.5 ;
        RECT  -7.35 266.4 -6.45 267.3 ;
        RECT  -7.35 266.4 -6.45 267.3 ;
        RECT  -7.35 271.2 -6.45 272.1 ;
        RECT  -7.35 271.2 -6.45 272.1 ;
        RECT  -7.35 276.0 -6.45 276.9 ;
        RECT  -7.35 276.0 -6.45 276.9 ;
        RECT  -7.35 280.8 -6.45 281.7 ;
        RECT  -7.35 280.8 -6.45 281.7 ;
        RECT  -7.35 285.6 -6.45 286.5 ;
        RECT  -7.35 285.6 -6.45 286.5 ;
        RECT  -7.35 290.4 -6.45 291.3 ;
        RECT  -7.35 290.4 -6.45 291.3 ;
        RECT  -7.35 295.2 -6.45 296.1 ;
        RECT  -6.45 261.6 -5.55 262.5 ;
        RECT  -6.9 261.6 -6.45 262.5 ;
        RECT  -7.35 262.05 -6.45 266.85 ;
        RECT  -6.9 266.4 -5.55 267.3 ;
        RECT  -6.45 266.4 -5.55 267.3 ;
        RECT  -6.9 266.4 -6.45 267.3 ;
        RECT  -7.35 266.85 -6.45 271.65 ;
        RECT  -6.9 271.2 -5.55 272.1 ;
        RECT  -6.45 271.2 -5.55 272.1 ;
        RECT  -6.9 271.2 -6.45 272.1 ;
        RECT  -7.35 271.65 -6.45 276.45 ;
        RECT  -6.9 276.0 -5.55 276.9 ;
        RECT  -6.45 276.0 -5.55 276.9 ;
        RECT  -6.9 276.0 -6.45 276.9 ;
        RECT  -7.35 276.45 -6.45 281.25 ;
        RECT  -6.9 280.8 -5.55 281.7 ;
        RECT  -6.45 280.8 -5.55 281.7 ;
        RECT  -6.9 280.8 -6.45 281.7 ;
        RECT  -7.35 281.25 -6.45 286.05 ;
        RECT  -6.9 285.6 -5.55 286.5 ;
        RECT  -6.45 285.6 -5.55 286.5 ;
        RECT  -6.9 285.6 -6.45 286.5 ;
        RECT  -7.35 286.05 -6.45 290.85 ;
        RECT  -6.9 290.4 -5.55 291.3 ;
        RECT  -6.45 290.4 -5.55 291.3 ;
        RECT  -6.9 290.4 -6.45 291.3 ;
        RECT  -7.35 290.85 -6.45 295.65 ;
        RECT  -6.9 295.2 -5.55 296.1 ;
        RECT  -3.45 259.2 -2.55 298.5 ;
        RECT  -7.35 261.6 -6.45 296.1 ;
        RECT  -6.75 259.2 -5.55 260.4 ;
        RECT  -6.75 261.6 -5.55 262.8 ;
        RECT  -6.75 264.0 -5.55 265.2 ;
        RECT  -6.75 266.4 -5.55 267.6 ;
        RECT  -6.75 268.8 -5.55 270.0 ;
        RECT  -6.75 271.2 -5.55 272.4 ;
        RECT  -6.75 273.6 -5.55 274.8 ;
        RECT  -6.75 276.0 -5.55 277.2 ;
        RECT  -6.75 278.4 -5.55 279.6 ;
        RECT  -6.75 280.8 -5.55 282.0 ;
        RECT  -6.75 283.2 -5.55 284.4 ;
        RECT  -6.75 285.6 -5.55 286.8 ;
        RECT  -6.75 288.0 -5.55 289.2 ;
        RECT  -6.75 290.4 -5.55 291.6 ;
        RECT  -6.75 292.8 -5.55 294.0 ;
        RECT  -6.75 295.2 -5.55 296.4 ;
        RECT  -6.75 297.6 -5.55 298.8 ;
        RECT  -15.45 259.2 -14.25 260.4 ;
        RECT  -15.45 261.6 -14.25 262.8 ;
        RECT  -15.45 264.0 -14.25 265.2 ;
        RECT  -15.45 266.4 -14.25 267.6 ;
        RECT  -15.45 268.8 -14.25 270.0 ;
        RECT  -15.45 271.2 -14.25 272.4 ;
        RECT  -15.45 273.6 -14.25 274.8 ;
        RECT  -15.45 276.0 -14.25 277.2 ;
        RECT  -15.45 278.4 -14.25 279.6 ;
        RECT  -15.45 280.8 -14.25 282.0 ;
        RECT  -15.45 283.2 -14.25 284.4 ;
        RECT  -15.45 285.6 -14.25 286.8 ;
        RECT  -15.45 288.0 -14.25 289.2 ;
        RECT  -15.45 290.4 -14.25 291.6 ;
        RECT  -15.45 292.8 -14.25 294.0 ;
        RECT  -15.45 295.2 -14.25 296.4 ;
        RECT  -15.45 297.6 -14.25 298.8 ;
        RECT  -17.25 259.2 -16.35 260.1 ;
        RECT  -17.25 264.0 -16.35 264.9 ;
        RECT  -17.25 264.0 -16.35 264.9 ;
        RECT  -17.25 268.8 -16.35 269.7 ;
        RECT  -17.25 268.8 -16.35 269.7 ;
        RECT  -17.25 273.6 -16.35 274.5 ;
        RECT  -17.25 273.6 -16.35 274.5 ;
        RECT  -17.25 278.4 -16.35 279.3 ;
        RECT  -17.25 278.4 -16.35 279.3 ;
        RECT  -17.25 283.2 -16.35 284.1 ;
        RECT  -17.25 283.2 -16.35 284.1 ;
        RECT  -17.25 288.0 -16.35 288.9 ;
        RECT  -17.25 288.0 -16.35 288.9 ;
        RECT  -17.25 292.8 -16.35 293.7 ;
        RECT  -17.25 292.8 -16.35 293.7 ;
        RECT  -17.25 297.6 -16.35 298.5 ;
        RECT  -16.35 259.2 -14.25 260.1 ;
        RECT  -16.8 259.2 -16.35 260.1 ;
        RECT  -17.25 259.65 -16.35 264.45 ;
        RECT  -16.8 264.0 -14.25 264.9 ;
        RECT  -16.35 264.0 -14.25 264.9 ;
        RECT  -16.8 264.0 -16.35 264.9 ;
        RECT  -17.25 264.45 -16.35 269.25 ;
        RECT  -16.8 268.8 -14.25 269.7 ;
        RECT  -16.35 268.8 -14.25 269.7 ;
        RECT  -16.8 268.8 -16.35 269.7 ;
        RECT  -17.25 269.25 -16.35 274.05 ;
        RECT  -16.8 273.6 -14.25 274.5 ;
        RECT  -16.35 273.6 -14.25 274.5 ;
        RECT  -16.8 273.6 -16.35 274.5 ;
        RECT  -17.25 274.05 -16.35 278.85 ;
        RECT  -16.8 278.4 -14.25 279.3 ;
        RECT  -16.35 278.4 -14.25 279.3 ;
        RECT  -16.8 278.4 -16.35 279.3 ;
        RECT  -17.25 278.85 -16.35 283.65 ;
        RECT  -16.8 283.2 -14.25 284.1 ;
        RECT  -16.35 283.2 -14.25 284.1 ;
        RECT  -16.8 283.2 -16.35 284.1 ;
        RECT  -17.25 283.65 -16.35 288.45 ;
        RECT  -16.8 288.0 -14.25 288.9 ;
        RECT  -16.35 288.0 -14.25 288.9 ;
        RECT  -16.8 288.0 -16.35 288.9 ;
        RECT  -17.25 288.45 -16.35 293.25 ;
        RECT  -16.8 292.8 -14.25 293.7 ;
        RECT  -16.35 292.8 -14.25 293.7 ;
        RECT  -16.8 292.8 -16.35 293.7 ;
        RECT  -17.25 293.25 -16.35 298.05 ;
        RECT  -16.8 297.6 -14.25 298.5 ;
        RECT  -13.35 261.6 -12.45 262.5 ;
        RECT  -13.35 266.4 -12.45 267.3 ;
        RECT  -13.35 266.4 -12.45 267.3 ;
        RECT  -13.35 271.2 -12.45 272.1 ;
        RECT  -13.35 271.2 -12.45 272.1 ;
        RECT  -13.35 276.0 -12.45 276.9 ;
        RECT  -13.35 276.0 -12.45 276.9 ;
        RECT  -13.35 280.8 -12.45 281.7 ;
        RECT  -13.35 280.8 -12.45 281.7 ;
        RECT  -13.35 285.6 -12.45 286.5 ;
        RECT  -13.35 285.6 -12.45 286.5 ;
        RECT  -13.35 290.4 -12.45 291.3 ;
        RECT  -13.35 290.4 -12.45 291.3 ;
        RECT  -13.35 295.2 -12.45 296.1 ;
        RECT  -14.25 261.6 -13.35 262.5 ;
        RECT  -13.35 261.6 -12.9 262.5 ;
        RECT  -13.35 262.05 -12.45 266.85 ;
        RECT  -14.25 266.4 -12.9 267.3 ;
        RECT  -14.25 266.4 -13.35 267.3 ;
        RECT  -13.35 266.4 -12.9 267.3 ;
        RECT  -13.35 266.85 -12.45 271.65 ;
        RECT  -14.25 271.2 -12.9 272.1 ;
        RECT  -14.25 271.2 -13.35 272.1 ;
        RECT  -13.35 271.2 -12.9 272.1 ;
        RECT  -13.35 271.65 -12.45 276.45 ;
        RECT  -14.25 276.0 -12.9 276.9 ;
        RECT  -14.25 276.0 -13.35 276.9 ;
        RECT  -13.35 276.0 -12.9 276.9 ;
        RECT  -13.35 276.45 -12.45 281.25 ;
        RECT  -14.25 280.8 -12.9 281.7 ;
        RECT  -14.25 280.8 -13.35 281.7 ;
        RECT  -13.35 280.8 -12.9 281.7 ;
        RECT  -13.35 281.25 -12.45 286.05 ;
        RECT  -14.25 285.6 -12.9 286.5 ;
        RECT  -14.25 285.6 -13.35 286.5 ;
        RECT  -13.35 285.6 -12.9 286.5 ;
        RECT  -13.35 286.05 -12.45 290.85 ;
        RECT  -14.25 290.4 -12.9 291.3 ;
        RECT  -14.25 290.4 -13.35 291.3 ;
        RECT  -13.35 290.4 -12.9 291.3 ;
        RECT  -13.35 290.85 -12.45 295.65 ;
        RECT  -14.25 295.2 -12.9 296.1 ;
        RECT  -17.25 259.2 -16.35 298.5 ;
        RECT  -13.35 261.6 -12.45 296.1 ;
        RECT  -15.45 259.2 -14.25 260.4 ;
        RECT  -15.45 261.6 -14.25 262.8 ;
        RECT  -15.45 264.0 -14.25 265.2 ;
        RECT  -15.45 266.4 -14.25 267.6 ;
        RECT  -15.45 268.8 -14.25 270.0 ;
        RECT  -15.45 271.2 -14.25 272.4 ;
        RECT  -15.45 273.6 -14.25 274.8 ;
        RECT  -15.45 276.0 -14.25 277.2 ;
        RECT  -15.45 278.4 -14.25 279.6 ;
        RECT  -15.45 280.8 -14.25 282.0 ;
        RECT  -15.45 283.2 -14.25 284.4 ;
        RECT  -15.45 285.6 -14.25 286.8 ;
        RECT  -15.45 288.0 -14.25 289.2 ;
        RECT  -15.45 290.4 -14.25 291.6 ;
        RECT  -15.45 292.8 -14.25 294.0 ;
        RECT  -15.45 295.2 -14.25 296.4 ;
        RECT  -15.45 297.6 -14.25 298.8 ;
        RECT  -15.45 300.0 -14.25 301.2 ;
        RECT  -5.55 300.0 -4.35 301.2 ;
        RECT  -10.05 259.5 -8.85 260.7 ;
        RECT  -15.3 340.8 -4.8 341.7 ;
        RECT  -17.1 342.6 -14.25 343.5 ;
        RECT  -6.6 342.6 -3.0 343.5 ;
        RECT  -17.1 333.15 -14.25 334.05 ;
        RECT  -17.1 337.95 -14.25 338.85 ;
        RECT  -5.85 333.15 -3.0 334.05 ;
        RECT  -12.75 330.0 -11.85 334.5 ;
        RECT  -8.55 330.0 -7.65 339.3 ;
        RECT  -10.65 330.0 -9.75 336.9 ;
        RECT  -17.55 330.0 -16.65 345.6 ;
        RECT  -3.45 330.0 -2.55 345.6 ;
        RECT  -10.65 340.8 -9.75 345.6 ;
        RECT  -6.45 333.0 -5.25 334.2 ;
        RECT  -6.45 335.4 -5.25 336.6 ;
        RECT  -7.65 333.0 -6.45 334.2 ;
        RECT  -7.65 335.4 -6.45 336.6 ;
        RECT  -6.45 335.4 -5.25 336.6 ;
        RECT  -6.45 337.8 -5.25 339.0 ;
        RECT  -7.65 335.4 -6.45 336.6 ;
        RECT  -7.65 337.8 -6.45 339.0 ;
        RECT  -6.45 337.8 -5.25 339.0 ;
        RECT  -6.45 340.2 -5.25 341.4 ;
        RECT  -7.65 337.8 -6.45 339.0 ;
        RECT  -7.65 340.2 -6.45 341.4 ;
        RECT  -15.45 333.0 -14.25 334.2 ;
        RECT  -15.45 335.4 -14.25 336.6 ;
        RECT  -15.45 333.0 -14.25 334.2 ;
        RECT  -15.45 335.4 -14.25 336.6 ;
        RECT  -15.45 335.4 -14.25 336.6 ;
        RECT  -15.45 337.8 -14.25 339.0 ;
        RECT  -15.45 335.4 -14.25 336.6 ;
        RECT  -15.45 337.8 -14.25 339.0 ;
        RECT  -15.45 337.8 -14.25 339.0 ;
        RECT  -15.45 340.2 -14.25 341.4 ;
        RECT  -15.45 337.8 -14.25 339.0 ;
        RECT  -15.45 340.2 -14.25 341.4 ;
        RECT  -15.45 342.6 -14.25 343.8 ;
        RECT  -6.45 342.6 -5.25 343.8 ;
        RECT  -15.45 335.4 -14.25 336.6 ;
        RECT  -15.45 340.2 -14.25 341.4 ;
        RECT  -13.05 333.9 -11.85 335.1 ;
        RECT  -10.95 336.3 -9.75 337.5 ;
        RECT  -8.85 338.7 -7.65 339.9 ;
        RECT  -16.65 352.2 -14.25 353.4 ;
        RECT  -5.25 352.2 -3.45 353.4 ;
        RECT  -4.35 347.4 -3.45 348.6 ;
        RECT  -16.65 347.4 -15.45 348.6 ;
        RECT  -14.4 349.8 -5.55 351.0 ;
        RECT  -9.9 345.6 -9.0 347.7 ;
        RECT  -9.9 351.0 -9.0 355.2 ;
        RECT  -17.55 345.6 -16.65 355.2 ;
        RECT  -3.45 345.6 -2.55 355.2 ;
        RECT  -5.55 347.4 -4.35 348.6 ;
        RECT  -5.55 349.8 -4.35 351.0 ;
        RECT  -6.75 347.4 -5.55 348.6 ;
        RECT  -6.75 349.8 -5.55 351.0 ;
        RECT  -15.45 347.4 -14.25 348.6 ;
        RECT  -15.45 349.8 -14.25 351.0 ;
        RECT  -15.45 347.4 -14.25 348.6 ;
        RECT  -15.45 349.8 -14.25 351.0 ;
        RECT  -15.45 352.2 -14.25 353.4 ;
        RECT  -5.55 352.2 -4.35 353.4 ;
        RECT  -10.05 347.7 -8.85 348.9 ;
        RECT  -27.3 334.35 -26.4 335.25 ;
        RECT  -27.3 334.8 -26.4 346.8 ;
        RECT  -29.85 334.35 -26.85 335.25 ;
        RECT  -27.3 342.0 -26.4 346.8 ;
        RECT  -21.3 343.8 -17.1 344.7 ;
        RECT  -31.2 339.0 -29.85 339.9 ;
        RECT  -21.3 331.8 -17.55 332.7 ;
        RECT  -23.1 334.35 -22.2 335.25 ;
        RECT  -22.65 334.35 -21.3 335.25 ;
        RECT  -23.1 334.8 -22.2 337.2 ;
        RECT  -23.1 339.15 -22.2 340.05 ;
        RECT  -22.65 339.15 -21.3 340.05 ;
        RECT  -23.1 337.2 -22.2 339.6 ;
        RECT  -31.65 331.8 -29.85 332.7 ;
        RECT  -31.65 336.6 -29.85 337.5 ;
        RECT  -27.3 330.0 -26.4 333.3 ;
        RECT  -27.3 342.0 -26.4 346.8 ;
        RECT  -25.2 330.0 -24.3 340.5 ;
        RECT  -17.55 330.0 -16.65 346.8 ;
        RECT  -31.65 330.0 -30.75 346.8 ;
        RECT  -25.05 331.8 -23.85 333.0 ;
        RECT  -25.05 334.2 -23.85 335.4 ;
        RECT  -26.25 331.8 -25.05 333.0 ;
        RECT  -26.25 334.2 -25.05 335.4 ;
        RECT  -25.05 334.2 -23.85 335.4 ;
        RECT  -25.05 336.6 -23.85 337.8 ;
        RECT  -26.25 334.2 -25.05 335.4 ;
        RECT  -26.25 336.6 -25.05 337.8 ;
        RECT  -28.5 331.8 -25.8 333.0 ;
        RECT  -28.5 334.2 -25.8 335.4 ;
        RECT  -28.5 331.8 -25.8 333.0 ;
        RECT  -28.5 334.2 -25.8 335.4 ;
        RECT  -28.5 339.0 -25.8 340.2 ;
        RECT  -28.5 341.4 -25.8 342.6 ;
        RECT  -28.5 339.0 -25.8 340.2 ;
        RECT  -28.5 341.4 -25.8 342.6 ;
        RECT  -24.0 343.8 -21.3 345.0 ;
        RECT  -31.05 339.0 -29.85 340.2 ;
        RECT  -28.65 332.1 -27.45 333.3 ;
        RECT  -26.55 339.3 -25.35 340.5 ;
        RECT  -22.5 341.4 -21.3 342.6 ;
        RECT  -28.65 341.4 -27.45 342.6 ;
        RECT  -19.95 358.5 -17.1 359.4 ;
        RECT  -31.2 358.5 -28.8 359.4 ;
        RECT  -19.95 351.45 -17.1 352.35 ;
        RECT  -19.95 356.25 -17.1 357.15 ;
        RECT  -31.2 351.45 -28.35 352.35 ;
        RECT  -23.1 356.7 -22.2 357.6 ;
        RECT  -23.1 353.7 -22.2 354.6 ;
        RECT  -29.55 356.7 -22.65 357.6 ;
        RECT  -23.1 354.15 -22.2 357.15 ;
        RECT  -22.65 353.7 -19.95 354.6 ;
        RECT  -23.1 349.5 -22.2 351.6 ;
        RECT  -25.2 357.15 -24.3 361.5 ;
        RECT  -25.8 349.5 -24.9 354.6 ;
        RECT  -17.55 349.5 -16.65 361.5 ;
        RECT  -31.65 349.5 -30.75 361.5 ;
        RECT  -23.55 351.3 -22.35 352.5 ;
        RECT  -23.55 353.7 -22.35 354.9 ;
        RECT  -24.75 351.3 -23.55 352.5 ;
        RECT  -24.75 353.7 -23.55 354.9 ;
        RECT  -23.55 353.7 -22.35 354.9 ;
        RECT  -23.55 356.1 -22.35 357.3 ;
        RECT  -24.75 353.7 -23.55 354.9 ;
        RECT  -24.75 356.1 -23.55 357.3 ;
        RECT  -25.95 351.3 -24.75 352.5 ;
        RECT  -25.95 353.7 -24.75 354.9 ;
        RECT  -25.95 351.3 -24.75 352.5 ;
        RECT  -25.95 353.7 -24.75 354.9 ;
        RECT  -25.95 353.7 -24.75 354.9 ;
        RECT  -25.95 356.1 -24.75 357.3 ;
        RECT  -25.95 353.7 -24.75 354.9 ;
        RECT  -25.95 356.1 -24.75 357.3 ;
        RECT  -21.15 358.5 -19.95 359.7 ;
        RECT  -30.75 358.5 -29.55 359.7 ;
        RECT  -24.6 351.6 -23.4 352.8 ;
        RECT  -27.3 354.6 -26.1 355.8 ;
        RECT  -19.95 366.0 -17.55 367.2 ;
        RECT  -30.75 366.0 -28.95 367.2 ;
        RECT  -30.75 370.8 -29.85 372.0 ;
        RECT  -18.75 370.8 -17.55 372.0 ;
        RECT  -28.65 368.4 -19.8 369.6 ;
        RECT  -25.2 371.7 -24.3 373.8 ;
        RECT  -25.2 364.2 -24.3 368.4 ;
        RECT  -17.55 364.2 -16.65 373.8 ;
        RECT  -31.65 364.2 -30.75 373.8 ;
        RECT  -29.85 370.8 -28.65 372.0 ;
        RECT  -29.85 368.4 -28.65 369.6 ;
        RECT  -28.65 370.8 -27.45 372.0 ;
        RECT  -28.65 368.4 -27.45 369.6 ;
        RECT  -19.95 370.8 -18.75 372.0 ;
        RECT  -19.95 368.4 -18.75 369.6 ;
        RECT  -19.95 370.8 -18.75 372.0 ;
        RECT  -19.95 368.4 -18.75 369.6 ;
        RECT  -19.95 366.0 -18.75 367.2 ;
        RECT  -29.85 366.0 -28.65 367.2 ;
        RECT  -25.35 370.5 -24.15 371.7 ;
        RECT  -19.95 375.6 -17.55 376.8 ;
        RECT  -30.75 375.6 -28.95 376.8 ;
        RECT  -30.75 380.4 -29.85 381.6 ;
        RECT  -18.75 380.4 -17.55 381.6 ;
        RECT  -28.65 378.0 -19.8 379.2 ;
        RECT  -25.2 381.3 -24.3 383.4 ;
        RECT  -25.2 373.8 -24.3 378.0 ;
        RECT  -17.55 373.8 -16.65 383.4 ;
        RECT  -31.65 373.8 -30.75 383.4 ;
        RECT  -29.85 380.4 -28.65 381.6 ;
        RECT  -29.85 378.0 -28.65 379.2 ;
        RECT  -28.65 380.4 -27.45 381.6 ;
        RECT  -28.65 378.0 -27.45 379.2 ;
        RECT  -19.95 380.4 -18.75 381.6 ;
        RECT  -19.95 378.0 -18.75 379.2 ;
        RECT  -19.95 380.4 -18.75 381.6 ;
        RECT  -19.95 378.0 -18.75 379.2 ;
        RECT  -19.95 375.6 -18.75 376.8 ;
        RECT  -29.85 375.6 -28.65 376.8 ;
        RECT  -25.35 380.1 -24.15 381.3 ;
        RECT  -43.5 350.4 -33.0 351.3 ;
        RECT  -45.3 352.2 -42.45 353.1 ;
        RECT  -34.8 352.2 -31.2 353.1 ;
        RECT  -45.3 342.75 -42.45 343.65 ;
        RECT  -45.3 347.55 -42.45 348.45 ;
        RECT  -34.05 342.75 -31.2 343.65 ;
        RECT  -40.95 339.6 -40.05 344.1 ;
        RECT  -36.75 339.6 -35.85 348.9 ;
        RECT  -38.85 339.6 -37.95 346.5 ;
        RECT  -45.75 339.6 -44.85 355.2 ;
        RECT  -31.65 339.6 -30.75 355.2 ;
        RECT  -38.85 350.4 -37.95 355.2 ;
        RECT  -34.65 342.6 -33.45 343.8 ;
        RECT  -34.65 345.0 -33.45 346.2 ;
        RECT  -35.85 342.6 -34.65 343.8 ;
        RECT  -35.85 345.0 -34.65 346.2 ;
        RECT  -34.65 345.0 -33.45 346.2 ;
        RECT  -34.65 347.4 -33.45 348.6 ;
        RECT  -35.85 345.0 -34.65 346.2 ;
        RECT  -35.85 347.4 -34.65 348.6 ;
        RECT  -34.65 347.4 -33.45 348.6 ;
        RECT  -34.65 349.8 -33.45 351.0 ;
        RECT  -35.85 347.4 -34.65 348.6 ;
        RECT  -35.85 349.8 -34.65 351.0 ;
        RECT  -43.65 342.6 -42.45 343.8 ;
        RECT  -43.65 345.0 -42.45 346.2 ;
        RECT  -43.65 342.6 -42.45 343.8 ;
        RECT  -43.65 345.0 -42.45 346.2 ;
        RECT  -43.65 345.0 -42.45 346.2 ;
        RECT  -43.65 347.4 -42.45 348.6 ;
        RECT  -43.65 345.0 -42.45 346.2 ;
        RECT  -43.65 347.4 -42.45 348.6 ;
        RECT  -43.65 347.4 -42.45 348.6 ;
        RECT  -43.65 349.8 -42.45 351.0 ;
        RECT  -43.65 347.4 -42.45 348.6 ;
        RECT  -43.65 349.8 -42.45 351.0 ;
        RECT  -43.65 352.2 -42.45 353.4 ;
        RECT  -34.65 352.2 -33.45 353.4 ;
        RECT  -43.65 345.0 -42.45 346.2 ;
        RECT  -43.65 349.8 -42.45 351.0 ;
        RECT  -41.25 343.5 -40.05 344.7 ;
        RECT  -39.15 345.9 -37.95 347.1 ;
        RECT  -37.05 348.3 -35.85 349.5 ;
        RECT  -44.85 361.8 -42.45 363.0 ;
        RECT  -33.45 361.8 -31.65 363.0 ;
        RECT  -32.55 357.0 -31.65 358.2 ;
        RECT  -44.85 357.0 -43.65 358.2 ;
        RECT  -42.6 359.4 -33.75 360.6 ;
        RECT  -38.1 355.2 -37.2 357.3 ;
        RECT  -38.1 360.6 -37.2 364.8 ;
        RECT  -45.75 355.2 -44.85 364.8 ;
        RECT  -31.65 355.2 -30.75 364.8 ;
        RECT  -33.75 357.0 -32.55 358.2 ;
        RECT  -33.75 359.4 -32.55 360.6 ;
        RECT  -34.95 357.0 -33.75 358.2 ;
        RECT  -34.95 359.4 -33.75 360.6 ;
        RECT  -43.65 357.0 -42.45 358.2 ;
        RECT  -43.65 359.4 -42.45 360.6 ;
        RECT  -43.65 357.0 -42.45 358.2 ;
        RECT  -43.65 359.4 -42.45 360.6 ;
        RECT  -43.65 361.8 -42.45 363.0 ;
        RECT  -33.75 361.8 -32.55 363.0 ;
        RECT  -38.25 357.3 -37.05 358.5 ;
        RECT  -44.85 371.4 -42.45 372.6 ;
        RECT  -33.45 371.4 -31.65 372.6 ;
        RECT  -32.55 366.6 -31.65 367.8 ;
        RECT  -44.85 366.6 -43.65 367.8 ;
        RECT  -42.6 369.0 -33.75 370.2 ;
        RECT  -38.1 364.8 -37.2 366.9 ;
        RECT  -38.1 370.2 -37.2 374.4 ;
        RECT  -45.75 364.8 -44.85 374.4 ;
        RECT  -31.65 364.8 -30.75 374.4 ;
        RECT  -33.75 366.6 -32.55 367.8 ;
        RECT  -33.75 369.0 -32.55 370.2 ;
        RECT  -34.95 366.6 -33.75 367.8 ;
        RECT  -34.95 369.0 -33.75 370.2 ;
        RECT  -43.65 366.6 -42.45 367.8 ;
        RECT  -43.65 369.0 -42.45 370.2 ;
        RECT  -43.65 366.6 -42.45 367.8 ;
        RECT  -43.65 369.0 -42.45 370.2 ;
        RECT  -43.65 371.4 -42.45 372.6 ;
        RECT  -33.75 371.4 -32.55 372.6 ;
        RECT  -38.25 366.9 -37.05 368.1 ;
        RECT  -44.85 381.0 -42.45 382.2 ;
        RECT  -33.45 381.0 -31.65 382.2 ;
        RECT  -32.55 376.2 -31.65 377.4 ;
        RECT  -44.85 376.2 -43.65 377.4 ;
        RECT  -42.6 378.6 -33.75 379.8 ;
        RECT  -38.1 374.4 -37.2 376.5 ;
        RECT  -38.1 379.8 -37.2 384.0 ;
        RECT  -45.75 374.4 -44.85 384.0 ;
        RECT  -31.65 374.4 -30.75 384.0 ;
        RECT  -33.75 376.2 -32.55 377.4 ;
        RECT  -33.75 378.6 -32.55 379.8 ;
        RECT  -34.95 376.2 -33.75 377.4 ;
        RECT  -34.95 378.6 -33.75 379.8 ;
        RECT  -43.65 376.2 -42.45 377.4 ;
        RECT  -43.65 378.6 -42.45 379.8 ;
        RECT  -43.65 376.2 -42.45 377.4 ;
        RECT  -43.65 378.6 -42.45 379.8 ;
        RECT  -43.65 381.0 -42.45 382.2 ;
        RECT  -33.75 381.0 -32.55 382.2 ;
        RECT  -38.25 376.5 -37.05 377.7 ;
        RECT  -51.45 262.2 -50.25 263.4 ;
        RECT  -48.75 262.2 -47.55 263.4 ;
        RECT  -35.85 262.2 -34.65 263.4 ;
        RECT  -31.05 262.2 -29.85 263.4 ;
        RECT  -36.6 422.1 -30.75 423.0 ;
        RECT  -36.6 444.9 -30.75 445.8 ;
        RECT  -46.8 450.45 -31.2 451.35 ;
        RECT  -48.9 433.5 -36.6 434.4 ;
        RECT  -48.9 405.3 -36.6 406.2 ;
        RECT  -25.2 420.45 -24.3 421.35 ;
        RECT  -25.2 420.9 -24.3 434.1 ;
        RECT  -24.75 420.45 -24.6 421.35 ;
        RECT  -25.05 416.85 -24.15 417.75 ;
        RECT  -25.05 417.3 -24.15 420.9 ;
        RECT  -36.6 416.85 -24.6 417.75 ;
        RECT  -21.75 421.65 -17.1 422.55 ;
        RECT  -22.2 407.55 -21.3 408.45 ;
        RECT  -25.2 407.55 -24.3 408.45 ;
        RECT  -22.2 408.0 -21.3 419.7 ;
        RECT  -24.75 407.55 -21.75 408.45 ;
        RECT  -25.2 405.3 -24.3 408.0 ;
        RECT  -33.45 407.55 -24.75 408.45 ;
        RECT  -40.2 400.05 -33.45 400.95 ;
        RECT  -9.9 386.1 -9.0 435.0 ;
        RECT  -49.8 386.1 -48.9 448.65 ;
        RECT  -17.55 386.1 -16.65 434.1 ;
        RECT  -31.65 386.1 -30.75 405.3 ;
        RECT  -3.45 386.1 -2.55 434.1 ;
        RECT  -25.2 386.1 -24.3 395.7 ;
        RECT  -19.95 411.9 -17.55 413.1 ;
        RECT  -30.75 411.9 -28.95 413.1 ;
        RECT  -30.75 407.1 -29.85 408.3 ;
        RECT  -18.75 407.1 -17.55 408.3 ;
        RECT  -28.65 409.5 -19.8 410.7 ;
        RECT  -25.2 405.3 -24.3 407.4 ;
        RECT  -25.2 410.7 -24.3 414.9 ;
        RECT  -17.55 405.3 -16.65 414.9 ;
        RECT  -31.65 405.3 -30.75 414.9 ;
        RECT  -25.05 407.1 -23.85 408.3 ;
        RECT  -25.05 409.5 -23.85 410.7 ;
        RECT  -26.25 407.1 -25.05 408.3 ;
        RECT  -26.25 409.5 -25.05 410.7 ;
        RECT  -25.95 407.1 -24.75 408.3 ;
        RECT  -25.95 409.5 -24.75 410.7 ;
        RECT  -25.95 407.1 -24.75 408.3 ;
        RECT  -25.95 409.5 -24.75 410.7 ;
        RECT  -21.15 411.9 -19.95 413.1 ;
        RECT  -31.05 411.9 -29.85 413.1 ;
        RECT  -26.55 407.4 -25.35 408.6 ;
        RECT  -22.35 414.3 -21.15 415.5 ;
        RECT  -22.35 411.9 -21.15 413.1 ;
        RECT  -22.35 414.3 -21.15 415.5 ;
        RECT  -22.35 411.9 -21.15 413.1 ;
        RECT  -31.65 412.65 -30.75 413.55 ;
        RECT  -3.45 412.65 -2.55 413.55 ;
        RECT  -31.65 413.1 -30.75 414.9 ;
        RECT  -31.2 412.65 -3.0 413.55 ;
        RECT  -3.45 413.1 -2.55 414.9 ;
        RECT  -25.2 429.9 -24.3 434.1 ;
        RECT  -17.55 414.9 -16.65 434.1 ;
        RECT  -31.65 414.9 -30.75 434.1 ;
        RECT  -3.45 414.9 -2.55 434.1 ;
        RECT  -9.9 433.2 -9.0 434.1 ;
        RECT  -10.2 432.9 -9.0 434.1 ;
        RECT  -16.65 426.3 -14.25 427.5 ;
        RECT  -5.25 426.3 -3.45 427.5 ;
        RECT  -4.35 431.1 -3.45 432.3 ;
        RECT  -16.65 431.1 -15.45 432.3 ;
        RECT  -14.4 428.7 -5.55 429.9 ;
        RECT  -9.9 432.0 -9.0 434.1 ;
        RECT  -9.9 427.8 -9.0 428.7 ;
        RECT  -17.55 424.5 -16.65 434.1 ;
        RECT  -3.45 424.5 -2.55 434.1 ;
        RECT  -10.35 431.1 -9.15 432.3 ;
        RECT  -10.35 428.7 -9.15 429.9 ;
        RECT  -9.15 431.1 -7.95 432.3 ;
        RECT  -9.15 428.7 -7.95 429.9 ;
        RECT  -9.45 431.1 -8.25 432.3 ;
        RECT  -9.45 428.7 -8.25 429.9 ;
        RECT  -9.45 431.1 -8.25 432.3 ;
        RECT  -9.45 428.7 -8.25 429.9 ;
        RECT  -14.25 426.3 -13.05 427.5 ;
        RECT  -4.35 426.3 -3.15 427.5 ;
        RECT  -8.85 430.8 -7.65 432.0 ;
        RECT  -10.2 423.3 -9.0 424.5 ;
        RECT  -16.65 416.7 -14.25 417.9 ;
        RECT  -5.25 416.7 -3.45 417.9 ;
        RECT  -4.35 421.5 -3.45 422.7 ;
        RECT  -16.65 421.5 -15.45 422.7 ;
        RECT  -14.4 419.1 -5.55 420.3 ;
        RECT  -9.9 422.4 -9.0 424.5 ;
        RECT  -9.9 418.2 -9.0 419.1 ;
        RECT  -17.55 414.9 -16.65 424.5 ;
        RECT  -3.45 414.9 -2.55 424.5 ;
        RECT  -10.35 421.5 -9.15 422.7 ;
        RECT  -10.35 419.1 -9.15 420.3 ;
        RECT  -9.15 421.5 -7.95 422.7 ;
        RECT  -9.15 419.1 -7.95 420.3 ;
        RECT  -9.45 421.5 -8.25 422.7 ;
        RECT  -9.45 419.1 -8.25 420.3 ;
        RECT  -9.45 421.5 -8.25 422.7 ;
        RECT  -9.45 419.1 -8.25 420.3 ;
        RECT  -14.25 416.7 -13.05 417.9 ;
        RECT  -4.35 416.7 -3.15 417.9 ;
        RECT  -8.85 421.2 -7.65 422.4 ;
        RECT  -25.2 414.9 -24.0 416.1 ;
        RECT  -19.95 421.5 -17.55 422.7 ;
        RECT  -30.75 421.5 -28.95 422.7 ;
        RECT  -30.75 416.7 -29.85 417.9 ;
        RECT  -18.75 416.7 -17.55 417.9 ;
        RECT  -28.65 419.1 -19.8 420.3 ;
        RECT  -25.2 414.9 -24.3 417.0 ;
        RECT  -25.2 420.3 -24.3 421.2 ;
        RECT  -17.55 414.9 -16.65 424.5 ;
        RECT  -31.65 414.9 -30.75 424.5 ;
        RECT  -25.05 416.7 -23.85 417.9 ;
        RECT  -25.05 419.1 -23.85 420.3 ;
        RECT  -26.25 416.7 -25.05 417.9 ;
        RECT  -26.25 419.1 -25.05 420.3 ;
        RECT  -25.95 416.7 -24.75 417.9 ;
        RECT  -25.95 419.1 -24.75 420.3 ;
        RECT  -25.95 416.7 -24.75 417.9 ;
        RECT  -25.95 419.1 -24.75 420.3 ;
        RECT  -21.15 421.5 -19.95 422.7 ;
        RECT  -31.05 421.5 -29.85 422.7 ;
        RECT  -26.55 417.0 -25.35 418.2 ;
        RECT  -25.2 424.5 -24.0 425.7 ;
        RECT  -19.95 431.1 -17.55 432.3 ;
        RECT  -30.75 431.1 -28.95 432.3 ;
        RECT  -30.75 426.3 -29.85 427.5 ;
        RECT  -18.75 426.3 -17.55 427.5 ;
        RECT  -28.65 428.7 -19.8 429.9 ;
        RECT  -25.2 424.5 -24.3 426.6 ;
        RECT  -25.2 429.9 -24.3 430.8 ;
        RECT  -17.55 424.5 -16.65 434.1 ;
        RECT  -31.65 424.5 -30.75 434.1 ;
        RECT  -25.05 426.3 -23.85 427.5 ;
        RECT  -25.05 428.7 -23.85 429.9 ;
        RECT  -26.25 426.3 -25.05 427.5 ;
        RECT  -26.25 428.7 -25.05 429.9 ;
        RECT  -25.95 426.3 -24.75 427.5 ;
        RECT  -25.95 428.7 -24.75 429.9 ;
        RECT  -25.95 426.3 -24.75 427.5 ;
        RECT  -25.95 428.7 -24.75 429.9 ;
        RECT  -21.15 431.1 -19.95 432.3 ;
        RECT  -31.05 431.1 -29.85 432.3 ;
        RECT  -26.55 426.6 -25.35 427.8 ;
        RECT  -10.2 427.5 -9.0 428.7 ;
        RECT  -10.2 417.9 -9.0 419.1 ;
        RECT  -25.2 420.3 -24.0 421.5 ;
        RECT  -47.4 433.5 -36.6 434.7 ;
        RECT  -38.4 431.4 -37.2 433.5 ;
        RECT  -41.4 431.4 -40.2 432.6 ;
        RECT  -44.4 431.4 -43.2 432.6 ;
        RECT  -47.4 431.4 -46.2 433.5 ;
        RECT  -41.1 430.5 -39.9 431.4 ;
        RECT  -42.3 429.3 -37.2 430.5 ;
        RECT  -38.4 424.2 -37.2 429.3 ;
        RECT  -41.1 426.0 -39.9 429.3 ;
        RECT  -44.7 427.8 -43.5 431.4 ;
        RECT  -44.7 426.6 -42.9 427.8 ;
        RECT  -44.7 426.0 -43.5 426.6 ;
        RECT  -40.8 424.8 -39.6 426.0 ;
        RECT  -45.0 424.8 -43.8 426.0 ;
        RECT  -47.4 424.8 -46.2 430.5 ;
        RECT  -42.9 423.3 -41.7 423.6 ;
        RECT  -47.4 422.1 -36.6 423.3 ;
        RECT  -40.8 420.0 -38.1 421.2 ;
        RECT  -45.0 420.0 -42.3 421.2 ;
        RECT  -47.4 422.1 -36.6 423.3 ;
        RECT  -47.4 433.5 -36.6 434.7 ;
        RECT  -47.4 416.7 -36.0 417.9 ;
        RECT  -47.4 393.9 -36.0 395.1 ;
        RECT  -47.4 405.6 -36.0 406.5 ;
        RECT  -45.0 418.8 -42.3 420.0 ;
        RECT  -40.8 418.8 -38.1 420.0 ;
        RECT  -47.4 416.7 -36.0 417.9 ;
        RECT  -42.9 416.4 -41.7 416.7 ;
        RECT  -47.4 409.5 -46.2 415.2 ;
        RECT  -45.0 414.0 -43.8 415.2 ;
        RECT  -40.8 414.0 -39.6 415.2 ;
        RECT  -44.7 413.4 -43.5 414.0 ;
        RECT  -44.7 412.2 -42.9 413.4 ;
        RECT  -44.7 408.6 -43.5 412.2 ;
        RECT  -41.1 410.7 -39.9 414.0 ;
        RECT  -42.3 409.5 -39.9 410.7 ;
        RECT  -38.4 409.5 -37.2 415.2 ;
        RECT  -41.1 408.6 -39.9 409.5 ;
        RECT  -47.4 406.5 -46.2 408.6 ;
        RECT  -44.4 407.4 -43.2 408.6 ;
        RECT  -41.4 407.4 -40.2 408.6 ;
        RECT  -38.4 406.5 -37.2 408.6 ;
        RECT  -47.4 405.3 -36.0 406.5 ;
        RECT  -47.4 416.7 -36.0 417.9 ;
        RECT  -47.4 405.3 -36.0 406.5 ;
        RECT  -45.0 391.8 -42.3 393.0 ;
        RECT  -40.8 391.8 -38.1 393.0 ;
        RECT  -47.4 393.9 -36.0 395.1 ;
        RECT  -42.9 395.1 -41.7 395.4 ;
        RECT  -47.4 396.6 -46.2 402.3 ;
        RECT  -45.0 396.6 -43.8 397.8 ;
        RECT  -40.8 396.6 -39.6 397.8 ;
        RECT  -44.7 397.8 -43.5 398.4 ;
        RECT  -44.7 398.4 -42.9 399.6 ;
        RECT  -44.7 399.6 -43.5 403.2 ;
        RECT  -41.1 397.8 -39.9 401.1 ;
        RECT  -42.3 401.1 -39.9 402.3 ;
        RECT  -38.4 396.6 -37.2 402.3 ;
        RECT  -41.1 402.3 -39.9 403.2 ;
        RECT  -47.4 403.2 -46.2 405.3 ;
        RECT  -44.4 403.2 -43.2 404.4 ;
        RECT  -41.4 403.2 -40.2 404.4 ;
        RECT  -38.4 403.2 -37.2 405.3 ;
        RECT  -47.4 405.3 -36.0 406.5 ;
        RECT  -47.4 393.9 -36.0 395.1 ;
        RECT  -47.4 405.3 -36.0 406.5 ;
        RECT  -31.95 420.9 -30.75 422.1 ;
        RECT  -31.95 443.7 -30.75 444.9 ;
        RECT  -31.95 432.9 -30.75 434.1 ;
        RECT  -31.95 393.3 -30.75 394.5 ;
        RECT  -31.8 449.1 -30.6 450.3 ;
        RECT  -47.4 449.1 -46.2 450.3 ;
        RECT  -25.2 419.1 -24.0 420.3 ;
        RECT  -34.05 406.2 -32.85 407.4 ;
        RECT  -34.05 398.7 -32.85 399.9 ;
        RECT  -40.8 398.7 -39.6 399.9 ;
        RECT  -10.05 305.55 -8.85 306.75 ;
        RECT  -10.2 257.4 -9.0 258.6 ;
        RECT  -20.4 204.45 -19.2 205.65 ;
        RECT  -27.45 305.55 -26.25 306.75 ;
        RECT  -25.35 310.95 -24.15 312.15 ;
        RECT  -23.4 349.5 -22.2 350.7 ;
        RECT  -26.1 349.5 -24.9 350.7 ;
        RECT  -12.9 324.45 -11.7 325.65 ;
        RECT  -10.8 321.75 -9.6 322.95 ;
        RECT  -8.7 313.65 -7.5 314.85 ;
        RECT  -41.1 324.45 -39.9 325.65 ;
        RECT  -39.0 316.35 -37.8 317.55 ;
        RECT  -36.9 313.65 -35.7 314.85 ;
        RECT  -27.3 346.8 -26.1 348.0 ;
        RECT  -25.2 361.5 -24.0 362.7 ;
        RECT  -38.1 384.0 -36.9 385.2 ;
        RECT  -25.2 364.2 -24.0 365.4 ;
        RECT  -3.6 308.25 -2.4 309.45 ;
        RECT  -17.7 319.05 -16.5 320.25 ;
        RECT  -31.8 308.25 -30.6 309.45 ;
        RECT  -45.9 319.05 -44.7 320.25 ;
        RECT  1.65 319.05 2.85 320.25 ;
        LAYER  via1 ;
        RECT  126.3 199.5 126.9 200.1 ;
        RECT  122.1 199.5 122.7 200.1 ;
        RECT  130.2 208.8 130.8 209.4 ;
        RECT  121.2 208.8 121.8 209.4 ;
        RECT  126.3 226.5 126.9 227.1 ;
        RECT  122.1 226.5 122.7 227.1 ;
        RECT  130.2 217.2 130.8 217.8 ;
        RECT  121.2 217.2 121.8 217.8 ;
        RECT  126.3 227.7 126.9 228.3 ;
        RECT  122.1 227.7 122.7 228.3 ;
        RECT  130.2 237.0 130.8 237.6 ;
        RECT  121.2 237.0 121.8 237.6 ;
        RECT  126.3 254.7 126.9 255.3 ;
        RECT  122.1 254.7 122.7 255.3 ;
        RECT  130.2 245.4 130.8 246.0 ;
        RECT  121.2 245.4 121.8 246.0 ;
        RECT  126.3 255.9 126.9 256.5 ;
        RECT  122.1 255.9 122.7 256.5 ;
        RECT  130.2 265.2 130.8 265.8 ;
        RECT  121.2 265.2 121.8 265.8 ;
        RECT  126.3 282.9 126.9 283.5 ;
        RECT  122.1 282.9 122.7 283.5 ;
        RECT  130.2 273.6 130.8 274.2 ;
        RECT  121.2 273.6 121.8 274.2 ;
        RECT  126.3 284.1 126.9 284.7 ;
        RECT  122.1 284.1 122.7 284.7 ;
        RECT  130.2 293.4 130.8 294.0 ;
        RECT  121.2 293.4 121.8 294.0 ;
        RECT  126.3 311.1 126.9 311.7 ;
        RECT  122.1 311.1 122.7 311.7 ;
        RECT  130.2 301.8 130.8 302.4 ;
        RECT  121.2 301.8 121.8 302.4 ;
        RECT  126.3 312.3 126.9 312.9 ;
        RECT  122.1 312.3 122.7 312.9 ;
        RECT  130.2 321.6 130.8 322.2 ;
        RECT  121.2 321.6 121.8 322.2 ;
        RECT  126.3 339.3 126.9 339.9 ;
        RECT  122.1 339.3 122.7 339.9 ;
        RECT  130.2 330.0 130.8 330.6 ;
        RECT  121.2 330.0 121.8 330.6 ;
        RECT  126.3 340.5 126.9 341.1 ;
        RECT  122.1 340.5 122.7 341.1 ;
        RECT  130.2 349.8 130.8 350.4 ;
        RECT  121.2 349.8 121.8 350.4 ;
        RECT  126.3 367.5 126.9 368.1 ;
        RECT  122.1 367.5 122.7 368.1 ;
        RECT  130.2 358.2 130.8 358.8 ;
        RECT  121.2 358.2 121.8 358.8 ;
        RECT  126.3 368.7 126.9 369.3 ;
        RECT  122.1 368.7 122.7 369.3 ;
        RECT  130.2 378.0 130.8 378.6 ;
        RECT  121.2 378.0 121.8 378.6 ;
        RECT  126.3 395.7 126.9 396.3 ;
        RECT  122.1 395.7 122.7 396.3 ;
        RECT  130.2 386.4 130.8 387.0 ;
        RECT  121.2 386.4 121.8 387.0 ;
        RECT  126.3 396.9 126.9 397.5 ;
        RECT  122.1 396.9 122.7 397.5 ;
        RECT  130.2 406.2 130.8 406.8 ;
        RECT  121.2 406.2 121.8 406.8 ;
        RECT  126.3 423.9 126.9 424.5 ;
        RECT  122.1 423.9 122.7 424.5 ;
        RECT  130.2 414.6 130.8 415.2 ;
        RECT  121.2 414.6 121.8 415.2 ;
        RECT  136.5 199.5 137.1 200.1 ;
        RECT  132.3 199.5 132.9 200.1 ;
        RECT  140.4 208.8 141.0 209.4 ;
        RECT  131.4 208.8 132.0 209.4 ;
        RECT  136.5 226.5 137.1 227.1 ;
        RECT  132.3 226.5 132.9 227.1 ;
        RECT  140.4 217.2 141.0 217.8 ;
        RECT  131.4 217.2 132.0 217.8 ;
        RECT  136.5 227.7 137.1 228.3 ;
        RECT  132.3 227.7 132.9 228.3 ;
        RECT  140.4 237.0 141.0 237.6 ;
        RECT  131.4 237.0 132.0 237.6 ;
        RECT  136.5 254.7 137.1 255.3 ;
        RECT  132.3 254.7 132.9 255.3 ;
        RECT  140.4 245.4 141.0 246.0 ;
        RECT  131.4 245.4 132.0 246.0 ;
        RECT  136.5 255.9 137.1 256.5 ;
        RECT  132.3 255.9 132.9 256.5 ;
        RECT  140.4 265.2 141.0 265.8 ;
        RECT  131.4 265.2 132.0 265.8 ;
        RECT  136.5 282.9 137.1 283.5 ;
        RECT  132.3 282.9 132.9 283.5 ;
        RECT  140.4 273.6 141.0 274.2 ;
        RECT  131.4 273.6 132.0 274.2 ;
        RECT  136.5 284.1 137.1 284.7 ;
        RECT  132.3 284.1 132.9 284.7 ;
        RECT  140.4 293.4 141.0 294.0 ;
        RECT  131.4 293.4 132.0 294.0 ;
        RECT  136.5 311.1 137.1 311.7 ;
        RECT  132.3 311.1 132.9 311.7 ;
        RECT  140.4 301.8 141.0 302.4 ;
        RECT  131.4 301.8 132.0 302.4 ;
        RECT  136.5 312.3 137.1 312.9 ;
        RECT  132.3 312.3 132.9 312.9 ;
        RECT  140.4 321.6 141.0 322.2 ;
        RECT  131.4 321.6 132.0 322.2 ;
        RECT  136.5 339.3 137.1 339.9 ;
        RECT  132.3 339.3 132.9 339.9 ;
        RECT  140.4 330.0 141.0 330.6 ;
        RECT  131.4 330.0 132.0 330.6 ;
        RECT  136.5 340.5 137.1 341.1 ;
        RECT  132.3 340.5 132.9 341.1 ;
        RECT  140.4 349.8 141.0 350.4 ;
        RECT  131.4 349.8 132.0 350.4 ;
        RECT  136.5 367.5 137.1 368.1 ;
        RECT  132.3 367.5 132.9 368.1 ;
        RECT  140.4 358.2 141.0 358.8 ;
        RECT  131.4 358.2 132.0 358.8 ;
        RECT  136.5 368.7 137.1 369.3 ;
        RECT  132.3 368.7 132.9 369.3 ;
        RECT  140.4 378.0 141.0 378.6 ;
        RECT  131.4 378.0 132.0 378.6 ;
        RECT  136.5 395.7 137.1 396.3 ;
        RECT  132.3 395.7 132.9 396.3 ;
        RECT  140.4 386.4 141.0 387.0 ;
        RECT  131.4 386.4 132.0 387.0 ;
        RECT  136.5 396.9 137.1 397.5 ;
        RECT  132.3 396.9 132.9 397.5 ;
        RECT  140.4 406.2 141.0 406.8 ;
        RECT  131.4 406.2 132.0 406.8 ;
        RECT  136.5 423.9 137.1 424.5 ;
        RECT  132.3 423.9 132.9 424.5 ;
        RECT  140.4 414.6 141.0 415.2 ;
        RECT  131.4 414.6 132.0 415.2 ;
        RECT  123.6 436.2 124.2 436.8 ;
        RECT  128.4 436.2 129.0 436.8 ;
        RECT  123.6 427.8 124.2 428.4 ;
        RECT  126.0 427.8 126.6 428.4 ;
        RECT  133.8 436.2 134.4 436.8 ;
        RECT  138.6 436.2 139.2 436.8 ;
        RECT  133.8 427.8 134.4 428.4 ;
        RECT  136.2 427.8 136.8 428.4 ;
        RECT  130.2 193.2 130.8 193.8 ;
        RECT  124.5 163.8 125.1 164.4 ;
        RECT  127.2 163.8 127.8 164.4 ;
        RECT  121.5 153.9 122.1 154.5 ;
        RECT  140.4 193.2 141.0 193.8 ;
        RECT  134.7 163.8 135.3 164.4 ;
        RECT  137.4 163.8 138.0 164.4 ;
        RECT  131.7 153.9 132.3 154.5 ;
        RECT  122.1 147.3 122.7 147.9 ;
        RECT  126.6 146.7 127.2 147.3 ;
        RECT  123.9 137.1 124.5 137.7 ;
        RECT  123.0 125.4 123.6 126.0 ;
        RECT  129.6 114.6 130.2 115.2 ;
        RECT  126.3 109.2 126.9 109.8 ;
        RECT  123.0 99.3 123.6 99.9 ;
        RECT  130.2 95.1 130.8 95.7 ;
        RECT  124.2 93.0 124.8 93.6 ;
        RECT  132.3 147.3 132.9 147.9 ;
        RECT  136.8 146.7 137.4 147.3 ;
        RECT  134.1 137.1 134.7 137.7 ;
        RECT  133.2 125.4 133.8 126.0 ;
        RECT  139.8 114.6 140.4 115.2 ;
        RECT  136.5 109.2 137.1 109.8 ;
        RECT  133.2 99.3 133.8 99.9 ;
        RECT  140.4 95.1 141.0 95.7 ;
        RECT  134.4 93.0 135.0 93.6 ;
        RECT  124.2 84.6 124.8 85.2 ;
        RECT  126.6 80.1 127.2 80.7 ;
        RECT  125.7 76.8 126.3 77.4 ;
        RECT  130.2 76.2 130.8 76.8 ;
        RECT  125.7 74.7 126.3 75.3 ;
        RECT  122.4 73.8 123.0 74.4 ;
        RECT  126.6 70.2 127.2 70.8 ;
        RECT  126.6 67.8 127.2 68.4 ;
        RECT  124.2 64.8 124.8 65.4 ;
        RECT  125.1 61.5 125.7 62.1 ;
        RECT  122.4 60.3 123.0 60.9 ;
        RECT  126.6 54.6 127.2 55.2 ;
        RECT  125.7 51.3 126.3 51.9 ;
        RECT  130.2 50.7 130.8 51.3 ;
        RECT  125.7 48.3 126.3 48.9 ;
        RECT  122.4 47.4 123.0 48.0 ;
        RECT  126.6 43.8 127.2 44.4 ;
        RECT  126.6 41.4 127.2 42.0 ;
        RECT  124.2 38.4 124.8 39.0 ;
        RECT  136.2 84.6 136.8 85.2 ;
        RECT  133.8 80.1 134.4 80.7 ;
        RECT  134.7 76.8 135.3 77.4 ;
        RECT  130.2 76.2 130.8 76.8 ;
        RECT  134.7 74.7 135.3 75.3 ;
        RECT  138.0 73.8 138.6 74.4 ;
        RECT  133.8 70.2 134.4 70.8 ;
        RECT  133.8 67.8 134.4 68.4 ;
        RECT  136.2 64.8 136.8 65.4 ;
        RECT  135.3 61.5 135.9 62.1 ;
        RECT  138.0 60.3 138.6 60.9 ;
        RECT  133.8 54.6 134.4 55.2 ;
        RECT  134.7 51.3 135.3 51.9 ;
        RECT  130.2 50.7 130.8 51.3 ;
        RECT  134.7 48.3 135.3 48.9 ;
        RECT  138.0 47.4 138.6 48.0 ;
        RECT  133.8 43.8 134.4 44.4 ;
        RECT  133.8 41.4 134.4 42.0 ;
        RECT  136.2 38.4 136.8 39.0 ;
        RECT  123.3 44.1 123.9 44.7 ;
        RECT  128.1 40.5 128.7 41.1 ;
        RECT  130.2 36.0 130.8 36.6 ;
        RECT  133.5 44.1 134.1 44.7 ;
        RECT  138.3 40.5 138.9 41.1 ;
        RECT  140.4 36.0 141.0 36.6 ;
        RECT  56.1 96.75 56.7 97.35 ;
        RECT  74.7 91.35 75.3 91.95 ;
        RECT  53.1 110.85 53.7 111.45 ;
        RECT  71.7 106.65 72.3 107.25 ;
        RECT  74.7 115.35 75.3 115.95 ;
        RECT  50.1 115.35 50.7 115.95 ;
        RECT  71.7 129.45 72.3 130.05 ;
        RECT  47.1 129.45 47.7 130.05 ;
        RECT  56.1 93.45 56.7 94.05 ;
        RECT  53.1 90.75 53.7 91.35 ;
        RECT  50.1 104.55 50.7 105.15 ;
        RECT  53.1 107.25 53.7 107.85 ;
        RECT  56.1 121.65 56.7 122.25 ;
        RECT  47.1 118.95 47.7 119.55 ;
        RECT  50.1 132.75 50.7 133.35 ;
        RECT  47.1 135.45 47.7 136.05 ;
        RECT  56.1 153.15 56.7 153.75 ;
        RECT  74.7 147.75 75.3 148.35 ;
        RECT  53.1 167.25 53.7 167.85 ;
        RECT  71.7 163.05 72.3 163.65 ;
        RECT  74.7 171.75 75.3 172.35 ;
        RECT  50.1 171.75 50.7 172.35 ;
        RECT  71.7 185.85 72.3 186.45 ;
        RECT  47.1 185.85 47.7 186.45 ;
        RECT  56.1 149.85 56.7 150.45 ;
        RECT  53.1 147.15 53.7 147.75 ;
        RECT  50.1 160.95 50.7 161.55 ;
        RECT  53.1 163.65 53.7 164.25 ;
        RECT  56.1 178.05 56.7 178.65 ;
        RECT  47.1 175.35 47.7 175.95 ;
        RECT  50.1 189.15 50.7 189.75 ;
        RECT  47.1 191.85 47.7 192.45 ;
        RECT  6.6 92.7 7.2 93.3 ;
        RECT  8.7 108.0 9.3 108.6 ;
        RECT  10.8 120.9 11.4 121.5 ;
        RECT  12.9 136.2 13.5 136.8 ;
        RECT  15.0 149.1 15.6 149.7 ;
        RECT  17.1 164.4 17.7 165.0 ;
        RECT  19.2 177.3 19.8 177.9 ;
        RECT  21.3 192.6 21.9 193.2 ;
        RECT  6.6 207.6 7.2 208.2 ;
        RECT  15.0 204.9 15.6 205.5 ;
        RECT  6.6 218.7 7.2 219.3 ;
        RECT  17.1 221.4 17.7 222.0 ;
        RECT  6.6 235.8 7.2 236.4 ;
        RECT  19.2 233.1 19.8 233.7 ;
        RECT  6.6 246.9 7.2 247.5 ;
        RECT  21.3 249.6 21.9 250.2 ;
        RECT  8.7 264.0 9.3 264.6 ;
        RECT  15.0 261.3 15.6 261.9 ;
        RECT  8.7 275.1 9.3 275.7 ;
        RECT  17.1 277.8 17.7 278.4 ;
        RECT  8.7 292.2 9.3 292.8 ;
        RECT  19.2 289.5 19.8 290.1 ;
        RECT  8.7 303.3 9.3 303.9 ;
        RECT  21.3 306.0 21.9 306.6 ;
        RECT  10.8 320.4 11.4 321.0 ;
        RECT  15.0 317.7 15.6 318.3 ;
        RECT  10.8 331.5 11.4 332.1 ;
        RECT  17.1 334.2 17.7 334.8 ;
        RECT  10.8 348.6 11.4 349.2 ;
        RECT  19.2 345.9 19.8 346.5 ;
        RECT  10.8 359.7 11.4 360.3 ;
        RECT  21.3 362.4 21.9 363.0 ;
        RECT  12.9 376.8 13.5 377.4 ;
        RECT  15.0 374.1 15.6 374.7 ;
        RECT  12.9 387.9 13.5 388.5 ;
        RECT  17.1 390.6 17.7 391.2 ;
        RECT  12.9 405.0 13.5 405.6 ;
        RECT  19.2 402.3 19.8 402.9 ;
        RECT  12.9 416.1 13.5 416.7 ;
        RECT  21.3 418.8 21.9 419.4 ;
        RECT  47.55 205.35 48.15 205.95 ;
        RECT  49.5 207.45 50.1 208.05 ;
        RECT  60.9 207.45 61.5 208.05 ;
        RECT  47.55 220.65 48.15 221.25 ;
        RECT  49.5 218.55 50.1 219.15 ;
        RECT  60.9 218.55 61.5 219.15 ;
        RECT  47.55 233.55 48.15 234.15 ;
        RECT  49.5 235.65 50.1 236.25 ;
        RECT  60.9 235.65 61.5 236.25 ;
        RECT  47.55 248.85 48.15 249.45 ;
        RECT  49.5 246.75 50.1 247.35 ;
        RECT  60.9 246.75 61.5 247.35 ;
        RECT  47.55 261.75 48.15 262.35 ;
        RECT  49.5 263.85 50.1 264.45 ;
        RECT  60.9 263.85 61.5 264.45 ;
        RECT  47.55 277.05 48.15 277.65 ;
        RECT  49.5 274.95 50.1 275.55 ;
        RECT  60.9 274.95 61.5 275.55 ;
        RECT  47.55 289.95 48.15 290.55 ;
        RECT  49.5 292.05 50.1 292.65 ;
        RECT  60.9 292.05 61.5 292.65 ;
        RECT  47.55 305.25 48.15 305.85 ;
        RECT  49.5 303.15 50.1 303.75 ;
        RECT  60.9 303.15 61.5 303.75 ;
        RECT  47.55 318.15 48.15 318.75 ;
        RECT  49.5 320.25 50.1 320.85 ;
        RECT  60.9 320.25 61.5 320.85 ;
        RECT  47.55 333.45 48.15 334.05 ;
        RECT  49.5 331.35 50.1 331.95 ;
        RECT  60.9 331.35 61.5 331.95 ;
        RECT  47.55 346.35 48.15 346.95 ;
        RECT  49.5 348.45 50.1 349.05 ;
        RECT  60.9 348.45 61.5 349.05 ;
        RECT  47.55 361.65 48.15 362.25 ;
        RECT  49.5 359.55 50.1 360.15 ;
        RECT  60.9 359.55 61.5 360.15 ;
        RECT  47.55 374.55 48.15 375.15 ;
        RECT  49.5 376.65 50.1 377.25 ;
        RECT  60.9 376.65 61.5 377.25 ;
        RECT  47.55 389.85 48.15 390.45 ;
        RECT  49.5 387.75 50.1 388.35 ;
        RECT  60.9 387.75 61.5 388.35 ;
        RECT  47.55 402.75 48.15 403.35 ;
        RECT  49.5 404.85 50.1 405.45 ;
        RECT  60.9 404.85 61.5 405.45 ;
        RECT  47.55 418.05 48.15 418.65 ;
        RECT  49.5 415.95 50.1 416.55 ;
        RECT  60.9 415.95 61.5 416.55 ;
        RECT  60.9 76.5 61.5 77.1 ;
        RECT  56.4 74.1 57.0 74.7 ;
        RECT  53.1 75.0 53.7 75.6 ;
        RECT  52.5 70.5 53.1 71.1 ;
        RECT  51.0 75.0 51.6 75.6 ;
        RECT  50.1 78.3 50.7 78.9 ;
        RECT  46.5 74.1 47.1 74.7 ;
        RECT  44.1 74.1 44.7 74.7 ;
        RECT  41.1 76.5 41.7 77.1 ;
        RECT  37.8 75.6 38.4 76.2 ;
        RECT  36.6 78.3 37.2 78.9 ;
        RECT  30.9 74.1 31.5 74.7 ;
        RECT  27.6 75.0 28.2 75.6 ;
        RECT  27.0 70.5 27.6 71.1 ;
        RECT  24.6 75.0 25.2 75.6 ;
        RECT  23.7 78.3 24.3 78.9 ;
        RECT  20.1 74.1 20.7 74.7 ;
        RECT  17.7 74.1 18.3 74.7 ;
        RECT  14.7 76.5 15.3 77.1 ;
        RECT  60.9 64.5 61.5 65.1 ;
        RECT  56.4 66.9 57.0 67.5 ;
        RECT  53.1 66.0 53.7 66.6 ;
        RECT  52.5 70.5 53.1 71.1 ;
        RECT  51.0 66.0 51.6 66.6 ;
        RECT  50.1 62.7 50.7 63.3 ;
        RECT  46.5 66.9 47.1 67.5 ;
        RECT  44.1 66.9 44.7 67.5 ;
        RECT  41.1 64.5 41.7 65.1 ;
        RECT  37.8 65.4 38.4 66.0 ;
        RECT  36.6 62.7 37.2 63.3 ;
        RECT  30.9 66.9 31.5 67.5 ;
        RECT  27.6 66.0 28.2 66.6 ;
        RECT  27.0 70.5 27.6 71.1 ;
        RECT  24.6 66.0 25.2 66.6 ;
        RECT  23.7 62.7 24.3 63.3 ;
        RECT  20.1 66.9 20.7 67.5 ;
        RECT  17.7 66.9 18.3 67.5 ;
        RECT  14.7 64.5 15.3 65.1 ;
        RECT  60.9 56.1 61.5 56.7 ;
        RECT  56.4 53.7 57.0 54.3 ;
        RECT  53.1 54.6 53.7 55.2 ;
        RECT  52.5 50.1 53.1 50.7 ;
        RECT  51.0 54.6 51.6 55.2 ;
        RECT  50.1 57.9 50.7 58.5 ;
        RECT  46.5 53.7 47.1 54.3 ;
        RECT  44.1 53.7 44.7 54.3 ;
        RECT  41.1 56.1 41.7 56.7 ;
        RECT  37.8 55.2 38.4 55.8 ;
        RECT  36.6 57.9 37.2 58.5 ;
        RECT  30.9 53.7 31.5 54.3 ;
        RECT  27.6 54.6 28.2 55.2 ;
        RECT  27.0 50.1 27.6 50.7 ;
        RECT  24.6 54.6 25.2 55.2 ;
        RECT  23.7 57.9 24.3 58.5 ;
        RECT  20.1 53.7 20.7 54.3 ;
        RECT  17.7 53.7 18.3 54.3 ;
        RECT  14.7 56.1 15.3 56.7 ;
        RECT  60.9 44.1 61.5 44.7 ;
        RECT  56.4 46.5 57.0 47.1 ;
        RECT  53.1 45.6 53.7 46.2 ;
        RECT  52.5 50.1 53.1 50.7 ;
        RECT  51.0 45.6 51.6 46.2 ;
        RECT  50.1 42.3 50.7 42.9 ;
        RECT  46.5 46.5 47.1 47.1 ;
        RECT  44.1 46.5 44.7 47.1 ;
        RECT  41.1 44.1 41.7 44.7 ;
        RECT  37.8 45.0 38.4 45.6 ;
        RECT  36.6 42.3 37.2 42.9 ;
        RECT  30.9 46.5 31.5 47.1 ;
        RECT  27.6 45.6 28.2 46.2 ;
        RECT  27.0 50.1 27.6 50.7 ;
        RECT  24.6 45.6 25.2 46.2 ;
        RECT  23.7 42.3 24.3 42.9 ;
        RECT  20.1 46.5 20.7 47.1 ;
        RECT  17.7 46.5 18.3 47.1 ;
        RECT  14.7 44.1 15.3 44.7 ;
        RECT  93.15 198.9 93.75 199.5 ;
        RECT  93.15 227.1 93.75 227.7 ;
        RECT  93.15 255.3 93.75 255.9 ;
        RECT  93.15 283.5 93.75 284.1 ;
        RECT  93.15 311.7 93.75 312.3 ;
        RECT  93.15 339.9 93.75 340.5 ;
        RECT  93.15 368.1 93.75 368.7 ;
        RECT  93.15 396.3 93.75 396.9 ;
        RECT  93.15 424.5 93.75 425.1 ;
        RECT  74.4 88.95 75.0 89.55 ;
        RECT  79.35 88.95 79.95 89.55 ;
        RECT  71.4 103.05 72.0 103.65 ;
        RECT  82.05 103.05 82.65 103.65 ;
        RECT  74.4 145.35 75.0 145.95 ;
        RECT  84.75 145.35 85.35 145.95 ;
        RECT  71.4 159.45 72.0 160.05 ;
        RECT  87.45 159.45 88.05 160.05 ;
        RECT  76.5 86.1 77.1 86.7 ;
        RECT  76.5 114.3 77.1 114.9 ;
        RECT  76.5 142.5 77.1 143.1 ;
        RECT  76.5 170.7 77.1 171.3 ;
        RECT  66.6 75.6 67.2 76.2 ;
        RECT  79.35 75.75 79.95 76.35 ;
        RECT  66.6 65.4 67.2 66.0 ;
        RECT  82.05 65.55 82.65 66.15 ;
        RECT  66.6 55.2 67.2 55.8 ;
        RECT  84.75 55.35 85.35 55.95 ;
        RECT  66.6 45.0 67.2 45.6 ;
        RECT  87.45 45.15 88.05 45.75 ;
        RECT  66.6 70.5 67.2 71.1 ;
        RECT  93.15 70.65 93.75 71.25 ;
        RECT  66.6 50.1 67.2 50.7 ;
        RECT  93.15 50.25 93.75 50.85 ;
        RECT  108.3 32.55 108.9 33.15 ;
        RECT  102.9 28.05 103.5 28.65 ;
        RECT  105.6 25.65 106.2 26.25 ;
        RECT  108.3 431.55 108.9 432.15 ;
        RECT  111.0 97.05 111.6 97.65 ;
        RECT  113.7 195.15 114.3 195.75 ;
        RECT  100.35 82.95 100.95 83.55 ;
        RECT  47.55 426.6 48.15 427.2 ;
        RECT  100.35 426.75 100.95 427.35 ;
        RECT  96.45 23.7 97.05 24.3 ;
        RECT  96.45 193.2 97.05 193.8 ;
        RECT  96.45 95.1 97.05 95.7 ;
        RECT  -49.2 256.8 -48.6 257.4 ;
        RECT  -46.8 252.3 -46.2 252.9 ;
        RECT  -47.7 249.0 -47.1 249.6 ;
        RECT  -43.2 248.4 -42.6 249.0 ;
        RECT  -47.7 246.9 -47.1 247.5 ;
        RECT  -51.0 246.0 -50.4 246.6 ;
        RECT  -46.8 242.4 -46.2 243.0 ;
        RECT  -46.8 240.0 -46.2 240.6 ;
        RECT  -49.2 237.0 -48.6 237.6 ;
        RECT  -48.3 233.7 -47.7 234.3 ;
        RECT  -51.0 232.5 -50.4 233.1 ;
        RECT  -46.8 226.8 -46.2 227.4 ;
        RECT  -47.7 223.5 -47.1 224.1 ;
        RECT  -43.2 222.9 -42.6 223.5 ;
        RECT  -47.7 220.5 -47.1 221.1 ;
        RECT  -51.0 219.6 -50.4 220.2 ;
        RECT  -46.8 216.0 -46.2 216.6 ;
        RECT  -46.8 213.6 -46.2 214.2 ;
        RECT  -49.2 210.6 -48.6 211.2 ;
        RECT  -37.2 256.8 -36.6 257.4 ;
        RECT  -39.6 252.3 -39.0 252.9 ;
        RECT  -38.7 249.0 -38.1 249.6 ;
        RECT  -43.2 248.4 -42.6 249.0 ;
        RECT  -38.7 246.9 -38.1 247.5 ;
        RECT  -35.4 246.0 -34.8 246.6 ;
        RECT  -39.6 242.4 -39.0 243.0 ;
        RECT  -39.6 240.0 -39.0 240.6 ;
        RECT  -37.2 237.0 -36.6 237.6 ;
        RECT  -38.1 233.7 -37.5 234.3 ;
        RECT  -35.4 232.5 -34.8 233.1 ;
        RECT  -39.6 226.8 -39.0 227.4 ;
        RECT  -38.7 223.5 -38.1 224.1 ;
        RECT  -43.2 222.9 -42.6 223.5 ;
        RECT  -38.7 220.5 -38.1 221.1 ;
        RECT  -35.4 219.6 -34.8 220.2 ;
        RECT  -39.6 216.0 -39.0 216.6 ;
        RECT  -39.6 213.6 -39.0 214.2 ;
        RECT  -37.2 210.6 -36.6 211.2 ;
        RECT  -28.8 256.8 -28.2 257.4 ;
        RECT  -26.4 252.3 -25.8 252.9 ;
        RECT  -27.3 249.0 -26.7 249.6 ;
        RECT  -22.8 248.4 -22.2 249.0 ;
        RECT  -27.3 246.9 -26.7 247.5 ;
        RECT  -30.6 246.0 -30.0 246.6 ;
        RECT  -26.4 242.4 -25.8 243.0 ;
        RECT  -26.4 240.0 -25.8 240.6 ;
        RECT  -28.8 237.0 -28.2 237.6 ;
        RECT  -27.9 233.7 -27.3 234.3 ;
        RECT  -30.6 232.5 -30.0 233.1 ;
        RECT  -26.4 226.8 -25.8 227.4 ;
        RECT  -27.3 223.5 -26.7 224.1 ;
        RECT  -22.8 222.9 -22.2 223.5 ;
        RECT  -27.3 220.5 -26.7 221.1 ;
        RECT  -30.6 219.6 -30.0 220.2 ;
        RECT  -26.4 216.0 -25.8 216.6 ;
        RECT  -26.4 213.6 -25.8 214.2 ;
        RECT  -28.8 210.6 -28.2 211.2 ;
        RECT  -15.15 335.7 -14.55 336.3 ;
        RECT  -15.15 340.5 -14.55 341.1 ;
        RECT  -22.2 341.7 -21.6 342.3 ;
        RECT  -28.35 341.7 -27.75 342.3 ;
        RECT  -43.35 345.3 -42.75 345.9 ;
        RECT  -43.35 350.1 -42.75 350.7 ;
        RECT  -51.15 262.5 -50.55 263.1 ;
        RECT  -48.45 262.5 -47.85 263.1 ;
        RECT  -35.55 262.5 -34.95 263.1 ;
        RECT  -30.75 262.5 -30.15 263.1 ;
        RECT  -9.9 433.2 -9.3 433.8 ;
        RECT  -9.9 423.6 -9.3 424.2 ;
        RECT  -24.9 415.2 -24.3 415.8 ;
        RECT  -24.9 424.8 -24.3 425.4 ;
        RECT  -9.9 427.8 -9.3 428.4 ;
        RECT  -9.9 418.2 -9.3 418.8 ;
        RECT  -24.9 420.6 -24.3 421.2 ;
        RECT  -38.1 429.6 -37.5 430.2 ;
        RECT  -47.1 429.6 -46.5 430.2 ;
        RECT  -39.0 420.3 -38.4 420.9 ;
        RECT  -43.2 420.3 -42.6 420.9 ;
        RECT  -43.2 419.1 -42.6 419.7 ;
        RECT  -39.0 419.1 -38.4 419.7 ;
        RECT  -47.1 409.8 -46.5 410.4 ;
        RECT  -38.1 409.8 -37.5 410.4 ;
        RECT  -43.2 392.1 -42.6 392.7 ;
        RECT  -39.0 392.1 -38.4 392.7 ;
        RECT  -47.1 401.4 -46.5 402.0 ;
        RECT  -38.1 401.4 -37.5 402.0 ;
        RECT  -31.65 421.2 -31.05 421.8 ;
        RECT  -31.65 444.0 -31.05 444.6 ;
        RECT  -31.65 433.2 -31.05 433.8 ;
        RECT  -31.65 393.6 -31.05 394.2 ;
        RECT  -31.5 449.4 -30.9 450.0 ;
        RECT  -47.1 449.4 -46.5 450.0 ;
        RECT  -33.75 406.5 -33.15 407.1 ;
        RECT  -33.75 399.0 -33.15 399.6 ;
        RECT  -40.5 399.0 -39.9 399.6 ;
        RECT  -9.75 305.85 -9.15 306.45 ;
        RECT  -9.9 257.7 -9.3 258.3 ;
        RECT  -20.1 204.75 -19.5 205.35 ;
        RECT  -27.15 305.85 -26.55 306.45 ;
        RECT  -25.05 311.25 -24.45 311.85 ;
        RECT  -23.1 349.8 -22.5 350.4 ;
        RECT  -25.8 349.8 -25.2 350.4 ;
        RECT  -12.6 324.75 -12.0 325.35 ;
        RECT  -10.5 322.05 -9.9 322.65 ;
        RECT  -8.4 313.95 -7.8 314.55 ;
        RECT  -40.8 324.75 -40.2 325.35 ;
        RECT  -38.7 316.65 -38.1 317.25 ;
        RECT  -36.6 313.95 -36.0 314.55 ;
        RECT  -27.0 347.1 -26.4 347.7 ;
        RECT  -24.9 361.8 -24.3 362.4 ;
        RECT  -37.8 384.3 -37.2 384.9 ;
        RECT  -24.9 364.5 -24.3 365.1 ;
        RECT  -3.3 308.55 -2.7 309.15 ;
        RECT  -17.4 319.35 -16.8 319.95 ;
        RECT  -31.5 308.55 -30.9 309.15 ;
        RECT  -45.6 319.35 -45.0 319.95 ;
        RECT  1.95 319.35 2.55 319.95 ;
        LAYER  metal2 ;
        RECT  113.55 361.95 114.45 364.65 ;
        RECT  110.85 381.75 111.75 384.45 ;
        RECT  105.45 344.55 106.35 347.25 ;
        RECT  102.75 359.25 103.65 361.95 ;
        RECT  108.15 322.35 109.05 325.05 ;
        RECT  100.05 303.45 100.95 306.15 ;
        RECT  -3.0 319.2 2.25 320.1 ;
        RECT  94.65 306.15 95.55 308.85 ;
        RECT  124.8 0.0 125.7 1.8 ;
        RECT  135.0 0.0 135.9 1.8 ;
        RECT  92.85 0.0 97.35 444.3 ;
        RECT  100.05 0.0 100.95 444.3 ;
        RECT  102.75 0.0 103.65 444.3 ;
        RECT  105.45 0.0 106.35 444.3 ;
        RECT  108.15 0.0 109.05 444.3 ;
        RECT  110.85 0.0 111.75 444.3 ;
        RECT  113.55 0.0 114.45 444.3 ;
        RECT  79.35 34.8 80.25 199.2 ;
        RECT  82.05 34.8 82.95 199.2 ;
        RECT  84.75 34.8 85.65 199.2 ;
        RECT  87.45 34.8 88.35 199.2 ;
        RECT  124.95 5.85 125.85 6.75 ;
        RECT  121.8 5.85 125.4 6.75 ;
        RECT  124.95 6.3 125.85 8.1 ;
        RECT  135.15 5.85 136.05 6.75 ;
        RECT  132.0 5.85 135.6 6.75 ;
        RECT  135.15 6.3 136.05 8.1 ;
        RECT  47.4 424.8 48.3 426.9 ;
        RECT  124.8 0.0 125.7 1.8 ;
        RECT  135.0 0.0 135.9 1.8 ;
        RECT  110.85 0.0 111.75 444.3 ;
        RECT  108.15 0.0 109.05 444.3 ;
        RECT  100.05 0.0 100.95 444.3 ;
        RECT  113.55 0.0 114.45 444.3 ;
        RECT  102.75 0.0 103.65 444.3 ;
        RECT  92.85 0.0 97.35 444.3 ;
        RECT  105.45 0.0 106.35 444.3 ;
        RECT  126.3 199.2 127.5 424.8 ;
        RECT  133.5 199.2 134.7 424.8 ;
        RECT  136.5 199.2 137.7 424.8 ;
        RECT  123.3 199.2 124.5 424.8 ;
        RECT  129.9 199.2 131.1 424.8 ;
        RECT  129.9 199.2 131.1 213.9 ;
        RECT  126.0 199.2 127.5 200.4 ;
        RECT  121.8 199.2 124.5 200.4 ;
        RECT  126.3 199.2 127.5 213.9 ;
        RECT  123.3 199.2 124.5 212.7 ;
        RECT  119.7 203.4 122.1 213.9 ;
        RECT  123.3 199.2 124.5 212.7 ;
        RECT  129.9 199.2 131.1 213.9 ;
        RECT  119.7 203.4 122.1 213.9 ;
        RECT  126.3 199.2 127.5 213.9 ;
        RECT  129.9 212.7 131.1 227.4 ;
        RECT  126.0 226.2 127.5 227.4 ;
        RECT  121.8 226.2 124.5 227.4 ;
        RECT  126.3 212.7 127.5 227.4 ;
        RECT  123.3 213.9 124.5 227.4 ;
        RECT  119.7 212.7 122.1 223.2 ;
        RECT  123.3 213.9 124.5 227.4 ;
        RECT  129.9 212.7 131.1 227.4 ;
        RECT  119.7 212.7 122.1 223.2 ;
        RECT  126.3 212.7 127.5 227.4 ;
        RECT  129.9 227.4 131.1 242.1 ;
        RECT  126.0 227.4 127.5 228.6 ;
        RECT  121.8 227.4 124.5 228.6 ;
        RECT  126.3 227.4 127.5 242.1 ;
        RECT  123.3 227.4 124.5 240.9 ;
        RECT  119.7 231.6 122.1 242.1 ;
        RECT  123.3 227.4 124.5 240.9 ;
        RECT  129.9 227.4 131.1 242.1 ;
        RECT  119.7 231.6 122.1 242.1 ;
        RECT  126.3 227.4 127.5 242.1 ;
        RECT  129.9 240.9 131.1 255.6 ;
        RECT  126.0 254.4 127.5 255.6 ;
        RECT  121.8 254.4 124.5 255.6 ;
        RECT  126.3 240.9 127.5 255.6 ;
        RECT  123.3 242.1 124.5 255.6 ;
        RECT  119.7 240.9 122.1 251.4 ;
        RECT  123.3 242.1 124.5 255.6 ;
        RECT  129.9 240.9 131.1 255.6 ;
        RECT  119.7 240.9 122.1 251.4 ;
        RECT  126.3 240.9 127.5 255.6 ;
        RECT  129.9 255.6 131.1 270.3 ;
        RECT  126.0 255.6 127.5 256.8 ;
        RECT  121.8 255.6 124.5 256.8 ;
        RECT  126.3 255.6 127.5 270.3 ;
        RECT  123.3 255.6 124.5 269.1 ;
        RECT  119.7 259.8 122.1 270.3 ;
        RECT  123.3 255.6 124.5 269.1 ;
        RECT  129.9 255.6 131.1 270.3 ;
        RECT  119.7 259.8 122.1 270.3 ;
        RECT  126.3 255.6 127.5 270.3 ;
        RECT  129.9 269.1 131.1 283.8 ;
        RECT  126.0 282.6 127.5 283.8 ;
        RECT  121.8 282.6 124.5 283.8 ;
        RECT  126.3 269.1 127.5 283.8 ;
        RECT  123.3 270.3 124.5 283.8 ;
        RECT  119.7 269.1 122.1 279.6 ;
        RECT  123.3 270.3 124.5 283.8 ;
        RECT  129.9 269.1 131.1 283.8 ;
        RECT  119.7 269.1 122.1 279.6 ;
        RECT  126.3 269.1 127.5 283.8 ;
        RECT  129.9 283.8 131.1 298.5 ;
        RECT  126.0 283.8 127.5 285.0 ;
        RECT  121.8 283.8 124.5 285.0 ;
        RECT  126.3 283.8 127.5 298.5 ;
        RECT  123.3 283.8 124.5 297.3 ;
        RECT  119.7 288.0 122.1 298.5 ;
        RECT  123.3 283.8 124.5 297.3 ;
        RECT  129.9 283.8 131.1 298.5 ;
        RECT  119.7 288.0 122.1 298.5 ;
        RECT  126.3 283.8 127.5 298.5 ;
        RECT  129.9 297.3 131.1 312.0 ;
        RECT  126.0 310.8 127.5 312.0 ;
        RECT  121.8 310.8 124.5 312.0 ;
        RECT  126.3 297.3 127.5 312.0 ;
        RECT  123.3 298.5 124.5 312.0 ;
        RECT  119.7 297.3 122.1 307.8 ;
        RECT  123.3 298.5 124.5 312.0 ;
        RECT  129.9 297.3 131.1 312.0 ;
        RECT  119.7 297.3 122.1 307.8 ;
        RECT  126.3 297.3 127.5 312.0 ;
        RECT  129.9 312.0 131.1 326.7 ;
        RECT  126.0 312.0 127.5 313.2 ;
        RECT  121.8 312.0 124.5 313.2 ;
        RECT  126.3 312.0 127.5 326.7 ;
        RECT  123.3 312.0 124.5 325.5 ;
        RECT  119.7 316.2 122.1 326.7 ;
        RECT  123.3 312.0 124.5 325.5 ;
        RECT  129.9 312.0 131.1 326.7 ;
        RECT  119.7 316.2 122.1 326.7 ;
        RECT  126.3 312.0 127.5 326.7 ;
        RECT  129.9 325.5 131.1 340.2 ;
        RECT  126.0 339.0 127.5 340.2 ;
        RECT  121.8 339.0 124.5 340.2 ;
        RECT  126.3 325.5 127.5 340.2 ;
        RECT  123.3 326.7 124.5 340.2 ;
        RECT  119.7 325.5 122.1 336.0 ;
        RECT  123.3 326.7 124.5 340.2 ;
        RECT  129.9 325.5 131.1 340.2 ;
        RECT  119.7 325.5 122.1 336.0 ;
        RECT  126.3 325.5 127.5 340.2 ;
        RECT  129.9 340.2 131.1 354.9 ;
        RECT  126.0 340.2 127.5 341.4 ;
        RECT  121.8 340.2 124.5 341.4 ;
        RECT  126.3 340.2 127.5 354.9 ;
        RECT  123.3 340.2 124.5 353.7 ;
        RECT  119.7 344.4 122.1 354.9 ;
        RECT  123.3 340.2 124.5 353.7 ;
        RECT  129.9 340.2 131.1 354.9 ;
        RECT  119.7 344.4 122.1 354.9 ;
        RECT  126.3 340.2 127.5 354.9 ;
        RECT  129.9 353.7 131.1 368.4 ;
        RECT  126.0 367.2 127.5 368.4 ;
        RECT  121.8 367.2 124.5 368.4 ;
        RECT  126.3 353.7 127.5 368.4 ;
        RECT  123.3 354.9 124.5 368.4 ;
        RECT  119.7 353.7 122.1 364.2 ;
        RECT  123.3 354.9 124.5 368.4 ;
        RECT  129.9 353.7 131.1 368.4 ;
        RECT  119.7 353.7 122.1 364.2 ;
        RECT  126.3 353.7 127.5 368.4 ;
        RECT  129.9 368.4 131.1 383.1 ;
        RECT  126.0 368.4 127.5 369.6 ;
        RECT  121.8 368.4 124.5 369.6 ;
        RECT  126.3 368.4 127.5 383.1 ;
        RECT  123.3 368.4 124.5 381.9 ;
        RECT  119.7 372.6 122.1 383.1 ;
        RECT  123.3 368.4 124.5 381.9 ;
        RECT  129.9 368.4 131.1 383.1 ;
        RECT  119.7 372.6 122.1 383.1 ;
        RECT  126.3 368.4 127.5 383.1 ;
        RECT  129.9 381.9 131.1 396.6 ;
        RECT  126.0 395.4 127.5 396.6 ;
        RECT  121.8 395.4 124.5 396.6 ;
        RECT  126.3 381.9 127.5 396.6 ;
        RECT  123.3 383.1 124.5 396.6 ;
        RECT  119.7 381.9 122.1 392.4 ;
        RECT  123.3 383.1 124.5 396.6 ;
        RECT  129.9 381.9 131.1 396.6 ;
        RECT  119.7 381.9 122.1 392.4 ;
        RECT  126.3 381.9 127.5 396.6 ;
        RECT  129.9 396.6 131.1 411.3 ;
        RECT  126.0 396.6 127.5 397.8 ;
        RECT  121.8 396.6 124.5 397.8 ;
        RECT  126.3 396.6 127.5 411.3 ;
        RECT  123.3 396.6 124.5 410.1 ;
        RECT  119.7 400.8 122.1 411.3 ;
        RECT  123.3 396.6 124.5 410.1 ;
        RECT  129.9 396.6 131.1 411.3 ;
        RECT  119.7 400.8 122.1 411.3 ;
        RECT  126.3 396.6 127.5 411.3 ;
        RECT  129.9 410.1 131.1 424.8 ;
        RECT  126.0 423.6 127.5 424.8 ;
        RECT  121.8 423.6 124.5 424.8 ;
        RECT  126.3 410.1 127.5 424.8 ;
        RECT  123.3 411.3 124.5 424.8 ;
        RECT  119.7 410.1 122.1 420.6 ;
        RECT  123.3 411.3 124.5 424.8 ;
        RECT  129.9 410.1 131.1 424.8 ;
        RECT  119.7 410.1 122.1 420.6 ;
        RECT  126.3 410.1 127.5 424.8 ;
        RECT  140.1 199.2 141.3 213.9 ;
        RECT  136.2 199.2 137.7 200.4 ;
        RECT  132.0 199.2 134.7 200.4 ;
        RECT  136.5 199.2 137.7 213.9 ;
        RECT  133.5 199.2 134.7 212.7 ;
        RECT  129.9 203.4 132.3 213.9 ;
        RECT  133.5 199.2 134.7 212.7 ;
        RECT  140.1 199.2 141.3 213.9 ;
        RECT  129.9 203.4 132.3 213.9 ;
        RECT  136.5 199.2 137.7 213.9 ;
        RECT  140.1 212.7 141.3 227.4 ;
        RECT  136.2 226.2 137.7 227.4 ;
        RECT  132.0 226.2 134.7 227.4 ;
        RECT  136.5 212.7 137.7 227.4 ;
        RECT  133.5 213.9 134.7 227.4 ;
        RECT  129.9 212.7 132.3 223.2 ;
        RECT  133.5 213.9 134.7 227.4 ;
        RECT  140.1 212.7 141.3 227.4 ;
        RECT  129.9 212.7 132.3 223.2 ;
        RECT  136.5 212.7 137.7 227.4 ;
        RECT  140.1 227.4 141.3 242.1 ;
        RECT  136.2 227.4 137.7 228.6 ;
        RECT  132.0 227.4 134.7 228.6 ;
        RECT  136.5 227.4 137.7 242.1 ;
        RECT  133.5 227.4 134.7 240.9 ;
        RECT  129.9 231.6 132.3 242.1 ;
        RECT  133.5 227.4 134.7 240.9 ;
        RECT  140.1 227.4 141.3 242.1 ;
        RECT  129.9 231.6 132.3 242.1 ;
        RECT  136.5 227.4 137.7 242.1 ;
        RECT  140.1 240.9 141.3 255.6 ;
        RECT  136.2 254.4 137.7 255.6 ;
        RECT  132.0 254.4 134.7 255.6 ;
        RECT  136.5 240.9 137.7 255.6 ;
        RECT  133.5 242.1 134.7 255.6 ;
        RECT  129.9 240.9 132.3 251.4 ;
        RECT  133.5 242.1 134.7 255.6 ;
        RECT  140.1 240.9 141.3 255.6 ;
        RECT  129.9 240.9 132.3 251.4 ;
        RECT  136.5 240.9 137.7 255.6 ;
        RECT  140.1 255.6 141.3 270.3 ;
        RECT  136.2 255.6 137.7 256.8 ;
        RECT  132.0 255.6 134.7 256.8 ;
        RECT  136.5 255.6 137.7 270.3 ;
        RECT  133.5 255.6 134.7 269.1 ;
        RECT  129.9 259.8 132.3 270.3 ;
        RECT  133.5 255.6 134.7 269.1 ;
        RECT  140.1 255.6 141.3 270.3 ;
        RECT  129.9 259.8 132.3 270.3 ;
        RECT  136.5 255.6 137.7 270.3 ;
        RECT  140.1 269.1 141.3 283.8 ;
        RECT  136.2 282.6 137.7 283.8 ;
        RECT  132.0 282.6 134.7 283.8 ;
        RECT  136.5 269.1 137.7 283.8 ;
        RECT  133.5 270.3 134.7 283.8 ;
        RECT  129.9 269.1 132.3 279.6 ;
        RECT  133.5 270.3 134.7 283.8 ;
        RECT  140.1 269.1 141.3 283.8 ;
        RECT  129.9 269.1 132.3 279.6 ;
        RECT  136.5 269.1 137.7 283.8 ;
        RECT  140.1 283.8 141.3 298.5 ;
        RECT  136.2 283.8 137.7 285.0 ;
        RECT  132.0 283.8 134.7 285.0 ;
        RECT  136.5 283.8 137.7 298.5 ;
        RECT  133.5 283.8 134.7 297.3 ;
        RECT  129.9 288.0 132.3 298.5 ;
        RECT  133.5 283.8 134.7 297.3 ;
        RECT  140.1 283.8 141.3 298.5 ;
        RECT  129.9 288.0 132.3 298.5 ;
        RECT  136.5 283.8 137.7 298.5 ;
        RECT  140.1 297.3 141.3 312.0 ;
        RECT  136.2 310.8 137.7 312.0 ;
        RECT  132.0 310.8 134.7 312.0 ;
        RECT  136.5 297.3 137.7 312.0 ;
        RECT  133.5 298.5 134.7 312.0 ;
        RECT  129.9 297.3 132.3 307.8 ;
        RECT  133.5 298.5 134.7 312.0 ;
        RECT  140.1 297.3 141.3 312.0 ;
        RECT  129.9 297.3 132.3 307.8 ;
        RECT  136.5 297.3 137.7 312.0 ;
        RECT  140.1 312.0 141.3 326.7 ;
        RECT  136.2 312.0 137.7 313.2 ;
        RECT  132.0 312.0 134.7 313.2 ;
        RECT  136.5 312.0 137.7 326.7 ;
        RECT  133.5 312.0 134.7 325.5 ;
        RECT  129.9 316.2 132.3 326.7 ;
        RECT  133.5 312.0 134.7 325.5 ;
        RECT  140.1 312.0 141.3 326.7 ;
        RECT  129.9 316.2 132.3 326.7 ;
        RECT  136.5 312.0 137.7 326.7 ;
        RECT  140.1 325.5 141.3 340.2 ;
        RECT  136.2 339.0 137.7 340.2 ;
        RECT  132.0 339.0 134.7 340.2 ;
        RECT  136.5 325.5 137.7 340.2 ;
        RECT  133.5 326.7 134.7 340.2 ;
        RECT  129.9 325.5 132.3 336.0 ;
        RECT  133.5 326.7 134.7 340.2 ;
        RECT  140.1 325.5 141.3 340.2 ;
        RECT  129.9 325.5 132.3 336.0 ;
        RECT  136.5 325.5 137.7 340.2 ;
        RECT  140.1 340.2 141.3 354.9 ;
        RECT  136.2 340.2 137.7 341.4 ;
        RECT  132.0 340.2 134.7 341.4 ;
        RECT  136.5 340.2 137.7 354.9 ;
        RECT  133.5 340.2 134.7 353.7 ;
        RECT  129.9 344.4 132.3 354.9 ;
        RECT  133.5 340.2 134.7 353.7 ;
        RECT  140.1 340.2 141.3 354.9 ;
        RECT  129.9 344.4 132.3 354.9 ;
        RECT  136.5 340.2 137.7 354.9 ;
        RECT  140.1 353.7 141.3 368.4 ;
        RECT  136.2 367.2 137.7 368.4 ;
        RECT  132.0 367.2 134.7 368.4 ;
        RECT  136.5 353.7 137.7 368.4 ;
        RECT  133.5 354.9 134.7 368.4 ;
        RECT  129.9 353.7 132.3 364.2 ;
        RECT  133.5 354.9 134.7 368.4 ;
        RECT  140.1 353.7 141.3 368.4 ;
        RECT  129.9 353.7 132.3 364.2 ;
        RECT  136.5 353.7 137.7 368.4 ;
        RECT  140.1 368.4 141.3 383.1 ;
        RECT  136.2 368.4 137.7 369.6 ;
        RECT  132.0 368.4 134.7 369.6 ;
        RECT  136.5 368.4 137.7 383.1 ;
        RECT  133.5 368.4 134.7 381.9 ;
        RECT  129.9 372.6 132.3 383.1 ;
        RECT  133.5 368.4 134.7 381.9 ;
        RECT  140.1 368.4 141.3 383.1 ;
        RECT  129.9 372.6 132.3 383.1 ;
        RECT  136.5 368.4 137.7 383.1 ;
        RECT  140.1 381.9 141.3 396.6 ;
        RECT  136.2 395.4 137.7 396.6 ;
        RECT  132.0 395.4 134.7 396.6 ;
        RECT  136.5 381.9 137.7 396.6 ;
        RECT  133.5 383.1 134.7 396.6 ;
        RECT  129.9 381.9 132.3 392.4 ;
        RECT  133.5 383.1 134.7 396.6 ;
        RECT  140.1 381.9 141.3 396.6 ;
        RECT  129.9 381.9 132.3 392.4 ;
        RECT  136.5 381.9 137.7 396.6 ;
        RECT  140.1 396.6 141.3 411.3 ;
        RECT  136.2 396.6 137.7 397.8 ;
        RECT  132.0 396.6 134.7 397.8 ;
        RECT  136.5 396.6 137.7 411.3 ;
        RECT  133.5 396.6 134.7 410.1 ;
        RECT  129.9 400.8 132.3 411.3 ;
        RECT  133.5 396.6 134.7 410.1 ;
        RECT  140.1 396.6 141.3 411.3 ;
        RECT  129.9 400.8 132.3 411.3 ;
        RECT  136.5 396.6 137.7 411.3 ;
        RECT  140.1 410.1 141.3 424.8 ;
        RECT  136.2 423.6 137.7 424.8 ;
        RECT  132.0 423.6 134.7 424.8 ;
        RECT  136.5 410.1 137.7 424.8 ;
        RECT  133.5 411.3 134.7 424.8 ;
        RECT  129.9 410.1 132.3 420.6 ;
        RECT  133.5 411.3 134.7 424.8 ;
        RECT  140.1 410.1 141.3 424.8 ;
        RECT  129.9 410.1 132.3 420.6 ;
        RECT  136.5 410.1 137.7 424.8 ;
        RECT  133.65 424.8 134.55 444.3 ;
        RECT  123.45 424.8 124.35 444.3 ;
        RECT  136.65 424.8 137.55 444.3 ;
        RECT  126.45 424.8 127.35 444.3 ;
        RECT  123.75 435.9 123.9 437.1 ;
        RECT  126.45 435.9 128.1 437.1 ;
        RECT  123.75 427.5 123.9 428.7 ;
        RECT  125.7 427.5 126.45 428.7 ;
        RECT  123.45 424.8 124.35 444.3 ;
        RECT  126.45 424.8 127.35 444.3 ;
        RECT  123.3 435.9 124.5 437.1 ;
        RECT  128.1 435.9 129.3 437.1 ;
        RECT  123.3 427.5 124.5 428.7 ;
        RECT  125.7 427.5 126.9 428.7 ;
        RECT  133.95 435.9 134.1 437.1 ;
        RECT  136.65 435.9 138.3 437.1 ;
        RECT  133.95 427.5 134.1 428.7 ;
        RECT  135.9 427.5 136.65 428.7 ;
        RECT  133.65 424.8 134.55 444.3 ;
        RECT  136.65 424.8 137.55 444.3 ;
        RECT  133.5 435.9 134.7 437.1 ;
        RECT  138.3 435.9 139.5 437.1 ;
        RECT  133.5 427.5 134.7 428.7 ;
        RECT  135.9 427.5 137.1 428.7 ;
        RECT  133.5 150.3 134.7 163.5 ;
        RECT  123.3 150.3 124.5 163.5 ;
        RECT  136.5 150.3 137.7 163.5 ;
        RECT  126.3 150.3 127.5 163.5 ;
        RECT  123.3 164.7 124.5 199.2 ;
        RECT  126.3 164.7 127.5 199.2 ;
        RECT  129.9 191.7 131.1 199.2 ;
        RECT  123.3 163.5 125.4 164.7 ;
        RECT  126.3 163.5 128.1 164.7 ;
        RECT  121.2 150.3 122.4 154.8 ;
        RECT  123.3 150.3 124.5 163.5 ;
        RECT  126.3 150.3 127.5 163.5 ;
        RECT  126.3 150.3 127.5 163.5 ;
        RECT  123.3 150.3 124.5 163.5 ;
        RECT  133.5 164.7 134.7 199.2 ;
        RECT  136.5 164.7 137.7 199.2 ;
        RECT  140.1 191.7 141.3 199.2 ;
        RECT  133.5 163.5 135.6 164.7 ;
        RECT  136.5 163.5 138.3 164.7 ;
        RECT  131.4 150.3 132.6 154.8 ;
        RECT  133.5 150.3 134.7 163.5 ;
        RECT  136.5 150.3 137.7 163.5 ;
        RECT  136.5 150.3 137.7 163.5 ;
        RECT  133.5 150.3 134.7 163.5 ;
        RECT  124.8 90.0 126.0 92.7 ;
        RECT  135.0 90.0 136.2 92.7 ;
        RECT  123.3 148.2 124.5 150.3 ;
        RECT  133.5 148.2 134.7 150.3 ;
        RECT  136.5 142.8 137.7 150.3 ;
        RECT  126.3 142.8 127.5 150.3 ;
        RECT  123.3 148.2 124.5 150.3 ;
        RECT  121.8 147.0 124.5 148.2 ;
        RECT  126.3 142.8 127.5 150.3 ;
        RECT  129.9 138.0 131.1 148.5 ;
        RECT  123.6 136.8 131.1 138.0 ;
        RECT  122.7 99.0 123.9 126.3 ;
        RECT  129.9 115.5 131.1 136.8 ;
        RECT  129.3 114.3 131.1 115.5 ;
        RECT  129.9 111.3 131.1 114.3 ;
        RECT  126.0 110.1 131.1 111.3 ;
        RECT  126.0 108.9 127.2 110.1 ;
        RECT  123.9 92.7 126.3 93.9 ;
        RECT  124.8 90.0 126.0 92.7 ;
        RECT  129.9 90.0 131.1 110.1 ;
        RECT  124.8 90.0 126.0 92.7 ;
        RECT  126.3 142.8 127.5 150.3 ;
        RECT  123.3 148.2 124.5 150.3 ;
        RECT  133.5 148.2 134.7 150.3 ;
        RECT  132.0 147.0 134.7 148.2 ;
        RECT  136.5 142.8 137.7 150.3 ;
        RECT  140.1 138.0 141.3 148.5 ;
        RECT  133.8 136.8 141.3 138.0 ;
        RECT  132.9 99.0 134.1 126.3 ;
        RECT  140.1 115.5 141.3 136.8 ;
        RECT  139.5 114.3 141.3 115.5 ;
        RECT  140.1 111.3 141.3 114.3 ;
        RECT  136.2 110.1 141.3 111.3 ;
        RECT  136.2 108.9 137.4 110.1 ;
        RECT  134.1 92.7 136.5 93.9 ;
        RECT  135.0 90.0 136.2 92.7 ;
        RECT  140.1 90.0 141.3 110.1 ;
        RECT  135.0 90.0 136.2 92.7 ;
        RECT  136.5 142.8 137.7 150.3 ;
        RECT  133.5 148.2 134.7 150.3 ;
        RECT  137.7 85.5 138.9 90.0 ;
        RECT  135.0 30.0 136.2 31.2 ;
        RECT  124.8 30.0 126.0 31.2 ;
        RECT  129.9 30.0 131.1 90.0 ;
        RECT  122.1 85.5 123.3 90.0 ;
        RECT  124.8 88.8 126.0 90.0 ;
        RECT  135.0 88.8 136.2 90.0 ;
        RECT  122.1 85.5 123.3 90.0 ;
        RECT  124.8 88.8 126.0 90.0 ;
        RECT  124.8 87.6 127.5 88.8 ;
        RECT  122.1 84.3 125.1 85.5 ;
        RECT  122.1 74.7 123.0 84.3 ;
        RECT  126.3 79.8 127.5 87.6 ;
        RECT  125.4 76.5 128.4 77.7 ;
        RECT  122.1 73.5 123.3 74.7 ;
        RECT  125.4 74.4 126.6 75.6 ;
        RECT  125.7 72.9 126.6 74.4 ;
        RECT  124.2 72.0 126.6 72.9 ;
        RECT  124.2 65.7 125.1 72.0 ;
        RECT  127.5 71.1 128.4 76.5 ;
        RECT  126.3 69.9 128.4 71.1 ;
        RECT  126.3 67.5 128.4 68.7 ;
        RECT  123.9 64.5 125.1 65.7 ;
        RECT  121.8 60.0 123.3 61.2 ;
        RECT  121.8 48.3 122.7 60.0 ;
        RECT  124.8 57.9 126.0 62.4 ;
        RECT  123.6 57.0 126.0 57.9 ;
        RECT  123.6 50.1 124.5 57.0 ;
        RECT  127.5 55.5 128.4 67.5 ;
        RECT  126.3 54.3 128.4 55.5 ;
        RECT  125.4 51.0 128.4 52.2 ;
        RECT  123.6 49.2 125.1 50.1 ;
        RECT  121.8 47.1 123.3 48.3 ;
        RECT  124.2 48.0 126.6 49.2 ;
        RECT  124.2 39.3 125.1 48.0 ;
        RECT  127.5 44.7 128.4 51.0 ;
        RECT  126.3 43.5 128.4 44.7 ;
        RECT  126.3 41.1 128.4 42.3 ;
        RECT  123.9 38.1 125.1 39.3 ;
        RECT  127.5 32.4 128.4 41.1 ;
        RECT  124.8 31.2 128.4 32.4 ;
        RECT  124.8 30.0 126.0 31.2 ;
        RECT  129.9 30.0 131.1 90.0 ;
        RECT  124.8 30.0 126.0 31.2 ;
        RECT  124.8 88.8 126.0 90.0 ;
        RECT  122.1 85.5 123.3 90.0 ;
        RECT  129.9 30.0 131.1 90.0 ;
        RECT  137.7 85.5 138.9 90.0 ;
        RECT  135.0 88.8 136.2 90.0 ;
        RECT  133.5 87.6 136.2 88.8 ;
        RECT  135.9 84.3 138.9 85.5 ;
        RECT  138.0 74.7 138.9 84.3 ;
        RECT  133.5 79.8 134.7 87.6 ;
        RECT  132.6 76.5 135.6 77.7 ;
        RECT  137.7 73.5 138.9 74.7 ;
        RECT  134.4 74.4 135.6 75.6 ;
        RECT  134.4 72.9 135.3 74.4 ;
        RECT  134.4 72.0 136.8 72.9 ;
        RECT  135.9 65.7 136.8 72.0 ;
        RECT  132.6 71.1 133.5 76.5 ;
        RECT  132.6 69.9 134.7 71.1 ;
        RECT  132.6 67.5 134.7 68.7 ;
        RECT  135.9 64.5 137.1 65.7 ;
        RECT  137.7 60.0 139.2 61.2 ;
        RECT  138.3 48.3 139.2 60.0 ;
        RECT  135.0 57.9 136.2 62.4 ;
        RECT  135.0 57.0 137.4 57.9 ;
        RECT  136.5 50.1 137.4 57.0 ;
        RECT  132.6 55.5 133.5 67.5 ;
        RECT  132.6 54.3 134.7 55.5 ;
        RECT  132.6 51.0 135.6 52.2 ;
        RECT  135.9 49.2 137.4 50.1 ;
        RECT  137.7 47.1 139.2 48.3 ;
        RECT  134.4 48.0 136.8 49.2 ;
        RECT  135.9 39.3 136.8 48.0 ;
        RECT  132.6 44.7 133.5 51.0 ;
        RECT  132.6 43.5 134.7 44.7 ;
        RECT  132.6 41.1 134.7 42.3 ;
        RECT  135.9 38.1 137.1 39.3 ;
        RECT  132.6 32.4 133.5 41.1 ;
        RECT  132.6 31.2 136.2 32.4 ;
        RECT  135.0 30.0 136.2 31.2 ;
        RECT  129.9 30.0 131.1 90.0 ;
        RECT  135.0 30.0 136.2 31.2 ;
        RECT  135.0 88.8 136.2 90.0 ;
        RECT  137.7 85.5 138.9 90.0 ;
        RECT  129.9 30.0 131.1 90.0 ;
        RECT  124.8 8.1 126.0 15.0 ;
        RECT  124.8 28.5 126.0 30.0 ;
        RECT  135.0 28.5 136.2 30.0 ;
        RECT  135.0 8.1 136.2 15.0 ;
        RECT  124.8 45.0 126.0 51.9 ;
        RECT  123.0 43.8 126.0 45.0 ;
        RECT  124.8 40.2 129.0 41.4 ;
        RECT  124.8 32.7 126.0 40.2 ;
        RECT  124.8 31.5 126.3 32.7 ;
        RECT  124.8 30.0 126.0 31.5 ;
        RECT  129.9 30.0 131.1 51.9 ;
        RECT  129.9 30.0 131.1 51.9 ;
        RECT  124.8 45.0 126.0 51.9 ;
        RECT  124.8 30.0 126.0 31.5 ;
        RECT  135.0 45.0 136.2 51.9 ;
        RECT  133.2 43.8 136.2 45.0 ;
        RECT  135.0 40.2 139.2 41.4 ;
        RECT  135.0 32.7 136.2 40.2 ;
        RECT  135.0 31.5 136.5 32.7 ;
        RECT  135.0 30.0 136.2 31.5 ;
        RECT  140.1 30.0 141.3 51.9 ;
        RECT  140.1 30.0 141.3 51.9 ;
        RECT  135.0 45.0 136.2 51.9 ;
        RECT  135.0 30.0 136.2 31.5 ;
        RECT  6.3 86.4 7.2 424.8 ;
        RECT  8.4 86.4 9.3 424.8 ;
        RECT  10.5 86.4 11.4 424.8 ;
        RECT  12.6 86.4 13.5 424.8 ;
        RECT  14.7 86.4 15.6 424.8 ;
        RECT  16.8 86.4 17.7 424.8 ;
        RECT  18.9 86.4 19.8 424.8 ;
        RECT  21.0 86.4 21.9 424.8 ;
        RECT  71.4 142.8 72.3 198.3 ;
        RECT  71.4 86.4 72.3 141.9 ;
        RECT  74.4 86.4 75.3 141.9 ;
        RECT  74.4 142.8 75.3 198.3 ;
        RECT  49.8 86.4 50.7 141.9 ;
        RECT  46.8 86.4 47.7 141.9 ;
        RECT  55.8 86.4 56.7 141.9 ;
        RECT  52.8 86.4 53.7 141.9 ;
        RECT  74.4 86.4 75.3 141.9 ;
        RECT  71.4 86.4 72.3 141.9 ;
        RECT  55.8 96.45 57.0 97.65 ;
        RECT  74.4 91.05 75.6 92.25 ;
        RECT  52.8 110.55 54.0 111.75 ;
        RECT  71.4 106.35 72.6 107.55 ;
        RECT  74.4 115.05 75.6 116.25 ;
        RECT  49.8 115.05 51.0 116.25 ;
        RECT  71.4 129.15 72.6 130.35 ;
        RECT  46.8 129.15 48.0 130.35 ;
        RECT  55.8 93.15 57.0 94.35 ;
        RECT  52.8 90.45 54.0 91.65 ;
        RECT  49.8 104.25 51.0 105.45 ;
        RECT  52.8 106.95 54.0 108.15 ;
        RECT  55.8 121.35 57.0 122.55 ;
        RECT  46.8 118.65 48.0 119.85 ;
        RECT  49.8 132.45 51.0 133.65 ;
        RECT  46.8 135.15 48.0 136.35 ;
        RECT  49.8 142.8 50.7 198.3 ;
        RECT  46.8 142.8 47.7 198.3 ;
        RECT  55.8 142.8 56.7 198.3 ;
        RECT  52.8 142.8 53.7 198.3 ;
        RECT  74.4 142.8 75.3 198.3 ;
        RECT  71.4 142.8 72.3 198.3 ;
        RECT  55.8 152.85 57.0 154.05 ;
        RECT  74.4 147.45 75.6 148.65 ;
        RECT  52.8 166.95 54.0 168.15 ;
        RECT  71.4 162.75 72.6 163.95 ;
        RECT  74.4 171.45 75.6 172.65 ;
        RECT  49.8 171.45 51.0 172.65 ;
        RECT  71.4 185.55 72.6 186.75 ;
        RECT  46.8 185.55 48.0 186.75 ;
        RECT  55.8 149.55 57.0 150.75 ;
        RECT  52.8 146.85 54.0 148.05 ;
        RECT  49.8 160.65 51.0 161.85 ;
        RECT  52.8 163.35 54.0 164.55 ;
        RECT  55.8 177.75 57.0 178.95 ;
        RECT  46.8 175.05 48.0 176.25 ;
        RECT  49.8 188.85 51.0 190.05 ;
        RECT  46.8 191.55 48.0 192.75 ;
        RECT  6.3 92.4 7.5 93.6 ;
        RECT  8.4 107.7 9.6 108.9 ;
        RECT  10.5 120.6 11.7 121.8 ;
        RECT  12.6 135.9 13.8 137.1 ;
        RECT  14.7 148.8 15.9 150.0 ;
        RECT  16.8 164.1 18.0 165.3 ;
        RECT  18.9 177.0 20.1 178.2 ;
        RECT  21.0 192.3 22.2 193.5 ;
        RECT  6.3 207.3 7.5 208.5 ;
        RECT  14.7 204.6 15.9 205.8 ;
        RECT  6.3 218.4 7.5 219.6 ;
        RECT  16.8 221.1 18.0 222.3 ;
        RECT  6.3 235.5 7.5 236.7 ;
        RECT  18.9 232.8 20.1 234.0 ;
        RECT  6.3 246.6 7.5 247.8 ;
        RECT  21.0 249.3 22.2 250.5 ;
        RECT  8.4 263.7 9.6 264.9 ;
        RECT  14.7 261.0 15.9 262.2 ;
        RECT  8.4 274.8 9.6 276.0 ;
        RECT  16.8 277.5 18.0 278.7 ;
        RECT  8.4 291.9 9.6 293.1 ;
        RECT  18.9 289.2 20.1 290.4 ;
        RECT  8.4 303.0 9.6 304.2 ;
        RECT  21.0 305.7 22.2 306.9 ;
        RECT  10.5 320.1 11.7 321.3 ;
        RECT  14.7 317.4 15.9 318.6 ;
        RECT  10.5 331.2 11.7 332.4 ;
        RECT  16.8 333.9 18.0 335.1 ;
        RECT  10.5 348.3 11.7 349.5 ;
        RECT  18.9 345.6 20.1 346.8 ;
        RECT  10.5 359.4 11.7 360.6 ;
        RECT  21.0 362.1 22.2 363.3 ;
        RECT  12.6 376.5 13.8 377.7 ;
        RECT  14.7 373.8 15.9 375.0 ;
        RECT  12.6 387.6 13.8 388.8 ;
        RECT  16.8 390.3 18.0 391.5 ;
        RECT  12.6 404.7 13.8 405.9 ;
        RECT  18.9 402.0 20.1 403.2 ;
        RECT  12.6 415.8 13.8 417.0 ;
        RECT  21.0 418.5 22.2 419.7 ;
        RECT  49.8 207.3 60.6 208.2 ;
        RECT  49.8 218.4 60.6 219.3 ;
        RECT  49.8 235.5 60.6 236.4 ;
        RECT  49.8 246.6 60.6 247.5 ;
        RECT  49.8 263.7 60.6 264.6 ;
        RECT  49.8 274.8 60.6 275.7 ;
        RECT  49.8 291.9 60.6 292.8 ;
        RECT  49.8 303.0 60.6 303.9 ;
        RECT  49.8 320.1 60.6 321.0 ;
        RECT  49.8 331.2 60.6 332.1 ;
        RECT  49.8 348.3 60.6 349.2 ;
        RECT  49.8 359.4 60.6 360.3 ;
        RECT  49.8 376.5 60.6 377.4 ;
        RECT  49.8 387.6 60.6 388.5 ;
        RECT  49.8 404.7 60.6 405.6 ;
        RECT  49.8 415.8 60.6 416.7 ;
        RECT  47.4 199.2 48.3 424.8 ;
        RECT  47.25 205.05 48.45 206.25 ;
        RECT  49.2 207.15 50.4 208.35 ;
        RECT  60.6 207.15 61.8 208.35 ;
        RECT  47.25 220.35 48.45 221.55 ;
        RECT  49.2 218.25 50.4 219.45 ;
        RECT  60.6 218.25 61.8 219.45 ;
        RECT  47.25 233.25 48.45 234.45 ;
        RECT  49.2 235.35 50.4 236.55 ;
        RECT  60.6 235.35 61.8 236.55 ;
        RECT  47.25 248.55 48.45 249.75 ;
        RECT  49.2 246.45 50.4 247.65 ;
        RECT  60.6 246.45 61.8 247.65 ;
        RECT  47.25 261.45 48.45 262.65 ;
        RECT  49.2 263.55 50.4 264.75 ;
        RECT  60.6 263.55 61.8 264.75 ;
        RECT  47.25 276.75 48.45 277.95 ;
        RECT  49.2 274.65 50.4 275.85 ;
        RECT  60.6 274.65 61.8 275.85 ;
        RECT  47.25 289.65 48.45 290.85 ;
        RECT  49.2 291.75 50.4 292.95 ;
        RECT  60.6 291.75 61.8 292.95 ;
        RECT  47.25 304.95 48.45 306.15 ;
        RECT  49.2 302.85 50.4 304.05 ;
        RECT  60.6 302.85 61.8 304.05 ;
        RECT  47.25 317.85 48.45 319.05 ;
        RECT  49.2 319.95 50.4 321.15 ;
        RECT  60.6 319.95 61.8 321.15 ;
        RECT  47.25 333.15 48.45 334.35 ;
        RECT  49.2 331.05 50.4 332.25 ;
        RECT  60.6 331.05 61.8 332.25 ;
        RECT  47.25 346.05 48.45 347.25 ;
        RECT  49.2 348.15 50.4 349.35 ;
        RECT  60.6 348.15 61.8 349.35 ;
        RECT  47.25 361.35 48.45 362.55 ;
        RECT  49.2 359.25 50.4 360.45 ;
        RECT  60.6 359.25 61.8 360.45 ;
        RECT  47.25 374.25 48.45 375.45 ;
        RECT  49.2 376.35 50.4 377.55 ;
        RECT  60.6 376.35 61.8 377.55 ;
        RECT  47.25 389.55 48.45 390.75 ;
        RECT  49.2 387.45 50.4 388.65 ;
        RECT  60.6 387.45 61.8 388.65 ;
        RECT  47.25 402.45 48.45 403.65 ;
        RECT  49.2 404.55 50.4 405.75 ;
        RECT  60.6 404.55 61.8 405.75 ;
        RECT  47.25 417.75 48.45 418.95 ;
        RECT  49.2 415.65 50.4 416.85 ;
        RECT  60.6 415.65 61.8 416.85 ;
        RECT  61.8 62.4 66.3 63.6 ;
        RECT  6.3 44.7 7.5 45.9 ;
        RECT  61.8 57.6 66.3 58.8 ;
        RECT  61.8 42.0 66.3 43.2 ;
        RECT  6.3 65.1 7.5 66.3 ;
        RECT  6.3 75.3 7.5 76.5 ;
        RECT  6.3 54.9 7.5 56.1 ;
        RECT  6.3 70.2 66.3 71.4 ;
        RECT  6.3 49.8 66.3 51.0 ;
        RECT  61.8 78.0 66.3 79.2 ;
        RECT  65.1 75.3 66.3 76.5 ;
        RECT  65.1 65.1 66.3 66.3 ;
        RECT  65.1 44.7 66.3 45.9 ;
        RECT  65.1 54.9 66.3 56.1 ;
        RECT  61.8 78.0 66.3 79.2 ;
        RECT  65.1 75.3 66.3 76.5 ;
        RECT  63.9 73.8 65.1 76.5 ;
        RECT  60.6 76.2 61.8 79.2 ;
        RECT  51.0 78.3 60.6 79.2 ;
        RECT  56.1 73.8 63.9 75.0 ;
        RECT  52.8 72.9 54.0 75.9 ;
        RECT  49.8 78.0 51.0 79.2 ;
        RECT  50.7 74.7 51.9 75.9 ;
        RECT  49.2 74.7 50.7 75.6 ;
        RECT  48.3 74.7 49.2 77.1 ;
        RECT  42.0 76.2 48.3 77.1 ;
        RECT  47.4 72.9 52.8 73.8 ;
        RECT  46.2 72.9 47.4 75.0 ;
        RECT  43.8 72.9 45.0 75.0 ;
        RECT  40.8 76.2 42.0 77.4 ;
        RECT  36.3 78.0 37.5 79.5 ;
        RECT  24.6 78.6 36.3 79.5 ;
        RECT  34.2 75.3 38.7 76.5 ;
        RECT  33.3 75.3 34.2 77.7 ;
        RECT  26.4 76.8 33.3 77.7 ;
        RECT  31.8 72.9 43.8 73.8 ;
        RECT  30.6 72.9 31.8 75.0 ;
        RECT  27.3 72.9 28.5 75.9 ;
        RECT  25.5 76.2 26.4 77.7 ;
        RECT  23.4 78.0 24.6 79.5 ;
        RECT  24.3 74.7 25.5 77.1 ;
        RECT  15.6 76.2 24.3 77.1 ;
        RECT  21.0 72.9 27.3 73.8 ;
        RECT  19.8 72.9 21.0 75.0 ;
        RECT  17.4 72.9 18.6 75.0 ;
        RECT  14.4 76.2 15.6 77.4 ;
        RECT  8.7 72.9 17.4 73.8 ;
        RECT  7.5 72.9 8.7 76.5 ;
        RECT  6.3 75.3 7.5 76.5 ;
        RECT  6.3 70.2 66.3 71.4 ;
        RECT  6.3 75.3 7.5 76.5 ;
        RECT  65.1 75.3 66.3 76.5 ;
        RECT  61.8 78.0 66.3 79.2 ;
        RECT  6.3 70.2 66.3 71.4 ;
        RECT  61.8 62.4 66.3 63.6 ;
        RECT  65.1 65.1 66.3 66.3 ;
        RECT  63.9 65.1 65.1 67.8 ;
        RECT  60.6 62.4 61.8 65.4 ;
        RECT  51.0 62.4 60.6 63.3 ;
        RECT  56.1 66.6 63.9 67.8 ;
        RECT  52.8 65.7 54.0 68.7 ;
        RECT  49.8 62.4 51.0 63.6 ;
        RECT  50.7 65.7 51.9 66.9 ;
        RECT  49.2 66.0 50.7 66.9 ;
        RECT  48.3 64.5 49.2 66.9 ;
        RECT  42.0 64.5 48.3 65.4 ;
        RECT  47.4 67.8 52.8 68.7 ;
        RECT  46.2 66.6 47.4 68.7 ;
        RECT  43.8 66.6 45.0 68.7 ;
        RECT  40.8 64.2 42.0 65.4 ;
        RECT  36.3 62.1 37.5 63.6 ;
        RECT  24.6 62.1 36.3 63.0 ;
        RECT  34.2 65.1 38.7 66.3 ;
        RECT  33.3 63.9 34.2 66.3 ;
        RECT  26.4 63.9 33.3 64.8 ;
        RECT  31.8 67.8 43.8 68.7 ;
        RECT  30.6 66.6 31.8 68.7 ;
        RECT  27.3 65.7 28.5 68.7 ;
        RECT  25.5 63.9 26.4 65.4 ;
        RECT  23.4 62.1 24.6 63.6 ;
        RECT  24.3 64.5 25.5 66.9 ;
        RECT  15.6 64.5 24.3 65.4 ;
        RECT  21.0 67.8 27.3 68.7 ;
        RECT  19.8 66.6 21.0 68.7 ;
        RECT  17.4 66.6 18.6 68.7 ;
        RECT  14.4 64.2 15.6 65.4 ;
        RECT  8.7 67.8 17.4 68.7 ;
        RECT  7.5 65.1 8.7 68.7 ;
        RECT  6.3 65.1 7.5 66.3 ;
        RECT  6.3 70.2 66.3 71.4 ;
        RECT  6.3 65.1 7.5 66.3 ;
        RECT  65.1 65.1 66.3 66.3 ;
        RECT  61.8 62.4 66.3 63.6 ;
        RECT  6.3 70.2 66.3 71.4 ;
        RECT  61.8 57.6 66.3 58.8 ;
        RECT  65.1 54.9 66.3 56.1 ;
        RECT  63.9 53.4 65.1 56.1 ;
        RECT  60.6 55.8 61.8 58.8 ;
        RECT  51.0 57.9 60.6 58.8 ;
        RECT  56.1 53.4 63.9 54.6 ;
        RECT  52.8 52.5 54.0 55.5 ;
        RECT  49.8 57.6 51.0 58.8 ;
        RECT  50.7 54.3 51.9 55.5 ;
        RECT  49.2 54.3 50.7 55.2 ;
        RECT  48.3 54.3 49.2 56.7 ;
        RECT  42.0 55.8 48.3 56.7 ;
        RECT  47.4 52.5 52.8 53.4 ;
        RECT  46.2 52.5 47.4 54.6 ;
        RECT  43.8 52.5 45.0 54.6 ;
        RECT  40.8 55.8 42.0 57.0 ;
        RECT  36.3 57.6 37.5 59.1 ;
        RECT  24.6 58.2 36.3 59.1 ;
        RECT  34.2 54.9 38.7 56.1 ;
        RECT  33.3 54.9 34.2 57.3 ;
        RECT  26.4 56.4 33.3 57.3 ;
        RECT  31.8 52.5 43.8 53.4 ;
        RECT  30.6 52.5 31.8 54.6 ;
        RECT  27.3 52.5 28.5 55.5 ;
        RECT  25.5 55.8 26.4 57.3 ;
        RECT  23.4 57.6 24.6 59.1 ;
        RECT  24.3 54.3 25.5 56.7 ;
        RECT  15.6 55.8 24.3 56.7 ;
        RECT  21.0 52.5 27.3 53.4 ;
        RECT  19.8 52.5 21.0 54.6 ;
        RECT  17.4 52.5 18.6 54.6 ;
        RECT  14.4 55.8 15.6 57.0 ;
        RECT  8.7 52.5 17.4 53.4 ;
        RECT  7.5 52.5 8.7 56.1 ;
        RECT  6.3 54.9 7.5 56.1 ;
        RECT  6.3 49.8 66.3 51.0 ;
        RECT  6.3 54.9 7.5 56.1 ;
        RECT  65.1 54.9 66.3 56.1 ;
        RECT  61.8 57.6 66.3 58.8 ;
        RECT  6.3 49.8 66.3 51.0 ;
        RECT  61.8 42.0 66.3 43.2 ;
        RECT  65.1 44.7 66.3 45.9 ;
        RECT  63.9 44.7 65.1 47.4 ;
        RECT  60.6 42.0 61.8 45.0 ;
        RECT  51.0 42.0 60.6 42.9 ;
        RECT  56.1 46.2 63.9 47.4 ;
        RECT  52.8 45.3 54.0 48.3 ;
        RECT  49.8 42.0 51.0 43.2 ;
        RECT  50.7 45.3 51.9 46.5 ;
        RECT  49.2 45.6 50.7 46.5 ;
        RECT  48.3 44.1 49.2 46.5 ;
        RECT  42.0 44.1 48.3 45.0 ;
        RECT  47.4 47.4 52.8 48.3 ;
        RECT  46.2 46.2 47.4 48.3 ;
        RECT  43.8 46.2 45.0 48.3 ;
        RECT  40.8 43.8 42.0 45.0 ;
        RECT  36.3 41.7 37.5 43.2 ;
        RECT  24.6 41.7 36.3 42.6 ;
        RECT  34.2 44.7 38.7 45.9 ;
        RECT  33.3 43.5 34.2 45.9 ;
        RECT  26.4 43.5 33.3 44.4 ;
        RECT  31.8 47.4 43.8 48.3 ;
        RECT  30.6 46.2 31.8 48.3 ;
        RECT  27.3 45.3 28.5 48.3 ;
        RECT  25.5 43.5 26.4 45.0 ;
        RECT  23.4 41.7 24.6 43.2 ;
        RECT  24.3 44.1 25.5 46.5 ;
        RECT  15.6 44.1 24.3 45.0 ;
        RECT  21.0 47.4 27.3 48.3 ;
        RECT  19.8 46.2 21.0 48.3 ;
        RECT  17.4 46.2 18.6 48.3 ;
        RECT  14.4 43.8 15.6 45.0 ;
        RECT  8.7 47.4 17.4 48.3 ;
        RECT  7.5 44.7 8.7 48.3 ;
        RECT  6.3 44.7 7.5 45.9 ;
        RECT  6.3 49.8 66.3 51.0 ;
        RECT  6.3 44.7 7.5 45.9 ;
        RECT  65.1 44.7 66.3 45.9 ;
        RECT  61.8 42.0 66.3 43.2 ;
        RECT  6.3 49.8 66.3 51.0 ;
        RECT  121.35 5.85 122.55 7.05 ;
        RECT  131.55 5.85 132.75 7.05 ;
        RECT  125.1 0.3 126.3 1.5 ;
        RECT  135.3 0.3 136.5 1.5 ;
        RECT  92.85 198.6 94.05 199.8 ;
        RECT  92.85 226.8 94.05 228.0 ;
        RECT  92.85 255.0 94.05 256.2 ;
        RECT  92.85 283.2 94.05 284.4 ;
        RECT  92.85 311.4 94.05 312.6 ;
        RECT  92.85 339.6 94.05 340.8 ;
        RECT  92.85 367.8 94.05 369.0 ;
        RECT  92.85 396.0 94.05 397.2 ;
        RECT  92.85 424.2 94.05 425.4 ;
        RECT  74.1 88.65 75.3 89.85 ;
        RECT  79.05 88.65 80.25 89.85 ;
        RECT  71.1 102.75 72.3 103.95 ;
        RECT  81.75 102.75 82.95 103.95 ;
        RECT  74.1 145.05 75.3 146.25 ;
        RECT  84.45 145.05 85.65 146.25 ;
        RECT  71.1 159.15 72.3 160.35 ;
        RECT  87.15 159.15 88.35 160.35 ;
        RECT  76.2 85.8 77.4 87.0 ;
        RECT  76.2 85.8 77.4 87.0 ;
        RECT  92.25 85.8 93.45 87.0 ;
        RECT  76.2 114.0 77.4 115.2 ;
        RECT  76.2 114.0 77.4 115.2 ;
        RECT  92.25 114.0 93.45 115.2 ;
        RECT  76.2 142.2 77.4 143.4 ;
        RECT  76.2 142.2 77.4 143.4 ;
        RECT  92.25 142.2 93.45 143.4 ;
        RECT  76.2 170.4 77.4 171.6 ;
        RECT  76.2 170.4 77.4 171.6 ;
        RECT  92.25 170.4 93.45 171.6 ;
        RECT  66.3 75.3 67.5 76.5 ;
        RECT  79.05 75.45 80.25 76.65 ;
        RECT  66.3 65.1 67.5 66.3 ;
        RECT  81.75 65.25 82.95 66.45 ;
        RECT  66.3 54.9 67.5 56.1 ;
        RECT  84.45 55.05 85.65 56.25 ;
        RECT  66.3 44.7 67.5 45.9 ;
        RECT  87.15 44.85 88.35 46.05 ;
        RECT  66.3 70.2 67.5 71.4 ;
        RECT  92.85 70.35 94.05 71.55 ;
        RECT  66.3 49.8 67.5 51.0 ;
        RECT  92.85 49.95 94.05 51.15 ;
        RECT  108.0 32.25 109.2 33.45 ;
        RECT  102.6 27.75 103.8 28.95 ;
        RECT  105.3 25.35 106.5 26.55 ;
        RECT  108.0 431.25 109.2 432.45 ;
        RECT  110.7 96.75 111.9 97.95 ;
        RECT  113.4 194.85 114.6 196.05 ;
        RECT  100.05 82.65 101.25 83.85 ;
        RECT  47.25 426.3 48.45 427.5 ;
        RECT  100.05 426.45 101.25 427.65 ;
        RECT  96.15 23.4 97.35 24.6 ;
        RECT  96.15 192.9 97.35 194.1 ;
        RECT  96.15 94.8 97.35 96.0 ;
        RECT  -53.1 311.1 -3.0 312.0 ;
        RECT  -53.1 313.8 -3.0 314.7 ;
        RECT  -53.1 316.5 -3.0 317.4 ;
        RECT  -53.1 321.9 -3.0 322.8 ;
        RECT  -50.7 321.9 -48.0 322.8 ;
        RECT  -48.0 311.1 -45.3 312.0 ;
        RECT  -35.1 313.8 -32.4 314.7 ;
        RECT  -30.3 316.5 -27.6 317.4 ;
        RECT  -42.9 308.4 -40.2 309.3 ;
        RECT  -22.5 308.4 -19.8 309.3 ;
        RECT  -9.45 305.7 -6.75 306.6 ;
        RECT  -9.45 324.6 -6.75 325.5 ;
        RECT  -20.25 205.05 -19.35 306.15 ;
        RECT  -26.85 305.7 -24.15 306.6 ;
        RECT  -24.75 311.1 -22.05 312.0 ;
        RECT  -22.65 324.6 -19.95 325.5 ;
        RECT  -25.35 321.9 -22.65 322.8 ;
        RECT  -12.3 324.6 -9.6 325.5 ;
        RECT  -10.2 321.9 -7.5 322.8 ;
        RECT  -8.1 313.8 -5.4 314.7 ;
        RECT  -40.5 324.6 -37.8 325.5 ;
        RECT  -38.4 316.5 -35.7 317.4 ;
        RECT  -36.3 313.8 -33.6 314.7 ;
        RECT  -5.7 308.4 -3.0 309.3 ;
        RECT  -17.1 319.2 -14.4 320.1 ;
        RECT  -31.2 308.4 -28.5 309.3 ;
        RECT  -45.3 319.2 -42.6 320.1 ;
        RECT  -53.1 324.6 -3.0 325.5 ;
        RECT  -38.1 384.0 -3.0 384.9 ;
        RECT  -53.1 305.7 -3.0 306.6 ;
        RECT  -25.2 361.5 -3.0 362.4 ;
        RECT  -53.1 319.2 -3.0 320.1 ;
        RECT  -53.1 308.4 -3.0 309.3 ;
        RECT  -25.2 364.2 -3.0 365.1 ;
        RECT  -27.3 346.8 -3.0 347.7 ;
        RECT  -35.7 257.7 -34.5 262.2 ;
        RECT  -30.9 257.7 -29.7 262.2 ;
        RECT  -38.4 202.2 -37.2 203.4 ;
        RECT  -48.6 202.2 -47.4 203.4 ;
        RECT  -28.2 202.2 -27.0 203.4 ;
        RECT  -43.5 202.2 -42.3 262.2 ;
        RECT  -23.1 202.2 -21.9 262.2 ;
        RECT  -51.3 257.7 -50.1 262.2 ;
        RECT  -48.6 261.0 -47.4 262.2 ;
        RECT  -38.4 261.0 -37.2 262.2 ;
        RECT  -28.2 261.0 -27.0 262.2 ;
        RECT  -51.3 257.7 -50.1 262.2 ;
        RECT  -48.6 261.0 -47.4 262.2 ;
        RECT  -48.6 259.8 -45.9 261.0 ;
        RECT  -51.3 256.5 -48.3 257.7 ;
        RECT  -51.3 246.9 -50.4 256.5 ;
        RECT  -47.1 252.0 -45.9 259.8 ;
        RECT  -48.0 248.7 -45.0 249.9 ;
        RECT  -51.3 245.7 -50.1 246.9 ;
        RECT  -48.0 246.6 -46.8 247.8 ;
        RECT  -47.7 245.1 -46.8 246.6 ;
        RECT  -49.2 244.2 -46.8 245.1 ;
        RECT  -49.2 237.9 -48.3 244.2 ;
        RECT  -45.9 243.3 -45.0 248.7 ;
        RECT  -47.1 242.1 -45.0 243.3 ;
        RECT  -47.1 239.7 -45.0 240.9 ;
        RECT  -49.5 236.7 -48.3 237.9 ;
        RECT  -51.6 232.2 -50.1 233.4 ;
        RECT  -51.6 220.5 -50.7 232.2 ;
        RECT  -48.6 230.1 -47.4 234.6 ;
        RECT  -49.8 229.2 -47.4 230.1 ;
        RECT  -49.8 222.3 -48.9 229.2 ;
        RECT  -45.9 227.7 -45.0 239.7 ;
        RECT  -47.1 226.5 -45.0 227.7 ;
        RECT  -48.0 223.2 -45.0 224.4 ;
        RECT  -49.8 221.4 -48.3 222.3 ;
        RECT  -51.6 219.3 -50.1 220.5 ;
        RECT  -49.2 220.2 -46.8 221.4 ;
        RECT  -49.2 211.5 -48.3 220.2 ;
        RECT  -45.9 216.9 -45.0 223.2 ;
        RECT  -47.1 215.7 -45.0 216.9 ;
        RECT  -47.1 213.3 -45.0 214.5 ;
        RECT  -49.5 210.3 -48.3 211.5 ;
        RECT  -45.9 204.6 -45.0 213.3 ;
        RECT  -48.6 203.4 -45.0 204.6 ;
        RECT  -48.6 202.2 -47.4 203.4 ;
        RECT  -43.5 202.2 -42.3 262.2 ;
        RECT  -48.6 202.2 -47.4 203.4 ;
        RECT  -48.6 261.0 -47.4 262.2 ;
        RECT  -51.3 257.7 -50.1 262.2 ;
        RECT  -43.5 202.2 -42.3 262.2 ;
        RECT  -35.7 257.7 -34.5 262.2 ;
        RECT  -38.4 261.0 -37.2 262.2 ;
        RECT  -39.9 259.8 -37.2 261.0 ;
        RECT  -37.5 256.5 -34.5 257.7 ;
        RECT  -35.4 246.9 -34.5 256.5 ;
        RECT  -39.9 252.0 -38.7 259.8 ;
        RECT  -40.8 248.7 -37.8 249.9 ;
        RECT  -35.7 245.7 -34.5 246.9 ;
        RECT  -39.0 246.6 -37.8 247.8 ;
        RECT  -39.0 245.1 -38.1 246.6 ;
        RECT  -39.0 244.2 -36.6 245.1 ;
        RECT  -37.5 237.9 -36.6 244.2 ;
        RECT  -40.8 243.3 -39.9 248.7 ;
        RECT  -40.8 242.1 -38.7 243.3 ;
        RECT  -40.8 239.7 -38.7 240.9 ;
        RECT  -37.5 236.7 -36.3 237.9 ;
        RECT  -35.7 232.2 -34.2 233.4 ;
        RECT  -35.1 220.5 -34.2 232.2 ;
        RECT  -38.4 230.1 -37.2 234.6 ;
        RECT  -38.4 229.2 -36.0 230.1 ;
        RECT  -36.9 222.3 -36.0 229.2 ;
        RECT  -40.8 227.7 -39.9 239.7 ;
        RECT  -40.8 226.5 -38.7 227.7 ;
        RECT  -40.8 223.2 -37.8 224.4 ;
        RECT  -37.5 221.4 -36.0 222.3 ;
        RECT  -35.7 219.3 -34.2 220.5 ;
        RECT  -39.0 220.2 -36.6 221.4 ;
        RECT  -37.5 211.5 -36.6 220.2 ;
        RECT  -40.8 216.9 -39.9 223.2 ;
        RECT  -40.8 215.7 -38.7 216.9 ;
        RECT  -40.8 213.3 -38.7 214.5 ;
        RECT  -37.5 210.3 -36.3 211.5 ;
        RECT  -40.8 204.6 -39.9 213.3 ;
        RECT  -40.8 203.4 -37.2 204.6 ;
        RECT  -38.4 202.2 -37.2 203.4 ;
        RECT  -43.5 202.2 -42.3 262.2 ;
        RECT  -38.4 202.2 -37.2 203.4 ;
        RECT  -38.4 261.0 -37.2 262.2 ;
        RECT  -35.7 257.7 -34.5 262.2 ;
        RECT  -43.5 202.2 -42.3 262.2 ;
        RECT  -30.9 257.7 -29.7 262.2 ;
        RECT  -28.2 261.0 -27.0 262.2 ;
        RECT  -28.2 259.8 -25.5 261.0 ;
        RECT  -30.9 256.5 -27.9 257.7 ;
        RECT  -30.9 246.9 -30.0 256.5 ;
        RECT  -26.7 252.0 -25.5 259.8 ;
        RECT  -27.6 248.7 -24.6 249.9 ;
        RECT  -30.9 245.7 -29.7 246.9 ;
        RECT  -27.6 246.6 -26.4 247.8 ;
        RECT  -27.3 245.1 -26.4 246.6 ;
        RECT  -28.8 244.2 -26.4 245.1 ;
        RECT  -28.8 237.9 -27.9 244.2 ;
        RECT  -25.5 243.3 -24.6 248.7 ;
        RECT  -26.7 242.1 -24.6 243.3 ;
        RECT  -26.7 239.7 -24.6 240.9 ;
        RECT  -29.1 236.7 -27.9 237.9 ;
        RECT  -31.2 232.2 -29.7 233.4 ;
        RECT  -31.2 220.5 -30.3 232.2 ;
        RECT  -28.2 230.1 -27.0 234.6 ;
        RECT  -29.4 229.2 -27.0 230.1 ;
        RECT  -29.4 222.3 -28.5 229.2 ;
        RECT  -25.5 227.7 -24.6 239.7 ;
        RECT  -26.7 226.5 -24.6 227.7 ;
        RECT  -27.6 223.2 -24.6 224.4 ;
        RECT  -29.4 221.4 -27.9 222.3 ;
        RECT  -31.2 219.3 -29.7 220.5 ;
        RECT  -28.8 220.2 -26.4 221.4 ;
        RECT  -28.8 211.5 -27.9 220.2 ;
        RECT  -25.5 216.9 -24.6 223.2 ;
        RECT  -26.7 215.7 -24.6 216.9 ;
        RECT  -26.7 213.3 -24.6 214.5 ;
        RECT  -29.1 210.3 -27.9 211.5 ;
        RECT  -25.5 204.6 -24.6 213.3 ;
        RECT  -28.2 203.4 -24.6 204.6 ;
        RECT  -28.2 202.2 -27.0 203.4 ;
        RECT  -23.1 202.2 -21.9 262.2 ;
        RECT  -28.2 202.2 -27.0 203.4 ;
        RECT  -28.2 261.0 -27.0 262.2 ;
        RECT  -30.9 257.7 -29.7 262.2 ;
        RECT  -23.1 202.2 -21.9 262.2 ;
        RECT  -15.45 335.4 -14.25 341.4 ;
        RECT  -15.45 335.4 -14.25 336.6 ;
        RECT  -15.45 340.2 -14.25 341.4 ;
        RECT  -26.85 341.55 -21.3 342.45 ;
        RECT  -22.5 341.4 -21.3 342.6 ;
        RECT  -28.65 341.4 -27.45 342.6 ;
        RECT  -43.65 345.0 -42.45 351.0 ;
        RECT  -43.65 345.0 -42.45 346.2 ;
        RECT  -43.65 349.8 -42.45 351.0 ;
        RECT  -51.3 321.75 -50.1 322.95 ;
        RECT  -51.45 262.2 -50.25 263.4 ;
        RECT  -51.45 261.9 -50.25 263.1 ;
        RECT  -48.6 310.95 -47.4 312.15 ;
        RECT  -48.75 262.2 -47.55 263.4 ;
        RECT  -48.75 261.9 -47.55 263.1 ;
        RECT  -35.7 313.65 -34.5 314.85 ;
        RECT  -35.85 262.2 -34.65 263.4 ;
        RECT  -35.85 261.9 -34.65 263.1 ;
        RECT  -30.9 316.35 -29.7 317.55 ;
        RECT  -31.05 262.2 -29.85 263.4 ;
        RECT  -31.05 261.9 -29.85 263.1 ;
        RECT  -43.5 308.25 -42.3 309.45 ;
        RECT  -43.65 261.9 -42.45 263.1 ;
        RECT  -23.1 308.25 -21.9 309.45 ;
        RECT  -23.25 261.9 -22.05 263.1 ;
        RECT  -31.65 395.7 -30.75 450.9 ;
        RECT  -31.65 405.3 -30.75 408.0 ;
        RECT  -31.65 408.0 -30.75 450.9 ;
        RECT  -47.25 448.2 -46.35 450.9 ;
        RECT  -33.9 400.5 -33.0 408.0 ;
        RECT  -40.65 400.5 -39.75 405.3 ;
        RECT  -9.9 424.5 -9.0 428.7 ;
        RECT  -9.9 415.35 -9.0 419.1 ;
        RECT  -25.2 414.9 -24.3 415.35 ;
        RECT  -25.2 420.3 -24.3 424.5 ;
        RECT  -10.2 432.9 -9.0 434.1 ;
        RECT  -10.2 423.3 -9.0 424.5 ;
        RECT  -25.2 414.9 -24.0 416.1 ;
        RECT  -25.2 424.5 -24.0 425.7 ;
        RECT  -10.2 427.5 -9.0 428.7 ;
        RECT  -10.2 417.9 -9.0 419.1 ;
        RECT  -10.05 414.75 -8.85 415.95 ;
        RECT  -25.35 414.75 -24.15 415.95 ;
        RECT  -25.2 420.3 -24.0 421.5 ;
        RECT  -38.4 424.2 -36.6 434.7 ;
        RECT  -40.8 421.2 -39.6 434.7 ;
        RECT  -43.8 421.2 -42.6 434.7 ;
        RECT  -40.8 420.0 -38.1 421.2 ;
        RECT  -43.8 420.0 -42.3 421.2 ;
        RECT  -47.4 420.0 -46.2 434.7 ;
        RECT  -40.8 421.2 -39.6 434.7 ;
        RECT  -38.4 424.2 -36.6 434.7 ;
        RECT  -47.4 420.0 -46.2 434.7 ;
        RECT  -43.8 421.2 -42.6 434.7 ;
        RECT  -40.8 391.8 -39.6 420.0 ;
        RECT  -47.4 391.8 -46.2 420.0 ;
        RECT  -43.8 391.8 -42.6 420.0 ;
        RECT  -47.4 405.3 -46.2 420.0 ;
        RECT  -43.8 418.8 -42.3 420.0 ;
        RECT  -40.8 418.8 -38.1 420.0 ;
        RECT  -43.8 405.3 -42.6 420.0 ;
        RECT  -40.8 406.5 -39.6 420.0 ;
        RECT  -38.4 405.3 -36.0 415.8 ;
        RECT  -40.8 406.5 -39.6 420.0 ;
        RECT  -47.4 405.3 -46.2 420.0 ;
        RECT  -38.4 405.3 -36.0 415.8 ;
        RECT  -43.8 405.3 -42.6 420.0 ;
        RECT  -47.4 391.8 -46.2 406.5 ;
        RECT  -43.8 391.8 -42.3 393.0 ;
        RECT  -40.8 391.8 -38.1 393.0 ;
        RECT  -43.8 391.8 -42.6 406.5 ;
        RECT  -40.8 391.8 -39.6 405.3 ;
        RECT  -38.4 396.0 -36.0 406.5 ;
        RECT  -40.8 391.8 -39.6 405.3 ;
        RECT  -47.4 391.8 -46.2 406.5 ;
        RECT  -38.4 396.0 -36.0 406.5 ;
        RECT  -43.8 391.8 -42.6 406.5 ;
        RECT  -31.95 420.9 -30.75 422.1 ;
        RECT  -31.95 443.7 -30.75 444.9 ;
        RECT  -31.95 432.9 -30.75 434.1 ;
        RECT  -31.95 393.3 -30.75 394.5 ;
        RECT  -31.8 449.1 -30.6 450.3 ;
        RECT  -47.4 449.1 -46.2 450.3 ;
        RECT  -34.05 406.2 -32.85 407.4 ;
        RECT  -34.05 398.7 -32.85 399.9 ;
        RECT  -40.8 398.7 -39.6 399.9 ;
        RECT  -10.05 305.55 -8.85 306.75 ;
        RECT  -10.05 324.45 -8.85 325.65 ;
        RECT  -10.2 257.4 -9.0 258.6 ;
        RECT  -10.2 257.1 -9.0 258.3 ;
        RECT  -20.4 204.45 -19.2 205.65 ;
        RECT  -27.45 305.55 -26.25 306.75 ;
        RECT  -25.35 310.95 -24.15 312.15 ;
        RECT  -23.25 324.45 -22.05 325.65 ;
        RECT  -23.4 349.5 -22.2 350.7 ;
        RECT  -23.4 349.2 -22.2 350.4 ;
        RECT  -25.95 321.75 -24.75 322.95 ;
        RECT  -26.1 349.5 -24.9 350.7 ;
        RECT  -26.1 349.2 -24.9 350.4 ;
        RECT  -12.9 324.45 -11.7 325.65 ;
        RECT  -10.8 321.75 -9.6 322.95 ;
        RECT  -8.7 313.65 -7.5 314.85 ;
        RECT  -41.1 324.45 -39.9 325.65 ;
        RECT  -39.0 316.35 -37.8 317.55 ;
        RECT  -36.9 313.65 -35.7 314.85 ;
        RECT  -27.3 346.8 -26.1 348.0 ;
        RECT  -25.2 361.5 -24.0 362.7 ;
        RECT  -38.1 384.0 -36.9 385.2 ;
        RECT  -25.2 364.2 -24.0 365.4 ;
        RECT  -3.6 308.25 -2.4 309.45 ;
        RECT  -17.7 319.05 -16.5 320.25 ;
        RECT  -31.8 308.25 -30.6 309.45 ;
        RECT  -45.9 319.05 -44.7 320.25 ;
        RECT  113.4 364.05 114.6 365.25 ;
        RECT  -4.5 364.2 -3.3 365.4 ;
        RECT  110.7 383.85 111.9 385.05 ;
        RECT  -4.5 384.0 -3.3 385.2 ;
        RECT  105.3 346.65 106.5 347.85 ;
        RECT  -4.5 346.8 -3.3 348.0 ;
        RECT  102.6 361.35 103.8 362.55 ;
        RECT  -4.5 361.5 -3.3 362.7 ;
        RECT  108.0 324.45 109.2 325.65 ;
        RECT  -4.5 324.6 -3.3 325.8 ;
        RECT  99.9 305.55 101.1 306.75 ;
        RECT  -4.5 305.7 -3.3 306.9 ;
        RECT  1.65 319.05 2.85 320.25 ;
        RECT  94.5 308.25 95.7 309.45 ;
        RECT  -4.5 308.4 -3.3 309.6 ;
        LAYER  via2 ;
        RECT  121.5 151.8 122.1 152.4 ;
        RECT  131.7 151.8 132.3 152.4 ;
        RECT  125.1 31.5 125.7 32.1 ;
        RECT  135.3 31.5 135.9 32.1 ;
        RECT  125.1 31.8 125.7 32.4 ;
        RECT  135.3 31.8 135.9 32.4 ;
        RECT  7.8 75.6 8.4 76.2 ;
        RECT  7.8 65.4 8.4 66.0 ;
        RECT  7.8 55.2 8.4 55.8 ;
        RECT  7.8 45.0 8.4 45.6 ;
        RECT  121.65 6.15 122.25 6.75 ;
        RECT  131.85 6.15 132.45 6.75 ;
        RECT  125.4 0.6 126.0 1.2 ;
        RECT  135.6 0.6 136.2 1.2 ;
        RECT  76.5 86.1 77.1 86.7 ;
        RECT  92.55 86.1 93.15 86.7 ;
        RECT  76.5 114.3 77.1 114.9 ;
        RECT  92.55 114.3 93.15 114.9 ;
        RECT  76.5 142.5 77.1 143.1 ;
        RECT  92.55 142.5 93.15 143.1 ;
        RECT  76.5 170.7 77.1 171.3 ;
        RECT  92.55 170.7 93.15 171.3 ;
        RECT  -48.3 203.7 -47.7 204.3 ;
        RECT  -38.1 203.7 -37.5 204.3 ;
        RECT  -27.9 203.7 -27.3 204.3 ;
        RECT  -51.0 322.05 -50.4 322.65 ;
        RECT  -51.15 262.2 -50.55 262.8 ;
        RECT  -48.3 311.25 -47.7 311.85 ;
        RECT  -48.45 262.2 -47.85 262.8 ;
        RECT  -35.4 313.95 -34.8 314.55 ;
        RECT  -35.55 262.2 -34.95 262.8 ;
        RECT  -30.6 316.65 -30.0 317.25 ;
        RECT  -30.75 262.2 -30.15 262.8 ;
        RECT  -43.2 308.55 -42.6 309.15 ;
        RECT  -43.35 262.2 -42.75 262.8 ;
        RECT  -22.8 308.55 -22.2 309.15 ;
        RECT  -22.95 262.2 -22.35 262.8 ;
        RECT  -9.75 415.05 -9.15 415.65 ;
        RECT  -25.05 415.05 -24.45 415.65 ;
        RECT  -9.75 324.75 -9.15 325.35 ;
        RECT  -9.9 257.4 -9.3 258.0 ;
        RECT  -22.95 324.75 -22.35 325.35 ;
        RECT  -23.1 349.5 -22.5 350.1 ;
        RECT  -25.65 322.05 -25.05 322.65 ;
        RECT  -25.8 349.5 -25.2 350.1 ;
        RECT  113.7 364.35 114.3 364.95 ;
        RECT  -4.2 364.5 -3.6 365.1 ;
        RECT  111.0 384.15 111.6 384.75 ;
        RECT  -4.2 384.3 -3.6 384.9 ;
        RECT  105.6 346.95 106.2 347.55 ;
        RECT  -4.2 347.1 -3.6 347.7 ;
        RECT  102.9 361.65 103.5 362.25 ;
        RECT  -4.2 361.8 -3.6 362.4 ;
        RECT  108.3 324.75 108.9 325.35 ;
        RECT  -4.2 324.9 -3.6 325.5 ;
        RECT  100.2 305.85 100.8 306.45 ;
        RECT  -4.2 306.0 -3.6 306.6 ;
        RECT  94.8 308.55 95.4 309.15 ;
        RECT  -4.2 308.7 -3.6 309.3 ;
        LAYER  metal3 ;
        RECT  -3.0 363.9 114.0 365.4 ;
        RECT  -3.0 383.7 111.3 385.2 ;
        RECT  -3.0 346.5 105.9 348.0 ;
        RECT  -3.0 361.2 103.2 362.7 ;
        RECT  -3.0 324.3 108.6 325.8 ;
        RECT  -3.0 305.4 100.5 306.9 ;
        RECT  -3.0 308.1 95.1 309.6 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  0.0 44.4 7.2 45.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  0.0 64.8 7.2 66.3 ;
        RECT  0.0 75.0 7.2 76.5 ;
        RECT  0.0 54.6 7.2 56.1 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  121.05 6.3 122.55 151.2 ;
        RECT  131.25 6.3 132.75 151.2 ;
        RECT  124.8 0.0 126.3 30.0 ;
        RECT  135.0 0.0 136.5 30.0 ;
        RECT  76.8 85.65 92.85 87.15 ;
        RECT  76.8 113.85 92.85 115.35 ;
        RECT  76.8 142.05 92.85 143.55 ;
        RECT  76.8 170.25 92.85 171.75 ;
        RECT  0.0 44.4 7.2 45.9 ;
        RECT  0.0 64.8 7.2 66.3 ;
        RECT  0.0 75.0 7.2 76.5 ;
        RECT  0.0 54.6 7.2 56.1 ;
        RECT  120.9 151.2 122.7 153.0 ;
        RECT  131.1 151.2 132.9 153.0 ;
        RECT  120.9 151.2 122.7 153.0 ;
        RECT  120.9 151.2 122.7 153.0 ;
        RECT  131.1 151.2 132.9 153.0 ;
        RECT  131.1 151.2 132.9 153.0 ;
        RECT  134.7 30.9 136.5 32.7 ;
        RECT  124.5 30.9 126.3 32.7 ;
        RECT  124.5 30.9 126.3 32.7 ;
        RECT  124.5 30.9 126.3 32.7 ;
        RECT  134.7 30.9 136.5 32.7 ;
        RECT  134.7 30.9 136.5 32.7 ;
        RECT  124.5 31.2 126.3 33.0 ;
        RECT  134.7 31.2 136.5 33.0 ;
        RECT  7.2 44.4 9.0 46.2 ;
        RECT  7.2 64.8 9.0 66.6 ;
        RECT  7.2 75.0 9.0 76.8 ;
        RECT  7.2 54.6 9.0 56.4 ;
        RECT  7.2 75.0 9.0 76.8 ;
        RECT  7.2 75.0 9.0 76.8 ;
        RECT  7.2 64.8 9.0 66.6 ;
        RECT  7.2 64.8 9.0 66.6 ;
        RECT  7.2 54.6 9.0 56.4 ;
        RECT  7.2 54.6 9.0 56.4 ;
        RECT  7.2 44.4 9.0 46.2 ;
        RECT  7.2 44.4 9.0 46.2 ;
        RECT  121.05 5.55 122.85 7.35 ;
        RECT  131.25 5.55 133.05 7.35 ;
        RECT  124.8 0.0 126.6 1.8 ;
        RECT  135.0 0.0 136.8 1.8 ;
        RECT  75.9 85.5 77.7 87.3 ;
        RECT  91.95 85.5 93.75 87.3 ;
        RECT  75.9 113.7 77.7 115.5 ;
        RECT  91.95 113.7 93.75 115.5 ;
        RECT  75.9 141.9 77.7 143.7 ;
        RECT  91.95 141.9 93.75 143.7 ;
        RECT  75.9 170.1 77.7 171.9 ;
        RECT  91.95 170.1 93.75 171.9 ;
        RECT  -51.45 262.2 -49.95 322.35 ;
        RECT  -48.75 262.2 -47.25 311.55 ;
        RECT  -35.85 262.2 -34.35 314.25 ;
        RECT  -31.05 262.2 -29.55 316.95 ;
        RECT  -43.65 262.2 -42.15 308.85 ;
        RECT  -23.25 262.2 -21.75 308.85 ;
        RECT  -10.2 257.4 -8.7 325.05 ;
        RECT  -23.4 325.05 -21.9 349.5 ;
        RECT  -26.1 322.35 -24.6 349.5 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -51.6 321.45 -49.8 323.25 ;
        RECT  -51.75 261.6 -49.95 263.4 ;
        RECT  -48.9 310.65 -47.1 312.45 ;
        RECT  -49.05 261.6 -47.25 263.4 ;
        RECT  -36.0 313.35 -34.2 315.15 ;
        RECT  -36.15 261.6 -34.35 263.4 ;
        RECT  -31.2 316.05 -29.4 317.85 ;
        RECT  -31.35 261.6 -29.55 263.4 ;
        RECT  -43.8 307.95 -42.0 309.75 ;
        RECT  -43.95 261.6 -42.15 263.4 ;
        RECT  -23.4 307.95 -21.6 309.75 ;
        RECT  -23.55 261.6 -21.75 263.4 ;
        RECT  -24.75 414.6 -9.45 416.1 ;
        RECT  -10.35 414.45 -8.55 416.25 ;
        RECT  -25.65 414.45 -23.85 416.25 ;
        RECT  -10.35 324.15 -8.55 325.95 ;
        RECT  -10.5 256.8 -8.7 258.6 ;
        RECT  -23.55 324.15 -21.75 325.95 ;
        RECT  -23.7 348.9 -21.9 350.7 ;
        RECT  -26.25 321.45 -24.45 323.25 ;
        RECT  -26.4 348.9 -24.6 350.7 ;
        RECT  113.1 363.75 114.9 365.55 ;
        RECT  -4.8 363.9 -3.0 365.7 ;
        RECT  110.4 383.55 112.2 385.35 ;
        RECT  -4.8 383.7 -3.0 385.5 ;
        RECT  105.0 346.35 106.8 348.15 ;
        RECT  -4.8 346.5 -3.0 348.3 ;
        RECT  102.3 361.05 104.1 362.85 ;
        RECT  -4.8 361.2 -3.0 363.0 ;
        RECT  107.7 324.15 109.5 325.95 ;
        RECT  -4.8 324.3 -3.0 326.1 ;
        RECT  99.6 305.25 101.4 307.05 ;
        RECT  -4.8 305.4 -3.0 307.2 ;
        RECT  94.2 307.95 96.0 309.75 ;
        RECT  -4.8 308.1 -3.0 309.9 ;
    END
END    sram_2_16_1_scn3me_subm
END    LIBRARY
