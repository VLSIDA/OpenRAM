magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1296 -1277 2424 2731
<< nwell >>
rect -36 679 1164 1471
<< poly >>
rect 114 740 144 907
rect 81 674 144 740
rect 114 507 144 674
<< locali >>
rect 0 1397 1128 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 64 674 98 740
rect 596 724 630 1096
rect 596 690 647 724
rect 596 318 630 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 0 -17 1128 17
use pmos_m9_w2_000_sli_dli_da_p  pmos_m9_w2_000_sli_dli_da_p_0
timestamp 1595931502
transform 1 0 54 0 1 963
box -59 -56 1073 454
use nmos_m9_w2_000_sli_dli_da_p  nmos_m9_w2_000_sli_dli_da_p_0
timestamp 1595931502
transform 1 0 54 0 1 51
box 0 -26 1014 456
use contact_12  contact_12_0
timestamp 1595931502
transform 1 0 48 0 1 674
box 0 0 66 66
<< labels >>
rlabel corelocali s 564 0 564 0 4 gnd
rlabel corelocali s 630 707 630 707 4 Z
rlabel corelocali s 564 1414 564 1414 4 vdd
rlabel corelocali s 81 707 81 707 4 A
<< properties >>
string FIXED_BBOX 0 0 1128 1414
<< end >>
