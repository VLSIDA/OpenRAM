MACRO sram_2_16_1_freepdk45
    CLASS RING ;
    ORIGIN 4.22 0.0 ;
    FOREIGN  sram 0.0 0.0 ;
    SIZE 16.475 BY 42.27 ;
    SYMMETRY X Y R90 ;
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  11.95 0.0 12.3 42.27 ;
        RECT  11.95 0.0 12.3 42.27 ;
        RECT  0.0 0.0 0.35 42.27 ;
        RECT  0.0 0.0 0.35 42.27 ;
        END
    END vdd
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal2 ;
        RECT  8.2525 0.0 8.6025 42.27 ;
        RECT  8.2525 0.0 8.6025 42.27 ;
        END
    END gnd
    PIN DATA[0]
        DIRECTION INOUT ;
        PORT
        LAYER metal2 ;
        RECT  10.6625 0.0 10.7325 0.14 ;
        RECT  10.6625 0.0 10.7325 0.14 ;
        RECT  10.6625 0.0 10.7325 0.135 ;
        END
    END DATA[0]
    PIN DATA[1]
        DIRECTION INOUT ;
        PORT
        LAYER metal2 ;
        RECT  11.3675 0.0 11.4375 0.14 ;
        RECT  11.3675 0.0 11.4375 0.14 ;
        RECT  11.3675 0.0 11.4375 0.135 ;
        END
    END DATA[1]
    PIN ADDR[0]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 7.5325 0.48 7.6025 ;
        RECT  0.0 7.5325 0.48 7.6025 ;
        END
    END ADDR[0]
    PIN ADDR[1]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 6.8275 0.48 6.8975 ;
        RECT  0.0 6.8275 0.48 6.8975 ;
        END
    END ADDR[1]
    PIN ADDR[2]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 6.1225 0.48 6.1925 ;
        RECT  0.0 6.1225 0.48 6.1925 ;
        END
    END ADDR[2]
    PIN ADDR[3]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 5.4175 0.48 5.4875 ;
        RECT  0.0 5.4175 0.48 5.4875 ;
        END
    END ADDR[3]
    PIN CSb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        END
    END CSb
    PIN OEb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        END
    END OEb
    PIN WEb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        END
    END WEb
    PIN clk
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.79 19.355 -0.655 19.42 ;
        RECT  -0.79 19.355 -0.655 19.42 ;
        RECT  -0.79 19.355 -0.655 19.42 ;
        RECT  -0.79 19.355 -0.655 19.42 ;
        END
    END clk
    OBS
        LAYER  metal1 ;
        RECT  0.1425 26.935 0.2075 27.14 ;
        RECT  -0.79 19.355 -0.655 19.42 ;
        RECT  11.95 0.0 12.3 42.27 ;
        RECT  0.0 0.0 0.35 42.27 ;
        RECT  4.3 19.64 4.365 19.705 ;
        RECT  4.3 19.4125 4.365 19.4775 ;
        RECT  4.23 19.64 4.3325 19.705 ;
        RECT  4.3 19.445 4.365 19.6725 ;
        RECT  4.3325 19.4125 4.435 19.4775 ;
        RECT  8.4575 19.64 8.5225 19.705 ;
        RECT  8.4575 19.1975 8.5225 19.2625 ;
        RECT  6.725 19.64 8.49 19.705 ;
        RECT  8.4575 19.23 8.5225 19.6725 ;
        RECT  8.49 19.1975 10.255 19.2625 ;
        RECT  4.3 21.165 4.365 21.23 ;
        RECT  4.3 21.3925 4.365 21.4575 ;
        RECT  4.23 21.165 4.3325 21.23 ;
        RECT  4.3 21.1975 4.365 21.425 ;
        RECT  4.3325 21.3925 4.435 21.4575 ;
        RECT  8.4575 21.165 8.5225 21.23 ;
        RECT  8.4575 21.6075 8.5225 21.6725 ;
        RECT  6.725 21.165 8.49 21.23 ;
        RECT  8.4575 21.1975 8.5225 21.64 ;
        RECT  8.49 21.6075 10.255 21.6725 ;
        RECT  4.3 22.33 4.365 22.395 ;
        RECT  4.3 22.1025 4.365 22.1675 ;
        RECT  4.23 22.33 4.3325 22.395 ;
        RECT  4.3 22.135 4.365 22.3625 ;
        RECT  4.3325 22.1025 4.435 22.1675 ;
        RECT  8.4575 22.33 8.5225 22.395 ;
        RECT  8.4575 21.8875 8.5225 21.9525 ;
        RECT  6.725 22.33 8.49 22.395 ;
        RECT  8.4575 21.92 8.5225 22.3625 ;
        RECT  8.49 21.8875 10.255 21.9525 ;
        RECT  4.3 23.855 4.365 23.92 ;
        RECT  4.3 24.0825 4.365 24.1475 ;
        RECT  4.23 23.855 4.3325 23.92 ;
        RECT  4.3 23.8875 4.365 24.115 ;
        RECT  4.3325 24.0825 4.435 24.1475 ;
        RECT  8.4575 23.855 8.5225 23.92 ;
        RECT  8.4575 24.2975 8.5225 24.3625 ;
        RECT  6.725 23.855 8.49 23.92 ;
        RECT  8.4575 23.8875 8.5225 24.33 ;
        RECT  8.49 24.2975 10.255 24.3625 ;
        RECT  4.3 25.02 4.365 25.085 ;
        RECT  4.3 24.7925 4.365 24.8575 ;
        RECT  4.23 25.02 4.3325 25.085 ;
        RECT  4.3 24.825 4.365 25.0525 ;
        RECT  4.3325 24.7925 4.435 24.8575 ;
        RECT  8.4575 25.02 8.5225 25.085 ;
        RECT  8.4575 24.5775 8.5225 24.6425 ;
        RECT  6.725 25.02 8.49 25.085 ;
        RECT  8.4575 24.61 8.5225 25.0525 ;
        RECT  8.49 24.5775 10.255 24.6425 ;
        RECT  4.3 26.545 4.365 26.61 ;
        RECT  4.3 26.7725 4.365 26.8375 ;
        RECT  4.23 26.545 4.3325 26.61 ;
        RECT  4.3 26.5775 4.365 26.805 ;
        RECT  4.3325 26.7725 4.435 26.8375 ;
        RECT  8.4575 26.545 8.5225 26.61 ;
        RECT  8.4575 26.9875 8.5225 27.0525 ;
        RECT  6.725 26.545 8.49 26.61 ;
        RECT  8.4575 26.5775 8.5225 27.02 ;
        RECT  8.49 26.9875 10.255 27.0525 ;
        RECT  4.3 27.71 4.365 27.775 ;
        RECT  4.3 27.4825 4.365 27.5475 ;
        RECT  4.23 27.71 4.3325 27.775 ;
        RECT  4.3 27.515 4.365 27.7425 ;
        RECT  4.3325 27.4825 4.435 27.5475 ;
        RECT  8.4575 27.71 8.5225 27.775 ;
        RECT  8.4575 27.2675 8.5225 27.3325 ;
        RECT  6.725 27.71 8.49 27.775 ;
        RECT  8.4575 27.3 8.5225 27.7425 ;
        RECT  8.49 27.2675 10.255 27.3325 ;
        RECT  4.3 29.235 4.365 29.3 ;
        RECT  4.3 29.4625 4.365 29.5275 ;
        RECT  4.23 29.235 4.3325 29.3 ;
        RECT  4.3 29.2675 4.365 29.495 ;
        RECT  4.3325 29.4625 4.435 29.5275 ;
        RECT  8.4575 29.235 8.5225 29.3 ;
        RECT  8.4575 29.6775 8.5225 29.7425 ;
        RECT  6.725 29.235 8.49 29.3 ;
        RECT  8.4575 29.2675 8.5225 29.71 ;
        RECT  8.49 29.6775 10.255 29.7425 ;
        RECT  4.3 30.4 4.365 30.465 ;
        RECT  4.3 30.1725 4.365 30.2375 ;
        RECT  4.23 30.4 4.3325 30.465 ;
        RECT  4.3 30.205 4.365 30.4325 ;
        RECT  4.3325 30.1725 4.435 30.2375 ;
        RECT  8.4575 30.4 8.5225 30.465 ;
        RECT  8.4575 29.9575 8.5225 30.0225 ;
        RECT  6.725 30.4 8.49 30.465 ;
        RECT  8.4575 29.99 8.5225 30.4325 ;
        RECT  8.49 29.9575 10.255 30.0225 ;
        RECT  4.3 31.925 4.365 31.99 ;
        RECT  4.3 32.1525 4.365 32.2175 ;
        RECT  4.23 31.925 4.3325 31.99 ;
        RECT  4.3 31.9575 4.365 32.185 ;
        RECT  4.3325 32.1525 4.435 32.2175 ;
        RECT  8.4575 31.925 8.5225 31.99 ;
        RECT  8.4575 32.3675 8.5225 32.4325 ;
        RECT  6.725 31.925 8.49 31.99 ;
        RECT  8.4575 31.9575 8.5225 32.4 ;
        RECT  8.49 32.3675 10.255 32.4325 ;
        RECT  4.3 33.09 4.365 33.155 ;
        RECT  4.3 32.8625 4.365 32.9275 ;
        RECT  4.23 33.09 4.3325 33.155 ;
        RECT  4.3 32.895 4.365 33.1225 ;
        RECT  4.3325 32.8625 4.435 32.9275 ;
        RECT  8.4575 33.09 8.5225 33.155 ;
        RECT  8.4575 32.6475 8.5225 32.7125 ;
        RECT  6.725 33.09 8.49 33.155 ;
        RECT  8.4575 32.68 8.5225 33.1225 ;
        RECT  8.49 32.6475 10.255 32.7125 ;
        RECT  4.3 34.615 4.365 34.68 ;
        RECT  4.3 34.8425 4.365 34.9075 ;
        RECT  4.23 34.615 4.3325 34.68 ;
        RECT  4.3 34.6475 4.365 34.875 ;
        RECT  4.3325 34.8425 4.435 34.9075 ;
        RECT  8.4575 34.615 8.5225 34.68 ;
        RECT  8.4575 35.0575 8.5225 35.1225 ;
        RECT  6.725 34.615 8.49 34.68 ;
        RECT  8.4575 34.6475 8.5225 35.09 ;
        RECT  8.49 35.0575 10.255 35.1225 ;
        RECT  4.3 35.78 4.365 35.845 ;
        RECT  4.3 35.5525 4.365 35.6175 ;
        RECT  4.23 35.78 4.3325 35.845 ;
        RECT  4.3 35.585 4.365 35.8125 ;
        RECT  4.3325 35.5525 4.435 35.6175 ;
        RECT  8.4575 35.78 8.5225 35.845 ;
        RECT  8.4575 35.3375 8.5225 35.4025 ;
        RECT  6.725 35.78 8.49 35.845 ;
        RECT  8.4575 35.37 8.5225 35.8125 ;
        RECT  8.49 35.3375 10.255 35.4025 ;
        RECT  4.3 37.305 4.365 37.37 ;
        RECT  4.3 37.5325 4.365 37.5975 ;
        RECT  4.23 37.305 4.3325 37.37 ;
        RECT  4.3 37.3375 4.365 37.565 ;
        RECT  4.3325 37.5325 4.435 37.5975 ;
        RECT  8.4575 37.305 8.5225 37.37 ;
        RECT  8.4575 37.7475 8.5225 37.8125 ;
        RECT  6.725 37.305 8.49 37.37 ;
        RECT  8.4575 37.3375 8.5225 37.78 ;
        RECT  8.49 37.7475 10.255 37.8125 ;
        RECT  4.3 38.47 4.365 38.535 ;
        RECT  4.3 38.2425 4.365 38.3075 ;
        RECT  4.23 38.47 4.3325 38.535 ;
        RECT  4.3 38.275 4.365 38.5025 ;
        RECT  4.3325 38.2425 4.435 38.3075 ;
        RECT  8.4575 38.47 8.5225 38.535 ;
        RECT  8.4575 38.0275 8.5225 38.0925 ;
        RECT  6.725 38.47 8.49 38.535 ;
        RECT  8.4575 38.06 8.5225 38.5025 ;
        RECT  8.49 38.0275 10.255 38.0925 ;
        RECT  4.3 39.995 4.365 40.06 ;
        RECT  4.3 40.2225 4.365 40.2875 ;
        RECT  4.23 39.995 4.3325 40.06 ;
        RECT  4.3 40.0275 4.365 40.255 ;
        RECT  4.3325 40.2225 4.435 40.2875 ;
        RECT  8.4575 39.995 8.5225 40.06 ;
        RECT  8.4575 40.4375 8.5225 40.5025 ;
        RECT  6.725 39.995 8.49 40.06 ;
        RECT  8.4575 40.0275 8.5225 40.47 ;
        RECT  8.49 40.4375 10.255 40.5025 ;
        RECT  4.89 19.0575 10.345 19.1225 ;
        RECT  4.89 21.7475 10.345 21.8125 ;
        RECT  4.89 24.4375 10.345 24.5025 ;
        RECT  4.89 27.1275 10.345 27.1925 ;
        RECT  4.89 29.8175 10.345 29.8825 ;
        RECT  4.89 32.5075 10.345 32.5725 ;
        RECT  4.89 35.1975 10.345 35.2625 ;
        RECT  4.89 37.8875 10.345 37.9525 ;
        RECT  4.89 40.5775 10.345 40.6425 ;
        RECT  0.0 20.4025 12.3 20.4675 ;
        RECT  0.0 23.0925 12.3 23.1575 ;
        RECT  0.0 25.7825 12.3 25.8475 ;
        RECT  0.0 28.4725 12.3 28.5375 ;
        RECT  0.0 31.1625 12.3 31.2275 ;
        RECT  0.0 33.8525 12.3 33.9175 ;
        RECT  0.0 36.5425 12.3 36.6075 ;
        RECT  0.0 39.2325 12.3 39.2975 ;
        RECT  6.92 8.5025 7.2625 8.5675 ;
        RECT  6.645 9.8475 7.4675 9.9125 ;
        RECT  6.92 13.8825 7.6725 13.9475 ;
        RECT  6.645 15.2275 7.8775 15.2925 ;
        RECT  6.92 8.2975 7.0575 8.3625 ;
        RECT  6.92 10.9875 7.0575 11.0525 ;
        RECT  6.92 13.6775 7.0575 13.7425 ;
        RECT  6.92 16.3675 7.0575 16.4325 ;
        RECT  0.0 9.6425 6.92 9.7075 ;
        RECT  0.0 12.3325 6.92 12.3975 ;
        RECT  0.0 15.0225 6.92 15.0875 ;
        RECT  0.0 17.7125 6.92 17.7775 ;
        RECT  6.92 7.535 7.2625 7.6 ;
        RECT  6.92 6.83 7.4675 6.895 ;
        RECT  6.92 6.125 7.6725 6.19 ;
        RECT  6.92 5.42 7.8775 5.485 ;
        RECT  6.92 7.8875 8.3875 7.9525 ;
        RECT  6.92 7.1825 8.3875 7.2475 ;
        RECT  6.92 6.4775 8.3875 6.5425 ;
        RECT  6.92 5.7725 8.3875 5.8375 ;
        RECT  6.92 5.0675 8.3875 5.1325 ;
        RECT  3.69 4.8625 3.755 4.9275 ;
        RECT  3.69 4.895 3.755 5.1 ;
        RECT  0.0 4.8625 3.7225 4.9275 ;
        RECT  6.65 4.8625 6.715 4.9275 ;
        RECT  6.65 4.895 6.715 5.1 ;
        RECT  0.0 4.8625 6.6825 4.9275 ;
        RECT  1.7 4.8625 1.765 4.9275 ;
        RECT  1.7 4.895 1.765 5.1 ;
        RECT  0.0 4.8625 1.7325 4.9275 ;
        RECT  4.66 4.8625 4.725 4.9275 ;
        RECT  4.66 4.895 4.725 5.1 ;
        RECT  0.0 4.8625 4.6925 4.9275 ;
        RECT  9.4575 3.795 10.345 3.86 ;
        RECT  9.0475 1.61 10.345 1.675 ;
        RECT  9.2525 3.1575 10.345 3.2225 ;
        RECT  9.4575 41.4775 10.345 41.5425 ;
        RECT  9.6625 10.2975 10.345 10.3625 ;
        RECT  9.8675 14.3225 10.345 14.3875 ;
        RECT  0.685 8.0925 0.75 8.1575 ;
        RECT  0.685 7.92 0.75 8.125 ;
        RECT  0.7175 8.0925 8.8425 8.1575 ;
        RECT  4.665 40.7825 8.9075 40.8475 ;
        RECT  10.345 42.205 11.95 42.27 ;
        RECT  10.345 18.895 11.95 18.96 ;
        RECT  10.345 10.4275 11.95 10.4925 ;
        RECT  10.345 6.8 11.95 6.865 ;
        RECT  10.345 9.76 11.95 9.825 ;
        RECT  10.345 4.81 11.95 4.875 ;
        RECT  10.345 7.77 11.95 7.835 ;
        RECT  10.345 1.74 11.95 1.805 ;
        RECT  8.6025 3.0275 10.345 3.0925 ;
        RECT  8.6025 14.4525 10.345 14.5175 ;
        RECT  8.6025 3.955 10.345 4.02 ;
        RECT  8.6025 11.23 10.345 11.295 ;
        RECT  11.95 0.0 12.3 42.27 ;
        RECT  0.0 0.0 0.35 42.27 ;
        RECT  10.255 24.5775 11.845 24.6425 ;
        RECT  10.255 19.1975 11.845 19.2625 ;
        RECT  10.255 21.8875 11.845 21.9525 ;
        RECT  10.255 40.4375 11.845 40.5025 ;
        RECT  10.255 29.9575 11.845 30.0225 ;
        RECT  10.255 27.2675 11.845 27.3325 ;
        RECT  10.255 37.7475 11.845 37.8125 ;
        RECT  10.255 35.0575 11.845 35.1225 ;
        RECT  10.255 24.2975 11.845 24.3625 ;
        RECT  10.255 26.9875 11.845 27.0525 ;
        RECT  10.255 21.6075 11.845 21.6725 ;
        RECT  10.255 38.0275 11.845 38.0925 ;
        RECT  10.255 32.6475 11.845 32.7125 ;
        RECT  10.255 32.3675 11.845 32.4325 ;
        RECT  10.255 20.4025 11.845 20.4675 ;
        RECT  10.255 23.0925 11.845 23.1575 ;
        RECT  10.255 25.7825 11.845 25.8475 ;
        RECT  10.255 28.4725 11.845 28.5375 ;
        RECT  10.255 31.1625 11.845 31.2275 ;
        RECT  10.255 33.8525 11.845 33.9175 ;
        RECT  10.255 36.5425 11.845 36.6075 ;
        RECT  10.255 39.2325 11.845 39.2975 ;
        RECT  10.255 19.0575 11.845 19.1225 ;
        RECT  10.255 21.7475 11.845 21.8125 ;
        RECT  10.255 24.4375 11.845 24.5025 ;
        RECT  10.255 27.1275 11.845 27.1925 ;
        RECT  10.255 29.8175 11.845 29.8825 ;
        RECT  10.255 32.5075 11.845 32.5725 ;
        RECT  10.255 35.1975 11.845 35.2625 ;
        RECT  10.255 37.8875 11.845 37.9525 ;
        RECT  10.255 40.5775 11.845 40.6425 ;
        RECT  10.255 35.3375 11.845 35.4025 ;
        RECT  10.255 29.6775 11.845 29.7425 ;
        RECT  11.015 20.2025 11.08 20.3375 ;
        RECT  10.83 20.2025 10.895 20.3375 ;
        RECT  10.315 20.2025 10.38 20.3375 ;
        RECT  10.5 20.2025 10.565 20.3375 ;
        RECT  10.83 19.7375 10.895 19.8725 ;
        RECT  11.015 19.7375 11.08 19.8725 ;
        RECT  10.5 19.7375 10.565 19.8725 ;
        RECT  10.315 19.7375 10.38 19.8725 ;
        RECT  10.935 19.3475 11.0 19.4825 ;
        RECT  10.75 19.3475 10.815 19.4825 ;
        RECT  10.58 19.3475 10.645 19.4825 ;
        RECT  10.395 19.3475 10.46 19.4825 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  10.625 20.4025 10.76 20.4675 ;
        RECT  10.2775 19.0575 10.4125 19.1225 ;
        RECT  10.9825 19.0575 11.1175 19.1225 ;
        RECT  10.6125 19.1975 10.7475 19.2625 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  10.5175 20.0875 10.6525 20.1525 ;
        RECT  10.5175 20.0875 10.6525 20.1525 ;
        RECT  10.7425 19.9375 10.8775 20.0025 ;
        RECT  10.7425 19.9375 10.8775 20.0025 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  10.5675 19.3475 10.6325 19.4825 ;
        RECT  10.3125 19.84 10.3775 19.975 ;
        RECT  10.3125 19.84 10.3775 19.975 ;
        RECT  10.3125 19.84 10.3775 19.975 ;
        RECT  10.3125 19.84 10.3775 19.975 ;
        RECT  10.3125 19.84 10.3775 19.975 ;
        RECT  10.3125 19.84 10.3775 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  10.7625 19.3475 10.8275 19.4825 ;
        RECT  10.63 19.0575 10.765 19.1225 ;
        RECT  10.63 19.0575 10.765 19.1225 ;
        RECT  10.9825 19.0575 11.1175 19.1225 ;
        RECT  10.625 20.4025 10.76 20.4675 ;
        RECT  10.9825 19.0575 11.1175 19.1225 ;
        RECT  10.9825 19.0575 11.1175 19.1225 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  10.2775 19.0575 10.4125 19.1225 ;
        RECT  10.6375 20.4025 10.7375 20.465 ;
        RECT  10.6375 20.405 10.7375 20.4675 ;
        RECT  10.965 19.2 11.0175 19.2625 ;
        RECT  10.6375 20.4025 10.7375 20.465 ;
        RECT  11.015 20.2025 11.085 20.4025 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  10.255 19.0575 11.14 19.1225 ;
        RECT  10.83 19.5725 11.005 19.6375 ;
        RECT  10.31 19.7375 10.38 19.8725 ;
        RECT  10.5 19.5725 10.565 20.3125 ;
        RECT  10.6375 20.405 10.7375 20.4675 ;
        RECT  10.26 19.2 10.3125 19.2625 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  10.255 20.4025 11.14 20.4675 ;
        RECT  10.83 19.5725 10.895 20.2025 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  10.395 19.3475 10.465 19.6375 ;
        RECT  10.31 19.7375 10.38 19.8725 ;
        RECT  10.255 19.1975 11.14 19.2625 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  11.015 20.2025 11.085 20.4025 ;
        RECT  10.31 20.2025 10.38 20.4025 ;
        RECT  10.935 19.3475 11.005 19.6375 ;
        RECT  10.395 19.5725 10.565 19.6375 ;
        RECT  10.255 19.1975 11.14 19.2625 ;
        RECT  10.255 19.0575 11.14 19.1225 ;
        RECT  10.255 20.4025 11.14 20.4675 ;
        RECT  11.015 20.5325 11.08 20.6675 ;
        RECT  10.83 20.5325 10.895 20.6675 ;
        RECT  10.315 20.5325 10.38 20.6675 ;
        RECT  10.5 20.5325 10.565 20.6675 ;
        RECT  10.83 20.9975 10.895 21.1325 ;
        RECT  11.015 20.9975 11.08 21.1325 ;
        RECT  10.5 20.9975 10.565 21.1325 ;
        RECT  10.315 20.9975 10.38 21.1325 ;
        RECT  10.935 21.3875 11.0 21.5225 ;
        RECT  10.75 21.3875 10.815 21.5225 ;
        RECT  10.58 21.3875 10.645 21.5225 ;
        RECT  10.395 21.3875 10.46 21.5225 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  10.625 20.4025 10.76 20.4675 ;
        RECT  10.2775 21.7475 10.4125 21.8125 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  10.6125 21.6075 10.7475 21.6725 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  10.5175 20.7175 10.6525 20.7825 ;
        RECT  10.5175 20.7175 10.6525 20.7825 ;
        RECT  10.7425 20.8675 10.8775 20.9325 ;
        RECT  10.7425 20.8675 10.8775 20.9325 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  10.5675 21.3875 10.6325 21.5225 ;
        RECT  10.3125 20.895 10.3775 21.03 ;
        RECT  10.3125 20.895 10.3775 21.03 ;
        RECT  10.3125 20.895 10.3775 21.03 ;
        RECT  10.3125 20.895 10.3775 21.03 ;
        RECT  10.3125 20.895 10.3775 21.03 ;
        RECT  10.3125 20.895 10.3775 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  10.7625 21.3875 10.8275 21.5225 ;
        RECT  10.63 21.7475 10.765 21.8125 ;
        RECT  10.63 21.7475 10.765 21.8125 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  10.625 20.4025 10.76 20.4675 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  10.2775 21.7475 10.4125 21.8125 ;
        RECT  10.6375 20.405 10.7375 20.4675 ;
        RECT  10.6375 20.4025 10.7375 20.465 ;
        RECT  10.965 21.6075 11.0175 21.67 ;
        RECT  10.6375 20.405 10.7375 20.4675 ;
        RECT  11.015 20.4675 11.085 20.6675 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  10.255 21.7475 11.14 21.8125 ;
        RECT  10.83 21.2325 11.005 21.2975 ;
        RECT  10.31 20.9975 10.38 21.1325 ;
        RECT  10.5 20.5575 10.565 21.2975 ;
        RECT  10.6375 20.4025 10.7375 20.465 ;
        RECT  10.26 21.6075 10.3125 21.67 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  10.255 20.4025 11.14 20.4675 ;
        RECT  10.83 20.6675 10.895 21.2975 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  10.395 21.2325 10.465 21.5225 ;
        RECT  10.31 20.9975 10.38 21.1325 ;
        RECT  10.255 21.6075 11.14 21.6725 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  11.015 20.4675 11.085 20.6675 ;
        RECT  10.31 20.4675 10.38 20.6675 ;
        RECT  10.935 21.2325 11.005 21.5225 ;
        RECT  10.395 21.2325 10.565 21.2975 ;
        RECT  10.255 21.6075 11.14 21.6725 ;
        RECT  10.255 21.7475 11.14 21.8125 ;
        RECT  10.255 20.4025 11.14 20.4675 ;
        RECT  11.015 22.8925 11.08 23.0275 ;
        RECT  10.83 22.8925 10.895 23.0275 ;
        RECT  10.315 22.8925 10.38 23.0275 ;
        RECT  10.5 22.8925 10.565 23.0275 ;
        RECT  10.83 22.4275 10.895 22.5625 ;
        RECT  11.015 22.4275 11.08 22.5625 ;
        RECT  10.5 22.4275 10.565 22.5625 ;
        RECT  10.315 22.4275 10.38 22.5625 ;
        RECT  10.935 22.0375 11.0 22.1725 ;
        RECT  10.75 22.0375 10.815 22.1725 ;
        RECT  10.58 22.0375 10.645 22.1725 ;
        RECT  10.395 22.0375 10.46 22.1725 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  10.625 23.0925 10.76 23.1575 ;
        RECT  10.2775 21.7475 10.4125 21.8125 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  10.6125 21.8875 10.7475 21.9525 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  10.5175 22.7775 10.6525 22.8425 ;
        RECT  10.5175 22.7775 10.6525 22.8425 ;
        RECT  10.7425 22.6275 10.8775 22.6925 ;
        RECT  10.7425 22.6275 10.8775 22.6925 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  10.5675 22.0375 10.6325 22.1725 ;
        RECT  10.3125 22.53 10.3775 22.665 ;
        RECT  10.3125 22.53 10.3775 22.665 ;
        RECT  10.3125 22.53 10.3775 22.665 ;
        RECT  10.3125 22.53 10.3775 22.665 ;
        RECT  10.3125 22.53 10.3775 22.665 ;
        RECT  10.3125 22.53 10.3775 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  10.7625 22.0375 10.8275 22.1725 ;
        RECT  10.63 21.7475 10.765 21.8125 ;
        RECT  10.63 21.7475 10.765 21.8125 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  10.625 23.0925 10.76 23.1575 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  10.2775 21.7475 10.4125 21.8125 ;
        RECT  10.6375 23.0925 10.7375 23.155 ;
        RECT  10.6375 23.095 10.7375 23.1575 ;
        RECT  10.965 21.89 11.0175 21.9525 ;
        RECT  10.6375 23.0925 10.7375 23.155 ;
        RECT  11.015 22.8925 11.085 23.0925 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  10.255 21.7475 11.14 21.8125 ;
        RECT  10.83 22.2625 11.005 22.3275 ;
        RECT  10.31 22.4275 10.38 22.5625 ;
        RECT  10.5 22.2625 10.565 23.0025 ;
        RECT  10.6375 23.095 10.7375 23.1575 ;
        RECT  10.26 21.89 10.3125 21.9525 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  10.255 23.0925 11.14 23.1575 ;
        RECT  10.83 22.2625 10.895 22.8925 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  10.395 22.0375 10.465 22.3275 ;
        RECT  10.31 22.4275 10.38 22.5625 ;
        RECT  10.255 21.8875 11.14 21.9525 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  11.015 22.8925 11.085 23.0925 ;
        RECT  10.31 22.8925 10.38 23.0925 ;
        RECT  10.935 22.0375 11.005 22.3275 ;
        RECT  10.395 22.2625 10.565 22.3275 ;
        RECT  10.255 21.8875 11.14 21.9525 ;
        RECT  10.255 21.7475 11.14 21.8125 ;
        RECT  10.255 23.0925 11.14 23.1575 ;
        RECT  11.015 23.2225 11.08 23.3575 ;
        RECT  10.83 23.2225 10.895 23.3575 ;
        RECT  10.315 23.2225 10.38 23.3575 ;
        RECT  10.5 23.2225 10.565 23.3575 ;
        RECT  10.83 23.6875 10.895 23.8225 ;
        RECT  11.015 23.6875 11.08 23.8225 ;
        RECT  10.5 23.6875 10.565 23.8225 ;
        RECT  10.315 23.6875 10.38 23.8225 ;
        RECT  10.935 24.0775 11.0 24.2125 ;
        RECT  10.75 24.0775 10.815 24.2125 ;
        RECT  10.58 24.0775 10.645 24.2125 ;
        RECT  10.395 24.0775 10.46 24.2125 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  10.625 23.0925 10.76 23.1575 ;
        RECT  10.2775 24.4375 10.4125 24.5025 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  10.6125 24.2975 10.7475 24.3625 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  10.5175 23.4075 10.6525 23.4725 ;
        RECT  10.5175 23.4075 10.6525 23.4725 ;
        RECT  10.7425 23.5575 10.8775 23.6225 ;
        RECT  10.7425 23.5575 10.8775 23.6225 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  10.5675 24.0775 10.6325 24.2125 ;
        RECT  10.3125 23.585 10.3775 23.72 ;
        RECT  10.3125 23.585 10.3775 23.72 ;
        RECT  10.3125 23.585 10.3775 23.72 ;
        RECT  10.3125 23.585 10.3775 23.72 ;
        RECT  10.3125 23.585 10.3775 23.72 ;
        RECT  10.3125 23.585 10.3775 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  10.7625 24.0775 10.8275 24.2125 ;
        RECT  10.63 24.4375 10.765 24.5025 ;
        RECT  10.63 24.4375 10.765 24.5025 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  10.625 23.0925 10.76 23.1575 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  10.2775 24.4375 10.4125 24.5025 ;
        RECT  10.6375 23.095 10.7375 23.1575 ;
        RECT  10.6375 23.0925 10.7375 23.155 ;
        RECT  10.965 24.2975 11.0175 24.36 ;
        RECT  10.6375 23.095 10.7375 23.1575 ;
        RECT  11.015 23.1575 11.085 23.3575 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  10.255 24.4375 11.14 24.5025 ;
        RECT  10.83 23.9225 11.005 23.9875 ;
        RECT  10.31 23.6875 10.38 23.8225 ;
        RECT  10.5 23.2475 10.565 23.9875 ;
        RECT  10.6375 23.0925 10.7375 23.155 ;
        RECT  10.26 24.2975 10.3125 24.36 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  10.255 23.0925 11.14 23.1575 ;
        RECT  10.83 23.3575 10.895 23.9875 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  10.395 23.9225 10.465 24.2125 ;
        RECT  10.31 23.6875 10.38 23.8225 ;
        RECT  10.255 24.2975 11.14 24.3625 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  11.015 23.1575 11.085 23.3575 ;
        RECT  10.31 23.1575 10.38 23.3575 ;
        RECT  10.935 23.9225 11.005 24.2125 ;
        RECT  10.395 23.9225 10.565 23.9875 ;
        RECT  10.255 24.2975 11.14 24.3625 ;
        RECT  10.255 24.4375 11.14 24.5025 ;
        RECT  10.255 23.0925 11.14 23.1575 ;
        RECT  11.015 25.5825 11.08 25.7175 ;
        RECT  10.83 25.5825 10.895 25.7175 ;
        RECT  10.315 25.5825 10.38 25.7175 ;
        RECT  10.5 25.5825 10.565 25.7175 ;
        RECT  10.83 25.1175 10.895 25.2525 ;
        RECT  11.015 25.1175 11.08 25.2525 ;
        RECT  10.5 25.1175 10.565 25.2525 ;
        RECT  10.315 25.1175 10.38 25.2525 ;
        RECT  10.935 24.7275 11.0 24.8625 ;
        RECT  10.75 24.7275 10.815 24.8625 ;
        RECT  10.58 24.7275 10.645 24.8625 ;
        RECT  10.395 24.7275 10.46 24.8625 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  10.625 25.7825 10.76 25.8475 ;
        RECT  10.2775 24.4375 10.4125 24.5025 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  10.6125 24.5775 10.7475 24.6425 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  10.5175 25.4675 10.6525 25.5325 ;
        RECT  10.5175 25.4675 10.6525 25.5325 ;
        RECT  10.7425 25.3175 10.8775 25.3825 ;
        RECT  10.7425 25.3175 10.8775 25.3825 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  10.5675 24.7275 10.6325 24.8625 ;
        RECT  10.3125 25.22 10.3775 25.355 ;
        RECT  10.3125 25.22 10.3775 25.355 ;
        RECT  10.3125 25.22 10.3775 25.355 ;
        RECT  10.3125 25.22 10.3775 25.355 ;
        RECT  10.3125 25.22 10.3775 25.355 ;
        RECT  10.3125 25.22 10.3775 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  10.7625 24.7275 10.8275 24.8625 ;
        RECT  10.63 24.4375 10.765 24.5025 ;
        RECT  10.63 24.4375 10.765 24.5025 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  10.625 25.7825 10.76 25.8475 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  10.2775 24.4375 10.4125 24.5025 ;
        RECT  10.6375 25.7825 10.7375 25.845 ;
        RECT  10.6375 25.785 10.7375 25.8475 ;
        RECT  10.965 24.58 11.0175 24.6425 ;
        RECT  10.6375 25.7825 10.7375 25.845 ;
        RECT  11.015 25.5825 11.085 25.7825 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  10.255 24.4375 11.14 24.5025 ;
        RECT  10.83 24.9525 11.005 25.0175 ;
        RECT  10.31 25.1175 10.38 25.2525 ;
        RECT  10.5 24.9525 10.565 25.6925 ;
        RECT  10.6375 25.785 10.7375 25.8475 ;
        RECT  10.26 24.58 10.3125 24.6425 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  10.255 25.7825 11.14 25.8475 ;
        RECT  10.83 24.9525 10.895 25.5825 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  10.395 24.7275 10.465 25.0175 ;
        RECT  10.31 25.1175 10.38 25.2525 ;
        RECT  10.255 24.5775 11.14 24.6425 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  11.015 25.5825 11.085 25.7825 ;
        RECT  10.31 25.5825 10.38 25.7825 ;
        RECT  10.935 24.7275 11.005 25.0175 ;
        RECT  10.395 24.9525 10.565 25.0175 ;
        RECT  10.255 24.5775 11.14 24.6425 ;
        RECT  10.255 24.4375 11.14 24.5025 ;
        RECT  10.255 25.7825 11.14 25.8475 ;
        RECT  11.015 25.9125 11.08 26.0475 ;
        RECT  10.83 25.9125 10.895 26.0475 ;
        RECT  10.315 25.9125 10.38 26.0475 ;
        RECT  10.5 25.9125 10.565 26.0475 ;
        RECT  10.83 26.3775 10.895 26.5125 ;
        RECT  11.015 26.3775 11.08 26.5125 ;
        RECT  10.5 26.3775 10.565 26.5125 ;
        RECT  10.315 26.3775 10.38 26.5125 ;
        RECT  10.935 26.7675 11.0 26.9025 ;
        RECT  10.75 26.7675 10.815 26.9025 ;
        RECT  10.58 26.7675 10.645 26.9025 ;
        RECT  10.395 26.7675 10.46 26.9025 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  10.625 25.7825 10.76 25.8475 ;
        RECT  10.2775 27.1275 10.4125 27.1925 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  10.6125 26.9875 10.7475 27.0525 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  10.5175 26.0975 10.6525 26.1625 ;
        RECT  10.5175 26.0975 10.6525 26.1625 ;
        RECT  10.7425 26.2475 10.8775 26.3125 ;
        RECT  10.7425 26.2475 10.8775 26.3125 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  10.5675 26.7675 10.6325 26.9025 ;
        RECT  10.3125 26.275 10.3775 26.41 ;
        RECT  10.3125 26.275 10.3775 26.41 ;
        RECT  10.3125 26.275 10.3775 26.41 ;
        RECT  10.3125 26.275 10.3775 26.41 ;
        RECT  10.3125 26.275 10.3775 26.41 ;
        RECT  10.3125 26.275 10.3775 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  10.7625 26.7675 10.8275 26.9025 ;
        RECT  10.63 27.1275 10.765 27.1925 ;
        RECT  10.63 27.1275 10.765 27.1925 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  10.625 25.7825 10.76 25.8475 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  10.2775 27.1275 10.4125 27.1925 ;
        RECT  10.6375 25.785 10.7375 25.8475 ;
        RECT  10.6375 25.7825 10.7375 25.845 ;
        RECT  10.965 26.9875 11.0175 27.05 ;
        RECT  10.6375 25.785 10.7375 25.8475 ;
        RECT  11.015 25.8475 11.085 26.0475 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  10.255 27.1275 11.14 27.1925 ;
        RECT  10.83 26.6125 11.005 26.6775 ;
        RECT  10.31 26.3775 10.38 26.5125 ;
        RECT  10.5 25.9375 10.565 26.6775 ;
        RECT  10.6375 25.7825 10.7375 25.845 ;
        RECT  10.26 26.9875 10.3125 27.05 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  10.255 25.7825 11.14 25.8475 ;
        RECT  10.83 26.0475 10.895 26.6775 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  10.395 26.6125 10.465 26.9025 ;
        RECT  10.31 26.3775 10.38 26.5125 ;
        RECT  10.255 26.9875 11.14 27.0525 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  11.015 25.8475 11.085 26.0475 ;
        RECT  10.31 25.8475 10.38 26.0475 ;
        RECT  10.935 26.6125 11.005 26.9025 ;
        RECT  10.395 26.6125 10.565 26.6775 ;
        RECT  10.255 26.9875 11.14 27.0525 ;
        RECT  10.255 27.1275 11.14 27.1925 ;
        RECT  10.255 25.7825 11.14 25.8475 ;
        RECT  11.015 28.2725 11.08 28.4075 ;
        RECT  10.83 28.2725 10.895 28.4075 ;
        RECT  10.315 28.2725 10.38 28.4075 ;
        RECT  10.5 28.2725 10.565 28.4075 ;
        RECT  10.83 27.8075 10.895 27.9425 ;
        RECT  11.015 27.8075 11.08 27.9425 ;
        RECT  10.5 27.8075 10.565 27.9425 ;
        RECT  10.315 27.8075 10.38 27.9425 ;
        RECT  10.935 27.4175 11.0 27.5525 ;
        RECT  10.75 27.4175 10.815 27.5525 ;
        RECT  10.58 27.4175 10.645 27.5525 ;
        RECT  10.395 27.4175 10.46 27.5525 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  10.625 28.4725 10.76 28.5375 ;
        RECT  10.2775 27.1275 10.4125 27.1925 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  10.6125 27.2675 10.7475 27.3325 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  10.5175 28.1575 10.6525 28.2225 ;
        RECT  10.5175 28.1575 10.6525 28.2225 ;
        RECT  10.7425 28.0075 10.8775 28.0725 ;
        RECT  10.7425 28.0075 10.8775 28.0725 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  10.5675 27.4175 10.6325 27.5525 ;
        RECT  10.3125 27.91 10.3775 28.045 ;
        RECT  10.3125 27.91 10.3775 28.045 ;
        RECT  10.3125 27.91 10.3775 28.045 ;
        RECT  10.3125 27.91 10.3775 28.045 ;
        RECT  10.3125 27.91 10.3775 28.045 ;
        RECT  10.3125 27.91 10.3775 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  10.7625 27.4175 10.8275 27.5525 ;
        RECT  10.63 27.1275 10.765 27.1925 ;
        RECT  10.63 27.1275 10.765 27.1925 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  10.625 28.4725 10.76 28.5375 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  10.2775 27.1275 10.4125 27.1925 ;
        RECT  10.6375 28.4725 10.7375 28.535 ;
        RECT  10.6375 28.475 10.7375 28.5375 ;
        RECT  10.965 27.27 11.0175 27.3325 ;
        RECT  10.6375 28.4725 10.7375 28.535 ;
        RECT  11.015 28.2725 11.085 28.4725 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  10.255 27.1275 11.14 27.1925 ;
        RECT  10.83 27.6425 11.005 27.7075 ;
        RECT  10.31 27.8075 10.38 27.9425 ;
        RECT  10.5 27.6425 10.565 28.3825 ;
        RECT  10.6375 28.475 10.7375 28.5375 ;
        RECT  10.26 27.27 10.3125 27.3325 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  10.255 28.4725 11.14 28.5375 ;
        RECT  10.83 27.6425 10.895 28.2725 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  10.395 27.4175 10.465 27.7075 ;
        RECT  10.31 27.8075 10.38 27.9425 ;
        RECT  10.255 27.2675 11.14 27.3325 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  11.015 28.2725 11.085 28.4725 ;
        RECT  10.31 28.2725 10.38 28.4725 ;
        RECT  10.935 27.4175 11.005 27.7075 ;
        RECT  10.395 27.6425 10.565 27.7075 ;
        RECT  10.255 27.2675 11.14 27.3325 ;
        RECT  10.255 27.1275 11.14 27.1925 ;
        RECT  10.255 28.4725 11.14 28.5375 ;
        RECT  11.015 28.6025 11.08 28.7375 ;
        RECT  10.83 28.6025 10.895 28.7375 ;
        RECT  10.315 28.6025 10.38 28.7375 ;
        RECT  10.5 28.6025 10.565 28.7375 ;
        RECT  10.83 29.0675 10.895 29.2025 ;
        RECT  11.015 29.0675 11.08 29.2025 ;
        RECT  10.5 29.0675 10.565 29.2025 ;
        RECT  10.315 29.0675 10.38 29.2025 ;
        RECT  10.935 29.4575 11.0 29.5925 ;
        RECT  10.75 29.4575 10.815 29.5925 ;
        RECT  10.58 29.4575 10.645 29.5925 ;
        RECT  10.395 29.4575 10.46 29.5925 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  10.625 28.4725 10.76 28.5375 ;
        RECT  10.2775 29.8175 10.4125 29.8825 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  10.6125 29.6775 10.7475 29.7425 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  10.5175 28.7875 10.6525 28.8525 ;
        RECT  10.5175 28.7875 10.6525 28.8525 ;
        RECT  10.7425 28.9375 10.8775 29.0025 ;
        RECT  10.7425 28.9375 10.8775 29.0025 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  10.5675 29.4575 10.6325 29.5925 ;
        RECT  10.3125 28.965 10.3775 29.1 ;
        RECT  10.3125 28.965 10.3775 29.1 ;
        RECT  10.3125 28.965 10.3775 29.1 ;
        RECT  10.3125 28.965 10.3775 29.1 ;
        RECT  10.3125 28.965 10.3775 29.1 ;
        RECT  10.3125 28.965 10.3775 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  10.7625 29.4575 10.8275 29.5925 ;
        RECT  10.63 29.8175 10.765 29.8825 ;
        RECT  10.63 29.8175 10.765 29.8825 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  10.625 28.4725 10.76 28.5375 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  10.2775 29.8175 10.4125 29.8825 ;
        RECT  10.6375 28.475 10.7375 28.5375 ;
        RECT  10.6375 28.4725 10.7375 28.535 ;
        RECT  10.965 29.6775 11.0175 29.74 ;
        RECT  10.6375 28.475 10.7375 28.5375 ;
        RECT  11.015 28.5375 11.085 28.7375 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  10.255 29.8175 11.14 29.8825 ;
        RECT  10.83 29.3025 11.005 29.3675 ;
        RECT  10.31 29.0675 10.38 29.2025 ;
        RECT  10.5 28.6275 10.565 29.3675 ;
        RECT  10.6375 28.4725 10.7375 28.535 ;
        RECT  10.26 29.6775 10.3125 29.74 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  10.255 28.4725 11.14 28.5375 ;
        RECT  10.83 28.7375 10.895 29.3675 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  10.395 29.3025 10.465 29.5925 ;
        RECT  10.31 29.0675 10.38 29.2025 ;
        RECT  10.255 29.6775 11.14 29.7425 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  11.015 28.5375 11.085 28.7375 ;
        RECT  10.31 28.5375 10.38 28.7375 ;
        RECT  10.935 29.3025 11.005 29.5925 ;
        RECT  10.395 29.3025 10.565 29.3675 ;
        RECT  10.255 29.6775 11.14 29.7425 ;
        RECT  10.255 29.8175 11.14 29.8825 ;
        RECT  10.255 28.4725 11.14 28.5375 ;
        RECT  11.015 30.9625 11.08 31.0975 ;
        RECT  10.83 30.9625 10.895 31.0975 ;
        RECT  10.315 30.9625 10.38 31.0975 ;
        RECT  10.5 30.9625 10.565 31.0975 ;
        RECT  10.83 30.4975 10.895 30.6325 ;
        RECT  11.015 30.4975 11.08 30.6325 ;
        RECT  10.5 30.4975 10.565 30.6325 ;
        RECT  10.315 30.4975 10.38 30.6325 ;
        RECT  10.935 30.1075 11.0 30.2425 ;
        RECT  10.75 30.1075 10.815 30.2425 ;
        RECT  10.58 30.1075 10.645 30.2425 ;
        RECT  10.395 30.1075 10.46 30.2425 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  10.625 31.1625 10.76 31.2275 ;
        RECT  10.2775 29.8175 10.4125 29.8825 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  10.6125 29.9575 10.7475 30.0225 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  10.5175 30.8475 10.6525 30.9125 ;
        RECT  10.5175 30.8475 10.6525 30.9125 ;
        RECT  10.7425 30.6975 10.8775 30.7625 ;
        RECT  10.7425 30.6975 10.8775 30.7625 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  10.5675 30.1075 10.6325 30.2425 ;
        RECT  10.3125 30.6 10.3775 30.735 ;
        RECT  10.3125 30.6 10.3775 30.735 ;
        RECT  10.3125 30.6 10.3775 30.735 ;
        RECT  10.3125 30.6 10.3775 30.735 ;
        RECT  10.3125 30.6 10.3775 30.735 ;
        RECT  10.3125 30.6 10.3775 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  10.7625 30.1075 10.8275 30.2425 ;
        RECT  10.63 29.8175 10.765 29.8825 ;
        RECT  10.63 29.8175 10.765 29.8825 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  10.625 31.1625 10.76 31.2275 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  10.2775 29.8175 10.4125 29.8825 ;
        RECT  10.6375 31.1625 10.7375 31.225 ;
        RECT  10.6375 31.165 10.7375 31.2275 ;
        RECT  10.965 29.96 11.0175 30.0225 ;
        RECT  10.6375 31.1625 10.7375 31.225 ;
        RECT  11.015 30.9625 11.085 31.1625 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  10.255 29.8175 11.14 29.8825 ;
        RECT  10.83 30.3325 11.005 30.3975 ;
        RECT  10.31 30.4975 10.38 30.6325 ;
        RECT  10.5 30.3325 10.565 31.0725 ;
        RECT  10.6375 31.165 10.7375 31.2275 ;
        RECT  10.26 29.96 10.3125 30.0225 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  10.255 31.1625 11.14 31.2275 ;
        RECT  10.83 30.3325 10.895 30.9625 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  10.395 30.1075 10.465 30.3975 ;
        RECT  10.31 30.4975 10.38 30.6325 ;
        RECT  10.255 29.9575 11.14 30.0225 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  11.015 30.9625 11.085 31.1625 ;
        RECT  10.31 30.9625 10.38 31.1625 ;
        RECT  10.935 30.1075 11.005 30.3975 ;
        RECT  10.395 30.3325 10.565 30.3975 ;
        RECT  10.255 29.9575 11.14 30.0225 ;
        RECT  10.255 29.8175 11.14 29.8825 ;
        RECT  10.255 31.1625 11.14 31.2275 ;
        RECT  11.015 31.2925 11.08 31.4275 ;
        RECT  10.83 31.2925 10.895 31.4275 ;
        RECT  10.315 31.2925 10.38 31.4275 ;
        RECT  10.5 31.2925 10.565 31.4275 ;
        RECT  10.83 31.7575 10.895 31.8925 ;
        RECT  11.015 31.7575 11.08 31.8925 ;
        RECT  10.5 31.7575 10.565 31.8925 ;
        RECT  10.315 31.7575 10.38 31.8925 ;
        RECT  10.935 32.1475 11.0 32.2825 ;
        RECT  10.75 32.1475 10.815 32.2825 ;
        RECT  10.58 32.1475 10.645 32.2825 ;
        RECT  10.395 32.1475 10.46 32.2825 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  10.625 31.1625 10.76 31.2275 ;
        RECT  10.2775 32.5075 10.4125 32.5725 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  10.6125 32.3675 10.7475 32.4325 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  10.5175 31.4775 10.6525 31.5425 ;
        RECT  10.5175 31.4775 10.6525 31.5425 ;
        RECT  10.7425 31.6275 10.8775 31.6925 ;
        RECT  10.7425 31.6275 10.8775 31.6925 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  10.5675 32.1475 10.6325 32.2825 ;
        RECT  10.3125 31.655 10.3775 31.79 ;
        RECT  10.3125 31.655 10.3775 31.79 ;
        RECT  10.3125 31.655 10.3775 31.79 ;
        RECT  10.3125 31.655 10.3775 31.79 ;
        RECT  10.3125 31.655 10.3775 31.79 ;
        RECT  10.3125 31.655 10.3775 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  10.7625 32.1475 10.8275 32.2825 ;
        RECT  10.63 32.5075 10.765 32.5725 ;
        RECT  10.63 32.5075 10.765 32.5725 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  10.625 31.1625 10.76 31.2275 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  10.2775 32.5075 10.4125 32.5725 ;
        RECT  10.6375 31.165 10.7375 31.2275 ;
        RECT  10.6375 31.1625 10.7375 31.225 ;
        RECT  10.965 32.3675 11.0175 32.43 ;
        RECT  10.6375 31.165 10.7375 31.2275 ;
        RECT  11.015 31.2275 11.085 31.4275 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  10.255 32.5075 11.14 32.5725 ;
        RECT  10.83 31.9925 11.005 32.0575 ;
        RECT  10.31 31.7575 10.38 31.8925 ;
        RECT  10.5 31.3175 10.565 32.0575 ;
        RECT  10.6375 31.1625 10.7375 31.225 ;
        RECT  10.26 32.3675 10.3125 32.43 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  10.255 31.1625 11.14 31.2275 ;
        RECT  10.83 31.4275 10.895 32.0575 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  10.395 31.9925 10.465 32.2825 ;
        RECT  10.31 31.7575 10.38 31.8925 ;
        RECT  10.255 32.3675 11.14 32.4325 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  11.015 31.2275 11.085 31.4275 ;
        RECT  10.31 31.2275 10.38 31.4275 ;
        RECT  10.935 31.9925 11.005 32.2825 ;
        RECT  10.395 31.9925 10.565 32.0575 ;
        RECT  10.255 32.3675 11.14 32.4325 ;
        RECT  10.255 32.5075 11.14 32.5725 ;
        RECT  10.255 31.1625 11.14 31.2275 ;
        RECT  11.015 33.6525 11.08 33.7875 ;
        RECT  10.83 33.6525 10.895 33.7875 ;
        RECT  10.315 33.6525 10.38 33.7875 ;
        RECT  10.5 33.6525 10.565 33.7875 ;
        RECT  10.83 33.1875 10.895 33.3225 ;
        RECT  11.015 33.1875 11.08 33.3225 ;
        RECT  10.5 33.1875 10.565 33.3225 ;
        RECT  10.315 33.1875 10.38 33.3225 ;
        RECT  10.935 32.7975 11.0 32.9325 ;
        RECT  10.75 32.7975 10.815 32.9325 ;
        RECT  10.58 32.7975 10.645 32.9325 ;
        RECT  10.395 32.7975 10.46 32.9325 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  10.625 33.8525 10.76 33.9175 ;
        RECT  10.2775 32.5075 10.4125 32.5725 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  10.6125 32.6475 10.7475 32.7125 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  10.5175 33.5375 10.6525 33.6025 ;
        RECT  10.5175 33.5375 10.6525 33.6025 ;
        RECT  10.7425 33.3875 10.8775 33.4525 ;
        RECT  10.7425 33.3875 10.8775 33.4525 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  10.5675 32.7975 10.6325 32.9325 ;
        RECT  10.3125 33.29 10.3775 33.425 ;
        RECT  10.3125 33.29 10.3775 33.425 ;
        RECT  10.3125 33.29 10.3775 33.425 ;
        RECT  10.3125 33.29 10.3775 33.425 ;
        RECT  10.3125 33.29 10.3775 33.425 ;
        RECT  10.3125 33.29 10.3775 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  10.7625 32.7975 10.8275 32.9325 ;
        RECT  10.63 32.5075 10.765 32.5725 ;
        RECT  10.63 32.5075 10.765 32.5725 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  10.625 33.8525 10.76 33.9175 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  10.2775 32.5075 10.4125 32.5725 ;
        RECT  10.6375 33.8525 10.7375 33.915 ;
        RECT  10.6375 33.855 10.7375 33.9175 ;
        RECT  10.965 32.65 11.0175 32.7125 ;
        RECT  10.6375 33.8525 10.7375 33.915 ;
        RECT  11.015 33.6525 11.085 33.8525 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  10.255 32.5075 11.14 32.5725 ;
        RECT  10.83 33.0225 11.005 33.0875 ;
        RECT  10.31 33.1875 10.38 33.3225 ;
        RECT  10.5 33.0225 10.565 33.7625 ;
        RECT  10.6375 33.855 10.7375 33.9175 ;
        RECT  10.26 32.65 10.3125 32.7125 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  10.255 33.8525 11.14 33.9175 ;
        RECT  10.83 33.0225 10.895 33.6525 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  10.395 32.7975 10.465 33.0875 ;
        RECT  10.31 33.1875 10.38 33.3225 ;
        RECT  10.255 32.6475 11.14 32.7125 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  11.015 33.6525 11.085 33.8525 ;
        RECT  10.31 33.6525 10.38 33.8525 ;
        RECT  10.935 32.7975 11.005 33.0875 ;
        RECT  10.395 33.0225 10.565 33.0875 ;
        RECT  10.255 32.6475 11.14 32.7125 ;
        RECT  10.255 32.5075 11.14 32.5725 ;
        RECT  10.255 33.8525 11.14 33.9175 ;
        RECT  11.015 33.9825 11.08 34.1175 ;
        RECT  10.83 33.9825 10.895 34.1175 ;
        RECT  10.315 33.9825 10.38 34.1175 ;
        RECT  10.5 33.9825 10.565 34.1175 ;
        RECT  10.83 34.4475 10.895 34.5825 ;
        RECT  11.015 34.4475 11.08 34.5825 ;
        RECT  10.5 34.4475 10.565 34.5825 ;
        RECT  10.315 34.4475 10.38 34.5825 ;
        RECT  10.935 34.8375 11.0 34.9725 ;
        RECT  10.75 34.8375 10.815 34.9725 ;
        RECT  10.58 34.8375 10.645 34.9725 ;
        RECT  10.395 34.8375 10.46 34.9725 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  10.625 33.8525 10.76 33.9175 ;
        RECT  10.2775 35.1975 10.4125 35.2625 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  10.6125 35.0575 10.7475 35.1225 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  10.5175 34.1675 10.6525 34.2325 ;
        RECT  10.5175 34.1675 10.6525 34.2325 ;
        RECT  10.7425 34.3175 10.8775 34.3825 ;
        RECT  10.7425 34.3175 10.8775 34.3825 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  10.5675 34.8375 10.6325 34.9725 ;
        RECT  10.3125 34.345 10.3775 34.48 ;
        RECT  10.3125 34.345 10.3775 34.48 ;
        RECT  10.3125 34.345 10.3775 34.48 ;
        RECT  10.3125 34.345 10.3775 34.48 ;
        RECT  10.3125 34.345 10.3775 34.48 ;
        RECT  10.3125 34.345 10.3775 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  10.7625 34.8375 10.8275 34.9725 ;
        RECT  10.63 35.1975 10.765 35.2625 ;
        RECT  10.63 35.1975 10.765 35.2625 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  10.625 33.8525 10.76 33.9175 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  10.2775 35.1975 10.4125 35.2625 ;
        RECT  10.6375 33.855 10.7375 33.9175 ;
        RECT  10.6375 33.8525 10.7375 33.915 ;
        RECT  10.965 35.0575 11.0175 35.12 ;
        RECT  10.6375 33.855 10.7375 33.9175 ;
        RECT  11.015 33.9175 11.085 34.1175 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  10.255 35.1975 11.14 35.2625 ;
        RECT  10.83 34.6825 11.005 34.7475 ;
        RECT  10.31 34.4475 10.38 34.5825 ;
        RECT  10.5 34.0075 10.565 34.7475 ;
        RECT  10.6375 33.8525 10.7375 33.915 ;
        RECT  10.26 35.0575 10.3125 35.12 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  10.255 33.8525 11.14 33.9175 ;
        RECT  10.83 34.1175 10.895 34.7475 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  10.395 34.6825 10.465 34.9725 ;
        RECT  10.31 34.4475 10.38 34.5825 ;
        RECT  10.255 35.0575 11.14 35.1225 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  11.015 33.9175 11.085 34.1175 ;
        RECT  10.31 33.9175 10.38 34.1175 ;
        RECT  10.935 34.6825 11.005 34.9725 ;
        RECT  10.395 34.6825 10.565 34.7475 ;
        RECT  10.255 35.0575 11.14 35.1225 ;
        RECT  10.255 35.1975 11.14 35.2625 ;
        RECT  10.255 33.8525 11.14 33.9175 ;
        RECT  11.015 36.3425 11.08 36.4775 ;
        RECT  10.83 36.3425 10.895 36.4775 ;
        RECT  10.315 36.3425 10.38 36.4775 ;
        RECT  10.5 36.3425 10.565 36.4775 ;
        RECT  10.83 35.8775 10.895 36.0125 ;
        RECT  11.015 35.8775 11.08 36.0125 ;
        RECT  10.5 35.8775 10.565 36.0125 ;
        RECT  10.315 35.8775 10.38 36.0125 ;
        RECT  10.935 35.4875 11.0 35.6225 ;
        RECT  10.75 35.4875 10.815 35.6225 ;
        RECT  10.58 35.4875 10.645 35.6225 ;
        RECT  10.395 35.4875 10.46 35.6225 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  10.625 36.5425 10.76 36.6075 ;
        RECT  10.2775 35.1975 10.4125 35.2625 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  10.6125 35.3375 10.7475 35.4025 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  10.5175 36.2275 10.6525 36.2925 ;
        RECT  10.5175 36.2275 10.6525 36.2925 ;
        RECT  10.7425 36.0775 10.8775 36.1425 ;
        RECT  10.7425 36.0775 10.8775 36.1425 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  10.5675 35.4875 10.6325 35.6225 ;
        RECT  10.3125 35.98 10.3775 36.115 ;
        RECT  10.3125 35.98 10.3775 36.115 ;
        RECT  10.3125 35.98 10.3775 36.115 ;
        RECT  10.3125 35.98 10.3775 36.115 ;
        RECT  10.3125 35.98 10.3775 36.115 ;
        RECT  10.3125 35.98 10.3775 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  10.7625 35.4875 10.8275 35.6225 ;
        RECT  10.63 35.1975 10.765 35.2625 ;
        RECT  10.63 35.1975 10.765 35.2625 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  10.625 36.5425 10.76 36.6075 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  10.2775 35.1975 10.4125 35.2625 ;
        RECT  10.6375 36.5425 10.7375 36.605 ;
        RECT  10.6375 36.545 10.7375 36.6075 ;
        RECT  10.965 35.34 11.0175 35.4025 ;
        RECT  10.6375 36.5425 10.7375 36.605 ;
        RECT  11.015 36.3425 11.085 36.5425 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  10.255 35.1975 11.14 35.2625 ;
        RECT  10.83 35.7125 11.005 35.7775 ;
        RECT  10.31 35.8775 10.38 36.0125 ;
        RECT  10.5 35.7125 10.565 36.4525 ;
        RECT  10.6375 36.545 10.7375 36.6075 ;
        RECT  10.26 35.34 10.3125 35.4025 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  10.255 36.5425 11.14 36.6075 ;
        RECT  10.83 35.7125 10.895 36.3425 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  10.395 35.4875 10.465 35.7775 ;
        RECT  10.31 35.8775 10.38 36.0125 ;
        RECT  10.255 35.3375 11.14 35.4025 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  11.015 36.3425 11.085 36.5425 ;
        RECT  10.31 36.3425 10.38 36.5425 ;
        RECT  10.935 35.4875 11.005 35.7775 ;
        RECT  10.395 35.7125 10.565 35.7775 ;
        RECT  10.255 35.3375 11.14 35.4025 ;
        RECT  10.255 35.1975 11.14 35.2625 ;
        RECT  10.255 36.5425 11.14 36.6075 ;
        RECT  11.015 36.6725 11.08 36.8075 ;
        RECT  10.83 36.6725 10.895 36.8075 ;
        RECT  10.315 36.6725 10.38 36.8075 ;
        RECT  10.5 36.6725 10.565 36.8075 ;
        RECT  10.83 37.1375 10.895 37.2725 ;
        RECT  11.015 37.1375 11.08 37.2725 ;
        RECT  10.5 37.1375 10.565 37.2725 ;
        RECT  10.315 37.1375 10.38 37.2725 ;
        RECT  10.935 37.5275 11.0 37.6625 ;
        RECT  10.75 37.5275 10.815 37.6625 ;
        RECT  10.58 37.5275 10.645 37.6625 ;
        RECT  10.395 37.5275 10.46 37.6625 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  10.625 36.5425 10.76 36.6075 ;
        RECT  10.2775 37.8875 10.4125 37.9525 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  10.6125 37.7475 10.7475 37.8125 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  10.5175 36.8575 10.6525 36.9225 ;
        RECT  10.5175 36.8575 10.6525 36.9225 ;
        RECT  10.7425 37.0075 10.8775 37.0725 ;
        RECT  10.7425 37.0075 10.8775 37.0725 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  10.5675 37.5275 10.6325 37.6625 ;
        RECT  10.3125 37.035 10.3775 37.17 ;
        RECT  10.3125 37.035 10.3775 37.17 ;
        RECT  10.3125 37.035 10.3775 37.17 ;
        RECT  10.3125 37.035 10.3775 37.17 ;
        RECT  10.3125 37.035 10.3775 37.17 ;
        RECT  10.3125 37.035 10.3775 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  10.7625 37.5275 10.8275 37.6625 ;
        RECT  10.63 37.8875 10.765 37.9525 ;
        RECT  10.63 37.8875 10.765 37.9525 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  10.625 36.5425 10.76 36.6075 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  10.2775 37.8875 10.4125 37.9525 ;
        RECT  10.6375 36.545 10.7375 36.6075 ;
        RECT  10.6375 36.5425 10.7375 36.605 ;
        RECT  10.965 37.7475 11.0175 37.81 ;
        RECT  10.6375 36.545 10.7375 36.6075 ;
        RECT  11.015 36.6075 11.085 36.8075 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  10.255 37.8875 11.14 37.9525 ;
        RECT  10.83 37.3725 11.005 37.4375 ;
        RECT  10.31 37.1375 10.38 37.2725 ;
        RECT  10.5 36.6975 10.565 37.4375 ;
        RECT  10.6375 36.5425 10.7375 36.605 ;
        RECT  10.26 37.7475 10.3125 37.81 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  10.255 36.5425 11.14 36.6075 ;
        RECT  10.83 36.8075 10.895 37.4375 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  10.395 37.3725 10.465 37.6625 ;
        RECT  10.31 37.1375 10.38 37.2725 ;
        RECT  10.255 37.7475 11.14 37.8125 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  11.015 36.6075 11.085 36.8075 ;
        RECT  10.31 36.6075 10.38 36.8075 ;
        RECT  10.935 37.3725 11.005 37.6625 ;
        RECT  10.395 37.3725 10.565 37.4375 ;
        RECT  10.255 37.7475 11.14 37.8125 ;
        RECT  10.255 37.8875 11.14 37.9525 ;
        RECT  10.255 36.5425 11.14 36.6075 ;
        RECT  11.015 39.0325 11.08 39.1675 ;
        RECT  10.83 39.0325 10.895 39.1675 ;
        RECT  10.315 39.0325 10.38 39.1675 ;
        RECT  10.5 39.0325 10.565 39.1675 ;
        RECT  10.83 38.5675 10.895 38.7025 ;
        RECT  11.015 38.5675 11.08 38.7025 ;
        RECT  10.5 38.5675 10.565 38.7025 ;
        RECT  10.315 38.5675 10.38 38.7025 ;
        RECT  10.935 38.1775 11.0 38.3125 ;
        RECT  10.75 38.1775 10.815 38.3125 ;
        RECT  10.58 38.1775 10.645 38.3125 ;
        RECT  10.395 38.1775 10.46 38.3125 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  10.625 39.2325 10.76 39.2975 ;
        RECT  10.2775 37.8875 10.4125 37.9525 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  10.6125 38.0275 10.7475 38.0925 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  10.5175 38.9175 10.6525 38.9825 ;
        RECT  10.5175 38.9175 10.6525 38.9825 ;
        RECT  10.7425 38.7675 10.8775 38.8325 ;
        RECT  10.7425 38.7675 10.8775 38.8325 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  10.5675 38.1775 10.6325 38.3125 ;
        RECT  10.3125 38.67 10.3775 38.805 ;
        RECT  10.3125 38.67 10.3775 38.805 ;
        RECT  10.3125 38.67 10.3775 38.805 ;
        RECT  10.3125 38.67 10.3775 38.805 ;
        RECT  10.3125 38.67 10.3775 38.805 ;
        RECT  10.3125 38.67 10.3775 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  10.7625 38.1775 10.8275 38.3125 ;
        RECT  10.63 37.8875 10.765 37.9525 ;
        RECT  10.63 37.8875 10.765 37.9525 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  10.625 39.2325 10.76 39.2975 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  10.2775 37.8875 10.4125 37.9525 ;
        RECT  10.6375 39.2325 10.7375 39.295 ;
        RECT  10.6375 39.235 10.7375 39.2975 ;
        RECT  10.965 38.03 11.0175 38.0925 ;
        RECT  10.6375 39.2325 10.7375 39.295 ;
        RECT  11.015 39.0325 11.085 39.2325 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  10.255 37.8875 11.14 37.9525 ;
        RECT  10.83 38.4025 11.005 38.4675 ;
        RECT  10.31 38.5675 10.38 38.7025 ;
        RECT  10.5 38.4025 10.565 39.1425 ;
        RECT  10.6375 39.235 10.7375 39.2975 ;
        RECT  10.26 38.03 10.3125 38.0925 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  10.255 39.2325 11.14 39.2975 ;
        RECT  10.83 38.4025 10.895 39.0325 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  10.395 38.1775 10.465 38.4675 ;
        RECT  10.31 38.5675 10.38 38.7025 ;
        RECT  10.255 38.0275 11.14 38.0925 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  11.015 39.0325 11.085 39.2325 ;
        RECT  10.31 39.0325 10.38 39.2325 ;
        RECT  10.935 38.1775 11.005 38.4675 ;
        RECT  10.395 38.4025 10.565 38.4675 ;
        RECT  10.255 38.0275 11.14 38.0925 ;
        RECT  10.255 37.8875 11.14 37.9525 ;
        RECT  10.255 39.2325 11.14 39.2975 ;
        RECT  11.015 39.3625 11.08 39.4975 ;
        RECT  10.83 39.3625 10.895 39.4975 ;
        RECT  10.315 39.3625 10.38 39.4975 ;
        RECT  10.5 39.3625 10.565 39.4975 ;
        RECT  10.83 39.8275 10.895 39.9625 ;
        RECT  11.015 39.8275 11.08 39.9625 ;
        RECT  10.5 39.8275 10.565 39.9625 ;
        RECT  10.315 39.8275 10.38 39.9625 ;
        RECT  10.935 40.2175 11.0 40.3525 ;
        RECT  10.75 40.2175 10.815 40.3525 ;
        RECT  10.58 40.2175 10.645 40.3525 ;
        RECT  10.395 40.2175 10.46 40.3525 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  10.625 39.2325 10.76 39.2975 ;
        RECT  10.2775 40.5775 10.4125 40.6425 ;
        RECT  10.9825 40.5775 11.1175 40.6425 ;
        RECT  10.6125 40.4375 10.7475 40.5025 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  10.5175 39.5475 10.6525 39.6125 ;
        RECT  10.5175 39.5475 10.6525 39.6125 ;
        RECT  10.7425 39.6975 10.8775 39.7625 ;
        RECT  10.7425 39.6975 10.8775 39.7625 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  10.5675 40.2175 10.6325 40.3525 ;
        RECT  10.3125 39.725 10.3775 39.86 ;
        RECT  10.3125 39.725 10.3775 39.86 ;
        RECT  10.3125 39.725 10.3775 39.86 ;
        RECT  10.3125 39.725 10.3775 39.86 ;
        RECT  10.3125 39.725 10.3775 39.86 ;
        RECT  10.3125 39.725 10.3775 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  10.7625 40.2175 10.8275 40.3525 ;
        RECT  10.63 40.5775 10.765 40.6425 ;
        RECT  10.63 40.5775 10.765 40.6425 ;
        RECT  10.9825 40.5775 11.1175 40.6425 ;
        RECT  10.625 39.2325 10.76 39.2975 ;
        RECT  10.9825 40.5775 11.1175 40.6425 ;
        RECT  10.9825 40.5775 11.1175 40.6425 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  10.2775 40.5775 10.4125 40.6425 ;
        RECT  10.6375 39.235 10.7375 39.2975 ;
        RECT  10.6375 39.2325 10.7375 39.295 ;
        RECT  10.965 40.4375 11.0175 40.5 ;
        RECT  10.6375 39.235 10.7375 39.2975 ;
        RECT  11.015 39.2975 11.085 39.4975 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  10.255 40.5775 11.14 40.6425 ;
        RECT  10.83 40.0625 11.005 40.1275 ;
        RECT  10.31 39.8275 10.38 39.9625 ;
        RECT  10.5 39.3875 10.565 40.1275 ;
        RECT  10.6375 39.2325 10.7375 39.295 ;
        RECT  10.26 40.4375 10.3125 40.5 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  10.255 39.2325 11.14 39.2975 ;
        RECT  10.83 39.4975 10.895 40.1275 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  10.395 40.0625 10.465 40.3525 ;
        RECT  10.31 39.8275 10.38 39.9625 ;
        RECT  10.255 40.4375 11.14 40.5025 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  11.015 39.2975 11.085 39.4975 ;
        RECT  10.31 39.2975 10.38 39.4975 ;
        RECT  10.935 40.0625 11.005 40.3525 ;
        RECT  10.395 40.0625 10.565 40.1275 ;
        RECT  10.255 40.4375 11.14 40.5025 ;
        RECT  10.255 40.5775 11.14 40.6425 ;
        RECT  10.255 39.2325 11.14 39.2975 ;
        RECT  11.72 20.2025 11.785 20.3375 ;
        RECT  11.535 20.2025 11.6 20.3375 ;
        RECT  11.02 20.2025 11.085 20.3375 ;
        RECT  11.205 20.2025 11.27 20.3375 ;
        RECT  11.535 19.7375 11.6 19.8725 ;
        RECT  11.72 19.7375 11.785 19.8725 ;
        RECT  11.205 19.7375 11.27 19.8725 ;
        RECT  11.02 19.7375 11.085 19.8725 ;
        RECT  11.64 19.3475 11.705 19.4825 ;
        RECT  11.455 19.3475 11.52 19.4825 ;
        RECT  11.285 19.3475 11.35 19.4825 ;
        RECT  11.1 19.3475 11.165 19.4825 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.33 20.4025 11.465 20.4675 ;
        RECT  10.9825 19.0575 11.1175 19.1225 ;
        RECT  11.6875 19.0575 11.8225 19.1225 ;
        RECT  11.3175 19.1975 11.4525 19.2625 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.2225 20.0875 11.3575 20.1525 ;
        RECT  11.2225 20.0875 11.3575 20.1525 ;
        RECT  11.4475 19.9375 11.5825 20.0025 ;
        RECT  11.4475 19.9375 11.5825 20.0025 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.2725 19.3475 11.3375 19.4825 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.4675 19.3475 11.5325 19.4825 ;
        RECT  11.335 19.0575 11.47 19.1225 ;
        RECT  11.335 19.0575 11.47 19.1225 ;
        RECT  11.6875 19.0575 11.8225 19.1225 ;
        RECT  11.33 20.4025 11.465 20.4675 ;
        RECT  11.6875 19.0575 11.8225 19.1225 ;
        RECT  11.6875 19.0575 11.8225 19.1225 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  10.9825 19.0575 11.1175 19.1225 ;
        RECT  11.3425 20.4025 11.4425 20.465 ;
        RECT  11.3425 20.405 11.4425 20.4675 ;
        RECT  11.67 19.2 11.7225 19.2625 ;
        RECT  11.3425 20.4025 11.4425 20.465 ;
        RECT  11.72 20.2025 11.79 20.4025 ;
        RECT  11.72 19.7375 11.79 19.8725 ;
        RECT  11.72 19.7375 11.79 19.8725 ;
        RECT  10.96 19.0575 11.845 19.1225 ;
        RECT  11.535 19.5725 11.71 19.6375 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  11.205 19.5725 11.27 20.3125 ;
        RECT  11.3425 20.405 11.4425 20.4675 ;
        RECT  10.965 19.2 11.0175 19.2625 ;
        RECT  11.72 19.7375 11.79 19.8725 ;
        RECT  10.96 20.4025 11.845 20.4675 ;
        RECT  11.535 19.5725 11.6 20.2025 ;
        RECT  11.72 19.7375 11.79 19.8725 ;
        RECT  11.72 19.7375 11.79 19.8725 ;
        RECT  11.1 19.3475 11.17 19.6375 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  10.96 19.1975 11.845 19.2625 ;
        RECT  11.72 19.7375 11.79 19.8725 ;
        RECT  11.72 20.2025 11.79 20.4025 ;
        RECT  11.015 20.2025 11.085 20.4025 ;
        RECT  11.64 19.3475 11.71 19.6375 ;
        RECT  11.1 19.5725 11.27 19.6375 ;
        RECT  10.96 19.1975 11.845 19.2625 ;
        RECT  10.96 19.0575 11.845 19.1225 ;
        RECT  10.96 20.4025 11.845 20.4675 ;
        RECT  11.72 20.5325 11.785 20.6675 ;
        RECT  11.535 20.5325 11.6 20.6675 ;
        RECT  11.02 20.5325 11.085 20.6675 ;
        RECT  11.205 20.5325 11.27 20.6675 ;
        RECT  11.535 20.9975 11.6 21.1325 ;
        RECT  11.72 20.9975 11.785 21.1325 ;
        RECT  11.205 20.9975 11.27 21.1325 ;
        RECT  11.02 20.9975 11.085 21.1325 ;
        RECT  11.64 21.3875 11.705 21.5225 ;
        RECT  11.455 21.3875 11.52 21.5225 ;
        RECT  11.285 21.3875 11.35 21.5225 ;
        RECT  11.1 21.3875 11.165 21.5225 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.33 20.4025 11.465 20.4675 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.3175 21.6075 11.4525 21.6725 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.2225 20.7175 11.3575 20.7825 ;
        RECT  11.2225 20.7175 11.3575 20.7825 ;
        RECT  11.4475 20.8675 11.5825 20.9325 ;
        RECT  11.4475 20.8675 11.5825 20.9325 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.2725 21.3875 11.3375 21.5225 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.4675 21.3875 11.5325 21.5225 ;
        RECT  11.335 21.7475 11.47 21.8125 ;
        RECT  11.335 21.7475 11.47 21.8125 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.33 20.4025 11.465 20.4675 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  11.3425 20.405 11.4425 20.4675 ;
        RECT  11.3425 20.4025 11.4425 20.465 ;
        RECT  11.67 21.6075 11.7225 21.67 ;
        RECT  11.3425 20.405 11.4425 20.4675 ;
        RECT  11.72 20.4675 11.79 20.6675 ;
        RECT  11.72 20.9975 11.79 21.1325 ;
        RECT  11.72 20.9975 11.79 21.1325 ;
        RECT  10.96 21.7475 11.845 21.8125 ;
        RECT  11.535 21.2325 11.71 21.2975 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  11.205 20.5575 11.27 21.2975 ;
        RECT  11.3425 20.4025 11.4425 20.465 ;
        RECT  10.965 21.6075 11.0175 21.67 ;
        RECT  11.72 20.9975 11.79 21.1325 ;
        RECT  10.96 20.4025 11.845 20.4675 ;
        RECT  11.535 20.6675 11.6 21.2975 ;
        RECT  11.72 20.9975 11.79 21.1325 ;
        RECT  11.72 20.9975 11.79 21.1325 ;
        RECT  11.1 21.2325 11.17 21.5225 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  10.96 21.6075 11.845 21.6725 ;
        RECT  11.72 20.9975 11.79 21.1325 ;
        RECT  11.72 20.4675 11.79 20.6675 ;
        RECT  11.015 20.4675 11.085 20.6675 ;
        RECT  11.64 21.2325 11.71 21.5225 ;
        RECT  11.1 21.2325 11.27 21.2975 ;
        RECT  10.96 21.6075 11.845 21.6725 ;
        RECT  10.96 21.7475 11.845 21.8125 ;
        RECT  10.96 20.4025 11.845 20.4675 ;
        RECT  11.72 22.8925 11.785 23.0275 ;
        RECT  11.535 22.8925 11.6 23.0275 ;
        RECT  11.02 22.8925 11.085 23.0275 ;
        RECT  11.205 22.8925 11.27 23.0275 ;
        RECT  11.535 22.4275 11.6 22.5625 ;
        RECT  11.72 22.4275 11.785 22.5625 ;
        RECT  11.205 22.4275 11.27 22.5625 ;
        RECT  11.02 22.4275 11.085 22.5625 ;
        RECT  11.64 22.0375 11.705 22.1725 ;
        RECT  11.455 22.0375 11.52 22.1725 ;
        RECT  11.285 22.0375 11.35 22.1725 ;
        RECT  11.1 22.0375 11.165 22.1725 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.33 23.0925 11.465 23.1575 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.3175 21.8875 11.4525 21.9525 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.2225 22.7775 11.3575 22.8425 ;
        RECT  11.2225 22.7775 11.3575 22.8425 ;
        RECT  11.4475 22.6275 11.5825 22.6925 ;
        RECT  11.4475 22.6275 11.5825 22.6925 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.2725 22.0375 11.3375 22.1725 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.4675 22.0375 11.5325 22.1725 ;
        RECT  11.335 21.7475 11.47 21.8125 ;
        RECT  11.335 21.7475 11.47 21.8125 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.33 23.0925 11.465 23.1575 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  11.3425 23.0925 11.4425 23.155 ;
        RECT  11.3425 23.095 11.4425 23.1575 ;
        RECT  11.67 21.89 11.7225 21.9525 ;
        RECT  11.3425 23.0925 11.4425 23.155 ;
        RECT  11.72 22.8925 11.79 23.0925 ;
        RECT  11.72 22.4275 11.79 22.5625 ;
        RECT  11.72 22.4275 11.79 22.5625 ;
        RECT  10.96 21.7475 11.845 21.8125 ;
        RECT  11.535 22.2625 11.71 22.3275 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  11.205 22.2625 11.27 23.0025 ;
        RECT  11.3425 23.095 11.4425 23.1575 ;
        RECT  10.965 21.89 11.0175 21.9525 ;
        RECT  11.72 22.4275 11.79 22.5625 ;
        RECT  10.96 23.0925 11.845 23.1575 ;
        RECT  11.535 22.2625 11.6 22.8925 ;
        RECT  11.72 22.4275 11.79 22.5625 ;
        RECT  11.72 22.4275 11.79 22.5625 ;
        RECT  11.1 22.0375 11.17 22.3275 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  10.96 21.8875 11.845 21.9525 ;
        RECT  11.72 22.4275 11.79 22.5625 ;
        RECT  11.72 22.8925 11.79 23.0925 ;
        RECT  11.015 22.8925 11.085 23.0925 ;
        RECT  11.64 22.0375 11.71 22.3275 ;
        RECT  11.1 22.2625 11.27 22.3275 ;
        RECT  10.96 21.8875 11.845 21.9525 ;
        RECT  10.96 21.7475 11.845 21.8125 ;
        RECT  10.96 23.0925 11.845 23.1575 ;
        RECT  11.72 23.2225 11.785 23.3575 ;
        RECT  11.535 23.2225 11.6 23.3575 ;
        RECT  11.02 23.2225 11.085 23.3575 ;
        RECT  11.205 23.2225 11.27 23.3575 ;
        RECT  11.535 23.6875 11.6 23.8225 ;
        RECT  11.72 23.6875 11.785 23.8225 ;
        RECT  11.205 23.6875 11.27 23.8225 ;
        RECT  11.02 23.6875 11.085 23.8225 ;
        RECT  11.64 24.0775 11.705 24.2125 ;
        RECT  11.455 24.0775 11.52 24.2125 ;
        RECT  11.285 24.0775 11.35 24.2125 ;
        RECT  11.1 24.0775 11.165 24.2125 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.33 23.0925 11.465 23.1575 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.3175 24.2975 11.4525 24.3625 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.2225 23.4075 11.3575 23.4725 ;
        RECT  11.2225 23.4075 11.3575 23.4725 ;
        RECT  11.4475 23.5575 11.5825 23.6225 ;
        RECT  11.4475 23.5575 11.5825 23.6225 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.2725 24.0775 11.3375 24.2125 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.4675 24.0775 11.5325 24.2125 ;
        RECT  11.335 24.4375 11.47 24.5025 ;
        RECT  11.335 24.4375 11.47 24.5025 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.33 23.0925 11.465 23.1575 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  11.3425 23.095 11.4425 23.1575 ;
        RECT  11.3425 23.0925 11.4425 23.155 ;
        RECT  11.67 24.2975 11.7225 24.36 ;
        RECT  11.3425 23.095 11.4425 23.1575 ;
        RECT  11.72 23.1575 11.79 23.3575 ;
        RECT  11.72 23.6875 11.79 23.8225 ;
        RECT  11.72 23.6875 11.79 23.8225 ;
        RECT  10.96 24.4375 11.845 24.5025 ;
        RECT  11.535 23.9225 11.71 23.9875 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  11.205 23.2475 11.27 23.9875 ;
        RECT  11.3425 23.0925 11.4425 23.155 ;
        RECT  10.965 24.2975 11.0175 24.36 ;
        RECT  11.72 23.6875 11.79 23.8225 ;
        RECT  10.96 23.0925 11.845 23.1575 ;
        RECT  11.535 23.3575 11.6 23.9875 ;
        RECT  11.72 23.6875 11.79 23.8225 ;
        RECT  11.72 23.6875 11.79 23.8225 ;
        RECT  11.1 23.9225 11.17 24.2125 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  10.96 24.2975 11.845 24.3625 ;
        RECT  11.72 23.6875 11.79 23.8225 ;
        RECT  11.72 23.1575 11.79 23.3575 ;
        RECT  11.015 23.1575 11.085 23.3575 ;
        RECT  11.64 23.9225 11.71 24.2125 ;
        RECT  11.1 23.9225 11.27 23.9875 ;
        RECT  10.96 24.2975 11.845 24.3625 ;
        RECT  10.96 24.4375 11.845 24.5025 ;
        RECT  10.96 23.0925 11.845 23.1575 ;
        RECT  11.72 25.5825 11.785 25.7175 ;
        RECT  11.535 25.5825 11.6 25.7175 ;
        RECT  11.02 25.5825 11.085 25.7175 ;
        RECT  11.205 25.5825 11.27 25.7175 ;
        RECT  11.535 25.1175 11.6 25.2525 ;
        RECT  11.72 25.1175 11.785 25.2525 ;
        RECT  11.205 25.1175 11.27 25.2525 ;
        RECT  11.02 25.1175 11.085 25.2525 ;
        RECT  11.64 24.7275 11.705 24.8625 ;
        RECT  11.455 24.7275 11.52 24.8625 ;
        RECT  11.285 24.7275 11.35 24.8625 ;
        RECT  11.1 24.7275 11.165 24.8625 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.33 25.7825 11.465 25.8475 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.3175 24.5775 11.4525 24.6425 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.2225 25.4675 11.3575 25.5325 ;
        RECT  11.2225 25.4675 11.3575 25.5325 ;
        RECT  11.4475 25.3175 11.5825 25.3825 ;
        RECT  11.4475 25.3175 11.5825 25.3825 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.2725 24.7275 11.3375 24.8625 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.4675 24.7275 11.5325 24.8625 ;
        RECT  11.335 24.4375 11.47 24.5025 ;
        RECT  11.335 24.4375 11.47 24.5025 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.33 25.7825 11.465 25.8475 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  11.3425 25.7825 11.4425 25.845 ;
        RECT  11.3425 25.785 11.4425 25.8475 ;
        RECT  11.67 24.58 11.7225 24.6425 ;
        RECT  11.3425 25.7825 11.4425 25.845 ;
        RECT  11.72 25.5825 11.79 25.7825 ;
        RECT  11.72 25.1175 11.79 25.2525 ;
        RECT  11.72 25.1175 11.79 25.2525 ;
        RECT  10.96 24.4375 11.845 24.5025 ;
        RECT  11.535 24.9525 11.71 25.0175 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  11.205 24.9525 11.27 25.6925 ;
        RECT  11.3425 25.785 11.4425 25.8475 ;
        RECT  10.965 24.58 11.0175 24.6425 ;
        RECT  11.72 25.1175 11.79 25.2525 ;
        RECT  10.96 25.7825 11.845 25.8475 ;
        RECT  11.535 24.9525 11.6 25.5825 ;
        RECT  11.72 25.1175 11.79 25.2525 ;
        RECT  11.72 25.1175 11.79 25.2525 ;
        RECT  11.1 24.7275 11.17 25.0175 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  10.96 24.5775 11.845 24.6425 ;
        RECT  11.72 25.1175 11.79 25.2525 ;
        RECT  11.72 25.5825 11.79 25.7825 ;
        RECT  11.015 25.5825 11.085 25.7825 ;
        RECT  11.64 24.7275 11.71 25.0175 ;
        RECT  11.1 24.9525 11.27 25.0175 ;
        RECT  10.96 24.5775 11.845 24.6425 ;
        RECT  10.96 24.4375 11.845 24.5025 ;
        RECT  10.96 25.7825 11.845 25.8475 ;
        RECT  11.72 25.9125 11.785 26.0475 ;
        RECT  11.535 25.9125 11.6 26.0475 ;
        RECT  11.02 25.9125 11.085 26.0475 ;
        RECT  11.205 25.9125 11.27 26.0475 ;
        RECT  11.535 26.3775 11.6 26.5125 ;
        RECT  11.72 26.3775 11.785 26.5125 ;
        RECT  11.205 26.3775 11.27 26.5125 ;
        RECT  11.02 26.3775 11.085 26.5125 ;
        RECT  11.64 26.7675 11.705 26.9025 ;
        RECT  11.455 26.7675 11.52 26.9025 ;
        RECT  11.285 26.7675 11.35 26.9025 ;
        RECT  11.1 26.7675 11.165 26.9025 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.33 25.7825 11.465 25.8475 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.3175 26.9875 11.4525 27.0525 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.2225 26.0975 11.3575 26.1625 ;
        RECT  11.2225 26.0975 11.3575 26.1625 ;
        RECT  11.4475 26.2475 11.5825 26.3125 ;
        RECT  11.4475 26.2475 11.5825 26.3125 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.2725 26.7675 11.3375 26.9025 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.4675 26.7675 11.5325 26.9025 ;
        RECT  11.335 27.1275 11.47 27.1925 ;
        RECT  11.335 27.1275 11.47 27.1925 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.33 25.7825 11.465 25.8475 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  11.3425 25.785 11.4425 25.8475 ;
        RECT  11.3425 25.7825 11.4425 25.845 ;
        RECT  11.67 26.9875 11.7225 27.05 ;
        RECT  11.3425 25.785 11.4425 25.8475 ;
        RECT  11.72 25.8475 11.79 26.0475 ;
        RECT  11.72 26.3775 11.79 26.5125 ;
        RECT  11.72 26.3775 11.79 26.5125 ;
        RECT  10.96 27.1275 11.845 27.1925 ;
        RECT  11.535 26.6125 11.71 26.6775 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  11.205 25.9375 11.27 26.6775 ;
        RECT  11.3425 25.7825 11.4425 25.845 ;
        RECT  10.965 26.9875 11.0175 27.05 ;
        RECT  11.72 26.3775 11.79 26.5125 ;
        RECT  10.96 25.7825 11.845 25.8475 ;
        RECT  11.535 26.0475 11.6 26.6775 ;
        RECT  11.72 26.3775 11.79 26.5125 ;
        RECT  11.72 26.3775 11.79 26.5125 ;
        RECT  11.1 26.6125 11.17 26.9025 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  10.96 26.9875 11.845 27.0525 ;
        RECT  11.72 26.3775 11.79 26.5125 ;
        RECT  11.72 25.8475 11.79 26.0475 ;
        RECT  11.015 25.8475 11.085 26.0475 ;
        RECT  11.64 26.6125 11.71 26.9025 ;
        RECT  11.1 26.6125 11.27 26.6775 ;
        RECT  10.96 26.9875 11.845 27.0525 ;
        RECT  10.96 27.1275 11.845 27.1925 ;
        RECT  10.96 25.7825 11.845 25.8475 ;
        RECT  11.72 28.2725 11.785 28.4075 ;
        RECT  11.535 28.2725 11.6 28.4075 ;
        RECT  11.02 28.2725 11.085 28.4075 ;
        RECT  11.205 28.2725 11.27 28.4075 ;
        RECT  11.535 27.8075 11.6 27.9425 ;
        RECT  11.72 27.8075 11.785 27.9425 ;
        RECT  11.205 27.8075 11.27 27.9425 ;
        RECT  11.02 27.8075 11.085 27.9425 ;
        RECT  11.64 27.4175 11.705 27.5525 ;
        RECT  11.455 27.4175 11.52 27.5525 ;
        RECT  11.285 27.4175 11.35 27.5525 ;
        RECT  11.1 27.4175 11.165 27.5525 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.33 28.4725 11.465 28.5375 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.3175 27.2675 11.4525 27.3325 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.2225 28.1575 11.3575 28.2225 ;
        RECT  11.2225 28.1575 11.3575 28.2225 ;
        RECT  11.4475 28.0075 11.5825 28.0725 ;
        RECT  11.4475 28.0075 11.5825 28.0725 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.2725 27.4175 11.3375 27.5525 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.4675 27.4175 11.5325 27.5525 ;
        RECT  11.335 27.1275 11.47 27.1925 ;
        RECT  11.335 27.1275 11.47 27.1925 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.33 28.4725 11.465 28.5375 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  11.3425 28.4725 11.4425 28.535 ;
        RECT  11.3425 28.475 11.4425 28.5375 ;
        RECT  11.67 27.27 11.7225 27.3325 ;
        RECT  11.3425 28.4725 11.4425 28.535 ;
        RECT  11.72 28.2725 11.79 28.4725 ;
        RECT  11.72 27.8075 11.79 27.9425 ;
        RECT  11.72 27.8075 11.79 27.9425 ;
        RECT  10.96 27.1275 11.845 27.1925 ;
        RECT  11.535 27.6425 11.71 27.7075 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  11.205 27.6425 11.27 28.3825 ;
        RECT  11.3425 28.475 11.4425 28.5375 ;
        RECT  10.965 27.27 11.0175 27.3325 ;
        RECT  11.72 27.8075 11.79 27.9425 ;
        RECT  10.96 28.4725 11.845 28.5375 ;
        RECT  11.535 27.6425 11.6 28.2725 ;
        RECT  11.72 27.8075 11.79 27.9425 ;
        RECT  11.72 27.8075 11.79 27.9425 ;
        RECT  11.1 27.4175 11.17 27.7075 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  10.96 27.2675 11.845 27.3325 ;
        RECT  11.72 27.8075 11.79 27.9425 ;
        RECT  11.72 28.2725 11.79 28.4725 ;
        RECT  11.015 28.2725 11.085 28.4725 ;
        RECT  11.64 27.4175 11.71 27.7075 ;
        RECT  11.1 27.6425 11.27 27.7075 ;
        RECT  10.96 27.2675 11.845 27.3325 ;
        RECT  10.96 27.1275 11.845 27.1925 ;
        RECT  10.96 28.4725 11.845 28.5375 ;
        RECT  11.72 28.6025 11.785 28.7375 ;
        RECT  11.535 28.6025 11.6 28.7375 ;
        RECT  11.02 28.6025 11.085 28.7375 ;
        RECT  11.205 28.6025 11.27 28.7375 ;
        RECT  11.535 29.0675 11.6 29.2025 ;
        RECT  11.72 29.0675 11.785 29.2025 ;
        RECT  11.205 29.0675 11.27 29.2025 ;
        RECT  11.02 29.0675 11.085 29.2025 ;
        RECT  11.64 29.4575 11.705 29.5925 ;
        RECT  11.455 29.4575 11.52 29.5925 ;
        RECT  11.285 29.4575 11.35 29.5925 ;
        RECT  11.1 29.4575 11.165 29.5925 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.33 28.4725 11.465 28.5375 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.3175 29.6775 11.4525 29.7425 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.2225 28.7875 11.3575 28.8525 ;
        RECT  11.2225 28.7875 11.3575 28.8525 ;
        RECT  11.4475 28.9375 11.5825 29.0025 ;
        RECT  11.4475 28.9375 11.5825 29.0025 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.2725 29.4575 11.3375 29.5925 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.4675 29.4575 11.5325 29.5925 ;
        RECT  11.335 29.8175 11.47 29.8825 ;
        RECT  11.335 29.8175 11.47 29.8825 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.33 28.4725 11.465 28.5375 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  11.3425 28.475 11.4425 28.5375 ;
        RECT  11.3425 28.4725 11.4425 28.535 ;
        RECT  11.67 29.6775 11.7225 29.74 ;
        RECT  11.3425 28.475 11.4425 28.5375 ;
        RECT  11.72 28.5375 11.79 28.7375 ;
        RECT  11.72 29.0675 11.79 29.2025 ;
        RECT  11.72 29.0675 11.79 29.2025 ;
        RECT  10.96 29.8175 11.845 29.8825 ;
        RECT  11.535 29.3025 11.71 29.3675 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  11.205 28.6275 11.27 29.3675 ;
        RECT  11.3425 28.4725 11.4425 28.535 ;
        RECT  10.965 29.6775 11.0175 29.74 ;
        RECT  11.72 29.0675 11.79 29.2025 ;
        RECT  10.96 28.4725 11.845 28.5375 ;
        RECT  11.535 28.7375 11.6 29.3675 ;
        RECT  11.72 29.0675 11.79 29.2025 ;
        RECT  11.72 29.0675 11.79 29.2025 ;
        RECT  11.1 29.3025 11.17 29.5925 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  10.96 29.6775 11.845 29.7425 ;
        RECT  11.72 29.0675 11.79 29.2025 ;
        RECT  11.72 28.5375 11.79 28.7375 ;
        RECT  11.015 28.5375 11.085 28.7375 ;
        RECT  11.64 29.3025 11.71 29.5925 ;
        RECT  11.1 29.3025 11.27 29.3675 ;
        RECT  10.96 29.6775 11.845 29.7425 ;
        RECT  10.96 29.8175 11.845 29.8825 ;
        RECT  10.96 28.4725 11.845 28.5375 ;
        RECT  11.72 30.9625 11.785 31.0975 ;
        RECT  11.535 30.9625 11.6 31.0975 ;
        RECT  11.02 30.9625 11.085 31.0975 ;
        RECT  11.205 30.9625 11.27 31.0975 ;
        RECT  11.535 30.4975 11.6 30.6325 ;
        RECT  11.72 30.4975 11.785 30.6325 ;
        RECT  11.205 30.4975 11.27 30.6325 ;
        RECT  11.02 30.4975 11.085 30.6325 ;
        RECT  11.64 30.1075 11.705 30.2425 ;
        RECT  11.455 30.1075 11.52 30.2425 ;
        RECT  11.285 30.1075 11.35 30.2425 ;
        RECT  11.1 30.1075 11.165 30.2425 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.33 31.1625 11.465 31.2275 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.3175 29.9575 11.4525 30.0225 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.2225 30.8475 11.3575 30.9125 ;
        RECT  11.2225 30.8475 11.3575 30.9125 ;
        RECT  11.4475 30.6975 11.5825 30.7625 ;
        RECT  11.4475 30.6975 11.5825 30.7625 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.2725 30.1075 11.3375 30.2425 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.4675 30.1075 11.5325 30.2425 ;
        RECT  11.335 29.8175 11.47 29.8825 ;
        RECT  11.335 29.8175 11.47 29.8825 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.33 31.1625 11.465 31.2275 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  11.3425 31.1625 11.4425 31.225 ;
        RECT  11.3425 31.165 11.4425 31.2275 ;
        RECT  11.67 29.96 11.7225 30.0225 ;
        RECT  11.3425 31.1625 11.4425 31.225 ;
        RECT  11.72 30.9625 11.79 31.1625 ;
        RECT  11.72 30.4975 11.79 30.6325 ;
        RECT  11.72 30.4975 11.79 30.6325 ;
        RECT  10.96 29.8175 11.845 29.8825 ;
        RECT  11.535 30.3325 11.71 30.3975 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  11.205 30.3325 11.27 31.0725 ;
        RECT  11.3425 31.165 11.4425 31.2275 ;
        RECT  10.965 29.96 11.0175 30.0225 ;
        RECT  11.72 30.4975 11.79 30.6325 ;
        RECT  10.96 31.1625 11.845 31.2275 ;
        RECT  11.535 30.3325 11.6 30.9625 ;
        RECT  11.72 30.4975 11.79 30.6325 ;
        RECT  11.72 30.4975 11.79 30.6325 ;
        RECT  11.1 30.1075 11.17 30.3975 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  10.96 29.9575 11.845 30.0225 ;
        RECT  11.72 30.4975 11.79 30.6325 ;
        RECT  11.72 30.9625 11.79 31.1625 ;
        RECT  11.015 30.9625 11.085 31.1625 ;
        RECT  11.64 30.1075 11.71 30.3975 ;
        RECT  11.1 30.3325 11.27 30.3975 ;
        RECT  10.96 29.9575 11.845 30.0225 ;
        RECT  10.96 29.8175 11.845 29.8825 ;
        RECT  10.96 31.1625 11.845 31.2275 ;
        RECT  11.72 31.2925 11.785 31.4275 ;
        RECT  11.535 31.2925 11.6 31.4275 ;
        RECT  11.02 31.2925 11.085 31.4275 ;
        RECT  11.205 31.2925 11.27 31.4275 ;
        RECT  11.535 31.7575 11.6 31.8925 ;
        RECT  11.72 31.7575 11.785 31.8925 ;
        RECT  11.205 31.7575 11.27 31.8925 ;
        RECT  11.02 31.7575 11.085 31.8925 ;
        RECT  11.64 32.1475 11.705 32.2825 ;
        RECT  11.455 32.1475 11.52 32.2825 ;
        RECT  11.285 32.1475 11.35 32.2825 ;
        RECT  11.1 32.1475 11.165 32.2825 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.33 31.1625 11.465 31.2275 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.3175 32.3675 11.4525 32.4325 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.2225 31.4775 11.3575 31.5425 ;
        RECT  11.2225 31.4775 11.3575 31.5425 ;
        RECT  11.4475 31.6275 11.5825 31.6925 ;
        RECT  11.4475 31.6275 11.5825 31.6925 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.2725 32.1475 11.3375 32.2825 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.4675 32.1475 11.5325 32.2825 ;
        RECT  11.335 32.5075 11.47 32.5725 ;
        RECT  11.335 32.5075 11.47 32.5725 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.33 31.1625 11.465 31.2275 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  11.3425 31.165 11.4425 31.2275 ;
        RECT  11.3425 31.1625 11.4425 31.225 ;
        RECT  11.67 32.3675 11.7225 32.43 ;
        RECT  11.3425 31.165 11.4425 31.2275 ;
        RECT  11.72 31.2275 11.79 31.4275 ;
        RECT  11.72 31.7575 11.79 31.8925 ;
        RECT  11.72 31.7575 11.79 31.8925 ;
        RECT  10.96 32.5075 11.845 32.5725 ;
        RECT  11.535 31.9925 11.71 32.0575 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  11.205 31.3175 11.27 32.0575 ;
        RECT  11.3425 31.1625 11.4425 31.225 ;
        RECT  10.965 32.3675 11.0175 32.43 ;
        RECT  11.72 31.7575 11.79 31.8925 ;
        RECT  10.96 31.1625 11.845 31.2275 ;
        RECT  11.535 31.4275 11.6 32.0575 ;
        RECT  11.72 31.7575 11.79 31.8925 ;
        RECT  11.72 31.7575 11.79 31.8925 ;
        RECT  11.1 31.9925 11.17 32.2825 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  10.96 32.3675 11.845 32.4325 ;
        RECT  11.72 31.7575 11.79 31.8925 ;
        RECT  11.72 31.2275 11.79 31.4275 ;
        RECT  11.015 31.2275 11.085 31.4275 ;
        RECT  11.64 31.9925 11.71 32.2825 ;
        RECT  11.1 31.9925 11.27 32.0575 ;
        RECT  10.96 32.3675 11.845 32.4325 ;
        RECT  10.96 32.5075 11.845 32.5725 ;
        RECT  10.96 31.1625 11.845 31.2275 ;
        RECT  11.72 33.6525 11.785 33.7875 ;
        RECT  11.535 33.6525 11.6 33.7875 ;
        RECT  11.02 33.6525 11.085 33.7875 ;
        RECT  11.205 33.6525 11.27 33.7875 ;
        RECT  11.535 33.1875 11.6 33.3225 ;
        RECT  11.72 33.1875 11.785 33.3225 ;
        RECT  11.205 33.1875 11.27 33.3225 ;
        RECT  11.02 33.1875 11.085 33.3225 ;
        RECT  11.64 32.7975 11.705 32.9325 ;
        RECT  11.455 32.7975 11.52 32.9325 ;
        RECT  11.285 32.7975 11.35 32.9325 ;
        RECT  11.1 32.7975 11.165 32.9325 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.33 33.8525 11.465 33.9175 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.3175 32.6475 11.4525 32.7125 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.2225 33.5375 11.3575 33.6025 ;
        RECT  11.2225 33.5375 11.3575 33.6025 ;
        RECT  11.4475 33.3875 11.5825 33.4525 ;
        RECT  11.4475 33.3875 11.5825 33.4525 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.2725 32.7975 11.3375 32.9325 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.4675 32.7975 11.5325 32.9325 ;
        RECT  11.335 32.5075 11.47 32.5725 ;
        RECT  11.335 32.5075 11.47 32.5725 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.33 33.8525 11.465 33.9175 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  11.3425 33.8525 11.4425 33.915 ;
        RECT  11.3425 33.855 11.4425 33.9175 ;
        RECT  11.67 32.65 11.7225 32.7125 ;
        RECT  11.3425 33.8525 11.4425 33.915 ;
        RECT  11.72 33.6525 11.79 33.8525 ;
        RECT  11.72 33.1875 11.79 33.3225 ;
        RECT  11.72 33.1875 11.79 33.3225 ;
        RECT  10.96 32.5075 11.845 32.5725 ;
        RECT  11.535 33.0225 11.71 33.0875 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  11.205 33.0225 11.27 33.7625 ;
        RECT  11.3425 33.855 11.4425 33.9175 ;
        RECT  10.965 32.65 11.0175 32.7125 ;
        RECT  11.72 33.1875 11.79 33.3225 ;
        RECT  10.96 33.8525 11.845 33.9175 ;
        RECT  11.535 33.0225 11.6 33.6525 ;
        RECT  11.72 33.1875 11.79 33.3225 ;
        RECT  11.72 33.1875 11.79 33.3225 ;
        RECT  11.1 32.7975 11.17 33.0875 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  10.96 32.6475 11.845 32.7125 ;
        RECT  11.72 33.1875 11.79 33.3225 ;
        RECT  11.72 33.6525 11.79 33.8525 ;
        RECT  11.015 33.6525 11.085 33.8525 ;
        RECT  11.64 32.7975 11.71 33.0875 ;
        RECT  11.1 33.0225 11.27 33.0875 ;
        RECT  10.96 32.6475 11.845 32.7125 ;
        RECT  10.96 32.5075 11.845 32.5725 ;
        RECT  10.96 33.8525 11.845 33.9175 ;
        RECT  11.72 33.9825 11.785 34.1175 ;
        RECT  11.535 33.9825 11.6 34.1175 ;
        RECT  11.02 33.9825 11.085 34.1175 ;
        RECT  11.205 33.9825 11.27 34.1175 ;
        RECT  11.535 34.4475 11.6 34.5825 ;
        RECT  11.72 34.4475 11.785 34.5825 ;
        RECT  11.205 34.4475 11.27 34.5825 ;
        RECT  11.02 34.4475 11.085 34.5825 ;
        RECT  11.64 34.8375 11.705 34.9725 ;
        RECT  11.455 34.8375 11.52 34.9725 ;
        RECT  11.285 34.8375 11.35 34.9725 ;
        RECT  11.1 34.8375 11.165 34.9725 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.33 33.8525 11.465 33.9175 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.3175 35.0575 11.4525 35.1225 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.2225 34.1675 11.3575 34.2325 ;
        RECT  11.2225 34.1675 11.3575 34.2325 ;
        RECT  11.4475 34.3175 11.5825 34.3825 ;
        RECT  11.4475 34.3175 11.5825 34.3825 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.2725 34.8375 11.3375 34.9725 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.4675 34.8375 11.5325 34.9725 ;
        RECT  11.335 35.1975 11.47 35.2625 ;
        RECT  11.335 35.1975 11.47 35.2625 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.33 33.8525 11.465 33.9175 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  11.3425 33.855 11.4425 33.9175 ;
        RECT  11.3425 33.8525 11.4425 33.915 ;
        RECT  11.67 35.0575 11.7225 35.12 ;
        RECT  11.3425 33.855 11.4425 33.9175 ;
        RECT  11.72 33.9175 11.79 34.1175 ;
        RECT  11.72 34.4475 11.79 34.5825 ;
        RECT  11.72 34.4475 11.79 34.5825 ;
        RECT  10.96 35.1975 11.845 35.2625 ;
        RECT  11.535 34.6825 11.71 34.7475 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  11.205 34.0075 11.27 34.7475 ;
        RECT  11.3425 33.8525 11.4425 33.915 ;
        RECT  10.965 35.0575 11.0175 35.12 ;
        RECT  11.72 34.4475 11.79 34.5825 ;
        RECT  10.96 33.8525 11.845 33.9175 ;
        RECT  11.535 34.1175 11.6 34.7475 ;
        RECT  11.72 34.4475 11.79 34.5825 ;
        RECT  11.72 34.4475 11.79 34.5825 ;
        RECT  11.1 34.6825 11.17 34.9725 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  10.96 35.0575 11.845 35.1225 ;
        RECT  11.72 34.4475 11.79 34.5825 ;
        RECT  11.72 33.9175 11.79 34.1175 ;
        RECT  11.015 33.9175 11.085 34.1175 ;
        RECT  11.64 34.6825 11.71 34.9725 ;
        RECT  11.1 34.6825 11.27 34.7475 ;
        RECT  10.96 35.0575 11.845 35.1225 ;
        RECT  10.96 35.1975 11.845 35.2625 ;
        RECT  10.96 33.8525 11.845 33.9175 ;
        RECT  11.72 36.3425 11.785 36.4775 ;
        RECT  11.535 36.3425 11.6 36.4775 ;
        RECT  11.02 36.3425 11.085 36.4775 ;
        RECT  11.205 36.3425 11.27 36.4775 ;
        RECT  11.535 35.8775 11.6 36.0125 ;
        RECT  11.72 35.8775 11.785 36.0125 ;
        RECT  11.205 35.8775 11.27 36.0125 ;
        RECT  11.02 35.8775 11.085 36.0125 ;
        RECT  11.64 35.4875 11.705 35.6225 ;
        RECT  11.455 35.4875 11.52 35.6225 ;
        RECT  11.285 35.4875 11.35 35.6225 ;
        RECT  11.1 35.4875 11.165 35.6225 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.33 36.5425 11.465 36.6075 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.3175 35.3375 11.4525 35.4025 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.2225 36.2275 11.3575 36.2925 ;
        RECT  11.2225 36.2275 11.3575 36.2925 ;
        RECT  11.4475 36.0775 11.5825 36.1425 ;
        RECT  11.4475 36.0775 11.5825 36.1425 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.2725 35.4875 11.3375 35.6225 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.4675 35.4875 11.5325 35.6225 ;
        RECT  11.335 35.1975 11.47 35.2625 ;
        RECT  11.335 35.1975 11.47 35.2625 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.33 36.5425 11.465 36.6075 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  11.3425 36.5425 11.4425 36.605 ;
        RECT  11.3425 36.545 11.4425 36.6075 ;
        RECT  11.67 35.34 11.7225 35.4025 ;
        RECT  11.3425 36.5425 11.4425 36.605 ;
        RECT  11.72 36.3425 11.79 36.5425 ;
        RECT  11.72 35.8775 11.79 36.0125 ;
        RECT  11.72 35.8775 11.79 36.0125 ;
        RECT  10.96 35.1975 11.845 35.2625 ;
        RECT  11.535 35.7125 11.71 35.7775 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  11.205 35.7125 11.27 36.4525 ;
        RECT  11.3425 36.545 11.4425 36.6075 ;
        RECT  10.965 35.34 11.0175 35.4025 ;
        RECT  11.72 35.8775 11.79 36.0125 ;
        RECT  10.96 36.5425 11.845 36.6075 ;
        RECT  11.535 35.7125 11.6 36.3425 ;
        RECT  11.72 35.8775 11.79 36.0125 ;
        RECT  11.72 35.8775 11.79 36.0125 ;
        RECT  11.1 35.4875 11.17 35.7775 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  10.96 35.3375 11.845 35.4025 ;
        RECT  11.72 35.8775 11.79 36.0125 ;
        RECT  11.72 36.3425 11.79 36.5425 ;
        RECT  11.015 36.3425 11.085 36.5425 ;
        RECT  11.64 35.4875 11.71 35.7775 ;
        RECT  11.1 35.7125 11.27 35.7775 ;
        RECT  10.96 35.3375 11.845 35.4025 ;
        RECT  10.96 35.1975 11.845 35.2625 ;
        RECT  10.96 36.5425 11.845 36.6075 ;
        RECT  11.72 36.6725 11.785 36.8075 ;
        RECT  11.535 36.6725 11.6 36.8075 ;
        RECT  11.02 36.6725 11.085 36.8075 ;
        RECT  11.205 36.6725 11.27 36.8075 ;
        RECT  11.535 37.1375 11.6 37.2725 ;
        RECT  11.72 37.1375 11.785 37.2725 ;
        RECT  11.205 37.1375 11.27 37.2725 ;
        RECT  11.02 37.1375 11.085 37.2725 ;
        RECT  11.64 37.5275 11.705 37.6625 ;
        RECT  11.455 37.5275 11.52 37.6625 ;
        RECT  11.285 37.5275 11.35 37.6625 ;
        RECT  11.1 37.5275 11.165 37.6625 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.33 36.5425 11.465 36.6075 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.3175 37.7475 11.4525 37.8125 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.2225 36.8575 11.3575 36.9225 ;
        RECT  11.2225 36.8575 11.3575 36.9225 ;
        RECT  11.4475 37.0075 11.5825 37.0725 ;
        RECT  11.4475 37.0075 11.5825 37.0725 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.2725 37.5275 11.3375 37.6625 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.4675 37.5275 11.5325 37.6625 ;
        RECT  11.335 37.8875 11.47 37.9525 ;
        RECT  11.335 37.8875 11.47 37.9525 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.33 36.5425 11.465 36.6075 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  11.3425 36.545 11.4425 36.6075 ;
        RECT  11.3425 36.5425 11.4425 36.605 ;
        RECT  11.67 37.7475 11.7225 37.81 ;
        RECT  11.3425 36.545 11.4425 36.6075 ;
        RECT  11.72 36.6075 11.79 36.8075 ;
        RECT  11.72 37.1375 11.79 37.2725 ;
        RECT  11.72 37.1375 11.79 37.2725 ;
        RECT  10.96 37.8875 11.845 37.9525 ;
        RECT  11.535 37.3725 11.71 37.4375 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  11.205 36.6975 11.27 37.4375 ;
        RECT  11.3425 36.5425 11.4425 36.605 ;
        RECT  10.965 37.7475 11.0175 37.81 ;
        RECT  11.72 37.1375 11.79 37.2725 ;
        RECT  10.96 36.5425 11.845 36.6075 ;
        RECT  11.535 36.8075 11.6 37.4375 ;
        RECT  11.72 37.1375 11.79 37.2725 ;
        RECT  11.72 37.1375 11.79 37.2725 ;
        RECT  11.1 37.3725 11.17 37.6625 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  10.96 37.7475 11.845 37.8125 ;
        RECT  11.72 37.1375 11.79 37.2725 ;
        RECT  11.72 36.6075 11.79 36.8075 ;
        RECT  11.015 36.6075 11.085 36.8075 ;
        RECT  11.64 37.3725 11.71 37.6625 ;
        RECT  11.1 37.3725 11.27 37.4375 ;
        RECT  10.96 37.7475 11.845 37.8125 ;
        RECT  10.96 37.8875 11.845 37.9525 ;
        RECT  10.96 36.5425 11.845 36.6075 ;
        RECT  11.72 39.0325 11.785 39.1675 ;
        RECT  11.535 39.0325 11.6 39.1675 ;
        RECT  11.02 39.0325 11.085 39.1675 ;
        RECT  11.205 39.0325 11.27 39.1675 ;
        RECT  11.535 38.5675 11.6 38.7025 ;
        RECT  11.72 38.5675 11.785 38.7025 ;
        RECT  11.205 38.5675 11.27 38.7025 ;
        RECT  11.02 38.5675 11.085 38.7025 ;
        RECT  11.64 38.1775 11.705 38.3125 ;
        RECT  11.455 38.1775 11.52 38.3125 ;
        RECT  11.285 38.1775 11.35 38.3125 ;
        RECT  11.1 38.1775 11.165 38.3125 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.33 39.2325 11.465 39.2975 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.3175 38.0275 11.4525 38.0925 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.2225 38.9175 11.3575 38.9825 ;
        RECT  11.2225 38.9175 11.3575 38.9825 ;
        RECT  11.4475 38.7675 11.5825 38.8325 ;
        RECT  11.4475 38.7675 11.5825 38.8325 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.2725 38.1775 11.3375 38.3125 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.4675 38.1775 11.5325 38.3125 ;
        RECT  11.335 37.8875 11.47 37.9525 ;
        RECT  11.335 37.8875 11.47 37.9525 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.33 39.2325 11.465 39.2975 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  11.3425 39.2325 11.4425 39.295 ;
        RECT  11.3425 39.235 11.4425 39.2975 ;
        RECT  11.67 38.03 11.7225 38.0925 ;
        RECT  11.3425 39.2325 11.4425 39.295 ;
        RECT  11.72 39.0325 11.79 39.2325 ;
        RECT  11.72 38.5675 11.79 38.7025 ;
        RECT  11.72 38.5675 11.79 38.7025 ;
        RECT  10.96 37.8875 11.845 37.9525 ;
        RECT  11.535 38.4025 11.71 38.4675 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  11.205 38.4025 11.27 39.1425 ;
        RECT  11.3425 39.235 11.4425 39.2975 ;
        RECT  10.965 38.03 11.0175 38.0925 ;
        RECT  11.72 38.5675 11.79 38.7025 ;
        RECT  10.96 39.2325 11.845 39.2975 ;
        RECT  11.535 38.4025 11.6 39.0325 ;
        RECT  11.72 38.5675 11.79 38.7025 ;
        RECT  11.72 38.5675 11.79 38.7025 ;
        RECT  11.1 38.1775 11.17 38.4675 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  10.96 38.0275 11.845 38.0925 ;
        RECT  11.72 38.5675 11.79 38.7025 ;
        RECT  11.72 39.0325 11.79 39.2325 ;
        RECT  11.015 39.0325 11.085 39.2325 ;
        RECT  11.64 38.1775 11.71 38.4675 ;
        RECT  11.1 38.4025 11.27 38.4675 ;
        RECT  10.96 38.0275 11.845 38.0925 ;
        RECT  10.96 37.8875 11.845 37.9525 ;
        RECT  10.96 39.2325 11.845 39.2975 ;
        RECT  11.72 39.3625 11.785 39.4975 ;
        RECT  11.535 39.3625 11.6 39.4975 ;
        RECT  11.02 39.3625 11.085 39.4975 ;
        RECT  11.205 39.3625 11.27 39.4975 ;
        RECT  11.535 39.8275 11.6 39.9625 ;
        RECT  11.72 39.8275 11.785 39.9625 ;
        RECT  11.205 39.8275 11.27 39.9625 ;
        RECT  11.02 39.8275 11.085 39.9625 ;
        RECT  11.64 40.2175 11.705 40.3525 ;
        RECT  11.455 40.2175 11.52 40.3525 ;
        RECT  11.285 40.2175 11.35 40.3525 ;
        RECT  11.1 40.2175 11.165 40.3525 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.33 39.2325 11.465 39.2975 ;
        RECT  10.9825 40.5775 11.1175 40.6425 ;
        RECT  11.6875 40.5775 11.8225 40.6425 ;
        RECT  11.3175 40.4375 11.4525 40.5025 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.2225 39.5475 11.3575 39.6125 ;
        RECT  11.2225 39.5475 11.3575 39.6125 ;
        RECT  11.4475 39.6975 11.5825 39.7625 ;
        RECT  11.4475 39.6975 11.5825 39.7625 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.2725 40.2175 11.3375 40.3525 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.4675 40.2175 11.5325 40.3525 ;
        RECT  11.335 40.5775 11.47 40.6425 ;
        RECT  11.335 40.5775 11.47 40.6425 ;
        RECT  11.6875 40.5775 11.8225 40.6425 ;
        RECT  11.33 39.2325 11.465 39.2975 ;
        RECT  11.6875 40.5775 11.8225 40.6425 ;
        RECT  11.6875 40.5775 11.8225 40.6425 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  10.9825 40.5775 11.1175 40.6425 ;
        RECT  11.3425 39.235 11.4425 39.2975 ;
        RECT  11.3425 39.2325 11.4425 39.295 ;
        RECT  11.67 40.4375 11.7225 40.5 ;
        RECT  11.3425 39.235 11.4425 39.2975 ;
        RECT  11.72 39.2975 11.79 39.4975 ;
        RECT  11.72 39.8275 11.79 39.9625 ;
        RECT  11.72 39.8275 11.79 39.9625 ;
        RECT  10.96 40.5775 11.845 40.6425 ;
        RECT  11.535 40.0625 11.71 40.1275 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  11.205 39.3875 11.27 40.1275 ;
        RECT  11.3425 39.2325 11.4425 39.295 ;
        RECT  10.965 40.4375 11.0175 40.5 ;
        RECT  11.72 39.8275 11.79 39.9625 ;
        RECT  10.96 39.2325 11.845 39.2975 ;
        RECT  11.535 39.4975 11.6 40.1275 ;
        RECT  11.72 39.8275 11.79 39.9625 ;
        RECT  11.72 39.8275 11.79 39.9625 ;
        RECT  11.1 40.0625 11.17 40.3525 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  10.96 40.4375 11.845 40.5025 ;
        RECT  11.72 39.8275 11.79 39.9625 ;
        RECT  11.72 39.2975 11.79 39.4975 ;
        RECT  11.015 39.2975 11.085 39.4975 ;
        RECT  11.64 40.0625 11.71 40.3525 ;
        RECT  11.1 40.0625 11.27 40.1275 ;
        RECT  10.96 40.4375 11.845 40.5025 ;
        RECT  10.96 40.5775 11.845 40.6425 ;
        RECT  10.96 39.2325 11.845 39.2975 ;
        RECT  10.345 41.4775 11.755 41.5425 ;
        RECT  10.345 42.205 11.755 42.27 ;
        RECT  10.6975 41.7675 10.7625 42.27 ;
        RECT  10.345 42.205 11.05 42.27 ;
        RECT  10.345 41.4775 11.05 41.5425 ;
        RECT  10.5075 41.1825 10.5725 41.3175 ;
        RECT  10.6975 41.1825 10.7625 41.3175 ;
        RECT  10.5075 41.1825 10.5725 41.3175 ;
        RECT  10.6975 41.1825 10.7625 41.3175 ;
        RECT  10.5075 41.7675 10.5725 41.9025 ;
        RECT  10.6975 41.7675 10.7625 41.9025 ;
        RECT  10.5075 41.7675 10.5725 41.9025 ;
        RECT  10.6975 41.7675 10.7625 41.9025 ;
        RECT  10.6975 41.7675 10.7625 41.9025 ;
        RECT  10.8875 41.7675 10.9525 41.9025 ;
        RECT  10.6975 41.7675 10.7625 41.9025 ;
        RECT  10.8875 41.7675 10.9525 41.9025 ;
        RECT  10.5425 41.4775 10.6775 41.5425 ;
        RECT  10.6975 42.0675 10.7625 42.2025 ;
        RECT  10.5075 41.1825 10.5725 41.3175 ;
        RECT  10.6975 41.1825 10.7625 41.3175 ;
        RECT  10.5075 41.7675 10.5725 41.9025 ;
        RECT  10.8875 41.7675 10.9525 41.9025 ;
        RECT  10.5075 41.1825 10.5725 41.3175 ;
        RECT  10.6975 41.1825 10.7625 41.3175 ;
        RECT  10.5075 41.7675 10.5725 41.9025 ;
        RECT  10.8875 41.7675 10.9525 41.9025 ;
        RECT  11.4025 41.7675 11.4675 42.27 ;
        RECT  11.05 42.205 11.755 42.27 ;
        RECT  11.05 41.4775 11.755 41.5425 ;
        RECT  11.2125 41.1825 11.2775 41.3175 ;
        RECT  11.4025 41.1825 11.4675 41.3175 ;
        RECT  11.2125 41.1825 11.2775 41.3175 ;
        RECT  11.4025 41.1825 11.4675 41.3175 ;
        RECT  11.2125 41.7675 11.2775 41.9025 ;
        RECT  11.4025 41.7675 11.4675 41.9025 ;
        RECT  11.2125 41.7675 11.2775 41.9025 ;
        RECT  11.4025 41.7675 11.4675 41.9025 ;
        RECT  11.4025 41.7675 11.4675 41.9025 ;
        RECT  11.5925 41.7675 11.6575 41.9025 ;
        RECT  11.4025 41.7675 11.4675 41.9025 ;
        RECT  11.5925 41.7675 11.6575 41.9025 ;
        RECT  11.2475 41.4775 11.3825 41.5425 ;
        RECT  11.4025 42.0675 11.4675 42.2025 ;
        RECT  11.2125 41.1825 11.2775 41.3175 ;
        RECT  11.4025 41.1825 11.4675 41.3175 ;
        RECT  11.2125 41.7675 11.2775 41.9025 ;
        RECT  11.5925 41.7675 11.6575 41.9025 ;
        RECT  11.2125 41.1825 11.2775 41.3175 ;
        RECT  11.4025 41.1825 11.4675 41.3175 ;
        RECT  11.2125 41.7675 11.2775 41.9025 ;
        RECT  11.5925 41.7675 11.6575 41.9025 ;
        RECT  10.345 14.3225 11.755 14.3875 ;
        RECT  10.345 18.895 11.755 18.96 ;
        RECT  10.345 14.4525 11.755 14.5175 ;
        RECT  10.31 14.3225 11.085 14.3875 ;
        RECT  10.8525 15.3925 10.9175 16.255 ;
        RECT  10.4775 15.3875 10.5425 16.255 ;
        RECT  10.4775 15.4925 10.7675 15.5575 ;
        RECT  10.6275 15.6925 10.9175 15.7575 ;
        RECT  10.31 18.895 11.085 18.96 ;
        RECT  10.4775 16.4175 10.5425 17.515 ;
        RECT  10.8525 16.415 10.9175 16.61 ;
        RECT  10.31 14.4525 11.085 14.5175 ;
        RECT  10.6275 14.8475 10.6975 15.175 ;
        RECT  10.6675 16.545 10.9175 16.61 ;
        RECT  10.6675 16.545 10.7325 16.74 ;
        RECT  10.4775 17.515 10.975 17.58 ;
        RECT  10.665 17.515 10.73 17.7125 ;
        RECT  10.6575 18.6925 10.975 18.7625 ;
        RECT  10.9375 14.4525 11.0025 14.6825 ;
        RECT  10.7625 14.5175 10.8275 14.67 ;
        RECT  10.4075 18.895 10.475 18.96 ;
        RECT  10.91 17.515 10.975 18.7625 ;
        RECT  10.4075 18.5575 10.765 18.6225 ;
        RECT  10.4075 18.6225 10.475 18.96 ;
        RECT  11.0025 14.5175 11.0175 14.5875 ;
        RECT  10.575 14.3225 10.64 14.3875 ;
        RECT  10.615 14.4525 10.675 14.5175 ;
        RECT  10.7225 15.4575 10.7875 15.5925 ;
        RECT  10.6075 15.6575 10.6725 15.7925 ;
        RECT  10.665 16.345 10.73 16.48 ;
        RECT  10.665 18.4875 10.73 18.6225 ;
        RECT  10.63 18.5575 10.765 18.6225 ;
        RECT  10.4725 17.645 10.5375 17.78 ;
        RECT  10.9375 14.6825 11.0025 14.8175 ;
        RECT  10.855 17.235 10.92 17.37 ;
        RECT  10.3125 14.4525 10.3775 14.5875 ;
        RECT  11.0175 14.4525 11.0825 14.5875 ;
        RECT  10.635 14.3225 10.77 14.3875 ;
        RECT  10.66 18.6925 10.725 18.8275 ;
        RECT  10.6675 16.675 10.7325 17.37 ;
        RECT  10.8525 16.675 10.9175 17.37 ;
        RECT  10.4775 17.645 10.5425 18.34 ;
        RECT  10.6625 17.645 10.7275 18.34 ;
        RECT  10.6675 15.8625 10.7325 16.4175 ;
        RECT  10.8525 15.8625 10.9175 16.4175 ;
        RECT  10.4775 15.8625 10.5425 16.4175 ;
        RECT  10.6625 15.8625 10.7275 16.4175 ;
        RECT  10.5775 14.66 10.6425 14.935 ;
        RECT  10.7625 14.66 10.8275 14.935 ;
        RECT  10.4775 15.1175 10.5425 15.3925 ;
        RECT  10.6625 15.1175 10.7275 15.3925 ;
        RECT  10.6675 15.1175 10.7325 15.3925 ;
        RECT  10.8525 15.1175 10.9175 15.3925 ;
        RECT  10.31 14.3225 11.085 14.3875 ;
        RECT  10.31 18.895 11.085 18.96 ;
        RECT  10.31 14.4525 11.085 14.5175 ;
        RECT  11.015 14.3225 11.79 14.3875 ;
        RECT  11.5575 15.3925 11.6225 16.255 ;
        RECT  11.1825 15.3875 11.2475 16.255 ;
        RECT  11.1825 15.4925 11.4725 15.5575 ;
        RECT  11.3325 15.6925 11.6225 15.7575 ;
        RECT  11.015 18.895 11.79 18.96 ;
        RECT  11.1825 16.4175 11.2475 17.515 ;
        RECT  11.5575 16.415 11.6225 16.61 ;
        RECT  11.015 14.4525 11.79 14.5175 ;
        RECT  11.3325 14.8475 11.4025 15.175 ;
        RECT  11.3725 16.545 11.6225 16.61 ;
        RECT  11.3725 16.545 11.4375 16.74 ;
        RECT  11.1825 17.515 11.68 17.58 ;
        RECT  11.37 17.515 11.435 17.7125 ;
        RECT  11.3625 18.6925 11.68 18.7625 ;
        RECT  11.6425 14.4525 11.7075 14.6825 ;
        RECT  11.4675 14.5175 11.5325 14.67 ;
        RECT  11.1125 18.895 11.18 18.96 ;
        RECT  11.615 17.515 11.68 18.7625 ;
        RECT  11.1125 18.5575 11.47 18.6225 ;
        RECT  11.1125 18.6225 11.18 18.96 ;
        RECT  11.7075 14.5175 11.7225 14.5875 ;
        RECT  11.28 14.3225 11.345 14.3875 ;
        RECT  11.32 14.4525 11.38 14.5175 ;
        RECT  11.4275 15.4575 11.4925 15.5925 ;
        RECT  11.3125 15.6575 11.3775 15.7925 ;
        RECT  11.37 16.345 11.435 16.48 ;
        RECT  11.37 18.4875 11.435 18.6225 ;
        RECT  11.335 18.5575 11.47 18.6225 ;
        RECT  11.1775 17.645 11.2425 17.78 ;
        RECT  11.6425 14.6825 11.7075 14.8175 ;
        RECT  11.56 17.235 11.625 17.37 ;
        RECT  11.0175 14.4525 11.0825 14.5875 ;
        RECT  11.7225 14.4525 11.7875 14.5875 ;
        RECT  11.34 14.3225 11.475 14.3875 ;
        RECT  11.365 18.6925 11.43 18.8275 ;
        RECT  11.3725 16.675 11.4375 17.37 ;
        RECT  11.5575 16.675 11.6225 17.37 ;
        RECT  11.1825 17.645 11.2475 18.34 ;
        RECT  11.3675 17.645 11.4325 18.34 ;
        RECT  11.3725 15.8625 11.4375 16.4175 ;
        RECT  11.5575 15.8625 11.6225 16.4175 ;
        RECT  11.1825 15.8625 11.2475 16.4175 ;
        RECT  11.3675 15.8625 11.4325 16.4175 ;
        RECT  11.2825 14.66 11.3475 14.935 ;
        RECT  11.4675 14.66 11.5325 14.935 ;
        RECT  11.1825 15.1175 11.2475 15.3925 ;
        RECT  11.3675 15.1175 11.4325 15.3925 ;
        RECT  11.3725 15.1175 11.4375 15.3925 ;
        RECT  11.5575 15.1175 11.6225 15.3925 ;
        RECT  11.015 14.3225 11.79 14.3875 ;
        RECT  11.015 18.895 11.79 18.96 ;
        RECT  11.015 14.4525 11.79 14.5175 ;
        RECT  10.345 10.2975 11.755 10.3625 ;
        RECT  10.345 10.4275 11.755 10.4925 ;
        RECT  10.345 11.23 11.755 11.295 ;
        RECT  10.765 13.6925 10.83 13.8275 ;
        RECT  10.39 13.6925 10.455 13.8275 ;
        RECT  10.39 11.765 10.455 11.9 ;
        RECT  10.765 11.765 10.83 11.9 ;
        RECT  10.765 12.8975 10.83 13.3125 ;
        RECT  10.39 12.8975 10.455 13.3125 ;
        RECT  10.39 12.28 10.455 12.695 ;
        RECT  10.765 12.28 10.83 12.695 ;
        RECT  10.575 10.71 10.64 11.125 ;
        RECT  10.39 10.71 10.455 11.125 ;
        RECT  10.73 10.71 10.795 11.125 ;
        RECT  10.915 10.71 10.98 11.125 ;
        RECT  10.575 11.4 10.64 11.535 ;
        RECT  10.39 11.4 10.455 11.535 ;
        RECT  10.73 11.4 10.795 11.535 ;
        RECT  10.915 11.4 10.98 11.535 ;
        RECT  10.5525 10.165 10.6875 10.23 ;
        RECT  10.6275 12.12 10.6925 12.255 ;
        RECT  11.0175 11.765 11.0825 11.9 ;
        RECT  10.93 11.765 10.995 11.9 ;
        RECT  10.3125 12.7275 10.3775 12.8625 ;
        RECT  11.0175 11.195 11.0825 11.33 ;
        RECT  10.3125 11.195 10.3775 11.33 ;
        RECT  10.7325 11.4 10.7975 11.535 ;
        RECT  11.0175 13.6925 11.0825 13.8275 ;
        RECT  10.9325 13.6925 10.9975 13.8275 ;
        RECT  10.7325 10.99 10.7975 11.125 ;
        RECT  10.5925 10.99 10.6575 11.125 ;
        RECT  10.615 10.5775 10.75 10.6425 ;
        RECT  10.4475 10.1675 10.5825 10.2325 ;
        RECT  10.7875 10.2975 10.9225 10.3625 ;
        RECT  11.0175 11.4 11.0825 11.535 ;
        RECT  10.3125 11.4 10.3775 11.535 ;
        RECT  10.45 10.4275 10.585 10.4925 ;
        RECT  10.5925 13.37 10.6575 13.505 ;
        RECT  10.7625 11.765 10.8275 11.9 ;
        RECT  10.4525 12.68 10.5175 12.815 ;
        RECT  10.5925 11.4 10.6575 11.535 ;
        RECT  10.53 13.37 10.595 13.505 ;
        RECT  10.3125 11.765 10.3775 11.9 ;
        RECT  10.7625 12.28 10.8275 12.415 ;
        RECT  10.4975 13.9025 10.5625 14.0375 ;
        RECT  10.3125 13.6925 10.3775 13.8275 ;
        RECT  10.9975 13.6925 11.0175 13.8275 ;
        RECT  10.995 11.765 11.0175 11.9 ;
        RECT  10.665 11.2325 10.7225 11.2925 ;
        RECT  10.64 10.2975 10.7125 10.3625 ;
        RECT  10.6425 10.4275 10.7125 10.4925 ;
        RECT  10.3725 13.6925 10.385 13.8275 ;
        RECT  10.3775 12.7275 10.52 12.8625 ;
        RECT  10.31 11.23 11.085 11.295 ;
        RECT  10.6475 10.4925 10.7125 10.6425 ;
        RECT  10.975 11.4 11.0175 11.535 ;
        RECT  10.915 10.4925 10.98 10.71 ;
        RECT  10.39 10.4925 10.455 10.71 ;
        RECT  10.31 10.4275 11.085 10.4925 ;
        RECT  10.31 10.2975 11.085 10.3625 ;
        RECT  10.3725 11.4 10.385 11.535 ;
        RECT  10.44 12.68 10.455 12.815 ;
        RECT  10.3725 11.765 10.385 11.9 ;
        RECT  10.39 12.695 10.455 12.8975 ;
        RECT  10.765 13.8275 10.83 13.9025 ;
        RECT  10.6275 11.6075 10.79 11.6725 ;
        RECT  10.38 13.6925 10.39 13.8275 ;
        RECT  10.38 11.765 10.39 11.9 ;
        RECT  10.725 11.4825 10.79 11.6075 ;
        RECT  10.6275 11.6075 10.6925 12.205 ;
        RECT  10.765 13.3125 10.83 13.6925 ;
        RECT  10.495 13.9025 10.83 13.9675 ;
        RECT  10.38 11.4 10.39 11.535 ;
        RECT  10.31 10.2975 11.085 10.3625 ;
        RECT  10.31 10.4275 11.085 10.4925 ;
        RECT  10.31 11.23 11.085 11.295 ;
        RECT  11.47 13.6925 11.535 13.8275 ;
        RECT  11.095 13.6925 11.16 13.8275 ;
        RECT  11.095 11.765 11.16 11.9 ;
        RECT  11.47 11.765 11.535 11.9 ;
        RECT  11.47 12.8975 11.535 13.3125 ;
        RECT  11.095 12.8975 11.16 13.3125 ;
        RECT  11.095 12.28 11.16 12.695 ;
        RECT  11.47 12.28 11.535 12.695 ;
        RECT  11.28 10.71 11.345 11.125 ;
        RECT  11.095 10.71 11.16 11.125 ;
        RECT  11.435 10.71 11.5 11.125 ;
        RECT  11.62 10.71 11.685 11.125 ;
        RECT  11.28 11.4 11.345 11.535 ;
        RECT  11.095 11.4 11.16 11.535 ;
        RECT  11.435 11.4 11.5 11.535 ;
        RECT  11.62 11.4 11.685 11.535 ;
        RECT  11.2575 10.165 11.3925 10.23 ;
        RECT  11.3325 12.12 11.3975 12.255 ;
        RECT  11.7225 11.765 11.7875 11.9 ;
        RECT  11.635 11.765 11.7 11.9 ;
        RECT  11.0175 12.7275 11.0825 12.8625 ;
        RECT  11.7225 11.195 11.7875 11.33 ;
        RECT  11.0175 11.195 11.0825 11.33 ;
        RECT  11.4375 11.4 11.5025 11.535 ;
        RECT  11.7225 13.6925 11.7875 13.8275 ;
        RECT  11.6375 13.6925 11.7025 13.8275 ;
        RECT  11.4375 10.99 11.5025 11.125 ;
        RECT  11.2975 10.99 11.3625 11.125 ;
        RECT  11.32 10.5775 11.455 10.6425 ;
        RECT  11.1525 10.1675 11.2875 10.2325 ;
        RECT  11.4925 10.2975 11.6275 10.3625 ;
        RECT  11.7225 11.4 11.7875 11.535 ;
        RECT  11.0175 11.4 11.0825 11.535 ;
        RECT  11.155 10.4275 11.29 10.4925 ;
        RECT  11.2975 13.37 11.3625 13.505 ;
        RECT  11.4675 11.765 11.5325 11.9 ;
        RECT  11.1575 12.68 11.2225 12.815 ;
        RECT  11.2975 11.4 11.3625 11.535 ;
        RECT  11.235 13.37 11.3 13.505 ;
        RECT  11.0175 11.765 11.0825 11.9 ;
        RECT  11.4675 12.28 11.5325 12.415 ;
        RECT  11.2025 13.9025 11.2675 14.0375 ;
        RECT  11.0175 13.6925 11.0825 13.8275 ;
        RECT  11.7025 13.6925 11.7225 13.8275 ;
        RECT  11.7 11.765 11.7225 11.9 ;
        RECT  11.37 11.2325 11.4275 11.2925 ;
        RECT  11.345 10.2975 11.4175 10.3625 ;
        RECT  11.3475 10.4275 11.4175 10.4925 ;
        RECT  11.0775 13.6925 11.09 13.8275 ;
        RECT  11.0825 12.7275 11.225 12.8625 ;
        RECT  11.015 11.23 11.79 11.295 ;
        RECT  11.3525 10.4925 11.4175 10.6425 ;
        RECT  11.68 11.4 11.7225 11.535 ;
        RECT  11.62 10.4925 11.685 10.71 ;
        RECT  11.095 10.4925 11.16 10.71 ;
        RECT  11.015 10.4275 11.79 10.4925 ;
        RECT  11.015 10.2975 11.79 10.3625 ;
        RECT  11.0775 11.4 11.09 11.535 ;
        RECT  11.145 12.68 11.16 12.815 ;
        RECT  11.0775 11.765 11.09 11.9 ;
        RECT  11.095 12.695 11.16 12.8975 ;
        RECT  11.47 13.8275 11.535 13.9025 ;
        RECT  11.3325 11.6075 11.495 11.6725 ;
        RECT  11.085 13.6925 11.095 13.8275 ;
        RECT  11.085 11.765 11.095 11.9 ;
        RECT  11.43 11.4825 11.495 11.6075 ;
        RECT  11.3325 11.6075 11.3975 12.205 ;
        RECT  11.47 13.3125 11.535 13.6925 ;
        RECT  11.2 13.9025 11.535 13.9675 ;
        RECT  11.085 11.4 11.095 11.535 ;
        RECT  11.015 10.2975 11.79 10.3625 ;
        RECT  11.015 10.4275 11.79 10.4925 ;
        RECT  11.015 11.23 11.79 11.295 ;
        RECT  10.345 3.795 11.755 3.86 ;
        RECT  10.345 6.8 11.755 6.865 ;
        RECT  10.345 9.76 11.755 9.825 ;
        RECT  10.345 4.81 11.755 4.875 ;
        RECT  10.345 7.77 11.755 7.835 ;
        RECT  10.345 3.955 11.755 4.02 ;
        RECT  10.885 6.28 10.95 6.415 ;
        RECT  10.7 6.28 10.765 6.415 ;
        RECT  10.885 5.045 10.95 5.18 ;
        RECT  10.7 5.045 10.765 5.18 ;
        RECT  10.695 6.28 10.76 6.415 ;
        RECT  10.51 6.28 10.575 6.415 ;
        RECT  10.695 9.24 10.76 9.375 ;
        RECT  10.51 9.24 10.575 9.375 ;
        RECT  10.695 5.045 10.76 5.18 ;
        RECT  10.51 5.045 10.575 5.18 ;
        RECT  10.885 9.24 10.95 9.375 ;
        RECT  10.7 9.24 10.765 9.375 ;
        RECT  10.695 4.51 10.76 4.645 ;
        RECT  10.51 4.51 10.575 4.645 ;
        RECT  10.835 7.47 10.9 7.605 ;
        RECT  10.65 7.47 10.715 7.605 ;
        RECT  10.885 8.005 10.95 8.14 ;
        RECT  10.7 8.005 10.765 8.14 ;
        RECT  10.695 8.005 10.76 8.14 ;
        RECT  10.51 8.005 10.575 8.14 ;
        RECT  10.885 8.43 10.95 8.565 ;
        RECT  10.7 8.43 10.765 8.565 ;
        RECT  10.885 5.47 10.95 5.605 ;
        RECT  10.7 5.47 10.765 5.605 ;
        RECT  10.885 8.815 10.95 8.95 ;
        RECT  10.7 8.815 10.765 8.95 ;
        RECT  10.695 8.815 10.76 8.95 ;
        RECT  10.51 8.815 10.575 8.95 ;
        RECT  10.695 5.47 10.76 5.605 ;
        RECT  10.51 5.47 10.575 5.605 ;
        RECT  10.695 8.43 10.76 8.565 ;
        RECT  10.51 8.43 10.575 8.565 ;
        RECT  10.695 5.855 10.76 5.99 ;
        RECT  10.51 5.855 10.575 5.99 ;
        RECT  10.885 5.855 10.95 5.99 ;
        RECT  10.7 5.855 10.765 5.99 ;
        RECT  10.695 4.085 10.76 4.22 ;
        RECT  10.51 4.085 10.575 4.22 ;
        RECT  10.77 7.06 10.835 7.195 ;
        RECT  10.585 7.06 10.65 7.195 ;
        RECT  10.5725 3.795 10.7075 3.86 ;
        RECT  10.51 9.2925 10.575 9.4275 ;
        RECT  10.4 7.4775 10.465 7.6125 ;
        RECT  10.51 6.5775 10.575 6.7125 ;
        RECT  10.9325 7.0525 10.9975 7.1875 ;
        RECT  10.51 9.6575 10.575 9.7925 ;
        RECT  11.0175 4.115 11.0825 4.25 ;
        RECT  10.875 8.1975 10.94 8.3325 ;
        RECT  10.8775 6.59 10.9425 6.725 ;
        RECT  10.8775 5.1925 10.9425 5.3275 ;
        RECT  10.3125 3.975 10.3775 4.11 ;
        RECT  10.8875 4.0925 10.9525 4.2275 ;
        RECT  10.8875 5.7025 11.0225 5.7675 ;
        RECT  10.9275 4.6175 10.9925 4.7525 ;
        RECT  10.8875 8.6625 11.0225 8.7275 ;
        RECT  10.835 9.55 10.9 9.685 ;
        RECT  10.755 6.08 10.82 6.215 ;
        RECT  10.745 9.04 10.81 9.175 ;
        RECT  10.5125 7.35 10.6475 7.415 ;
        RECT  11.0175 7.0525 11.0825 7.1875 ;
        RECT  10.4025 4.345 10.5375 4.41 ;
        RECT  10.5125 5.8575 10.5775 5.9925 ;
        RECT  10.8775 9.55 10.9425 9.685 ;
        RECT  10.7 9.04 10.765 9.175 ;
        RECT  11.0175 8.6275 11.0825 8.7625 ;
        RECT  11.0175 3.925 11.0825 4.06 ;
        RECT  10.8775 6.59 10.9425 6.725 ;
        RECT  11.0175 5.6675 11.0825 5.8025 ;
        RECT  10.5125 5.4675 10.5775 5.6025 ;
        RECT  10.7 5.4675 10.765 5.6025 ;
        RECT  10.7 6.08 10.765 6.215 ;
        RECT  10.51 8.4275 10.575 8.5625 ;
        RECT  10.7 8.4275 10.765 8.5625 ;
        RECT  10.31 3.795 11.085 3.86 ;
        RECT  10.38 6.865 10.445 9.76 ;
        RECT  10.885 9.375 10.95 9.685 ;
        RECT  10.51 8.95 10.575 9.24 ;
        RECT  10.51 8.14 10.575 8.43 ;
        RECT  10.65 9.7625 10.7225 9.825 ;
        RECT  10.695 9.375 10.765 9.76 ;
        RECT  10.695 8.14 10.765 8.43 ;
        RECT  10.695 8.66 10.765 8.8175 ;
        RECT  10.885 8.95 10.95 9.24 ;
        RECT  10.885 8.14 10.95 8.43 ;
        RECT  10.695 8.66 11.08 8.73 ;
        RECT  10.31 9.76 11.085 9.825 ;
        RECT  10.31 7.77 11.085 7.835 ;
        RECT  10.38 4.875 10.445 6.8 ;
        RECT  10.885 6.415 10.95 6.725 ;
        RECT  10.51 5.99 10.575 6.28 ;
        RECT  10.585 7.155 10.65 7.605 ;
        RECT  10.695 6.415 10.765 6.8 ;
        RECT  10.695 5.7 10.765 5.8575 ;
        RECT  10.51 6.7125 10.575 6.8 ;
        RECT  10.885 5.99 10.95 6.28 ;
        RECT  10.77 6.93 11.015 6.995 ;
        RECT  10.9325 6.93 11.015 7.0525 ;
        RECT  10.9525 7.0525 11.02 7.1875 ;
        RECT  10.31 6.8 11.085 6.865 ;
        RECT  10.51 5.18 10.575 5.47 ;
        RECT  10.695 4.6425 10.76 4.81 ;
        RECT  10.76 4.15 11.0175 4.22 ;
        RECT  10.51 4.085 10.575 4.51 ;
        RECT  10.695 5.18 10.765 5.47 ;
        RECT  10.4025 4.34 10.575 4.415 ;
        RECT  10.885 5.18 10.95 5.47 ;
        RECT  10.8875 4.02 10.9525 4.0925 ;
        RECT  10.695 5.7 11.08 5.77 ;
        RECT  10.9275 4.73 10.9925 4.845 ;
        RECT  10.31 3.955 11.085 4.02 ;
        RECT  10.31 4.81 11.085 4.875 ;
        RECT  10.45 3.8 10.515 3.8575 ;
        RECT  11.0175 4.04 11.0825 4.1625 ;
        RECT  10.835 7.6025 10.9 7.77 ;
        RECT  10.77 6.995 10.8375 7.0975 ;
        RECT  10.31 3.795 11.085 3.86 ;
        RECT  10.31 6.8 11.085 6.865 ;
        RECT  10.31 9.76 11.085 9.825 ;
        RECT  10.31 4.81 11.085 4.875 ;
        RECT  10.31 7.77 11.085 7.835 ;
        RECT  10.31 3.955 11.085 4.02 ;
        RECT  11.15 6.28 11.215 6.415 ;
        RECT  11.335 6.28 11.4 6.415 ;
        RECT  11.15 5.045 11.215 5.18 ;
        RECT  11.335 5.045 11.4 5.18 ;
        RECT  11.34 6.28 11.405 6.415 ;
        RECT  11.525 6.28 11.59 6.415 ;
        RECT  11.34 9.24 11.405 9.375 ;
        RECT  11.525 9.24 11.59 9.375 ;
        RECT  11.34 5.045 11.405 5.18 ;
        RECT  11.525 5.045 11.59 5.18 ;
        RECT  11.15 9.24 11.215 9.375 ;
        RECT  11.335 9.24 11.4 9.375 ;
        RECT  11.34 4.51 11.405 4.645 ;
        RECT  11.525 4.51 11.59 4.645 ;
        RECT  11.2 7.47 11.265 7.605 ;
        RECT  11.385 7.47 11.45 7.605 ;
        RECT  11.15 8.005 11.215 8.14 ;
        RECT  11.335 8.005 11.4 8.14 ;
        RECT  11.34 8.005 11.405 8.14 ;
        RECT  11.525 8.005 11.59 8.14 ;
        RECT  11.15 8.43 11.215 8.565 ;
        RECT  11.335 8.43 11.4 8.565 ;
        RECT  11.15 5.47 11.215 5.605 ;
        RECT  11.335 5.47 11.4 5.605 ;
        RECT  11.15 8.815 11.215 8.95 ;
        RECT  11.335 8.815 11.4 8.95 ;
        RECT  11.34 8.815 11.405 8.95 ;
        RECT  11.525 8.815 11.59 8.95 ;
        RECT  11.34 5.47 11.405 5.605 ;
        RECT  11.525 5.47 11.59 5.605 ;
        RECT  11.34 8.43 11.405 8.565 ;
        RECT  11.525 8.43 11.59 8.565 ;
        RECT  11.34 5.855 11.405 5.99 ;
        RECT  11.525 5.855 11.59 5.99 ;
        RECT  11.15 5.855 11.215 5.99 ;
        RECT  11.335 5.855 11.4 5.99 ;
        RECT  11.34 4.085 11.405 4.22 ;
        RECT  11.525 4.085 11.59 4.22 ;
        RECT  11.265 7.06 11.33 7.195 ;
        RECT  11.45 7.06 11.515 7.195 ;
        RECT  11.3925 3.795 11.5275 3.86 ;
        RECT  11.525 9.2925 11.59 9.4275 ;
        RECT  11.635 7.4775 11.7 7.6125 ;
        RECT  11.525 6.5775 11.59 6.7125 ;
        RECT  11.1025 7.0525 11.1675 7.1875 ;
        RECT  11.525 9.6575 11.59 9.7925 ;
        RECT  11.0175 4.115 11.0825 4.25 ;
        RECT  11.16 8.1975 11.225 8.3325 ;
        RECT  11.1575 6.59 11.2225 6.725 ;
        RECT  11.1575 5.1925 11.2225 5.3275 ;
        RECT  11.7225 3.975 11.7875 4.11 ;
        RECT  11.1475 4.0925 11.2125 4.2275 ;
        RECT  11.0775 5.7025 11.2125 5.7675 ;
        RECT  11.1075 4.6175 11.1725 4.7525 ;
        RECT  11.0775 8.6625 11.2125 8.7275 ;
        RECT  11.2 9.55 11.265 9.685 ;
        RECT  11.28 6.08 11.345 6.215 ;
        RECT  11.29 9.04 11.355 9.175 ;
        RECT  11.4525 7.35 11.5875 7.415 ;
        RECT  11.0175 7.0525 11.0825 7.1875 ;
        RECT  11.5625 4.345 11.6975 4.41 ;
        RECT  11.5225 5.8575 11.5875 5.9925 ;
        RECT  11.1575 9.55 11.2225 9.685 ;
        RECT  11.335 9.04 11.4 9.175 ;
        RECT  11.0175 8.6275 11.0825 8.7625 ;
        RECT  11.0175 3.925 11.0825 4.06 ;
        RECT  11.1575 6.59 11.2225 6.725 ;
        RECT  11.0175 5.6675 11.0825 5.8025 ;
        RECT  11.5225 5.4675 11.5875 5.6025 ;
        RECT  11.335 5.4675 11.4 5.6025 ;
        RECT  11.335 6.08 11.4 6.215 ;
        RECT  11.525 8.4275 11.59 8.5625 ;
        RECT  11.335 8.4275 11.4 8.5625 ;
        RECT  11.015 3.795 11.79 3.86 ;
        RECT  11.655 6.865 11.72 9.76 ;
        RECT  11.15 9.375 11.215 9.685 ;
        RECT  11.525 8.95 11.59 9.24 ;
        RECT  11.525 8.14 11.59 8.43 ;
        RECT  11.3775 9.7625 11.45 9.825 ;
        RECT  11.335 9.375 11.405 9.76 ;
        RECT  11.335 8.14 11.405 8.43 ;
        RECT  11.335 8.66 11.405 8.8175 ;
        RECT  11.15 8.95 11.215 9.24 ;
        RECT  11.15 8.14 11.215 8.43 ;
        RECT  11.02 8.66 11.405 8.73 ;
        RECT  11.015 9.76 11.79 9.825 ;
        RECT  11.015 7.77 11.79 7.835 ;
        RECT  11.655 4.875 11.72 6.8 ;
        RECT  11.15 6.415 11.215 6.725 ;
        RECT  11.525 5.99 11.59 6.28 ;
        RECT  11.45 7.155 11.515 7.605 ;
        RECT  11.335 6.415 11.405 6.8 ;
        RECT  11.335 5.7 11.405 5.8575 ;
        RECT  11.525 6.7125 11.59 6.8 ;
        RECT  11.15 5.99 11.215 6.28 ;
        RECT  11.085 6.93 11.33 6.995 ;
        RECT  11.085 6.93 11.1675 7.0525 ;
        RECT  11.08 7.0525 11.1475 7.1875 ;
        RECT  11.015 6.8 11.79 6.865 ;
        RECT  11.525 5.18 11.59 5.47 ;
        RECT  11.34 4.6425 11.405 4.81 ;
        RECT  11.0825 4.15 11.34 4.22 ;
        RECT  11.525 4.085 11.59 4.51 ;
        RECT  11.335 5.18 11.405 5.47 ;
        RECT  11.525 4.34 11.6975 4.415 ;
        RECT  11.15 5.18 11.215 5.47 ;
        RECT  11.1475 4.02 11.2125 4.0925 ;
        RECT  11.02 5.7 11.405 5.77 ;
        RECT  11.1075 4.73 11.1725 4.845 ;
        RECT  11.015 3.955 11.79 4.02 ;
        RECT  11.015 4.81 11.79 4.875 ;
        RECT  11.585 3.8 11.65 3.8575 ;
        RECT  11.0175 4.04 11.0825 4.1625 ;
        RECT  11.2 7.6025 11.265 7.77 ;
        RECT  11.2625 6.995 11.33 7.0975 ;
        RECT  11.015 3.795 11.79 3.86 ;
        RECT  11.015 6.8 11.79 6.865 ;
        RECT  11.015 9.76 11.79 9.825 ;
        RECT  11.015 4.81 11.79 4.875 ;
        RECT  11.015 7.77 11.79 7.835 ;
        RECT  11.015 3.955 11.79 4.02 ;
        RECT  10.345 3.1575 11.755 3.2225 ;
        RECT  10.345 1.74 11.755 1.805 ;
        RECT  10.345 3.0275 11.755 3.0925 ;
        RECT  10.345 1.61 11.755 1.675 ;
        RECT  10.4875 5.375 10.5525 5.44 ;
        RECT  10.8275 5.2825 10.8925 5.375 ;
        RECT  10.345 5.375 11.085 5.44 ;
        RECT  10.345 5.505 11.085 5.57 ;
        RECT  10.72 6.1475 11.0175 6.2825 ;
        RECT  10.8275 4.1525 10.8925 4.24 ;
        RECT  10.345 4.0875 11.085 4.1525 ;
        RECT  10.345 3.9575 11.085 4.0225 ;
        RECT  10.7625 4.5075 10.8975 4.5725 ;
        RECT  10.4525 4.3525 10.5175 4.8675 ;
        RECT  10.515 5.765 10.58 6.285 ;
        RECT  10.6225 5.505 10.685 5.57 ;
        RECT  10.67 3.9575 10.7275 4.0225 ;
        RECT  10.6975 5.68 10.7625 5.815 ;
        RECT  10.49 5.9575 10.555 6.0925 ;
        RECT  10.785 5.375 10.92 5.44 ;
        RECT  10.7625 5.975 10.8975 6.04 ;
        RECT  11.0175 6.1475 11.0825 6.2825 ;
        RECT  10.7625 6.015 10.8975 6.08 ;
        RECT  10.5075 3.9575 10.6425 4.0225 ;
        RECT  10.4025 5.505 10.5375 5.57 ;
        RECT  11.0175 4.0875 11.0825 4.2225 ;
        RECT  10.785 4.0875 10.92 4.1525 ;
        RECT  10.63 5.375 10.765 5.44 ;
        RECT  10.865 6.1575 10.93 6.2925 ;
        RECT  10.8425 4.5075 10.9775 4.5725 ;
        RECT  10.4525 4.8675 10.5175 5.2825 ;
        RECT  10.8275 4.8675 10.8925 5.2825 ;
        RECT  10.4525 4.24 10.5175 4.375 ;
        RECT  10.8275 4.24 10.8925 4.375 ;
        RECT  10.515 6.15 10.58 6.285 ;
        RECT  10.7 6.15 10.765 6.285 ;
        RECT  10.515 5.635 10.58 5.77 ;
        RECT  10.7 5.635 10.765 5.77 ;
        RECT  10.345 3.9575 11.085 4.0225 ;
        RECT  10.345 5.375 11.085 5.44 ;
        RECT  10.345 4.0875 11.085 4.1525 ;
        RECT  10.345 5.505 11.085 5.57 ;
        RECT  10.4525 4.24 10.5175 4.375 ;
        RECT  11.1925 5.375 11.2575 5.44 ;
        RECT  11.5325 5.2825 11.5975 5.375 ;
        RECT  11.05 5.375 11.79 5.44 ;
        RECT  11.05 5.505 11.79 5.57 ;
        RECT  11.425 6.1475 11.7225 6.2825 ;
        RECT  11.5325 4.1525 11.5975 4.24 ;
        RECT  11.05 4.0875 11.79 4.1525 ;
        RECT  11.05 3.9575 11.79 4.0225 ;
        RECT  11.4675 4.5075 11.6025 4.5725 ;
        RECT  11.1575 4.3525 11.2225 4.8675 ;
        RECT  11.22 5.765 11.285 6.285 ;
        RECT  11.3275 5.505 11.39 5.57 ;
        RECT  11.375 3.9575 11.4325 4.0225 ;
        RECT  11.4025 5.68 11.4675 5.815 ;
        RECT  11.195 5.9575 11.26 6.0925 ;
        RECT  11.49 5.375 11.625 5.44 ;
        RECT  11.4675 5.975 11.6025 6.04 ;
        RECT  11.7225 6.1475 11.7875 6.2825 ;
        RECT  11.4675 6.015 11.6025 6.08 ;
        RECT  11.2125 3.9575 11.3475 4.0225 ;
        RECT  11.1075 5.505 11.2425 5.57 ;
        RECT  11.7225 4.0875 11.7875 4.2225 ;
        RECT  11.49 4.0875 11.625 4.1525 ;
        RECT  11.335 5.375 11.47 5.44 ;
        RECT  11.57 6.1575 11.635 6.2925 ;
        RECT  11.5475 4.5075 11.6825 4.5725 ;
        RECT  11.1575 4.8675 11.2225 5.2825 ;
        RECT  11.5325 4.8675 11.5975 5.2825 ;
        RECT  11.1575 4.24 11.2225 4.375 ;
        RECT  11.5325 4.24 11.5975 4.375 ;
        RECT  11.22 6.15 11.285 6.285 ;
        RECT  11.405 6.15 11.47 6.285 ;
        RECT  11.22 5.635 11.285 5.77 ;
        RECT  11.405 5.635 11.47 5.77 ;
        RECT  11.05 3.9575 11.79 4.0225 ;
        RECT  11.05 5.375 11.79 5.44 ;
        RECT  11.05 4.0875 11.79 4.1525 ;
        RECT  11.05 5.505 11.79 5.57 ;
        RECT  11.1575 4.24 11.2225 4.375 ;
        RECT  3.72 19.6975 3.785 19.7625 ;
        RECT  3.72 19.64 3.785 19.705 ;
        RECT  3.5025 19.6975 3.7525 19.7625 ;
        RECT  3.72 19.6725 3.785 19.73 ;
        RECT  3.7525 19.64 4.0 19.705 ;
        RECT  3.72 21.1075 3.785 21.1725 ;
        RECT  3.72 21.165 3.785 21.23 ;
        RECT  3.5025 21.1075 3.7525 21.1725 ;
        RECT  3.72 21.14 3.785 21.1975 ;
        RECT  3.7525 21.165 4.0 21.23 ;
        RECT  3.72 22.3875 3.785 22.4525 ;
        RECT  3.72 22.33 3.785 22.395 ;
        RECT  3.5025 22.3875 3.7525 22.4525 ;
        RECT  3.72 22.3625 3.785 22.42 ;
        RECT  3.7525 22.33 4.0 22.395 ;
        RECT  3.72 23.7975 3.785 23.8625 ;
        RECT  3.72 23.855 3.785 23.92 ;
        RECT  3.5025 23.7975 3.7525 23.8625 ;
        RECT  3.72 23.83 3.785 23.8875 ;
        RECT  3.7525 23.855 4.0 23.92 ;
        RECT  3.72 25.0775 3.785 25.1425 ;
        RECT  3.72 25.02 3.785 25.085 ;
        RECT  3.5025 25.0775 3.7525 25.1425 ;
        RECT  3.72 25.0525 3.785 25.11 ;
        RECT  3.7525 25.02 4.0 25.085 ;
        RECT  3.72 26.4875 3.785 26.5525 ;
        RECT  3.72 26.545 3.785 26.61 ;
        RECT  3.5025 26.4875 3.7525 26.5525 ;
        RECT  3.72 26.52 3.785 26.5775 ;
        RECT  3.7525 26.545 4.0 26.61 ;
        RECT  3.72 27.7675 3.785 27.8325 ;
        RECT  3.72 27.71 3.785 27.775 ;
        RECT  3.5025 27.7675 3.7525 27.8325 ;
        RECT  3.72 27.7425 3.785 27.8 ;
        RECT  3.7525 27.71 4.0 27.775 ;
        RECT  3.72 29.1775 3.785 29.2425 ;
        RECT  3.72 29.235 3.785 29.3 ;
        RECT  3.5025 29.1775 3.7525 29.2425 ;
        RECT  3.72 29.21 3.785 29.2675 ;
        RECT  3.7525 29.235 4.0 29.3 ;
        RECT  3.72 30.4575 3.785 30.5225 ;
        RECT  3.72 30.4 3.785 30.465 ;
        RECT  3.5025 30.4575 3.7525 30.5225 ;
        RECT  3.72 30.4325 3.785 30.49 ;
        RECT  3.7525 30.4 4.0 30.465 ;
        RECT  3.72 31.8675 3.785 31.9325 ;
        RECT  3.72 31.925 3.785 31.99 ;
        RECT  3.5025 31.8675 3.7525 31.9325 ;
        RECT  3.72 31.9 3.785 31.9575 ;
        RECT  3.7525 31.925 4.0 31.99 ;
        RECT  3.72 33.1475 3.785 33.2125 ;
        RECT  3.72 33.09 3.785 33.155 ;
        RECT  3.5025 33.1475 3.7525 33.2125 ;
        RECT  3.72 33.1225 3.785 33.18 ;
        RECT  3.7525 33.09 4.0 33.155 ;
        RECT  3.72 34.5575 3.785 34.6225 ;
        RECT  3.72 34.615 3.785 34.68 ;
        RECT  3.5025 34.5575 3.7525 34.6225 ;
        RECT  3.72 34.59 3.785 34.6475 ;
        RECT  3.7525 34.615 4.0 34.68 ;
        RECT  3.72 35.8375 3.785 35.9025 ;
        RECT  3.72 35.78 3.785 35.845 ;
        RECT  3.5025 35.8375 3.7525 35.9025 ;
        RECT  3.72 35.8125 3.785 35.87 ;
        RECT  3.7525 35.78 4.0 35.845 ;
        RECT  3.72 37.2475 3.785 37.3125 ;
        RECT  3.72 37.305 3.785 37.37 ;
        RECT  3.5025 37.2475 3.7525 37.3125 ;
        RECT  3.72 37.28 3.785 37.3375 ;
        RECT  3.7525 37.305 4.0 37.37 ;
        RECT  3.72 38.5275 3.785 38.5925 ;
        RECT  3.72 38.47 3.785 38.535 ;
        RECT  3.5025 38.5275 3.7525 38.5925 ;
        RECT  3.72 38.5025 3.785 38.56 ;
        RECT  3.7525 38.47 4.0 38.535 ;
        RECT  3.72 39.9375 3.785 40.0025 ;
        RECT  3.72 39.995 3.785 40.06 ;
        RECT  3.5025 39.9375 3.7525 40.0025 ;
        RECT  3.72 39.97 3.785 40.0275 ;
        RECT  3.7525 39.995 4.0 40.06 ;
        RECT  1.59 8.88 2.955 8.945 ;
        RECT  1.765 10.405 2.955 10.47 ;
        RECT  1.94 11.57 2.955 11.635 ;
        RECT  2.115 13.095 2.955 13.16 ;
        RECT  2.29 14.26 2.955 14.325 ;
        RECT  2.465 15.785 2.955 15.85 ;
        RECT  2.64 16.95 2.955 17.015 ;
        RECT  2.815 18.475 2.955 18.54 ;
        RECT  1.59 19.6975 3.015 19.7625 ;
        RECT  2.29 19.4825 3.2725 19.5475 ;
        RECT  1.59 21.1075 3.015 21.1725 ;
        RECT  2.465 21.3225 3.2725 21.3875 ;
        RECT  1.59 22.3875 3.015 22.4525 ;
        RECT  2.64 22.1725 3.2725 22.2375 ;
        RECT  1.59 23.7975 3.015 23.8625 ;
        RECT  2.815 24.0125 3.2725 24.0775 ;
        RECT  1.765 25.0775 3.015 25.1425 ;
        RECT  2.29 24.8625 3.2725 24.9275 ;
        RECT  1.765 26.4875 3.015 26.5525 ;
        RECT  2.465 26.7025 3.2725 26.7675 ;
        RECT  1.765 27.7675 3.015 27.8325 ;
        RECT  2.64 27.5525 3.2725 27.6175 ;
        RECT  1.765 29.1775 3.015 29.2425 ;
        RECT  2.815 29.3925 3.2725 29.4575 ;
        RECT  1.94 30.4575 3.015 30.5225 ;
        RECT  2.29 30.2425 3.2725 30.3075 ;
        RECT  1.94 31.8675 3.015 31.9325 ;
        RECT  2.465 32.0825 3.2725 32.1475 ;
        RECT  1.94 33.1475 3.015 33.2125 ;
        RECT  2.64 32.9325 3.2725 32.9975 ;
        RECT  1.94 34.5575 3.015 34.6225 ;
        RECT  2.815 34.7725 3.2725 34.8375 ;
        RECT  2.115 35.8375 3.015 35.9025 ;
        RECT  2.29 35.6225 3.2725 35.6875 ;
        RECT  2.115 37.2475 3.015 37.3125 ;
        RECT  2.465 37.4625 3.2725 37.5275 ;
        RECT  2.115 38.5275 3.015 38.5925 ;
        RECT  2.64 38.3125 3.2725 38.3775 ;
        RECT  2.115 39.9375 3.015 40.0025 ;
        RECT  2.815 40.1525 3.2725 40.2175 ;
        RECT  4.165 29.235 4.23 29.3 ;
        RECT  4.165 26.545 4.23 26.61 ;
        RECT  4.165 33.09 4.23 33.155 ;
        RECT  4.165 21.165 4.23 21.23 ;
        RECT  4.165 23.855 4.23 23.92 ;
        RECT  4.165 35.78 4.23 35.845 ;
        RECT  4.165 30.4 4.23 30.465 ;
        RECT  4.165 38.47 4.23 38.535 ;
        RECT  4.165 27.71 4.23 27.775 ;
        RECT  4.165 19.64 4.23 19.705 ;
        RECT  4.165 25.02 4.23 25.085 ;
        RECT  4.165 22.33 4.23 22.395 ;
        RECT  4.165 37.305 4.23 37.37 ;
        RECT  4.165 31.925 4.23 31.99 ;
        RECT  4.165 39.995 4.23 40.06 ;
        RECT  4.165 34.615 4.23 34.68 ;
        RECT  1.555 9.6425 6.92 9.7075 ;
        RECT  1.555 12.3325 6.92 12.3975 ;
        RECT  1.555 15.0225 6.92 15.0875 ;
        RECT  1.555 17.7125 6.92 17.7775 ;
        RECT  1.555 20.4025 6.92 20.4675 ;
        RECT  1.555 23.0925 6.92 23.1575 ;
        RECT  1.555 25.7825 6.92 25.8475 ;
        RECT  1.555 28.4725 6.92 28.5375 ;
        RECT  1.555 31.1625 6.92 31.2275 ;
        RECT  1.555 33.8525 6.92 33.9175 ;
        RECT  1.555 36.5425 6.92 36.6075 ;
        RECT  1.555 39.2325 6.92 39.2975 ;
        RECT  1.555 8.2975 6.92 8.3625 ;
        RECT  1.555 10.9875 6.92 11.0525 ;
        RECT  1.555 13.6775 6.92 13.7425 ;
        RECT  1.555 16.3675 6.92 16.4325 ;
        RECT  1.555 19.0575 6.92 19.1225 ;
        RECT  1.555 21.7475 6.92 21.8125 ;
        RECT  1.555 24.4375 6.92 24.5025 ;
        RECT  1.555 27.1275 6.92 27.1925 ;
        RECT  1.555 29.8175 6.92 29.8825 ;
        RECT  1.555 32.5075 6.92 32.5725 ;
        RECT  1.555 35.1975 6.92 35.2625 ;
        RECT  1.555 37.8875 6.92 37.9525 ;
        RECT  1.555 40.5775 6.92 40.6425 ;
        RECT  5.7125 8.88 5.7775 8.945 ;
        RECT  5.7125 9.4475 5.7775 9.5125 ;
        RECT  5.745 8.88 6.015 8.945 ;
        RECT  5.7125 8.9125 5.7775 9.48 ;
        RECT  5.5 9.4475 5.745 9.5125 ;
        RECT  6.245 8.88 6.885 8.945 ;
        RECT  5.7125 10.405 5.7775 10.47 ;
        RECT  5.7125 10.7925 5.7775 10.8575 ;
        RECT  5.745 10.405 6.015 10.47 ;
        RECT  5.7125 10.4375 5.7775 10.825 ;
        RECT  5.225 10.7925 5.745 10.8575 ;
        RECT  6.245 10.405 6.61 10.47 ;
        RECT  4.95 11.1225 6.885 11.1875 ;
        RECT  4.675 12.4675 6.61 12.5325 ;
        RECT  4.375 8.9375 5.5 9.0025 ;
        RECT  4.1175 8.7225 5.225 8.7875 ;
        RECT  4.375 10.3475 4.95 10.4125 ;
        RECT  4.1175 10.5625 5.225 10.6275 ;
        RECT  4.375 11.6275 5.5 11.6925 ;
        RECT  4.1175 11.4125 4.675 11.4775 ;
        RECT  4.375 13.0375 4.95 13.1025 ;
        RECT  4.1175 13.2525 4.675 13.3175 ;
        RECT  3.605 8.9375 3.67 9.0025 ;
        RECT  3.605 8.88 3.67 8.945 ;
        RECT  3.6375 8.9375 3.8875 9.0025 ;
        RECT  3.605 8.9125 3.67 8.97 ;
        RECT  3.39 8.88 3.6375 8.945 ;
        RECT  3.605 10.3475 3.67 10.4125 ;
        RECT  3.605 10.405 3.67 10.47 ;
        RECT  3.6375 10.3475 3.8875 10.4125 ;
        RECT  3.605 10.38 3.67 10.4375 ;
        RECT  3.39 10.405 3.6375 10.47 ;
        RECT  3.605 11.6275 3.67 11.6925 ;
        RECT  3.605 11.57 3.67 11.635 ;
        RECT  3.6375 11.6275 3.8875 11.6925 ;
        RECT  3.605 11.6025 3.67 11.66 ;
        RECT  3.39 11.57 3.6375 11.635 ;
        RECT  3.605 13.0375 3.67 13.1025 ;
        RECT  3.605 13.095 3.67 13.16 ;
        RECT  3.6375 13.0375 3.8875 13.1025 ;
        RECT  3.605 13.07 3.67 13.1275 ;
        RECT  3.39 13.095 3.6375 13.16 ;
        RECT  2.955 13.095 3.16 13.16 ;
        RECT  2.955 11.57 3.16 11.635 ;
        RECT  2.955 8.88 3.16 8.945 ;
        RECT  2.955 10.405 3.16 10.47 ;
        RECT  2.955 9.6425 6.92 9.7075 ;
        RECT  2.955 12.3325 6.92 12.3975 ;
        RECT  2.955 8.2975 6.92 8.3625 ;
        RECT  2.955 10.9875 6.92 11.0525 ;
        RECT  2.955 13.6775 6.92 13.7425 ;
        RECT  5.8775 8.145 5.9425 8.33 ;
        RECT  5.8775 6.985 5.9425 7.215 ;
        RECT  6.2375 8.2125 6.3025 8.3625 ;
        RECT  6.2375 6.9525 6.3025 7.3275 ;
        RECT  6.0475 7.3275 6.1125 8.0775 ;
        RECT  6.18 7.68 6.245 7.815 ;
        RECT  6.015 7.715 6.08 7.78 ;
        RECT  5.81 6.9525 6.37 7.0175 ;
        RECT  5.81 8.2975 6.37 8.3625 ;
        RECT  6.2375 7.1925 6.3025 7.3275 ;
        RECT  6.0475 7.1925 6.1125 7.3275 ;
        RECT  6.2375 7.1925 6.3025 7.3275 ;
        RECT  6.0475 7.1925 6.1125 7.3275 ;
        RECT  6.2375 8.0775 6.3025 8.2125 ;
        RECT  6.0475 8.0775 6.1125 8.2125 ;
        RECT  6.2375 8.0775 6.3025 8.2125 ;
        RECT  6.0475 8.0775 6.1125 8.2125 ;
        RECT  5.8775 8.0775 5.9425 8.2125 ;
        RECT  5.8775 7.1475 5.9425 7.2825 ;
        RECT  6.18 7.68 6.245 7.815 ;
        RECT  5.8775 11.02 5.9425 11.205 ;
        RECT  5.8775 12.135 5.9425 12.365 ;
        RECT  6.2375 10.9875 6.3025 11.1375 ;
        RECT  6.2375 12.0225 6.3025 12.3975 ;
        RECT  6.0475 11.2725 6.1125 12.0225 ;
        RECT  6.18 11.535 6.245 11.67 ;
        RECT  6.015 11.57 6.08 11.635 ;
        RECT  5.81 12.3325 6.37 12.3975 ;
        RECT  5.81 10.9875 6.37 11.0525 ;
        RECT  6.2375 11.7525 6.3025 11.8875 ;
        RECT  6.0475 11.7525 6.1125 11.8875 ;
        RECT  6.2375 11.7525 6.3025 11.8875 ;
        RECT  6.0475 11.7525 6.1125 11.8875 ;
        RECT  6.2375 11.0475 6.3025 11.1825 ;
        RECT  6.0475 11.0475 6.1125 11.1825 ;
        RECT  6.2375 11.0475 6.3025 11.1825 ;
        RECT  6.0475 11.0475 6.1125 11.1825 ;
        RECT  5.8775 11.0025 5.9425 11.1375 ;
        RECT  5.8775 11.9325 5.9425 12.0675 ;
        RECT  6.18 11.4 6.245 11.535 ;
        RECT  3.0225 8.145 3.0875 8.33 ;
        RECT  3.0225 6.985 3.0875 7.215 ;
        RECT  3.3825 8.2125 3.4475 8.3625 ;
        RECT  3.3825 6.9525 3.4475 7.3275 ;
        RECT  3.1925 7.3275 3.2575 8.0775 ;
        RECT  3.325 7.68 3.39 7.815 ;
        RECT  3.16 7.715 3.225 7.78 ;
        RECT  2.955 6.9525 3.515 7.0175 ;
        RECT  2.955 8.2975 3.515 8.3625 ;
        RECT  3.3825 7.1925 3.4475 7.3275 ;
        RECT  3.1925 7.1925 3.2575 7.3275 ;
        RECT  3.3825 7.1925 3.4475 7.3275 ;
        RECT  3.1925 7.1925 3.2575 7.3275 ;
        RECT  3.3825 8.0775 3.4475 8.2125 ;
        RECT  3.1925 8.0775 3.2575 8.2125 ;
        RECT  3.3825 8.0775 3.4475 8.2125 ;
        RECT  3.1925 8.0775 3.2575 8.2125 ;
        RECT  3.0225 8.0775 3.0875 8.2125 ;
        RECT  3.0225 7.1475 3.0875 7.2825 ;
        RECT  3.325 7.68 3.39 7.815 ;
        RECT  3.0225 11.02 3.0875 11.205 ;
        RECT  3.0225 12.135 3.0875 12.365 ;
        RECT  3.3825 10.9875 3.4475 11.1375 ;
        RECT  3.3825 12.0225 3.4475 12.3975 ;
        RECT  3.1925 11.2725 3.2575 12.0225 ;
        RECT  3.325 11.535 3.39 11.67 ;
        RECT  3.16 11.57 3.225 11.635 ;
        RECT  2.955 12.3325 3.515 12.3975 ;
        RECT  2.955 10.9875 3.515 11.0525 ;
        RECT  3.3825 11.7525 3.4475 11.8875 ;
        RECT  3.1925 11.7525 3.2575 11.8875 ;
        RECT  3.3825 11.7525 3.4475 11.8875 ;
        RECT  3.1925 11.7525 3.2575 11.8875 ;
        RECT  3.3825 11.0475 3.4475 11.1825 ;
        RECT  3.1925 11.0475 3.2575 11.1825 ;
        RECT  3.3825 11.0475 3.4475 11.1825 ;
        RECT  3.1925 11.0475 3.2575 11.1825 ;
        RECT  3.0225 11.0025 3.0875 11.1375 ;
        RECT  3.0225 11.9325 3.0875 12.0675 ;
        RECT  3.325 11.4 3.39 11.535 ;
        RECT  3.0225 10.835 3.0875 11.02 ;
        RECT  3.0225 9.675 3.0875 9.905 ;
        RECT  3.3825 10.9025 3.4475 11.0525 ;
        RECT  3.3825 9.6425 3.4475 10.0175 ;
        RECT  3.1925 10.0175 3.2575 10.7675 ;
        RECT  3.325 10.37 3.39 10.505 ;
        RECT  3.16 10.405 3.225 10.47 ;
        RECT  2.955 9.6425 3.515 9.7075 ;
        RECT  2.955 10.9875 3.515 11.0525 ;
        RECT  3.3825 9.8825 3.4475 10.0175 ;
        RECT  3.1925 9.8825 3.2575 10.0175 ;
        RECT  3.3825 9.8825 3.4475 10.0175 ;
        RECT  3.1925 9.8825 3.2575 10.0175 ;
        RECT  3.3825 10.7675 3.4475 10.9025 ;
        RECT  3.1925 10.7675 3.2575 10.9025 ;
        RECT  3.3825 10.7675 3.4475 10.9025 ;
        RECT  3.1925 10.7675 3.2575 10.9025 ;
        RECT  3.0225 10.7675 3.0875 10.9025 ;
        RECT  3.0225 9.8375 3.0875 9.9725 ;
        RECT  3.325 10.37 3.39 10.505 ;
        RECT  3.0225 13.71 3.0875 13.895 ;
        RECT  3.0225 14.825 3.0875 15.055 ;
        RECT  3.3825 13.6775 3.4475 13.8275 ;
        RECT  3.3825 14.7125 3.4475 15.0875 ;
        RECT  3.1925 13.9625 3.2575 14.7125 ;
        RECT  3.325 14.225 3.39 14.36 ;
        RECT  3.16 14.26 3.225 14.325 ;
        RECT  2.955 15.0225 3.515 15.0875 ;
        RECT  2.955 13.6775 3.515 13.7425 ;
        RECT  3.3825 14.4425 3.4475 14.5775 ;
        RECT  3.1925 14.4425 3.2575 14.5775 ;
        RECT  3.3825 14.4425 3.4475 14.5775 ;
        RECT  3.1925 14.4425 3.2575 14.5775 ;
        RECT  3.3825 13.7375 3.4475 13.8725 ;
        RECT  3.1925 13.7375 3.2575 13.8725 ;
        RECT  3.3825 13.7375 3.4475 13.8725 ;
        RECT  3.1925 13.7375 3.2575 13.8725 ;
        RECT  3.0225 13.6925 3.0875 13.8275 ;
        RECT  3.0225 14.6225 3.0875 14.7575 ;
        RECT  3.325 14.09 3.39 14.225 ;
        RECT  3.7525 8.145 3.8175 8.33 ;
        RECT  3.7525 6.985 3.8175 7.215 ;
        RECT  4.3025 8.1675 4.3675 8.3625 ;
        RECT  4.3025 6.9525 4.3675 7.3275 ;
        RECT  3.9225 6.9525 3.9875 7.3275 ;
        RECT  4.24 7.6575 4.375 7.7225 ;
        RECT  3.8875 7.6575 4.0225 7.7225 ;
        RECT  3.9825 7.8725 4.1175 7.9375 ;
        RECT  3.515 6.9525 4.435 7.0175 ;
        RECT  3.515 8.2975 4.435 8.3625 ;
        RECT  4.3025 7.1925 4.3675 7.3275 ;
        RECT  4.1125 7.1925 4.1775 7.3275 ;
        RECT  4.3025 7.1925 4.3675 7.3275 ;
        RECT  4.1125 7.1925 4.1775 7.3275 ;
        RECT  4.1125 7.1925 4.1775 7.3275 ;
        RECT  3.9225 7.1925 3.9875 7.3275 ;
        RECT  4.1125 7.1925 4.1775 7.3275 ;
        RECT  3.9225 7.1925 3.9875 7.3275 ;
        RECT  4.3025 8.0325 4.3675 8.1675 ;
        RECT  4.1125 8.0325 4.1775 8.1675 ;
        RECT  4.3025 8.0325 4.3675 8.1675 ;
        RECT  4.1125 8.0325 4.1775 8.1675 ;
        RECT  4.1125 8.0325 4.1775 8.1675 ;
        RECT  3.9225 8.0325 3.9875 8.1675 ;
        RECT  4.1125 8.0325 4.1775 8.1675 ;
        RECT  3.9225 8.0325 3.9875 8.1675 ;
        RECT  3.7525 8.0775 3.8175 8.2125 ;
        RECT  3.7525 7.1475 3.8175 7.2825 ;
        RECT  3.9825 7.8725 4.1175 7.9375 ;
        RECT  4.24 7.6575 4.375 7.7225 ;
        RECT  4.1125 7.1925 4.1775 7.3275 ;
        RECT  3.9225 8.0325 3.9875 8.1675 ;
        RECT  3.8875 7.6575 4.0225 7.7225 ;
        RECT  3.7525 11.02 3.8175 11.205 ;
        RECT  3.7525 12.135 3.8175 12.365 ;
        RECT  4.3025 10.9875 4.3675 11.1825 ;
        RECT  4.3025 12.0225 4.3675 12.3975 ;
        RECT  3.9225 12.0225 3.9875 12.3975 ;
        RECT  4.24 11.6275 4.375 11.6925 ;
        RECT  3.8875 11.6275 4.0225 11.6925 ;
        RECT  3.9825 11.4125 4.1175 11.4775 ;
        RECT  3.515 12.3325 4.435 12.3975 ;
        RECT  3.515 10.9875 4.435 11.0525 ;
        RECT  4.3025 11.7525 4.3675 11.8875 ;
        RECT  4.1125 11.7525 4.1775 11.8875 ;
        RECT  4.3025 11.7525 4.3675 11.8875 ;
        RECT  4.1125 11.7525 4.1775 11.8875 ;
        RECT  4.1125 11.7525 4.1775 11.8875 ;
        RECT  3.9225 11.7525 3.9875 11.8875 ;
        RECT  4.1125 11.7525 4.1775 11.8875 ;
        RECT  3.9225 11.7525 3.9875 11.8875 ;
        RECT  4.3025 11.0025 4.3675 11.1375 ;
        RECT  4.1125 11.0025 4.1775 11.1375 ;
        RECT  4.3025 11.0025 4.3675 11.1375 ;
        RECT  4.1125 11.0025 4.1775 11.1375 ;
        RECT  4.1125 11.0025 4.1775 11.1375 ;
        RECT  3.9225 11.0025 3.9875 11.1375 ;
        RECT  4.1125 11.0025 4.1775 11.1375 ;
        RECT  3.9225 11.0025 3.9875 11.1375 ;
        RECT  3.7525 11.0025 3.8175 11.1375 ;
        RECT  3.7525 11.9325 3.8175 12.0675 ;
        RECT  3.9825 11.3375 4.1175 11.4025 ;
        RECT  4.24 11.5525 4.375 11.6175 ;
        RECT  4.1125 11.8875 4.1775 12.0225 ;
        RECT  3.9225 11.0475 3.9875 11.1825 ;
        RECT  3.8875 11.5575 4.0225 11.6225 ;
        RECT  3.7525 10.835 3.8175 11.02 ;
        RECT  3.7525 9.675 3.8175 9.905 ;
        RECT  4.3025 10.8575 4.3675 11.0525 ;
        RECT  4.3025 9.6425 4.3675 10.0175 ;
        RECT  3.9225 9.6425 3.9875 10.0175 ;
        RECT  4.24 10.3475 4.375 10.4125 ;
        RECT  3.8875 10.3475 4.0225 10.4125 ;
        RECT  3.9825 10.5625 4.1175 10.6275 ;
        RECT  3.515 9.6425 4.435 9.7075 ;
        RECT  3.515 10.9875 4.435 11.0525 ;
        RECT  4.3025 9.8825 4.3675 10.0175 ;
        RECT  4.1125 9.8825 4.1775 10.0175 ;
        RECT  4.3025 9.8825 4.3675 10.0175 ;
        RECT  4.1125 9.8825 4.1775 10.0175 ;
        RECT  4.1125 9.8825 4.1775 10.0175 ;
        RECT  3.9225 9.8825 3.9875 10.0175 ;
        RECT  4.1125 9.8825 4.1775 10.0175 ;
        RECT  3.9225 9.8825 3.9875 10.0175 ;
        RECT  4.3025 10.7225 4.3675 10.8575 ;
        RECT  4.1125 10.7225 4.1775 10.8575 ;
        RECT  4.3025 10.7225 4.3675 10.8575 ;
        RECT  4.1125 10.7225 4.1775 10.8575 ;
        RECT  4.1125 10.7225 4.1775 10.8575 ;
        RECT  3.9225 10.7225 3.9875 10.8575 ;
        RECT  4.1125 10.7225 4.1775 10.8575 ;
        RECT  3.9225 10.7225 3.9875 10.8575 ;
        RECT  3.7525 10.7675 3.8175 10.9025 ;
        RECT  3.7525 9.8375 3.8175 9.9725 ;
        RECT  3.9825 10.5625 4.1175 10.6275 ;
        RECT  4.24 10.3475 4.375 10.4125 ;
        RECT  4.1125 9.8825 4.1775 10.0175 ;
        RECT  3.9225 10.7225 3.9875 10.8575 ;
        RECT  3.8875 10.3475 4.0225 10.4125 ;
        RECT  3.7525 13.71 3.8175 13.895 ;
        RECT  3.7525 14.825 3.8175 15.055 ;
        RECT  4.3025 13.6775 4.3675 13.8725 ;
        RECT  4.3025 14.7125 4.3675 15.0875 ;
        RECT  3.9225 14.7125 3.9875 15.0875 ;
        RECT  4.24 14.3175 4.375 14.3825 ;
        RECT  3.8875 14.3175 4.0225 14.3825 ;
        RECT  3.9825 14.1025 4.1175 14.1675 ;
        RECT  3.515 15.0225 4.435 15.0875 ;
        RECT  3.515 13.6775 4.435 13.7425 ;
        RECT  4.3025 14.4425 4.3675 14.5775 ;
        RECT  4.1125 14.4425 4.1775 14.5775 ;
        RECT  4.3025 14.4425 4.3675 14.5775 ;
        RECT  4.1125 14.4425 4.1775 14.5775 ;
        RECT  4.1125 14.4425 4.1775 14.5775 ;
        RECT  3.9225 14.4425 3.9875 14.5775 ;
        RECT  4.1125 14.4425 4.1775 14.5775 ;
        RECT  3.9225 14.4425 3.9875 14.5775 ;
        RECT  4.3025 13.6925 4.3675 13.8275 ;
        RECT  4.1125 13.6925 4.1775 13.8275 ;
        RECT  4.3025 13.6925 4.3675 13.8275 ;
        RECT  4.1125 13.6925 4.1775 13.8275 ;
        RECT  4.1125 13.6925 4.1775 13.8275 ;
        RECT  3.9225 13.6925 3.9875 13.8275 ;
        RECT  4.1125 13.6925 4.1775 13.8275 ;
        RECT  3.9225 13.6925 3.9875 13.8275 ;
        RECT  3.7525 13.6925 3.8175 13.8275 ;
        RECT  3.7525 14.6225 3.8175 14.7575 ;
        RECT  3.9825 14.0275 4.1175 14.0925 ;
        RECT  4.24 14.2425 4.375 14.3075 ;
        RECT  4.1125 14.5775 4.1775 14.7125 ;
        RECT  3.9225 13.7375 3.9875 13.8725 ;
        RECT  3.8875 14.2475 4.0225 14.3125 ;
        RECT  5.4325 9.3775 5.5675 9.4425 ;
        RECT  6.8175 8.81 6.9525 8.875 ;
        RECT  5.1575 10.7225 5.2925 10.7875 ;
        RECT  6.5425 10.335 6.6775 10.4 ;
        RECT  6.8175 11.0525 6.9525 11.1175 ;
        RECT  4.8825 11.0525 5.0175 11.1175 ;
        RECT  6.5425 12.3975 6.6775 12.4625 ;
        RECT  4.6075 12.3975 4.7425 12.4625 ;
        RECT  5.4325 8.8675 5.5675 8.9325 ;
        RECT  5.1575 8.6525 5.2925 8.7175 ;
        RECT  4.8825 10.2775 5.0175 10.3425 ;
        RECT  5.1575 10.4925 5.2925 10.5575 ;
        RECT  5.4325 11.5575 5.5675 11.6225 ;
        RECT  4.6075 11.3425 4.7425 11.4075 ;
        RECT  4.8825 12.9675 5.0175 13.0325 ;
        RECT  4.6075 13.1825 4.7425 13.2475 ;
        RECT  5.7125 14.26 5.7775 14.325 ;
        RECT  5.7125 14.8275 5.7775 14.8925 ;
        RECT  5.745 14.26 6.015 14.325 ;
        RECT  5.7125 14.2925 5.7775 14.86 ;
        RECT  5.5 14.8275 5.745 14.8925 ;
        RECT  6.245 14.26 6.885 14.325 ;
        RECT  5.7125 15.785 5.7775 15.85 ;
        RECT  5.7125 16.1725 5.7775 16.2375 ;
        RECT  5.745 15.785 6.015 15.85 ;
        RECT  5.7125 15.8175 5.7775 16.205 ;
        RECT  5.225 16.1725 5.745 16.2375 ;
        RECT  6.245 15.785 6.61 15.85 ;
        RECT  4.95 16.5025 6.885 16.5675 ;
        RECT  4.675 17.8475 6.61 17.9125 ;
        RECT  4.375 14.3175 5.5 14.3825 ;
        RECT  4.1175 14.1025 5.225 14.1675 ;
        RECT  4.375 15.7275 4.95 15.7925 ;
        RECT  4.1175 15.9425 5.225 16.0075 ;
        RECT  4.375 17.0075 5.5 17.0725 ;
        RECT  4.1175 16.7925 4.675 16.8575 ;
        RECT  4.375 18.4175 4.95 18.4825 ;
        RECT  4.1175 18.6325 4.675 18.6975 ;
        RECT  3.605 14.3175 3.67 14.3825 ;
        RECT  3.605 14.26 3.67 14.325 ;
        RECT  3.6375 14.3175 3.8875 14.3825 ;
        RECT  3.605 14.2925 3.67 14.35 ;
        RECT  3.39 14.26 3.6375 14.325 ;
        RECT  3.605 15.7275 3.67 15.7925 ;
        RECT  3.605 15.785 3.67 15.85 ;
        RECT  3.6375 15.7275 3.8875 15.7925 ;
        RECT  3.605 15.76 3.67 15.8175 ;
        RECT  3.39 15.785 3.6375 15.85 ;
        RECT  3.605 17.0075 3.67 17.0725 ;
        RECT  3.605 16.95 3.67 17.015 ;
        RECT  3.6375 17.0075 3.8875 17.0725 ;
        RECT  3.605 16.9825 3.67 17.04 ;
        RECT  3.39 16.95 3.6375 17.015 ;
        RECT  3.605 18.4175 3.67 18.4825 ;
        RECT  3.605 18.475 3.67 18.54 ;
        RECT  3.6375 18.4175 3.8875 18.4825 ;
        RECT  3.605 18.45 3.67 18.5075 ;
        RECT  3.39 18.475 3.6375 18.54 ;
        RECT  2.955 18.475 3.16 18.54 ;
        RECT  2.955 16.95 3.16 17.015 ;
        RECT  2.955 14.26 3.16 14.325 ;
        RECT  2.955 15.785 3.16 15.85 ;
        RECT  2.955 15.0225 6.92 15.0875 ;
        RECT  2.955 17.7125 6.92 17.7775 ;
        RECT  2.955 13.6775 6.92 13.7425 ;
        RECT  2.955 16.3675 6.92 16.4325 ;
        RECT  2.955 19.0575 6.92 19.1225 ;
        RECT  5.8775 13.525 5.9425 13.71 ;
        RECT  5.8775 12.365 5.9425 12.595 ;
        RECT  6.2375 13.5925 6.3025 13.7425 ;
        RECT  6.2375 12.3325 6.3025 12.7075 ;
        RECT  6.0475 12.7075 6.1125 13.4575 ;
        RECT  6.18 13.06 6.245 13.195 ;
        RECT  6.015 13.095 6.08 13.16 ;
        RECT  5.81 12.3325 6.37 12.3975 ;
        RECT  5.81 13.6775 6.37 13.7425 ;
        RECT  6.2375 12.5725 6.3025 12.7075 ;
        RECT  6.0475 12.5725 6.1125 12.7075 ;
        RECT  6.2375 12.5725 6.3025 12.7075 ;
        RECT  6.0475 12.5725 6.1125 12.7075 ;
        RECT  6.2375 13.4575 6.3025 13.5925 ;
        RECT  6.0475 13.4575 6.1125 13.5925 ;
        RECT  6.2375 13.4575 6.3025 13.5925 ;
        RECT  6.0475 13.4575 6.1125 13.5925 ;
        RECT  5.8775 13.4575 5.9425 13.5925 ;
        RECT  5.8775 12.5275 5.9425 12.6625 ;
        RECT  6.18 13.06 6.245 13.195 ;
        RECT  5.8775 16.4 5.9425 16.585 ;
        RECT  5.8775 17.515 5.9425 17.745 ;
        RECT  6.2375 16.3675 6.3025 16.5175 ;
        RECT  6.2375 17.4025 6.3025 17.7775 ;
        RECT  6.0475 16.6525 6.1125 17.4025 ;
        RECT  6.18 16.915 6.245 17.05 ;
        RECT  6.015 16.95 6.08 17.015 ;
        RECT  5.81 17.7125 6.37 17.7775 ;
        RECT  5.81 16.3675 6.37 16.4325 ;
        RECT  6.2375 17.1325 6.3025 17.2675 ;
        RECT  6.0475 17.1325 6.1125 17.2675 ;
        RECT  6.2375 17.1325 6.3025 17.2675 ;
        RECT  6.0475 17.1325 6.1125 17.2675 ;
        RECT  6.2375 16.4275 6.3025 16.5625 ;
        RECT  6.0475 16.4275 6.1125 16.5625 ;
        RECT  6.2375 16.4275 6.3025 16.5625 ;
        RECT  6.0475 16.4275 6.1125 16.5625 ;
        RECT  5.8775 16.3825 5.9425 16.5175 ;
        RECT  5.8775 17.3125 5.9425 17.4475 ;
        RECT  6.18 16.78 6.245 16.915 ;
        RECT  3.0225 13.525 3.0875 13.71 ;
        RECT  3.0225 12.365 3.0875 12.595 ;
        RECT  3.3825 13.5925 3.4475 13.7425 ;
        RECT  3.3825 12.3325 3.4475 12.7075 ;
        RECT  3.1925 12.7075 3.2575 13.4575 ;
        RECT  3.325 13.06 3.39 13.195 ;
        RECT  3.16 13.095 3.225 13.16 ;
        RECT  2.955 12.3325 3.515 12.3975 ;
        RECT  2.955 13.6775 3.515 13.7425 ;
        RECT  3.3825 12.5725 3.4475 12.7075 ;
        RECT  3.1925 12.5725 3.2575 12.7075 ;
        RECT  3.3825 12.5725 3.4475 12.7075 ;
        RECT  3.1925 12.5725 3.2575 12.7075 ;
        RECT  3.3825 13.4575 3.4475 13.5925 ;
        RECT  3.1925 13.4575 3.2575 13.5925 ;
        RECT  3.3825 13.4575 3.4475 13.5925 ;
        RECT  3.1925 13.4575 3.2575 13.5925 ;
        RECT  3.0225 13.4575 3.0875 13.5925 ;
        RECT  3.0225 12.5275 3.0875 12.6625 ;
        RECT  3.325 13.06 3.39 13.195 ;
        RECT  3.0225 16.4 3.0875 16.585 ;
        RECT  3.0225 17.515 3.0875 17.745 ;
        RECT  3.3825 16.3675 3.4475 16.5175 ;
        RECT  3.3825 17.4025 3.4475 17.7775 ;
        RECT  3.1925 16.6525 3.2575 17.4025 ;
        RECT  3.325 16.915 3.39 17.05 ;
        RECT  3.16 16.95 3.225 17.015 ;
        RECT  2.955 17.7125 3.515 17.7775 ;
        RECT  2.955 16.3675 3.515 16.4325 ;
        RECT  3.3825 17.1325 3.4475 17.2675 ;
        RECT  3.1925 17.1325 3.2575 17.2675 ;
        RECT  3.3825 17.1325 3.4475 17.2675 ;
        RECT  3.1925 17.1325 3.2575 17.2675 ;
        RECT  3.3825 16.4275 3.4475 16.5625 ;
        RECT  3.1925 16.4275 3.2575 16.5625 ;
        RECT  3.3825 16.4275 3.4475 16.5625 ;
        RECT  3.1925 16.4275 3.2575 16.5625 ;
        RECT  3.0225 16.3825 3.0875 16.5175 ;
        RECT  3.0225 17.3125 3.0875 17.4475 ;
        RECT  3.325 16.78 3.39 16.915 ;
        RECT  3.0225 16.215 3.0875 16.4 ;
        RECT  3.0225 15.055 3.0875 15.285 ;
        RECT  3.3825 16.2825 3.4475 16.4325 ;
        RECT  3.3825 15.0225 3.4475 15.3975 ;
        RECT  3.1925 15.3975 3.2575 16.1475 ;
        RECT  3.325 15.75 3.39 15.885 ;
        RECT  3.16 15.785 3.225 15.85 ;
        RECT  2.955 15.0225 3.515 15.0875 ;
        RECT  2.955 16.3675 3.515 16.4325 ;
        RECT  3.3825 15.2625 3.4475 15.3975 ;
        RECT  3.1925 15.2625 3.2575 15.3975 ;
        RECT  3.3825 15.2625 3.4475 15.3975 ;
        RECT  3.1925 15.2625 3.2575 15.3975 ;
        RECT  3.3825 16.1475 3.4475 16.2825 ;
        RECT  3.1925 16.1475 3.2575 16.2825 ;
        RECT  3.3825 16.1475 3.4475 16.2825 ;
        RECT  3.1925 16.1475 3.2575 16.2825 ;
        RECT  3.0225 16.1475 3.0875 16.2825 ;
        RECT  3.0225 15.2175 3.0875 15.3525 ;
        RECT  3.325 15.75 3.39 15.885 ;
        RECT  3.0225 19.09 3.0875 19.275 ;
        RECT  3.0225 20.205 3.0875 20.435 ;
        RECT  3.3825 19.0575 3.4475 19.2075 ;
        RECT  3.3825 20.0925 3.4475 20.4675 ;
        RECT  3.1925 19.3425 3.2575 20.0925 ;
        RECT  3.325 19.605 3.39 19.74 ;
        RECT  3.16 19.64 3.225 19.705 ;
        RECT  2.955 20.4025 3.515 20.4675 ;
        RECT  2.955 19.0575 3.515 19.1225 ;
        RECT  3.3825 19.8225 3.4475 19.9575 ;
        RECT  3.1925 19.8225 3.2575 19.9575 ;
        RECT  3.3825 19.8225 3.4475 19.9575 ;
        RECT  3.1925 19.8225 3.2575 19.9575 ;
        RECT  3.3825 19.1175 3.4475 19.2525 ;
        RECT  3.1925 19.1175 3.2575 19.2525 ;
        RECT  3.3825 19.1175 3.4475 19.2525 ;
        RECT  3.1925 19.1175 3.2575 19.2525 ;
        RECT  3.0225 19.0725 3.0875 19.2075 ;
        RECT  3.0225 20.0025 3.0875 20.1375 ;
        RECT  3.325 19.47 3.39 19.605 ;
        RECT  3.7525 13.525 3.8175 13.71 ;
        RECT  3.7525 12.365 3.8175 12.595 ;
        RECT  4.3025 13.5475 4.3675 13.7425 ;
        RECT  4.3025 12.3325 4.3675 12.7075 ;
        RECT  3.9225 12.3325 3.9875 12.7075 ;
        RECT  4.24 13.0375 4.375 13.1025 ;
        RECT  3.8875 13.0375 4.0225 13.1025 ;
        RECT  3.9825 13.2525 4.1175 13.3175 ;
        RECT  3.515 12.3325 4.435 12.3975 ;
        RECT  3.515 13.6775 4.435 13.7425 ;
        RECT  4.3025 12.5725 4.3675 12.7075 ;
        RECT  4.1125 12.5725 4.1775 12.7075 ;
        RECT  4.3025 12.5725 4.3675 12.7075 ;
        RECT  4.1125 12.5725 4.1775 12.7075 ;
        RECT  4.1125 12.5725 4.1775 12.7075 ;
        RECT  3.9225 12.5725 3.9875 12.7075 ;
        RECT  4.1125 12.5725 4.1775 12.7075 ;
        RECT  3.9225 12.5725 3.9875 12.7075 ;
        RECT  4.3025 13.4125 4.3675 13.5475 ;
        RECT  4.1125 13.4125 4.1775 13.5475 ;
        RECT  4.3025 13.4125 4.3675 13.5475 ;
        RECT  4.1125 13.4125 4.1775 13.5475 ;
        RECT  4.1125 13.4125 4.1775 13.5475 ;
        RECT  3.9225 13.4125 3.9875 13.5475 ;
        RECT  4.1125 13.4125 4.1775 13.5475 ;
        RECT  3.9225 13.4125 3.9875 13.5475 ;
        RECT  3.7525 13.4575 3.8175 13.5925 ;
        RECT  3.7525 12.5275 3.8175 12.6625 ;
        RECT  3.9825 13.2525 4.1175 13.3175 ;
        RECT  4.24 13.0375 4.375 13.1025 ;
        RECT  4.1125 12.5725 4.1775 12.7075 ;
        RECT  3.9225 13.4125 3.9875 13.5475 ;
        RECT  3.8875 13.0375 4.0225 13.1025 ;
        RECT  3.7525 16.4 3.8175 16.585 ;
        RECT  3.7525 17.515 3.8175 17.745 ;
        RECT  4.3025 16.3675 4.3675 16.5625 ;
        RECT  4.3025 17.4025 4.3675 17.7775 ;
        RECT  3.9225 17.4025 3.9875 17.7775 ;
        RECT  4.24 17.0075 4.375 17.0725 ;
        RECT  3.8875 17.0075 4.0225 17.0725 ;
        RECT  3.9825 16.7925 4.1175 16.8575 ;
        RECT  3.515 17.7125 4.435 17.7775 ;
        RECT  3.515 16.3675 4.435 16.4325 ;
        RECT  4.3025 17.1325 4.3675 17.2675 ;
        RECT  4.1125 17.1325 4.1775 17.2675 ;
        RECT  4.3025 17.1325 4.3675 17.2675 ;
        RECT  4.1125 17.1325 4.1775 17.2675 ;
        RECT  4.1125 17.1325 4.1775 17.2675 ;
        RECT  3.9225 17.1325 3.9875 17.2675 ;
        RECT  4.1125 17.1325 4.1775 17.2675 ;
        RECT  3.9225 17.1325 3.9875 17.2675 ;
        RECT  4.3025 16.3825 4.3675 16.5175 ;
        RECT  4.1125 16.3825 4.1775 16.5175 ;
        RECT  4.3025 16.3825 4.3675 16.5175 ;
        RECT  4.1125 16.3825 4.1775 16.5175 ;
        RECT  4.1125 16.3825 4.1775 16.5175 ;
        RECT  3.9225 16.3825 3.9875 16.5175 ;
        RECT  4.1125 16.3825 4.1775 16.5175 ;
        RECT  3.9225 16.3825 3.9875 16.5175 ;
        RECT  3.7525 16.3825 3.8175 16.5175 ;
        RECT  3.7525 17.3125 3.8175 17.4475 ;
        RECT  3.9825 16.7175 4.1175 16.7825 ;
        RECT  4.24 16.9325 4.375 16.9975 ;
        RECT  4.1125 17.2675 4.1775 17.4025 ;
        RECT  3.9225 16.4275 3.9875 16.5625 ;
        RECT  3.8875 16.9375 4.0225 17.0025 ;
        RECT  3.7525 16.215 3.8175 16.4 ;
        RECT  3.7525 15.055 3.8175 15.285 ;
        RECT  4.3025 16.2375 4.3675 16.4325 ;
        RECT  4.3025 15.0225 4.3675 15.3975 ;
        RECT  3.9225 15.0225 3.9875 15.3975 ;
        RECT  4.24 15.7275 4.375 15.7925 ;
        RECT  3.8875 15.7275 4.0225 15.7925 ;
        RECT  3.9825 15.9425 4.1175 16.0075 ;
        RECT  3.515 15.0225 4.435 15.0875 ;
        RECT  3.515 16.3675 4.435 16.4325 ;
        RECT  4.3025 15.2625 4.3675 15.3975 ;
        RECT  4.1125 15.2625 4.1775 15.3975 ;
        RECT  4.3025 15.2625 4.3675 15.3975 ;
        RECT  4.1125 15.2625 4.1775 15.3975 ;
        RECT  4.1125 15.2625 4.1775 15.3975 ;
        RECT  3.9225 15.2625 3.9875 15.3975 ;
        RECT  4.1125 15.2625 4.1775 15.3975 ;
        RECT  3.9225 15.2625 3.9875 15.3975 ;
        RECT  4.3025 16.1025 4.3675 16.2375 ;
        RECT  4.1125 16.1025 4.1775 16.2375 ;
        RECT  4.3025 16.1025 4.3675 16.2375 ;
        RECT  4.1125 16.1025 4.1775 16.2375 ;
        RECT  4.1125 16.1025 4.1775 16.2375 ;
        RECT  3.9225 16.1025 3.9875 16.2375 ;
        RECT  4.1125 16.1025 4.1775 16.2375 ;
        RECT  3.9225 16.1025 3.9875 16.2375 ;
        RECT  3.7525 16.1475 3.8175 16.2825 ;
        RECT  3.7525 15.2175 3.8175 15.3525 ;
        RECT  3.9825 15.9425 4.1175 16.0075 ;
        RECT  4.24 15.7275 4.375 15.7925 ;
        RECT  4.1125 15.2625 4.1775 15.3975 ;
        RECT  3.9225 16.1025 3.9875 16.2375 ;
        RECT  3.8875 15.7275 4.0225 15.7925 ;
        RECT  3.7525 19.09 3.8175 19.275 ;
        RECT  3.7525 20.205 3.8175 20.435 ;
        RECT  4.3025 19.0575 4.3675 19.2525 ;
        RECT  4.3025 20.0925 4.3675 20.4675 ;
        RECT  3.9225 20.0925 3.9875 20.4675 ;
        RECT  4.24 19.6975 4.375 19.7625 ;
        RECT  3.8875 19.6975 4.0225 19.7625 ;
        RECT  3.9825 19.4825 4.1175 19.5475 ;
        RECT  3.515 20.4025 4.435 20.4675 ;
        RECT  3.515 19.0575 4.435 19.1225 ;
        RECT  4.3025 19.8225 4.3675 19.9575 ;
        RECT  4.1125 19.8225 4.1775 19.9575 ;
        RECT  4.3025 19.8225 4.3675 19.9575 ;
        RECT  4.1125 19.8225 4.1775 19.9575 ;
        RECT  4.1125 19.8225 4.1775 19.9575 ;
        RECT  3.9225 19.8225 3.9875 19.9575 ;
        RECT  4.1125 19.8225 4.1775 19.9575 ;
        RECT  3.9225 19.8225 3.9875 19.9575 ;
        RECT  4.3025 19.0725 4.3675 19.2075 ;
        RECT  4.1125 19.0725 4.1775 19.2075 ;
        RECT  4.3025 19.0725 4.3675 19.2075 ;
        RECT  4.1125 19.0725 4.1775 19.2075 ;
        RECT  4.1125 19.0725 4.1775 19.2075 ;
        RECT  3.9225 19.0725 3.9875 19.2075 ;
        RECT  4.1125 19.0725 4.1775 19.2075 ;
        RECT  3.9225 19.0725 3.9875 19.2075 ;
        RECT  3.7525 19.0725 3.8175 19.2075 ;
        RECT  3.7525 20.0025 3.8175 20.1375 ;
        RECT  3.9825 19.4075 4.1175 19.4725 ;
        RECT  4.24 19.6225 4.375 19.6875 ;
        RECT  4.1125 19.9575 4.1775 20.0925 ;
        RECT  3.9225 19.1175 3.9875 19.2525 ;
        RECT  3.8875 19.6275 4.0225 19.6925 ;
        RECT  5.4325 14.7575 5.5675 14.8225 ;
        RECT  6.8175 14.19 6.9525 14.255 ;
        RECT  5.1575 16.1025 5.2925 16.1675 ;
        RECT  6.5425 15.715 6.6775 15.78 ;
        RECT  6.8175 16.4325 6.9525 16.4975 ;
        RECT  4.8825 16.4325 5.0175 16.4975 ;
        RECT  6.5425 17.7775 6.6775 17.8425 ;
        RECT  4.6075 17.7775 4.7425 17.8425 ;
        RECT  5.4325 14.2475 5.5675 14.3125 ;
        RECT  5.1575 14.0325 5.2925 14.0975 ;
        RECT  4.8825 15.6575 5.0175 15.7225 ;
        RECT  5.1575 15.8725 5.2925 15.9375 ;
        RECT  5.4325 16.9375 5.5675 17.0025 ;
        RECT  4.6075 16.7225 4.7425 16.7875 ;
        RECT  4.8825 18.3475 5.0175 18.4125 ;
        RECT  4.6075 18.5625 4.7425 18.6275 ;
        RECT  3.5725 19.09 3.6375 19.275 ;
        RECT  3.5725 20.205 3.6375 20.435 ;
        RECT  3.0225 19.0575 3.0875 19.2525 ;
        RECT  3.0225 20.0925 3.0875 20.4675 ;
        RECT  3.4025 20.0925 3.4675 20.4675 ;
        RECT  3.015 19.6975 3.15 19.7625 ;
        RECT  3.3675 19.6975 3.5025 19.7625 ;
        RECT  3.2725 19.4825 3.4075 19.5475 ;
        RECT  2.955 20.4025 3.875 20.4675 ;
        RECT  2.955 19.0575 3.875 19.1225 ;
        RECT  3.0225 20.0925 3.0875 20.2275 ;
        RECT  3.2125 20.0925 3.2775 20.2275 ;
        RECT  3.0225 20.0925 3.0875 20.2275 ;
        RECT  3.2125 20.0925 3.2775 20.2275 ;
        RECT  3.2125 20.0925 3.2775 20.2275 ;
        RECT  3.4025 20.0925 3.4675 20.2275 ;
        RECT  3.2125 20.0925 3.2775 20.2275 ;
        RECT  3.4025 20.0925 3.4675 20.2275 ;
        RECT  3.0225 19.2525 3.0875 19.3875 ;
        RECT  3.2125 19.2525 3.2775 19.3875 ;
        RECT  3.0225 19.2525 3.0875 19.3875 ;
        RECT  3.2125 19.2525 3.2775 19.3875 ;
        RECT  3.2125 19.2525 3.2775 19.3875 ;
        RECT  3.4025 19.2525 3.4675 19.3875 ;
        RECT  3.2125 19.2525 3.2775 19.3875 ;
        RECT  3.4025 19.2525 3.4675 19.3875 ;
        RECT  3.5725 19.2075 3.6375 19.3425 ;
        RECT  3.5725 20.1375 3.6375 20.2725 ;
        RECT  3.2725 19.4825 3.4075 19.5475 ;
        RECT  3.015 19.6975 3.15 19.7625 ;
        RECT  3.2125 20.0925 3.2775 20.2275 ;
        RECT  3.4025 19.2525 3.4675 19.3875 ;
        RECT  3.3675 19.6975 3.5025 19.7625 ;
        RECT  3.5725 21.595 3.6375 21.78 ;
        RECT  3.5725 20.435 3.6375 20.665 ;
        RECT  3.0225 21.6175 3.0875 21.8125 ;
        RECT  3.0225 20.4025 3.0875 20.7775 ;
        RECT  3.4025 20.4025 3.4675 20.7775 ;
        RECT  3.015 21.1075 3.15 21.1725 ;
        RECT  3.3675 21.1075 3.5025 21.1725 ;
        RECT  3.2725 21.3225 3.4075 21.3875 ;
        RECT  2.955 20.4025 3.875 20.4675 ;
        RECT  2.955 21.7475 3.875 21.8125 ;
        RECT  3.0225 20.9125 3.0875 21.0475 ;
        RECT  3.2125 20.9125 3.2775 21.0475 ;
        RECT  3.0225 20.9125 3.0875 21.0475 ;
        RECT  3.2125 20.9125 3.2775 21.0475 ;
        RECT  3.2125 20.9125 3.2775 21.0475 ;
        RECT  3.4025 20.9125 3.4675 21.0475 ;
        RECT  3.2125 20.9125 3.2775 21.0475 ;
        RECT  3.4025 20.9125 3.4675 21.0475 ;
        RECT  3.0225 21.6625 3.0875 21.7975 ;
        RECT  3.2125 21.6625 3.2775 21.7975 ;
        RECT  3.0225 21.6625 3.0875 21.7975 ;
        RECT  3.2125 21.6625 3.2775 21.7975 ;
        RECT  3.2125 21.6625 3.2775 21.7975 ;
        RECT  3.4025 21.6625 3.4675 21.7975 ;
        RECT  3.2125 21.6625 3.2775 21.7975 ;
        RECT  3.4025 21.6625 3.4675 21.7975 ;
        RECT  3.5725 21.6625 3.6375 21.7975 ;
        RECT  3.5725 20.7325 3.6375 20.8675 ;
        RECT  3.2725 21.3975 3.4075 21.4625 ;
        RECT  3.015 21.1825 3.15 21.2475 ;
        RECT  3.2125 20.7775 3.2775 20.9125 ;
        RECT  3.4025 21.6175 3.4675 21.7525 ;
        RECT  3.3675 21.1775 3.5025 21.2425 ;
        RECT  3.5725 21.78 3.6375 21.965 ;
        RECT  3.5725 22.895 3.6375 23.125 ;
        RECT  3.0225 21.7475 3.0875 21.9425 ;
        RECT  3.0225 22.7825 3.0875 23.1575 ;
        RECT  3.4025 22.7825 3.4675 23.1575 ;
        RECT  3.015 22.3875 3.15 22.4525 ;
        RECT  3.3675 22.3875 3.5025 22.4525 ;
        RECT  3.2725 22.1725 3.4075 22.2375 ;
        RECT  2.955 23.0925 3.875 23.1575 ;
        RECT  2.955 21.7475 3.875 21.8125 ;
        RECT  3.0225 22.7825 3.0875 22.9175 ;
        RECT  3.2125 22.7825 3.2775 22.9175 ;
        RECT  3.0225 22.7825 3.0875 22.9175 ;
        RECT  3.2125 22.7825 3.2775 22.9175 ;
        RECT  3.2125 22.7825 3.2775 22.9175 ;
        RECT  3.4025 22.7825 3.4675 22.9175 ;
        RECT  3.2125 22.7825 3.2775 22.9175 ;
        RECT  3.4025 22.7825 3.4675 22.9175 ;
        RECT  3.0225 21.9425 3.0875 22.0775 ;
        RECT  3.2125 21.9425 3.2775 22.0775 ;
        RECT  3.0225 21.9425 3.0875 22.0775 ;
        RECT  3.2125 21.9425 3.2775 22.0775 ;
        RECT  3.2125 21.9425 3.2775 22.0775 ;
        RECT  3.4025 21.9425 3.4675 22.0775 ;
        RECT  3.2125 21.9425 3.2775 22.0775 ;
        RECT  3.4025 21.9425 3.4675 22.0775 ;
        RECT  3.5725 21.8975 3.6375 22.0325 ;
        RECT  3.5725 22.8275 3.6375 22.9625 ;
        RECT  3.2725 22.1725 3.4075 22.2375 ;
        RECT  3.015 22.3875 3.15 22.4525 ;
        RECT  3.2125 22.7825 3.2775 22.9175 ;
        RECT  3.4025 21.9425 3.4675 22.0775 ;
        RECT  3.3675 22.3875 3.5025 22.4525 ;
        RECT  3.5725 24.285 3.6375 24.47 ;
        RECT  3.5725 23.125 3.6375 23.355 ;
        RECT  3.0225 24.3075 3.0875 24.5025 ;
        RECT  3.0225 23.0925 3.0875 23.4675 ;
        RECT  3.4025 23.0925 3.4675 23.4675 ;
        RECT  3.015 23.7975 3.15 23.8625 ;
        RECT  3.3675 23.7975 3.5025 23.8625 ;
        RECT  3.2725 24.0125 3.4075 24.0775 ;
        RECT  2.955 23.0925 3.875 23.1575 ;
        RECT  2.955 24.4375 3.875 24.5025 ;
        RECT  3.0225 23.6025 3.0875 23.7375 ;
        RECT  3.2125 23.6025 3.2775 23.7375 ;
        RECT  3.0225 23.6025 3.0875 23.7375 ;
        RECT  3.2125 23.6025 3.2775 23.7375 ;
        RECT  3.2125 23.6025 3.2775 23.7375 ;
        RECT  3.4025 23.6025 3.4675 23.7375 ;
        RECT  3.2125 23.6025 3.2775 23.7375 ;
        RECT  3.4025 23.6025 3.4675 23.7375 ;
        RECT  3.0225 24.3525 3.0875 24.4875 ;
        RECT  3.2125 24.3525 3.2775 24.4875 ;
        RECT  3.0225 24.3525 3.0875 24.4875 ;
        RECT  3.2125 24.3525 3.2775 24.4875 ;
        RECT  3.2125 24.3525 3.2775 24.4875 ;
        RECT  3.4025 24.3525 3.4675 24.4875 ;
        RECT  3.2125 24.3525 3.2775 24.4875 ;
        RECT  3.4025 24.3525 3.4675 24.4875 ;
        RECT  3.5725 24.3525 3.6375 24.4875 ;
        RECT  3.5725 23.4225 3.6375 23.5575 ;
        RECT  3.2725 24.0875 3.4075 24.1525 ;
        RECT  3.015 23.8725 3.15 23.9375 ;
        RECT  3.2125 23.4675 3.2775 23.6025 ;
        RECT  3.4025 24.3075 3.4675 24.4425 ;
        RECT  3.3675 23.8675 3.5025 23.9325 ;
        RECT  3.5725 24.47 3.6375 24.655 ;
        RECT  3.5725 25.585 3.6375 25.815 ;
        RECT  3.0225 24.4375 3.0875 24.6325 ;
        RECT  3.0225 25.4725 3.0875 25.8475 ;
        RECT  3.4025 25.4725 3.4675 25.8475 ;
        RECT  3.015 25.0775 3.15 25.1425 ;
        RECT  3.3675 25.0775 3.5025 25.1425 ;
        RECT  3.2725 24.8625 3.4075 24.9275 ;
        RECT  2.955 25.7825 3.875 25.8475 ;
        RECT  2.955 24.4375 3.875 24.5025 ;
        RECT  3.0225 25.4725 3.0875 25.6075 ;
        RECT  3.2125 25.4725 3.2775 25.6075 ;
        RECT  3.0225 25.4725 3.0875 25.6075 ;
        RECT  3.2125 25.4725 3.2775 25.6075 ;
        RECT  3.2125 25.4725 3.2775 25.6075 ;
        RECT  3.4025 25.4725 3.4675 25.6075 ;
        RECT  3.2125 25.4725 3.2775 25.6075 ;
        RECT  3.4025 25.4725 3.4675 25.6075 ;
        RECT  3.0225 24.6325 3.0875 24.7675 ;
        RECT  3.2125 24.6325 3.2775 24.7675 ;
        RECT  3.0225 24.6325 3.0875 24.7675 ;
        RECT  3.2125 24.6325 3.2775 24.7675 ;
        RECT  3.2125 24.6325 3.2775 24.7675 ;
        RECT  3.4025 24.6325 3.4675 24.7675 ;
        RECT  3.2125 24.6325 3.2775 24.7675 ;
        RECT  3.4025 24.6325 3.4675 24.7675 ;
        RECT  3.5725 24.5875 3.6375 24.7225 ;
        RECT  3.5725 25.5175 3.6375 25.6525 ;
        RECT  3.2725 24.8625 3.4075 24.9275 ;
        RECT  3.015 25.0775 3.15 25.1425 ;
        RECT  3.2125 25.4725 3.2775 25.6075 ;
        RECT  3.4025 24.6325 3.4675 24.7675 ;
        RECT  3.3675 25.0775 3.5025 25.1425 ;
        RECT  3.5725 26.975 3.6375 27.16 ;
        RECT  3.5725 25.815 3.6375 26.045 ;
        RECT  3.0225 26.9975 3.0875 27.1925 ;
        RECT  3.0225 25.7825 3.0875 26.1575 ;
        RECT  3.4025 25.7825 3.4675 26.1575 ;
        RECT  3.015 26.4875 3.15 26.5525 ;
        RECT  3.3675 26.4875 3.5025 26.5525 ;
        RECT  3.2725 26.7025 3.4075 26.7675 ;
        RECT  2.955 25.7825 3.875 25.8475 ;
        RECT  2.955 27.1275 3.875 27.1925 ;
        RECT  3.0225 26.2925 3.0875 26.4275 ;
        RECT  3.2125 26.2925 3.2775 26.4275 ;
        RECT  3.0225 26.2925 3.0875 26.4275 ;
        RECT  3.2125 26.2925 3.2775 26.4275 ;
        RECT  3.2125 26.2925 3.2775 26.4275 ;
        RECT  3.4025 26.2925 3.4675 26.4275 ;
        RECT  3.2125 26.2925 3.2775 26.4275 ;
        RECT  3.4025 26.2925 3.4675 26.4275 ;
        RECT  3.0225 27.0425 3.0875 27.1775 ;
        RECT  3.2125 27.0425 3.2775 27.1775 ;
        RECT  3.0225 27.0425 3.0875 27.1775 ;
        RECT  3.2125 27.0425 3.2775 27.1775 ;
        RECT  3.2125 27.0425 3.2775 27.1775 ;
        RECT  3.4025 27.0425 3.4675 27.1775 ;
        RECT  3.2125 27.0425 3.2775 27.1775 ;
        RECT  3.4025 27.0425 3.4675 27.1775 ;
        RECT  3.5725 27.0425 3.6375 27.1775 ;
        RECT  3.5725 26.1125 3.6375 26.2475 ;
        RECT  3.2725 26.7775 3.4075 26.8425 ;
        RECT  3.015 26.5625 3.15 26.6275 ;
        RECT  3.2125 26.1575 3.2775 26.2925 ;
        RECT  3.4025 26.9975 3.4675 27.1325 ;
        RECT  3.3675 26.5575 3.5025 26.6225 ;
        RECT  3.5725 27.16 3.6375 27.345 ;
        RECT  3.5725 28.275 3.6375 28.505 ;
        RECT  3.0225 27.1275 3.0875 27.3225 ;
        RECT  3.0225 28.1625 3.0875 28.5375 ;
        RECT  3.4025 28.1625 3.4675 28.5375 ;
        RECT  3.015 27.7675 3.15 27.8325 ;
        RECT  3.3675 27.7675 3.5025 27.8325 ;
        RECT  3.2725 27.5525 3.4075 27.6175 ;
        RECT  2.955 28.4725 3.875 28.5375 ;
        RECT  2.955 27.1275 3.875 27.1925 ;
        RECT  3.0225 28.1625 3.0875 28.2975 ;
        RECT  3.2125 28.1625 3.2775 28.2975 ;
        RECT  3.0225 28.1625 3.0875 28.2975 ;
        RECT  3.2125 28.1625 3.2775 28.2975 ;
        RECT  3.2125 28.1625 3.2775 28.2975 ;
        RECT  3.4025 28.1625 3.4675 28.2975 ;
        RECT  3.2125 28.1625 3.2775 28.2975 ;
        RECT  3.4025 28.1625 3.4675 28.2975 ;
        RECT  3.0225 27.3225 3.0875 27.4575 ;
        RECT  3.2125 27.3225 3.2775 27.4575 ;
        RECT  3.0225 27.3225 3.0875 27.4575 ;
        RECT  3.2125 27.3225 3.2775 27.4575 ;
        RECT  3.2125 27.3225 3.2775 27.4575 ;
        RECT  3.4025 27.3225 3.4675 27.4575 ;
        RECT  3.2125 27.3225 3.2775 27.4575 ;
        RECT  3.4025 27.3225 3.4675 27.4575 ;
        RECT  3.5725 27.2775 3.6375 27.4125 ;
        RECT  3.5725 28.2075 3.6375 28.3425 ;
        RECT  3.2725 27.5525 3.4075 27.6175 ;
        RECT  3.015 27.7675 3.15 27.8325 ;
        RECT  3.2125 28.1625 3.2775 28.2975 ;
        RECT  3.4025 27.3225 3.4675 27.4575 ;
        RECT  3.3675 27.7675 3.5025 27.8325 ;
        RECT  3.5725 29.665 3.6375 29.85 ;
        RECT  3.5725 28.505 3.6375 28.735 ;
        RECT  3.0225 29.6875 3.0875 29.8825 ;
        RECT  3.0225 28.4725 3.0875 28.8475 ;
        RECT  3.4025 28.4725 3.4675 28.8475 ;
        RECT  3.015 29.1775 3.15 29.2425 ;
        RECT  3.3675 29.1775 3.5025 29.2425 ;
        RECT  3.2725 29.3925 3.4075 29.4575 ;
        RECT  2.955 28.4725 3.875 28.5375 ;
        RECT  2.955 29.8175 3.875 29.8825 ;
        RECT  3.0225 28.9825 3.0875 29.1175 ;
        RECT  3.2125 28.9825 3.2775 29.1175 ;
        RECT  3.0225 28.9825 3.0875 29.1175 ;
        RECT  3.2125 28.9825 3.2775 29.1175 ;
        RECT  3.2125 28.9825 3.2775 29.1175 ;
        RECT  3.4025 28.9825 3.4675 29.1175 ;
        RECT  3.2125 28.9825 3.2775 29.1175 ;
        RECT  3.4025 28.9825 3.4675 29.1175 ;
        RECT  3.0225 29.7325 3.0875 29.8675 ;
        RECT  3.2125 29.7325 3.2775 29.8675 ;
        RECT  3.0225 29.7325 3.0875 29.8675 ;
        RECT  3.2125 29.7325 3.2775 29.8675 ;
        RECT  3.2125 29.7325 3.2775 29.8675 ;
        RECT  3.4025 29.7325 3.4675 29.8675 ;
        RECT  3.2125 29.7325 3.2775 29.8675 ;
        RECT  3.4025 29.7325 3.4675 29.8675 ;
        RECT  3.5725 29.7325 3.6375 29.8675 ;
        RECT  3.5725 28.8025 3.6375 28.9375 ;
        RECT  3.2725 29.4675 3.4075 29.5325 ;
        RECT  3.015 29.2525 3.15 29.3175 ;
        RECT  3.2125 28.8475 3.2775 28.9825 ;
        RECT  3.4025 29.6875 3.4675 29.8225 ;
        RECT  3.3675 29.2475 3.5025 29.3125 ;
        RECT  3.5725 29.85 3.6375 30.035 ;
        RECT  3.5725 30.965 3.6375 31.195 ;
        RECT  3.0225 29.8175 3.0875 30.0125 ;
        RECT  3.0225 30.8525 3.0875 31.2275 ;
        RECT  3.4025 30.8525 3.4675 31.2275 ;
        RECT  3.015 30.4575 3.15 30.5225 ;
        RECT  3.3675 30.4575 3.5025 30.5225 ;
        RECT  3.2725 30.2425 3.4075 30.3075 ;
        RECT  2.955 31.1625 3.875 31.2275 ;
        RECT  2.955 29.8175 3.875 29.8825 ;
        RECT  3.0225 30.8525 3.0875 30.9875 ;
        RECT  3.2125 30.8525 3.2775 30.9875 ;
        RECT  3.0225 30.8525 3.0875 30.9875 ;
        RECT  3.2125 30.8525 3.2775 30.9875 ;
        RECT  3.2125 30.8525 3.2775 30.9875 ;
        RECT  3.4025 30.8525 3.4675 30.9875 ;
        RECT  3.2125 30.8525 3.2775 30.9875 ;
        RECT  3.4025 30.8525 3.4675 30.9875 ;
        RECT  3.0225 30.0125 3.0875 30.1475 ;
        RECT  3.2125 30.0125 3.2775 30.1475 ;
        RECT  3.0225 30.0125 3.0875 30.1475 ;
        RECT  3.2125 30.0125 3.2775 30.1475 ;
        RECT  3.2125 30.0125 3.2775 30.1475 ;
        RECT  3.4025 30.0125 3.4675 30.1475 ;
        RECT  3.2125 30.0125 3.2775 30.1475 ;
        RECT  3.4025 30.0125 3.4675 30.1475 ;
        RECT  3.5725 29.9675 3.6375 30.1025 ;
        RECT  3.5725 30.8975 3.6375 31.0325 ;
        RECT  3.2725 30.2425 3.4075 30.3075 ;
        RECT  3.015 30.4575 3.15 30.5225 ;
        RECT  3.2125 30.8525 3.2775 30.9875 ;
        RECT  3.4025 30.0125 3.4675 30.1475 ;
        RECT  3.3675 30.4575 3.5025 30.5225 ;
        RECT  3.5725 32.355 3.6375 32.54 ;
        RECT  3.5725 31.195 3.6375 31.425 ;
        RECT  3.0225 32.3775 3.0875 32.5725 ;
        RECT  3.0225 31.1625 3.0875 31.5375 ;
        RECT  3.4025 31.1625 3.4675 31.5375 ;
        RECT  3.015 31.8675 3.15 31.9325 ;
        RECT  3.3675 31.8675 3.5025 31.9325 ;
        RECT  3.2725 32.0825 3.4075 32.1475 ;
        RECT  2.955 31.1625 3.875 31.2275 ;
        RECT  2.955 32.5075 3.875 32.5725 ;
        RECT  3.0225 31.6725 3.0875 31.8075 ;
        RECT  3.2125 31.6725 3.2775 31.8075 ;
        RECT  3.0225 31.6725 3.0875 31.8075 ;
        RECT  3.2125 31.6725 3.2775 31.8075 ;
        RECT  3.2125 31.6725 3.2775 31.8075 ;
        RECT  3.4025 31.6725 3.4675 31.8075 ;
        RECT  3.2125 31.6725 3.2775 31.8075 ;
        RECT  3.4025 31.6725 3.4675 31.8075 ;
        RECT  3.0225 32.4225 3.0875 32.5575 ;
        RECT  3.2125 32.4225 3.2775 32.5575 ;
        RECT  3.0225 32.4225 3.0875 32.5575 ;
        RECT  3.2125 32.4225 3.2775 32.5575 ;
        RECT  3.2125 32.4225 3.2775 32.5575 ;
        RECT  3.4025 32.4225 3.4675 32.5575 ;
        RECT  3.2125 32.4225 3.2775 32.5575 ;
        RECT  3.4025 32.4225 3.4675 32.5575 ;
        RECT  3.5725 32.4225 3.6375 32.5575 ;
        RECT  3.5725 31.4925 3.6375 31.6275 ;
        RECT  3.2725 32.1575 3.4075 32.2225 ;
        RECT  3.015 31.9425 3.15 32.0075 ;
        RECT  3.2125 31.5375 3.2775 31.6725 ;
        RECT  3.4025 32.3775 3.4675 32.5125 ;
        RECT  3.3675 31.9375 3.5025 32.0025 ;
        RECT  3.5725 32.54 3.6375 32.725 ;
        RECT  3.5725 33.655 3.6375 33.885 ;
        RECT  3.0225 32.5075 3.0875 32.7025 ;
        RECT  3.0225 33.5425 3.0875 33.9175 ;
        RECT  3.4025 33.5425 3.4675 33.9175 ;
        RECT  3.015 33.1475 3.15 33.2125 ;
        RECT  3.3675 33.1475 3.5025 33.2125 ;
        RECT  3.2725 32.9325 3.4075 32.9975 ;
        RECT  2.955 33.8525 3.875 33.9175 ;
        RECT  2.955 32.5075 3.875 32.5725 ;
        RECT  3.0225 33.5425 3.0875 33.6775 ;
        RECT  3.2125 33.5425 3.2775 33.6775 ;
        RECT  3.0225 33.5425 3.0875 33.6775 ;
        RECT  3.2125 33.5425 3.2775 33.6775 ;
        RECT  3.2125 33.5425 3.2775 33.6775 ;
        RECT  3.4025 33.5425 3.4675 33.6775 ;
        RECT  3.2125 33.5425 3.2775 33.6775 ;
        RECT  3.4025 33.5425 3.4675 33.6775 ;
        RECT  3.0225 32.7025 3.0875 32.8375 ;
        RECT  3.2125 32.7025 3.2775 32.8375 ;
        RECT  3.0225 32.7025 3.0875 32.8375 ;
        RECT  3.2125 32.7025 3.2775 32.8375 ;
        RECT  3.2125 32.7025 3.2775 32.8375 ;
        RECT  3.4025 32.7025 3.4675 32.8375 ;
        RECT  3.2125 32.7025 3.2775 32.8375 ;
        RECT  3.4025 32.7025 3.4675 32.8375 ;
        RECT  3.5725 32.6575 3.6375 32.7925 ;
        RECT  3.5725 33.5875 3.6375 33.7225 ;
        RECT  3.2725 32.9325 3.4075 32.9975 ;
        RECT  3.015 33.1475 3.15 33.2125 ;
        RECT  3.2125 33.5425 3.2775 33.6775 ;
        RECT  3.4025 32.7025 3.4675 32.8375 ;
        RECT  3.3675 33.1475 3.5025 33.2125 ;
        RECT  3.5725 35.045 3.6375 35.23 ;
        RECT  3.5725 33.885 3.6375 34.115 ;
        RECT  3.0225 35.0675 3.0875 35.2625 ;
        RECT  3.0225 33.8525 3.0875 34.2275 ;
        RECT  3.4025 33.8525 3.4675 34.2275 ;
        RECT  3.015 34.5575 3.15 34.6225 ;
        RECT  3.3675 34.5575 3.5025 34.6225 ;
        RECT  3.2725 34.7725 3.4075 34.8375 ;
        RECT  2.955 33.8525 3.875 33.9175 ;
        RECT  2.955 35.1975 3.875 35.2625 ;
        RECT  3.0225 34.3625 3.0875 34.4975 ;
        RECT  3.2125 34.3625 3.2775 34.4975 ;
        RECT  3.0225 34.3625 3.0875 34.4975 ;
        RECT  3.2125 34.3625 3.2775 34.4975 ;
        RECT  3.2125 34.3625 3.2775 34.4975 ;
        RECT  3.4025 34.3625 3.4675 34.4975 ;
        RECT  3.2125 34.3625 3.2775 34.4975 ;
        RECT  3.4025 34.3625 3.4675 34.4975 ;
        RECT  3.0225 35.1125 3.0875 35.2475 ;
        RECT  3.2125 35.1125 3.2775 35.2475 ;
        RECT  3.0225 35.1125 3.0875 35.2475 ;
        RECT  3.2125 35.1125 3.2775 35.2475 ;
        RECT  3.2125 35.1125 3.2775 35.2475 ;
        RECT  3.4025 35.1125 3.4675 35.2475 ;
        RECT  3.2125 35.1125 3.2775 35.2475 ;
        RECT  3.4025 35.1125 3.4675 35.2475 ;
        RECT  3.5725 35.1125 3.6375 35.2475 ;
        RECT  3.5725 34.1825 3.6375 34.3175 ;
        RECT  3.2725 34.8475 3.4075 34.9125 ;
        RECT  3.015 34.6325 3.15 34.6975 ;
        RECT  3.2125 34.2275 3.2775 34.3625 ;
        RECT  3.4025 35.0675 3.4675 35.2025 ;
        RECT  3.3675 34.6275 3.5025 34.6925 ;
        RECT  3.5725 35.23 3.6375 35.415 ;
        RECT  3.5725 36.345 3.6375 36.575 ;
        RECT  3.0225 35.1975 3.0875 35.3925 ;
        RECT  3.0225 36.2325 3.0875 36.6075 ;
        RECT  3.4025 36.2325 3.4675 36.6075 ;
        RECT  3.015 35.8375 3.15 35.9025 ;
        RECT  3.3675 35.8375 3.5025 35.9025 ;
        RECT  3.2725 35.6225 3.4075 35.6875 ;
        RECT  2.955 36.5425 3.875 36.6075 ;
        RECT  2.955 35.1975 3.875 35.2625 ;
        RECT  3.0225 36.2325 3.0875 36.3675 ;
        RECT  3.2125 36.2325 3.2775 36.3675 ;
        RECT  3.0225 36.2325 3.0875 36.3675 ;
        RECT  3.2125 36.2325 3.2775 36.3675 ;
        RECT  3.2125 36.2325 3.2775 36.3675 ;
        RECT  3.4025 36.2325 3.4675 36.3675 ;
        RECT  3.2125 36.2325 3.2775 36.3675 ;
        RECT  3.4025 36.2325 3.4675 36.3675 ;
        RECT  3.0225 35.3925 3.0875 35.5275 ;
        RECT  3.2125 35.3925 3.2775 35.5275 ;
        RECT  3.0225 35.3925 3.0875 35.5275 ;
        RECT  3.2125 35.3925 3.2775 35.5275 ;
        RECT  3.2125 35.3925 3.2775 35.5275 ;
        RECT  3.4025 35.3925 3.4675 35.5275 ;
        RECT  3.2125 35.3925 3.2775 35.5275 ;
        RECT  3.4025 35.3925 3.4675 35.5275 ;
        RECT  3.5725 35.3475 3.6375 35.4825 ;
        RECT  3.5725 36.2775 3.6375 36.4125 ;
        RECT  3.2725 35.6225 3.4075 35.6875 ;
        RECT  3.015 35.8375 3.15 35.9025 ;
        RECT  3.2125 36.2325 3.2775 36.3675 ;
        RECT  3.4025 35.3925 3.4675 35.5275 ;
        RECT  3.3675 35.8375 3.5025 35.9025 ;
        RECT  3.5725 37.735 3.6375 37.92 ;
        RECT  3.5725 36.575 3.6375 36.805 ;
        RECT  3.0225 37.7575 3.0875 37.9525 ;
        RECT  3.0225 36.5425 3.0875 36.9175 ;
        RECT  3.4025 36.5425 3.4675 36.9175 ;
        RECT  3.015 37.2475 3.15 37.3125 ;
        RECT  3.3675 37.2475 3.5025 37.3125 ;
        RECT  3.2725 37.4625 3.4075 37.5275 ;
        RECT  2.955 36.5425 3.875 36.6075 ;
        RECT  2.955 37.8875 3.875 37.9525 ;
        RECT  3.0225 37.0525 3.0875 37.1875 ;
        RECT  3.2125 37.0525 3.2775 37.1875 ;
        RECT  3.0225 37.0525 3.0875 37.1875 ;
        RECT  3.2125 37.0525 3.2775 37.1875 ;
        RECT  3.2125 37.0525 3.2775 37.1875 ;
        RECT  3.4025 37.0525 3.4675 37.1875 ;
        RECT  3.2125 37.0525 3.2775 37.1875 ;
        RECT  3.4025 37.0525 3.4675 37.1875 ;
        RECT  3.0225 37.8025 3.0875 37.9375 ;
        RECT  3.2125 37.8025 3.2775 37.9375 ;
        RECT  3.0225 37.8025 3.0875 37.9375 ;
        RECT  3.2125 37.8025 3.2775 37.9375 ;
        RECT  3.2125 37.8025 3.2775 37.9375 ;
        RECT  3.4025 37.8025 3.4675 37.9375 ;
        RECT  3.2125 37.8025 3.2775 37.9375 ;
        RECT  3.4025 37.8025 3.4675 37.9375 ;
        RECT  3.5725 37.8025 3.6375 37.9375 ;
        RECT  3.5725 36.8725 3.6375 37.0075 ;
        RECT  3.2725 37.5375 3.4075 37.6025 ;
        RECT  3.015 37.3225 3.15 37.3875 ;
        RECT  3.2125 36.9175 3.2775 37.0525 ;
        RECT  3.4025 37.7575 3.4675 37.8925 ;
        RECT  3.3675 37.3175 3.5025 37.3825 ;
        RECT  3.5725 37.92 3.6375 38.105 ;
        RECT  3.5725 39.035 3.6375 39.265 ;
        RECT  3.0225 37.8875 3.0875 38.0825 ;
        RECT  3.0225 38.9225 3.0875 39.2975 ;
        RECT  3.4025 38.9225 3.4675 39.2975 ;
        RECT  3.015 38.5275 3.15 38.5925 ;
        RECT  3.3675 38.5275 3.5025 38.5925 ;
        RECT  3.2725 38.3125 3.4075 38.3775 ;
        RECT  2.955 39.2325 3.875 39.2975 ;
        RECT  2.955 37.8875 3.875 37.9525 ;
        RECT  3.0225 38.9225 3.0875 39.0575 ;
        RECT  3.2125 38.9225 3.2775 39.0575 ;
        RECT  3.0225 38.9225 3.0875 39.0575 ;
        RECT  3.2125 38.9225 3.2775 39.0575 ;
        RECT  3.2125 38.9225 3.2775 39.0575 ;
        RECT  3.4025 38.9225 3.4675 39.0575 ;
        RECT  3.2125 38.9225 3.2775 39.0575 ;
        RECT  3.4025 38.9225 3.4675 39.0575 ;
        RECT  3.0225 38.0825 3.0875 38.2175 ;
        RECT  3.2125 38.0825 3.2775 38.2175 ;
        RECT  3.0225 38.0825 3.0875 38.2175 ;
        RECT  3.2125 38.0825 3.2775 38.2175 ;
        RECT  3.2125 38.0825 3.2775 38.2175 ;
        RECT  3.4025 38.0825 3.4675 38.2175 ;
        RECT  3.2125 38.0825 3.2775 38.2175 ;
        RECT  3.4025 38.0825 3.4675 38.2175 ;
        RECT  3.5725 38.0375 3.6375 38.1725 ;
        RECT  3.5725 38.9675 3.6375 39.1025 ;
        RECT  3.2725 38.3125 3.4075 38.3775 ;
        RECT  3.015 38.5275 3.15 38.5925 ;
        RECT  3.2125 38.9225 3.2775 39.0575 ;
        RECT  3.4025 38.0825 3.4675 38.2175 ;
        RECT  3.3675 38.5275 3.5025 38.5925 ;
        RECT  3.5725 40.425 3.6375 40.61 ;
        RECT  3.5725 39.265 3.6375 39.495 ;
        RECT  3.0225 40.4475 3.0875 40.6425 ;
        RECT  3.0225 39.2325 3.0875 39.6075 ;
        RECT  3.4025 39.2325 3.4675 39.6075 ;
        RECT  3.015 39.9375 3.15 40.0025 ;
        RECT  3.3675 39.9375 3.5025 40.0025 ;
        RECT  3.2725 40.1525 3.4075 40.2175 ;
        RECT  2.955 39.2325 3.875 39.2975 ;
        RECT  2.955 40.5775 3.875 40.6425 ;
        RECT  3.0225 39.7425 3.0875 39.8775 ;
        RECT  3.2125 39.7425 3.2775 39.8775 ;
        RECT  3.0225 39.7425 3.0875 39.8775 ;
        RECT  3.2125 39.7425 3.2775 39.8775 ;
        RECT  3.2125 39.7425 3.2775 39.8775 ;
        RECT  3.4025 39.7425 3.4675 39.8775 ;
        RECT  3.2125 39.7425 3.2775 39.8775 ;
        RECT  3.4025 39.7425 3.4675 39.8775 ;
        RECT  3.0225 40.4925 3.0875 40.6275 ;
        RECT  3.2125 40.4925 3.2775 40.6275 ;
        RECT  3.0225 40.4925 3.0875 40.6275 ;
        RECT  3.2125 40.4925 3.2775 40.6275 ;
        RECT  3.2125 40.4925 3.2775 40.6275 ;
        RECT  3.4025 40.4925 3.4675 40.6275 ;
        RECT  3.2125 40.4925 3.2775 40.6275 ;
        RECT  3.4025 40.4925 3.4675 40.6275 ;
        RECT  3.5725 40.4925 3.6375 40.6275 ;
        RECT  3.5725 39.5625 3.6375 39.6975 ;
        RECT  3.2725 40.2275 3.4075 40.2925 ;
        RECT  3.015 40.0125 3.15 40.0775 ;
        RECT  3.2125 39.6075 3.2775 39.7425 ;
        RECT  3.4025 40.4475 3.4675 40.5825 ;
        RECT  3.3675 40.0075 3.5025 40.0725 ;
        RECT  4.3025 19.09 4.3675 19.275 ;
        RECT  4.3025 20.205 4.3675 20.435 ;
        RECT  3.9425 19.0575 4.0075 19.2075 ;
        RECT  3.9425 20.0925 4.0075 20.4675 ;
        RECT  4.1325 19.3425 4.1975 20.0925 ;
        RECT  4.0 19.605 4.065 19.74 ;
        RECT  4.165 19.64 4.23 19.705 ;
        RECT  3.875 20.4025 4.435 20.4675 ;
        RECT  3.875 19.0575 4.435 19.1225 ;
        RECT  3.9425 20.0925 4.0075 20.2275 ;
        RECT  4.1325 20.0925 4.1975 20.2275 ;
        RECT  3.9425 20.0925 4.0075 20.2275 ;
        RECT  4.1325 20.0925 4.1975 20.2275 ;
        RECT  3.9425 19.2075 4.0075 19.3425 ;
        RECT  4.1325 19.2075 4.1975 19.3425 ;
        RECT  3.9425 19.2075 4.0075 19.3425 ;
        RECT  4.1325 19.2075 4.1975 19.3425 ;
        RECT  4.3025 19.2075 4.3675 19.3425 ;
        RECT  4.3025 20.1375 4.3675 20.2725 ;
        RECT  4.0 19.605 4.065 19.74 ;
        RECT  4.3025 21.595 4.3675 21.78 ;
        RECT  4.3025 20.435 4.3675 20.665 ;
        RECT  3.9425 21.6625 4.0075 21.8125 ;
        RECT  3.9425 20.4025 4.0075 20.7775 ;
        RECT  4.1325 20.7775 4.1975 21.5275 ;
        RECT  4.0 21.13 4.065 21.265 ;
        RECT  4.165 21.165 4.23 21.23 ;
        RECT  3.875 20.4025 4.435 20.4675 ;
        RECT  3.875 21.7475 4.435 21.8125 ;
        RECT  3.9425 20.9125 4.0075 21.0475 ;
        RECT  4.1325 20.9125 4.1975 21.0475 ;
        RECT  3.9425 20.9125 4.0075 21.0475 ;
        RECT  4.1325 20.9125 4.1975 21.0475 ;
        RECT  3.9425 21.6175 4.0075 21.7525 ;
        RECT  4.1325 21.6175 4.1975 21.7525 ;
        RECT  3.9425 21.6175 4.0075 21.7525 ;
        RECT  4.1325 21.6175 4.1975 21.7525 ;
        RECT  4.3025 21.6625 4.3675 21.7975 ;
        RECT  4.3025 20.7325 4.3675 20.8675 ;
        RECT  4.0 21.265 4.065 21.4 ;
        RECT  4.3025 21.78 4.3675 21.965 ;
        RECT  4.3025 22.895 4.3675 23.125 ;
        RECT  3.9425 21.7475 4.0075 21.8975 ;
        RECT  3.9425 22.7825 4.0075 23.1575 ;
        RECT  4.1325 22.0325 4.1975 22.7825 ;
        RECT  4.0 22.295 4.065 22.43 ;
        RECT  4.165 22.33 4.23 22.395 ;
        RECT  3.875 23.0925 4.435 23.1575 ;
        RECT  3.875 21.7475 4.435 21.8125 ;
        RECT  3.9425 22.7825 4.0075 22.9175 ;
        RECT  4.1325 22.7825 4.1975 22.9175 ;
        RECT  3.9425 22.7825 4.0075 22.9175 ;
        RECT  4.1325 22.7825 4.1975 22.9175 ;
        RECT  3.9425 21.8975 4.0075 22.0325 ;
        RECT  4.1325 21.8975 4.1975 22.0325 ;
        RECT  3.9425 21.8975 4.0075 22.0325 ;
        RECT  4.1325 21.8975 4.1975 22.0325 ;
        RECT  4.3025 21.8975 4.3675 22.0325 ;
        RECT  4.3025 22.8275 4.3675 22.9625 ;
        RECT  4.0 22.295 4.065 22.43 ;
        RECT  4.3025 24.285 4.3675 24.47 ;
        RECT  4.3025 23.125 4.3675 23.355 ;
        RECT  3.9425 24.3525 4.0075 24.5025 ;
        RECT  3.9425 23.0925 4.0075 23.4675 ;
        RECT  4.1325 23.4675 4.1975 24.2175 ;
        RECT  4.0 23.82 4.065 23.955 ;
        RECT  4.165 23.855 4.23 23.92 ;
        RECT  3.875 23.0925 4.435 23.1575 ;
        RECT  3.875 24.4375 4.435 24.5025 ;
        RECT  3.9425 23.6025 4.0075 23.7375 ;
        RECT  4.1325 23.6025 4.1975 23.7375 ;
        RECT  3.9425 23.6025 4.0075 23.7375 ;
        RECT  4.1325 23.6025 4.1975 23.7375 ;
        RECT  3.9425 24.3075 4.0075 24.4425 ;
        RECT  4.1325 24.3075 4.1975 24.4425 ;
        RECT  3.9425 24.3075 4.0075 24.4425 ;
        RECT  4.1325 24.3075 4.1975 24.4425 ;
        RECT  4.3025 24.3525 4.3675 24.4875 ;
        RECT  4.3025 23.4225 4.3675 23.5575 ;
        RECT  4.0 23.955 4.065 24.09 ;
        RECT  4.3025 24.47 4.3675 24.655 ;
        RECT  4.3025 25.585 4.3675 25.815 ;
        RECT  3.9425 24.4375 4.0075 24.5875 ;
        RECT  3.9425 25.4725 4.0075 25.8475 ;
        RECT  4.1325 24.7225 4.1975 25.4725 ;
        RECT  4.0 24.985 4.065 25.12 ;
        RECT  4.165 25.02 4.23 25.085 ;
        RECT  3.875 25.7825 4.435 25.8475 ;
        RECT  3.875 24.4375 4.435 24.5025 ;
        RECT  3.9425 25.4725 4.0075 25.6075 ;
        RECT  4.1325 25.4725 4.1975 25.6075 ;
        RECT  3.9425 25.4725 4.0075 25.6075 ;
        RECT  4.1325 25.4725 4.1975 25.6075 ;
        RECT  3.9425 24.5875 4.0075 24.7225 ;
        RECT  4.1325 24.5875 4.1975 24.7225 ;
        RECT  3.9425 24.5875 4.0075 24.7225 ;
        RECT  4.1325 24.5875 4.1975 24.7225 ;
        RECT  4.3025 24.5875 4.3675 24.7225 ;
        RECT  4.3025 25.5175 4.3675 25.6525 ;
        RECT  4.0 24.985 4.065 25.12 ;
        RECT  4.3025 26.975 4.3675 27.16 ;
        RECT  4.3025 25.815 4.3675 26.045 ;
        RECT  3.9425 27.0425 4.0075 27.1925 ;
        RECT  3.9425 25.7825 4.0075 26.1575 ;
        RECT  4.1325 26.1575 4.1975 26.9075 ;
        RECT  4.0 26.51 4.065 26.645 ;
        RECT  4.165 26.545 4.23 26.61 ;
        RECT  3.875 25.7825 4.435 25.8475 ;
        RECT  3.875 27.1275 4.435 27.1925 ;
        RECT  3.9425 26.2925 4.0075 26.4275 ;
        RECT  4.1325 26.2925 4.1975 26.4275 ;
        RECT  3.9425 26.2925 4.0075 26.4275 ;
        RECT  4.1325 26.2925 4.1975 26.4275 ;
        RECT  3.9425 26.9975 4.0075 27.1325 ;
        RECT  4.1325 26.9975 4.1975 27.1325 ;
        RECT  3.9425 26.9975 4.0075 27.1325 ;
        RECT  4.1325 26.9975 4.1975 27.1325 ;
        RECT  4.3025 27.0425 4.3675 27.1775 ;
        RECT  4.3025 26.1125 4.3675 26.2475 ;
        RECT  4.0 26.645 4.065 26.78 ;
        RECT  4.3025 27.16 4.3675 27.345 ;
        RECT  4.3025 28.275 4.3675 28.505 ;
        RECT  3.9425 27.1275 4.0075 27.2775 ;
        RECT  3.9425 28.1625 4.0075 28.5375 ;
        RECT  4.1325 27.4125 4.1975 28.1625 ;
        RECT  4.0 27.675 4.065 27.81 ;
        RECT  4.165 27.71 4.23 27.775 ;
        RECT  3.875 28.4725 4.435 28.5375 ;
        RECT  3.875 27.1275 4.435 27.1925 ;
        RECT  3.9425 28.1625 4.0075 28.2975 ;
        RECT  4.1325 28.1625 4.1975 28.2975 ;
        RECT  3.9425 28.1625 4.0075 28.2975 ;
        RECT  4.1325 28.1625 4.1975 28.2975 ;
        RECT  3.9425 27.2775 4.0075 27.4125 ;
        RECT  4.1325 27.2775 4.1975 27.4125 ;
        RECT  3.9425 27.2775 4.0075 27.4125 ;
        RECT  4.1325 27.2775 4.1975 27.4125 ;
        RECT  4.3025 27.2775 4.3675 27.4125 ;
        RECT  4.3025 28.2075 4.3675 28.3425 ;
        RECT  4.0 27.675 4.065 27.81 ;
        RECT  4.3025 29.665 4.3675 29.85 ;
        RECT  4.3025 28.505 4.3675 28.735 ;
        RECT  3.9425 29.7325 4.0075 29.8825 ;
        RECT  3.9425 28.4725 4.0075 28.8475 ;
        RECT  4.1325 28.8475 4.1975 29.5975 ;
        RECT  4.0 29.2 4.065 29.335 ;
        RECT  4.165 29.235 4.23 29.3 ;
        RECT  3.875 28.4725 4.435 28.5375 ;
        RECT  3.875 29.8175 4.435 29.8825 ;
        RECT  3.9425 28.9825 4.0075 29.1175 ;
        RECT  4.1325 28.9825 4.1975 29.1175 ;
        RECT  3.9425 28.9825 4.0075 29.1175 ;
        RECT  4.1325 28.9825 4.1975 29.1175 ;
        RECT  3.9425 29.6875 4.0075 29.8225 ;
        RECT  4.1325 29.6875 4.1975 29.8225 ;
        RECT  3.9425 29.6875 4.0075 29.8225 ;
        RECT  4.1325 29.6875 4.1975 29.8225 ;
        RECT  4.3025 29.7325 4.3675 29.8675 ;
        RECT  4.3025 28.8025 4.3675 28.9375 ;
        RECT  4.0 29.335 4.065 29.47 ;
        RECT  4.3025 29.85 4.3675 30.035 ;
        RECT  4.3025 30.965 4.3675 31.195 ;
        RECT  3.9425 29.8175 4.0075 29.9675 ;
        RECT  3.9425 30.8525 4.0075 31.2275 ;
        RECT  4.1325 30.1025 4.1975 30.8525 ;
        RECT  4.0 30.365 4.065 30.5 ;
        RECT  4.165 30.4 4.23 30.465 ;
        RECT  3.875 31.1625 4.435 31.2275 ;
        RECT  3.875 29.8175 4.435 29.8825 ;
        RECT  3.9425 30.8525 4.0075 30.9875 ;
        RECT  4.1325 30.8525 4.1975 30.9875 ;
        RECT  3.9425 30.8525 4.0075 30.9875 ;
        RECT  4.1325 30.8525 4.1975 30.9875 ;
        RECT  3.9425 29.9675 4.0075 30.1025 ;
        RECT  4.1325 29.9675 4.1975 30.1025 ;
        RECT  3.9425 29.9675 4.0075 30.1025 ;
        RECT  4.1325 29.9675 4.1975 30.1025 ;
        RECT  4.3025 29.9675 4.3675 30.1025 ;
        RECT  4.3025 30.8975 4.3675 31.0325 ;
        RECT  4.0 30.365 4.065 30.5 ;
        RECT  4.3025 32.355 4.3675 32.54 ;
        RECT  4.3025 31.195 4.3675 31.425 ;
        RECT  3.9425 32.4225 4.0075 32.5725 ;
        RECT  3.9425 31.1625 4.0075 31.5375 ;
        RECT  4.1325 31.5375 4.1975 32.2875 ;
        RECT  4.0 31.89 4.065 32.025 ;
        RECT  4.165 31.925 4.23 31.99 ;
        RECT  3.875 31.1625 4.435 31.2275 ;
        RECT  3.875 32.5075 4.435 32.5725 ;
        RECT  3.9425 31.6725 4.0075 31.8075 ;
        RECT  4.1325 31.6725 4.1975 31.8075 ;
        RECT  3.9425 31.6725 4.0075 31.8075 ;
        RECT  4.1325 31.6725 4.1975 31.8075 ;
        RECT  3.9425 32.3775 4.0075 32.5125 ;
        RECT  4.1325 32.3775 4.1975 32.5125 ;
        RECT  3.9425 32.3775 4.0075 32.5125 ;
        RECT  4.1325 32.3775 4.1975 32.5125 ;
        RECT  4.3025 32.4225 4.3675 32.5575 ;
        RECT  4.3025 31.4925 4.3675 31.6275 ;
        RECT  4.0 32.025 4.065 32.16 ;
        RECT  4.3025 32.54 4.3675 32.725 ;
        RECT  4.3025 33.655 4.3675 33.885 ;
        RECT  3.9425 32.5075 4.0075 32.6575 ;
        RECT  3.9425 33.5425 4.0075 33.9175 ;
        RECT  4.1325 32.7925 4.1975 33.5425 ;
        RECT  4.0 33.055 4.065 33.19 ;
        RECT  4.165 33.09 4.23 33.155 ;
        RECT  3.875 33.8525 4.435 33.9175 ;
        RECT  3.875 32.5075 4.435 32.5725 ;
        RECT  3.9425 33.5425 4.0075 33.6775 ;
        RECT  4.1325 33.5425 4.1975 33.6775 ;
        RECT  3.9425 33.5425 4.0075 33.6775 ;
        RECT  4.1325 33.5425 4.1975 33.6775 ;
        RECT  3.9425 32.6575 4.0075 32.7925 ;
        RECT  4.1325 32.6575 4.1975 32.7925 ;
        RECT  3.9425 32.6575 4.0075 32.7925 ;
        RECT  4.1325 32.6575 4.1975 32.7925 ;
        RECT  4.3025 32.6575 4.3675 32.7925 ;
        RECT  4.3025 33.5875 4.3675 33.7225 ;
        RECT  4.0 33.055 4.065 33.19 ;
        RECT  4.3025 35.045 4.3675 35.23 ;
        RECT  4.3025 33.885 4.3675 34.115 ;
        RECT  3.9425 35.1125 4.0075 35.2625 ;
        RECT  3.9425 33.8525 4.0075 34.2275 ;
        RECT  4.1325 34.2275 4.1975 34.9775 ;
        RECT  4.0 34.58 4.065 34.715 ;
        RECT  4.165 34.615 4.23 34.68 ;
        RECT  3.875 33.8525 4.435 33.9175 ;
        RECT  3.875 35.1975 4.435 35.2625 ;
        RECT  3.9425 34.3625 4.0075 34.4975 ;
        RECT  4.1325 34.3625 4.1975 34.4975 ;
        RECT  3.9425 34.3625 4.0075 34.4975 ;
        RECT  4.1325 34.3625 4.1975 34.4975 ;
        RECT  3.9425 35.0675 4.0075 35.2025 ;
        RECT  4.1325 35.0675 4.1975 35.2025 ;
        RECT  3.9425 35.0675 4.0075 35.2025 ;
        RECT  4.1325 35.0675 4.1975 35.2025 ;
        RECT  4.3025 35.1125 4.3675 35.2475 ;
        RECT  4.3025 34.1825 4.3675 34.3175 ;
        RECT  4.0 34.715 4.065 34.85 ;
        RECT  4.3025 35.23 4.3675 35.415 ;
        RECT  4.3025 36.345 4.3675 36.575 ;
        RECT  3.9425 35.1975 4.0075 35.3475 ;
        RECT  3.9425 36.2325 4.0075 36.6075 ;
        RECT  4.1325 35.4825 4.1975 36.2325 ;
        RECT  4.0 35.745 4.065 35.88 ;
        RECT  4.165 35.78 4.23 35.845 ;
        RECT  3.875 36.5425 4.435 36.6075 ;
        RECT  3.875 35.1975 4.435 35.2625 ;
        RECT  3.9425 36.2325 4.0075 36.3675 ;
        RECT  4.1325 36.2325 4.1975 36.3675 ;
        RECT  3.9425 36.2325 4.0075 36.3675 ;
        RECT  4.1325 36.2325 4.1975 36.3675 ;
        RECT  3.9425 35.3475 4.0075 35.4825 ;
        RECT  4.1325 35.3475 4.1975 35.4825 ;
        RECT  3.9425 35.3475 4.0075 35.4825 ;
        RECT  4.1325 35.3475 4.1975 35.4825 ;
        RECT  4.3025 35.3475 4.3675 35.4825 ;
        RECT  4.3025 36.2775 4.3675 36.4125 ;
        RECT  4.0 35.745 4.065 35.88 ;
        RECT  4.3025 37.735 4.3675 37.92 ;
        RECT  4.3025 36.575 4.3675 36.805 ;
        RECT  3.9425 37.8025 4.0075 37.9525 ;
        RECT  3.9425 36.5425 4.0075 36.9175 ;
        RECT  4.1325 36.9175 4.1975 37.6675 ;
        RECT  4.0 37.27 4.065 37.405 ;
        RECT  4.165 37.305 4.23 37.37 ;
        RECT  3.875 36.5425 4.435 36.6075 ;
        RECT  3.875 37.8875 4.435 37.9525 ;
        RECT  3.9425 37.0525 4.0075 37.1875 ;
        RECT  4.1325 37.0525 4.1975 37.1875 ;
        RECT  3.9425 37.0525 4.0075 37.1875 ;
        RECT  4.1325 37.0525 4.1975 37.1875 ;
        RECT  3.9425 37.7575 4.0075 37.8925 ;
        RECT  4.1325 37.7575 4.1975 37.8925 ;
        RECT  3.9425 37.7575 4.0075 37.8925 ;
        RECT  4.1325 37.7575 4.1975 37.8925 ;
        RECT  4.3025 37.8025 4.3675 37.9375 ;
        RECT  4.3025 36.8725 4.3675 37.0075 ;
        RECT  4.0 37.405 4.065 37.54 ;
        RECT  4.3025 37.92 4.3675 38.105 ;
        RECT  4.3025 39.035 4.3675 39.265 ;
        RECT  3.9425 37.8875 4.0075 38.0375 ;
        RECT  3.9425 38.9225 4.0075 39.2975 ;
        RECT  4.1325 38.1725 4.1975 38.9225 ;
        RECT  4.0 38.435 4.065 38.57 ;
        RECT  4.165 38.47 4.23 38.535 ;
        RECT  3.875 39.2325 4.435 39.2975 ;
        RECT  3.875 37.8875 4.435 37.9525 ;
        RECT  3.9425 38.9225 4.0075 39.0575 ;
        RECT  4.1325 38.9225 4.1975 39.0575 ;
        RECT  3.9425 38.9225 4.0075 39.0575 ;
        RECT  4.1325 38.9225 4.1975 39.0575 ;
        RECT  3.9425 38.0375 4.0075 38.1725 ;
        RECT  4.1325 38.0375 4.1975 38.1725 ;
        RECT  3.9425 38.0375 4.0075 38.1725 ;
        RECT  4.1325 38.0375 4.1975 38.1725 ;
        RECT  4.3025 38.0375 4.3675 38.1725 ;
        RECT  4.3025 38.9675 4.3675 39.1025 ;
        RECT  4.0 38.435 4.065 38.57 ;
        RECT  4.3025 40.425 4.3675 40.61 ;
        RECT  4.3025 39.265 4.3675 39.495 ;
        RECT  3.9425 40.4925 4.0075 40.6425 ;
        RECT  3.9425 39.2325 4.0075 39.6075 ;
        RECT  4.1325 39.6075 4.1975 40.3575 ;
        RECT  4.0 39.96 4.065 40.095 ;
        RECT  4.165 39.995 4.23 40.06 ;
        RECT  3.875 39.2325 4.435 39.2975 ;
        RECT  3.875 40.5775 4.435 40.6425 ;
        RECT  3.9425 39.7425 4.0075 39.8775 ;
        RECT  4.1325 39.7425 4.1975 39.8775 ;
        RECT  3.9425 39.7425 4.0075 39.8775 ;
        RECT  4.1325 39.7425 4.1975 39.8775 ;
        RECT  3.9425 40.4475 4.0075 40.5825 ;
        RECT  4.1325 40.4475 4.1975 40.5825 ;
        RECT  3.9425 40.4475 4.0075 40.5825 ;
        RECT  4.1325 40.4475 4.1975 40.5825 ;
        RECT  4.3025 40.4925 4.3675 40.6275 ;
        RECT  4.3025 39.5625 4.3675 39.6975 ;
        RECT  4.0 40.095 4.065 40.23 ;
        RECT  1.5225 8.88 1.6575 8.945 ;
        RECT  1.6975 10.405 1.8325 10.47 ;
        RECT  1.8725 11.57 2.0075 11.635 ;
        RECT  2.0475 13.095 2.1825 13.16 ;
        RECT  2.2225 14.26 2.3575 14.325 ;
        RECT  2.3975 15.785 2.5325 15.85 ;
        RECT  2.5725 16.95 2.7075 17.015 ;
        RECT  2.7475 18.475 2.8825 18.54 ;
        RECT  1.5225 19.6975 1.6575 19.7625 ;
        RECT  2.2225 19.4825 2.3575 19.5475 ;
        RECT  1.5225 21.1075 1.6575 21.1725 ;
        RECT  2.3975 21.3225 2.5325 21.3875 ;
        RECT  1.5225 22.3875 1.6575 22.4525 ;
        RECT  2.5725 22.1725 2.7075 22.2375 ;
        RECT  1.5225 23.7975 1.6575 23.8625 ;
        RECT  2.7475 24.0125 2.8825 24.0775 ;
        RECT  1.6975 25.0775 1.8325 25.1425 ;
        RECT  2.2225 24.8625 2.3575 24.9275 ;
        RECT  1.6975 26.4875 1.8325 26.5525 ;
        RECT  2.3975 26.7025 2.5325 26.7675 ;
        RECT  1.6975 27.7675 1.8325 27.8325 ;
        RECT  2.5725 27.5525 2.7075 27.6175 ;
        RECT  1.6975 29.1775 1.8325 29.2425 ;
        RECT  2.7475 29.3925 2.8825 29.4575 ;
        RECT  1.8725 30.4575 2.0075 30.5225 ;
        RECT  2.2225 30.2425 2.3575 30.3075 ;
        RECT  1.8725 31.8675 2.0075 31.9325 ;
        RECT  2.3975 32.0825 2.5325 32.1475 ;
        RECT  1.8725 33.1475 2.0075 33.2125 ;
        RECT  2.5725 32.9325 2.7075 32.9975 ;
        RECT  1.8725 34.5575 2.0075 34.6225 ;
        RECT  2.7475 34.7725 2.8825 34.8375 ;
        RECT  2.0475 35.8375 2.1825 35.9025 ;
        RECT  2.2225 35.6225 2.3575 35.6875 ;
        RECT  2.0475 37.2475 2.1825 37.3125 ;
        RECT  2.3975 37.4625 2.5325 37.5275 ;
        RECT  2.0475 38.5275 2.1825 38.5925 ;
        RECT  2.5725 38.3125 2.7075 38.3775 ;
        RECT  2.0475 39.9375 2.1825 40.0025 ;
        RECT  2.7475 40.1525 2.8825 40.2175 ;
        RECT  4.665 19.64 5.015 19.705 ;
        RECT  5.18 19.6975 5.245 19.7625 ;
        RECT  5.18 19.64 5.245 19.705 ;
        RECT  5.18 19.705 5.245 19.73 ;
        RECT  5.2125 19.6975 5.51 19.7625 ;
        RECT  5.51 19.6975 5.645 19.7625 ;
        RECT  6.215 19.6975 6.28 19.7625 ;
        RECT  6.215 19.64 6.28 19.705 ;
        RECT  5.9975 19.6975 6.2475 19.7625 ;
        RECT  6.215 19.6725 6.28 19.73 ;
        RECT  6.2475 19.64 6.495 19.705 ;
        RECT  4.665 21.165 5.015 21.23 ;
        RECT  5.18 21.1075 5.245 21.1725 ;
        RECT  5.18 21.165 5.245 21.23 ;
        RECT  5.18 21.14 5.245 21.23 ;
        RECT  5.2125 21.1075 5.51 21.1725 ;
        RECT  5.51 21.1075 5.645 21.1725 ;
        RECT  6.215 21.1075 6.28 21.1725 ;
        RECT  6.215 21.165 6.28 21.23 ;
        RECT  5.9975 21.1075 6.2475 21.1725 ;
        RECT  6.215 21.14 6.28 21.1975 ;
        RECT  6.2475 21.165 6.495 21.23 ;
        RECT  4.665 22.33 5.015 22.395 ;
        RECT  5.18 22.3875 5.245 22.4525 ;
        RECT  5.18 22.33 5.245 22.395 ;
        RECT  5.18 22.395 5.245 22.42 ;
        RECT  5.2125 22.3875 5.51 22.4525 ;
        RECT  5.51 22.3875 5.645 22.4525 ;
        RECT  6.215 22.3875 6.28 22.4525 ;
        RECT  6.215 22.33 6.28 22.395 ;
        RECT  5.9975 22.3875 6.2475 22.4525 ;
        RECT  6.215 22.3625 6.28 22.42 ;
        RECT  6.2475 22.33 6.495 22.395 ;
        RECT  4.665 23.855 5.015 23.92 ;
        RECT  5.18 23.7975 5.245 23.8625 ;
        RECT  5.18 23.855 5.245 23.92 ;
        RECT  5.18 23.83 5.245 23.92 ;
        RECT  5.2125 23.7975 5.51 23.8625 ;
        RECT  5.51 23.7975 5.645 23.8625 ;
        RECT  6.215 23.7975 6.28 23.8625 ;
        RECT  6.215 23.855 6.28 23.92 ;
        RECT  5.9975 23.7975 6.2475 23.8625 ;
        RECT  6.215 23.83 6.28 23.8875 ;
        RECT  6.2475 23.855 6.495 23.92 ;
        RECT  4.665 25.02 5.015 25.085 ;
        RECT  5.18 25.0775 5.245 25.1425 ;
        RECT  5.18 25.02 5.245 25.085 ;
        RECT  5.18 25.085 5.245 25.11 ;
        RECT  5.2125 25.0775 5.51 25.1425 ;
        RECT  5.51 25.0775 5.645 25.1425 ;
        RECT  6.215 25.0775 6.28 25.1425 ;
        RECT  6.215 25.02 6.28 25.085 ;
        RECT  5.9975 25.0775 6.2475 25.1425 ;
        RECT  6.215 25.0525 6.28 25.11 ;
        RECT  6.2475 25.02 6.495 25.085 ;
        RECT  4.665 26.545 5.015 26.61 ;
        RECT  5.18 26.4875 5.245 26.5525 ;
        RECT  5.18 26.545 5.245 26.61 ;
        RECT  5.18 26.52 5.245 26.61 ;
        RECT  5.2125 26.4875 5.51 26.5525 ;
        RECT  5.51 26.4875 5.645 26.5525 ;
        RECT  6.215 26.4875 6.28 26.5525 ;
        RECT  6.215 26.545 6.28 26.61 ;
        RECT  5.9975 26.4875 6.2475 26.5525 ;
        RECT  6.215 26.52 6.28 26.5775 ;
        RECT  6.2475 26.545 6.495 26.61 ;
        RECT  4.665 27.71 5.015 27.775 ;
        RECT  5.18 27.7675 5.245 27.8325 ;
        RECT  5.18 27.71 5.245 27.775 ;
        RECT  5.18 27.775 5.245 27.8 ;
        RECT  5.2125 27.7675 5.51 27.8325 ;
        RECT  5.51 27.7675 5.645 27.8325 ;
        RECT  6.215 27.7675 6.28 27.8325 ;
        RECT  6.215 27.71 6.28 27.775 ;
        RECT  5.9975 27.7675 6.2475 27.8325 ;
        RECT  6.215 27.7425 6.28 27.8 ;
        RECT  6.2475 27.71 6.495 27.775 ;
        RECT  4.665 29.235 5.015 29.3 ;
        RECT  5.18 29.1775 5.245 29.2425 ;
        RECT  5.18 29.235 5.245 29.3 ;
        RECT  5.18 29.21 5.245 29.3 ;
        RECT  5.2125 29.1775 5.51 29.2425 ;
        RECT  5.51 29.1775 5.645 29.2425 ;
        RECT  6.215 29.1775 6.28 29.2425 ;
        RECT  6.215 29.235 6.28 29.3 ;
        RECT  5.9975 29.1775 6.2475 29.2425 ;
        RECT  6.215 29.21 6.28 29.2675 ;
        RECT  6.2475 29.235 6.495 29.3 ;
        RECT  4.665 30.4 5.015 30.465 ;
        RECT  5.18 30.4575 5.245 30.5225 ;
        RECT  5.18 30.4 5.245 30.465 ;
        RECT  5.18 30.465 5.245 30.49 ;
        RECT  5.2125 30.4575 5.51 30.5225 ;
        RECT  5.51 30.4575 5.645 30.5225 ;
        RECT  6.215 30.4575 6.28 30.5225 ;
        RECT  6.215 30.4 6.28 30.465 ;
        RECT  5.9975 30.4575 6.2475 30.5225 ;
        RECT  6.215 30.4325 6.28 30.49 ;
        RECT  6.2475 30.4 6.495 30.465 ;
        RECT  4.665 31.925 5.015 31.99 ;
        RECT  5.18 31.8675 5.245 31.9325 ;
        RECT  5.18 31.925 5.245 31.99 ;
        RECT  5.18 31.9 5.245 31.99 ;
        RECT  5.2125 31.8675 5.51 31.9325 ;
        RECT  5.51 31.8675 5.645 31.9325 ;
        RECT  6.215 31.8675 6.28 31.9325 ;
        RECT  6.215 31.925 6.28 31.99 ;
        RECT  5.9975 31.8675 6.2475 31.9325 ;
        RECT  6.215 31.9 6.28 31.9575 ;
        RECT  6.2475 31.925 6.495 31.99 ;
        RECT  4.665 33.09 5.015 33.155 ;
        RECT  5.18 33.1475 5.245 33.2125 ;
        RECT  5.18 33.09 5.245 33.155 ;
        RECT  5.18 33.155 5.245 33.18 ;
        RECT  5.2125 33.1475 5.51 33.2125 ;
        RECT  5.51 33.1475 5.645 33.2125 ;
        RECT  6.215 33.1475 6.28 33.2125 ;
        RECT  6.215 33.09 6.28 33.155 ;
        RECT  5.9975 33.1475 6.2475 33.2125 ;
        RECT  6.215 33.1225 6.28 33.18 ;
        RECT  6.2475 33.09 6.495 33.155 ;
        RECT  4.665 34.615 5.015 34.68 ;
        RECT  5.18 34.5575 5.245 34.6225 ;
        RECT  5.18 34.615 5.245 34.68 ;
        RECT  5.18 34.59 5.245 34.68 ;
        RECT  5.2125 34.5575 5.51 34.6225 ;
        RECT  5.51 34.5575 5.645 34.6225 ;
        RECT  6.215 34.5575 6.28 34.6225 ;
        RECT  6.215 34.615 6.28 34.68 ;
        RECT  5.9975 34.5575 6.2475 34.6225 ;
        RECT  6.215 34.59 6.28 34.6475 ;
        RECT  6.2475 34.615 6.495 34.68 ;
        RECT  4.665 35.78 5.015 35.845 ;
        RECT  5.18 35.8375 5.245 35.9025 ;
        RECT  5.18 35.78 5.245 35.845 ;
        RECT  5.18 35.845 5.245 35.87 ;
        RECT  5.2125 35.8375 5.51 35.9025 ;
        RECT  5.51 35.8375 5.645 35.9025 ;
        RECT  6.215 35.8375 6.28 35.9025 ;
        RECT  6.215 35.78 6.28 35.845 ;
        RECT  5.9975 35.8375 6.2475 35.9025 ;
        RECT  6.215 35.8125 6.28 35.87 ;
        RECT  6.2475 35.78 6.495 35.845 ;
        RECT  4.665 37.305 5.015 37.37 ;
        RECT  5.18 37.2475 5.245 37.3125 ;
        RECT  5.18 37.305 5.245 37.37 ;
        RECT  5.18 37.28 5.245 37.37 ;
        RECT  5.2125 37.2475 5.51 37.3125 ;
        RECT  5.51 37.2475 5.645 37.3125 ;
        RECT  6.215 37.2475 6.28 37.3125 ;
        RECT  6.215 37.305 6.28 37.37 ;
        RECT  5.9975 37.2475 6.2475 37.3125 ;
        RECT  6.215 37.28 6.28 37.3375 ;
        RECT  6.2475 37.305 6.495 37.37 ;
        RECT  4.665 38.47 5.015 38.535 ;
        RECT  5.18 38.5275 5.245 38.5925 ;
        RECT  5.18 38.47 5.245 38.535 ;
        RECT  5.18 38.535 5.245 38.56 ;
        RECT  5.2125 38.5275 5.51 38.5925 ;
        RECT  5.51 38.5275 5.645 38.5925 ;
        RECT  6.215 38.5275 6.28 38.5925 ;
        RECT  6.215 38.47 6.28 38.535 ;
        RECT  5.9975 38.5275 6.2475 38.5925 ;
        RECT  6.215 38.5025 6.28 38.56 ;
        RECT  6.2475 38.47 6.495 38.535 ;
        RECT  4.665 39.995 5.015 40.06 ;
        RECT  5.18 39.9375 5.245 40.0025 ;
        RECT  5.18 39.995 5.245 40.06 ;
        RECT  5.18 39.97 5.245 40.06 ;
        RECT  5.2125 39.9375 5.51 40.0025 ;
        RECT  5.51 39.9375 5.645 40.0025 ;
        RECT  6.215 39.9375 6.28 40.0025 ;
        RECT  6.215 39.995 6.28 40.06 ;
        RECT  5.9975 39.9375 6.2475 40.0025 ;
        RECT  6.215 39.97 6.28 40.0275 ;
        RECT  6.2475 39.995 6.495 40.06 ;
        RECT  6.66 25.02 6.725 25.085 ;
        RECT  4.435 24.0825 4.805 24.1475 ;
        RECT  6.66 19.64 6.725 19.705 ;
        RECT  4.435 29.4625 4.805 29.5275 ;
        RECT  6.66 22.33 6.725 22.395 ;
        RECT  4.435 21.3925 4.805 21.4575 ;
        RECT  4.435 26.7725 4.805 26.8375 ;
        RECT  4.435 30.1725 4.805 30.2375 ;
        RECT  6.66 39.995 6.725 40.06 ;
        RECT  4.435 32.8625 4.805 32.9275 ;
        RECT  6.66 30.4 6.725 30.465 ;
        RECT  4.435 38.2425 4.805 38.3075 ;
        RECT  4.435 35.5525 4.805 35.6175 ;
        RECT  6.66 27.71 6.725 27.775 ;
        RECT  6.66 37.305 6.725 37.37 ;
        RECT  6.66 34.615 6.725 34.68 ;
        RECT  6.66 23.855 6.725 23.92 ;
        RECT  4.435 22.1025 4.805 22.1675 ;
        RECT  6.66 26.545 6.725 26.61 ;
        RECT  6.66 21.165 6.725 21.23 ;
        RECT  4.435 19.4125 4.805 19.4775 ;
        RECT  4.435 24.7925 4.805 24.8575 ;
        RECT  4.435 27.4825 4.805 27.5475 ;
        RECT  4.435 32.1525 4.805 32.2175 ;
        RECT  4.435 34.8425 4.805 34.9075 ;
        RECT  6.66 38.47 6.725 38.535 ;
        RECT  4.435 40.2225 4.805 40.2875 ;
        RECT  6.66 33.09 6.725 33.155 ;
        RECT  6.66 31.925 6.725 31.99 ;
        RECT  4.435 20.4025 4.89 20.4675 ;
        RECT  4.435 23.0925 4.89 23.1575 ;
        RECT  4.435 25.7825 4.89 25.8475 ;
        RECT  4.435 28.4725 4.89 28.5375 ;
        RECT  4.435 31.1625 4.89 31.2275 ;
        RECT  4.435 33.8525 4.89 33.9175 ;
        RECT  4.435 36.5425 4.89 36.6075 ;
        RECT  4.435 39.2325 4.89 39.2975 ;
        RECT  4.435 19.0575 4.89 19.1225 ;
        RECT  4.435 21.7475 4.89 21.8125 ;
        RECT  4.435 24.4375 4.89 24.5025 ;
        RECT  4.435 27.1275 4.89 27.1925 ;
        RECT  4.435 29.8175 4.89 29.8825 ;
        RECT  4.435 32.5075 4.89 32.5725 ;
        RECT  4.435 35.1975 4.89 35.2625 ;
        RECT  4.435 37.8875 4.89 37.9525 ;
        RECT  4.435 40.5775 4.89 40.6425 ;
        RECT  4.435 37.5325 4.805 37.5975 ;
        RECT  6.66 35.78 6.725 35.845 ;
        RECT  6.66 29.235 6.725 29.3 ;
        RECT  5.3175 19.09 5.3825 19.275 ;
        RECT  5.3175 20.205 5.3825 20.435 ;
        RECT  4.9575 19.0575 5.0225 19.2075 ;
        RECT  4.9575 20.0925 5.0225 20.4675 ;
        RECT  5.1475 19.3425 5.2125 20.0925 ;
        RECT  5.015 19.605 5.08 19.74 ;
        RECT  5.18 19.64 5.245 19.705 ;
        RECT  4.89 20.4025 5.45 20.4675 ;
        RECT  4.89 19.0575 5.45 19.1225 ;
        RECT  4.9575 20.0925 5.0225 20.2275 ;
        RECT  5.1475 20.0925 5.2125 20.2275 ;
        RECT  4.9575 20.0925 5.0225 20.2275 ;
        RECT  5.1475 20.0925 5.2125 20.2275 ;
        RECT  4.9575 19.2075 5.0225 19.3425 ;
        RECT  5.1475 19.2075 5.2125 19.3425 ;
        RECT  4.9575 19.2075 5.0225 19.3425 ;
        RECT  5.1475 19.2075 5.2125 19.3425 ;
        RECT  5.3175 19.2075 5.3825 19.3425 ;
        RECT  5.3175 20.1375 5.3825 20.2725 ;
        RECT  5.015 19.605 5.08 19.74 ;
        RECT  6.0675 19.09 6.1325 19.275 ;
        RECT  6.0675 20.205 6.1325 20.435 ;
        RECT  5.5175 19.0575 5.5825 19.2525 ;
        RECT  5.5175 20.0925 5.5825 20.4675 ;
        RECT  5.8975 20.0925 5.9625 20.4675 ;
        RECT  5.51 19.6975 5.645 19.7625 ;
        RECT  5.8625 19.6975 5.9975 19.7625 ;
        RECT  5.7675 19.4825 5.9025 19.5475 ;
        RECT  5.45 20.4025 6.37 20.4675 ;
        RECT  5.45 19.0575 6.37 19.1225 ;
        RECT  5.5175 20.0925 5.5825 20.2275 ;
        RECT  5.7075 20.0925 5.7725 20.2275 ;
        RECT  5.5175 20.0925 5.5825 20.2275 ;
        RECT  5.7075 20.0925 5.7725 20.2275 ;
        RECT  5.7075 20.0925 5.7725 20.2275 ;
        RECT  5.8975 20.0925 5.9625 20.2275 ;
        RECT  5.7075 20.0925 5.7725 20.2275 ;
        RECT  5.8975 20.0925 5.9625 20.2275 ;
        RECT  5.5175 19.2525 5.5825 19.3875 ;
        RECT  5.7075 19.2525 5.7725 19.3875 ;
        RECT  5.5175 19.2525 5.5825 19.3875 ;
        RECT  5.7075 19.2525 5.7725 19.3875 ;
        RECT  5.7075 19.2525 5.7725 19.3875 ;
        RECT  5.8975 19.2525 5.9625 19.3875 ;
        RECT  5.7075 19.2525 5.7725 19.3875 ;
        RECT  5.8975 19.2525 5.9625 19.3875 ;
        RECT  6.0675 19.2075 6.1325 19.3425 ;
        RECT  6.0675 20.1375 6.1325 20.2725 ;
        RECT  5.7675 19.4825 5.9025 19.5475 ;
        RECT  5.51 19.6975 5.645 19.7625 ;
        RECT  5.7075 20.0925 5.7725 20.2275 ;
        RECT  5.8975 19.2525 5.9625 19.3875 ;
        RECT  5.8625 19.6975 5.9975 19.7625 ;
        RECT  6.7975 19.09 6.8625 19.275 ;
        RECT  6.7975 20.205 6.8625 20.435 ;
        RECT  6.4375 19.0575 6.5025 19.2075 ;
        RECT  6.4375 20.0925 6.5025 20.4675 ;
        RECT  6.6275 19.3425 6.6925 20.0925 ;
        RECT  6.495 19.605 6.56 19.74 ;
        RECT  6.66 19.64 6.725 19.705 ;
        RECT  6.37 20.4025 6.93 20.4675 ;
        RECT  6.37 19.0575 6.93 19.1225 ;
        RECT  6.4375 20.0925 6.5025 20.2275 ;
        RECT  6.6275 20.0925 6.6925 20.2275 ;
        RECT  6.4375 20.0925 6.5025 20.2275 ;
        RECT  6.6275 20.0925 6.6925 20.2275 ;
        RECT  6.4375 19.2075 6.5025 19.3425 ;
        RECT  6.6275 19.2075 6.6925 19.3425 ;
        RECT  6.4375 19.2075 6.5025 19.3425 ;
        RECT  6.6275 19.2075 6.6925 19.3425 ;
        RECT  6.7975 19.2075 6.8625 19.3425 ;
        RECT  6.7975 20.1375 6.8625 20.2725 ;
        RECT  6.495 19.605 6.56 19.74 ;
        RECT  4.6325 19.605 4.6975 19.74 ;
        RECT  4.7725 19.3775 4.8375 19.5125 ;
        RECT  5.6325 19.4825 5.7675 19.5475 ;
        RECT  5.3175 21.595 5.3825 21.78 ;
        RECT  5.3175 20.435 5.3825 20.665 ;
        RECT  4.9575 21.6625 5.0225 21.8125 ;
        RECT  4.9575 20.4025 5.0225 20.7775 ;
        RECT  5.1475 20.7775 5.2125 21.5275 ;
        RECT  5.015 21.13 5.08 21.265 ;
        RECT  5.18 21.165 5.245 21.23 ;
        RECT  4.89 20.4025 5.45 20.4675 ;
        RECT  4.89 21.7475 5.45 21.8125 ;
        RECT  4.9575 20.9125 5.0225 21.0475 ;
        RECT  5.1475 20.9125 5.2125 21.0475 ;
        RECT  4.9575 20.9125 5.0225 21.0475 ;
        RECT  5.1475 20.9125 5.2125 21.0475 ;
        RECT  4.9575 21.6175 5.0225 21.7525 ;
        RECT  5.1475 21.6175 5.2125 21.7525 ;
        RECT  4.9575 21.6175 5.0225 21.7525 ;
        RECT  5.1475 21.6175 5.2125 21.7525 ;
        RECT  5.3175 21.6625 5.3825 21.7975 ;
        RECT  5.3175 20.7325 5.3825 20.8675 ;
        RECT  5.015 21.265 5.08 21.4 ;
        RECT  6.0675 21.595 6.1325 21.78 ;
        RECT  6.0675 20.435 6.1325 20.665 ;
        RECT  5.5175 21.6175 5.5825 21.8125 ;
        RECT  5.5175 20.4025 5.5825 20.7775 ;
        RECT  5.8975 20.4025 5.9625 20.7775 ;
        RECT  5.51 21.1075 5.645 21.1725 ;
        RECT  5.8625 21.1075 5.9975 21.1725 ;
        RECT  5.7675 21.3225 5.9025 21.3875 ;
        RECT  5.45 20.4025 6.37 20.4675 ;
        RECT  5.45 21.7475 6.37 21.8125 ;
        RECT  5.5175 20.9125 5.5825 21.0475 ;
        RECT  5.7075 20.9125 5.7725 21.0475 ;
        RECT  5.5175 20.9125 5.5825 21.0475 ;
        RECT  5.7075 20.9125 5.7725 21.0475 ;
        RECT  5.7075 20.9125 5.7725 21.0475 ;
        RECT  5.8975 20.9125 5.9625 21.0475 ;
        RECT  5.7075 20.9125 5.7725 21.0475 ;
        RECT  5.8975 20.9125 5.9625 21.0475 ;
        RECT  5.5175 21.6625 5.5825 21.7975 ;
        RECT  5.7075 21.6625 5.7725 21.7975 ;
        RECT  5.5175 21.6625 5.5825 21.7975 ;
        RECT  5.7075 21.6625 5.7725 21.7975 ;
        RECT  5.7075 21.6625 5.7725 21.7975 ;
        RECT  5.8975 21.6625 5.9625 21.7975 ;
        RECT  5.7075 21.6625 5.7725 21.7975 ;
        RECT  5.8975 21.6625 5.9625 21.7975 ;
        RECT  6.0675 21.6625 6.1325 21.7975 ;
        RECT  6.0675 20.7325 6.1325 20.8675 ;
        RECT  5.7675 21.3975 5.9025 21.4625 ;
        RECT  5.51 21.1825 5.645 21.2475 ;
        RECT  5.7075 20.7775 5.7725 20.9125 ;
        RECT  5.8975 21.6175 5.9625 21.7525 ;
        RECT  5.8625 21.1775 5.9975 21.2425 ;
        RECT  6.7975 21.595 6.8625 21.78 ;
        RECT  6.7975 20.435 6.8625 20.665 ;
        RECT  6.4375 21.6625 6.5025 21.8125 ;
        RECT  6.4375 20.4025 6.5025 20.7775 ;
        RECT  6.6275 20.7775 6.6925 21.5275 ;
        RECT  6.495 21.13 6.56 21.265 ;
        RECT  6.66 21.165 6.725 21.23 ;
        RECT  6.37 20.4025 6.93 20.4675 ;
        RECT  6.37 21.7475 6.93 21.8125 ;
        RECT  6.4375 20.9125 6.5025 21.0475 ;
        RECT  6.6275 20.9125 6.6925 21.0475 ;
        RECT  6.4375 20.9125 6.5025 21.0475 ;
        RECT  6.6275 20.9125 6.6925 21.0475 ;
        RECT  6.4375 21.6175 6.5025 21.7525 ;
        RECT  6.6275 21.6175 6.6925 21.7525 ;
        RECT  6.4375 21.6175 6.5025 21.7525 ;
        RECT  6.6275 21.6175 6.6925 21.7525 ;
        RECT  6.7975 21.6625 6.8625 21.7975 ;
        RECT  6.7975 20.7325 6.8625 20.8675 ;
        RECT  6.495 21.265 6.56 21.4 ;
        RECT  4.6325 21.13 4.6975 21.265 ;
        RECT  4.7725 21.3575 4.8375 21.4925 ;
        RECT  5.6325 21.3225 5.7675 21.3875 ;
        RECT  5.3175 21.78 5.3825 21.965 ;
        RECT  5.3175 22.895 5.3825 23.125 ;
        RECT  4.9575 21.7475 5.0225 21.8975 ;
        RECT  4.9575 22.7825 5.0225 23.1575 ;
        RECT  5.1475 22.0325 5.2125 22.7825 ;
        RECT  5.015 22.295 5.08 22.43 ;
        RECT  5.18 22.33 5.245 22.395 ;
        RECT  4.89 23.0925 5.45 23.1575 ;
        RECT  4.89 21.7475 5.45 21.8125 ;
        RECT  4.9575 22.7825 5.0225 22.9175 ;
        RECT  5.1475 22.7825 5.2125 22.9175 ;
        RECT  4.9575 22.7825 5.0225 22.9175 ;
        RECT  5.1475 22.7825 5.2125 22.9175 ;
        RECT  4.9575 21.8975 5.0225 22.0325 ;
        RECT  5.1475 21.8975 5.2125 22.0325 ;
        RECT  4.9575 21.8975 5.0225 22.0325 ;
        RECT  5.1475 21.8975 5.2125 22.0325 ;
        RECT  5.3175 21.8975 5.3825 22.0325 ;
        RECT  5.3175 22.8275 5.3825 22.9625 ;
        RECT  5.015 22.295 5.08 22.43 ;
        RECT  6.0675 21.78 6.1325 21.965 ;
        RECT  6.0675 22.895 6.1325 23.125 ;
        RECT  5.5175 21.7475 5.5825 21.9425 ;
        RECT  5.5175 22.7825 5.5825 23.1575 ;
        RECT  5.8975 22.7825 5.9625 23.1575 ;
        RECT  5.51 22.3875 5.645 22.4525 ;
        RECT  5.8625 22.3875 5.9975 22.4525 ;
        RECT  5.7675 22.1725 5.9025 22.2375 ;
        RECT  5.45 23.0925 6.37 23.1575 ;
        RECT  5.45 21.7475 6.37 21.8125 ;
        RECT  5.5175 22.7825 5.5825 22.9175 ;
        RECT  5.7075 22.7825 5.7725 22.9175 ;
        RECT  5.5175 22.7825 5.5825 22.9175 ;
        RECT  5.7075 22.7825 5.7725 22.9175 ;
        RECT  5.7075 22.7825 5.7725 22.9175 ;
        RECT  5.8975 22.7825 5.9625 22.9175 ;
        RECT  5.7075 22.7825 5.7725 22.9175 ;
        RECT  5.8975 22.7825 5.9625 22.9175 ;
        RECT  5.5175 21.9425 5.5825 22.0775 ;
        RECT  5.7075 21.9425 5.7725 22.0775 ;
        RECT  5.5175 21.9425 5.5825 22.0775 ;
        RECT  5.7075 21.9425 5.7725 22.0775 ;
        RECT  5.7075 21.9425 5.7725 22.0775 ;
        RECT  5.8975 21.9425 5.9625 22.0775 ;
        RECT  5.7075 21.9425 5.7725 22.0775 ;
        RECT  5.8975 21.9425 5.9625 22.0775 ;
        RECT  6.0675 21.8975 6.1325 22.0325 ;
        RECT  6.0675 22.8275 6.1325 22.9625 ;
        RECT  5.7675 22.1725 5.9025 22.2375 ;
        RECT  5.51 22.3875 5.645 22.4525 ;
        RECT  5.7075 22.7825 5.7725 22.9175 ;
        RECT  5.8975 21.9425 5.9625 22.0775 ;
        RECT  5.8625 22.3875 5.9975 22.4525 ;
        RECT  6.7975 21.78 6.8625 21.965 ;
        RECT  6.7975 22.895 6.8625 23.125 ;
        RECT  6.4375 21.7475 6.5025 21.8975 ;
        RECT  6.4375 22.7825 6.5025 23.1575 ;
        RECT  6.6275 22.0325 6.6925 22.7825 ;
        RECT  6.495 22.295 6.56 22.43 ;
        RECT  6.66 22.33 6.725 22.395 ;
        RECT  6.37 23.0925 6.93 23.1575 ;
        RECT  6.37 21.7475 6.93 21.8125 ;
        RECT  6.4375 22.7825 6.5025 22.9175 ;
        RECT  6.6275 22.7825 6.6925 22.9175 ;
        RECT  6.4375 22.7825 6.5025 22.9175 ;
        RECT  6.6275 22.7825 6.6925 22.9175 ;
        RECT  6.4375 21.8975 6.5025 22.0325 ;
        RECT  6.6275 21.8975 6.6925 22.0325 ;
        RECT  6.4375 21.8975 6.5025 22.0325 ;
        RECT  6.6275 21.8975 6.6925 22.0325 ;
        RECT  6.7975 21.8975 6.8625 22.0325 ;
        RECT  6.7975 22.8275 6.8625 22.9625 ;
        RECT  6.495 22.295 6.56 22.43 ;
        RECT  4.6325 22.295 4.6975 22.43 ;
        RECT  4.7725 22.0675 4.8375 22.2025 ;
        RECT  5.6325 22.1725 5.7675 22.2375 ;
        RECT  5.3175 24.285 5.3825 24.47 ;
        RECT  5.3175 23.125 5.3825 23.355 ;
        RECT  4.9575 24.3525 5.0225 24.5025 ;
        RECT  4.9575 23.0925 5.0225 23.4675 ;
        RECT  5.1475 23.4675 5.2125 24.2175 ;
        RECT  5.015 23.82 5.08 23.955 ;
        RECT  5.18 23.855 5.245 23.92 ;
        RECT  4.89 23.0925 5.45 23.1575 ;
        RECT  4.89 24.4375 5.45 24.5025 ;
        RECT  4.9575 23.6025 5.0225 23.7375 ;
        RECT  5.1475 23.6025 5.2125 23.7375 ;
        RECT  4.9575 23.6025 5.0225 23.7375 ;
        RECT  5.1475 23.6025 5.2125 23.7375 ;
        RECT  4.9575 24.3075 5.0225 24.4425 ;
        RECT  5.1475 24.3075 5.2125 24.4425 ;
        RECT  4.9575 24.3075 5.0225 24.4425 ;
        RECT  5.1475 24.3075 5.2125 24.4425 ;
        RECT  5.3175 24.3525 5.3825 24.4875 ;
        RECT  5.3175 23.4225 5.3825 23.5575 ;
        RECT  5.015 23.955 5.08 24.09 ;
        RECT  6.0675 24.285 6.1325 24.47 ;
        RECT  6.0675 23.125 6.1325 23.355 ;
        RECT  5.5175 24.3075 5.5825 24.5025 ;
        RECT  5.5175 23.0925 5.5825 23.4675 ;
        RECT  5.8975 23.0925 5.9625 23.4675 ;
        RECT  5.51 23.7975 5.645 23.8625 ;
        RECT  5.8625 23.7975 5.9975 23.8625 ;
        RECT  5.7675 24.0125 5.9025 24.0775 ;
        RECT  5.45 23.0925 6.37 23.1575 ;
        RECT  5.45 24.4375 6.37 24.5025 ;
        RECT  5.5175 23.6025 5.5825 23.7375 ;
        RECT  5.7075 23.6025 5.7725 23.7375 ;
        RECT  5.5175 23.6025 5.5825 23.7375 ;
        RECT  5.7075 23.6025 5.7725 23.7375 ;
        RECT  5.7075 23.6025 5.7725 23.7375 ;
        RECT  5.8975 23.6025 5.9625 23.7375 ;
        RECT  5.7075 23.6025 5.7725 23.7375 ;
        RECT  5.8975 23.6025 5.9625 23.7375 ;
        RECT  5.5175 24.3525 5.5825 24.4875 ;
        RECT  5.7075 24.3525 5.7725 24.4875 ;
        RECT  5.5175 24.3525 5.5825 24.4875 ;
        RECT  5.7075 24.3525 5.7725 24.4875 ;
        RECT  5.7075 24.3525 5.7725 24.4875 ;
        RECT  5.8975 24.3525 5.9625 24.4875 ;
        RECT  5.7075 24.3525 5.7725 24.4875 ;
        RECT  5.8975 24.3525 5.9625 24.4875 ;
        RECT  6.0675 24.3525 6.1325 24.4875 ;
        RECT  6.0675 23.4225 6.1325 23.5575 ;
        RECT  5.7675 24.0875 5.9025 24.1525 ;
        RECT  5.51 23.8725 5.645 23.9375 ;
        RECT  5.7075 23.4675 5.7725 23.6025 ;
        RECT  5.8975 24.3075 5.9625 24.4425 ;
        RECT  5.8625 23.8675 5.9975 23.9325 ;
        RECT  6.7975 24.285 6.8625 24.47 ;
        RECT  6.7975 23.125 6.8625 23.355 ;
        RECT  6.4375 24.3525 6.5025 24.5025 ;
        RECT  6.4375 23.0925 6.5025 23.4675 ;
        RECT  6.6275 23.4675 6.6925 24.2175 ;
        RECT  6.495 23.82 6.56 23.955 ;
        RECT  6.66 23.855 6.725 23.92 ;
        RECT  6.37 23.0925 6.93 23.1575 ;
        RECT  6.37 24.4375 6.93 24.5025 ;
        RECT  6.4375 23.6025 6.5025 23.7375 ;
        RECT  6.6275 23.6025 6.6925 23.7375 ;
        RECT  6.4375 23.6025 6.5025 23.7375 ;
        RECT  6.6275 23.6025 6.6925 23.7375 ;
        RECT  6.4375 24.3075 6.5025 24.4425 ;
        RECT  6.6275 24.3075 6.6925 24.4425 ;
        RECT  6.4375 24.3075 6.5025 24.4425 ;
        RECT  6.6275 24.3075 6.6925 24.4425 ;
        RECT  6.7975 24.3525 6.8625 24.4875 ;
        RECT  6.7975 23.4225 6.8625 23.5575 ;
        RECT  6.495 23.955 6.56 24.09 ;
        RECT  4.6325 23.82 4.6975 23.955 ;
        RECT  4.7725 24.0475 4.8375 24.1825 ;
        RECT  5.6325 24.0125 5.7675 24.0775 ;
        RECT  5.3175 24.47 5.3825 24.655 ;
        RECT  5.3175 25.585 5.3825 25.815 ;
        RECT  4.9575 24.4375 5.0225 24.5875 ;
        RECT  4.9575 25.4725 5.0225 25.8475 ;
        RECT  5.1475 24.7225 5.2125 25.4725 ;
        RECT  5.015 24.985 5.08 25.12 ;
        RECT  5.18 25.02 5.245 25.085 ;
        RECT  4.89 25.7825 5.45 25.8475 ;
        RECT  4.89 24.4375 5.45 24.5025 ;
        RECT  4.9575 25.4725 5.0225 25.6075 ;
        RECT  5.1475 25.4725 5.2125 25.6075 ;
        RECT  4.9575 25.4725 5.0225 25.6075 ;
        RECT  5.1475 25.4725 5.2125 25.6075 ;
        RECT  4.9575 24.5875 5.0225 24.7225 ;
        RECT  5.1475 24.5875 5.2125 24.7225 ;
        RECT  4.9575 24.5875 5.0225 24.7225 ;
        RECT  5.1475 24.5875 5.2125 24.7225 ;
        RECT  5.3175 24.5875 5.3825 24.7225 ;
        RECT  5.3175 25.5175 5.3825 25.6525 ;
        RECT  5.015 24.985 5.08 25.12 ;
        RECT  6.0675 24.47 6.1325 24.655 ;
        RECT  6.0675 25.585 6.1325 25.815 ;
        RECT  5.5175 24.4375 5.5825 24.6325 ;
        RECT  5.5175 25.4725 5.5825 25.8475 ;
        RECT  5.8975 25.4725 5.9625 25.8475 ;
        RECT  5.51 25.0775 5.645 25.1425 ;
        RECT  5.8625 25.0775 5.9975 25.1425 ;
        RECT  5.7675 24.8625 5.9025 24.9275 ;
        RECT  5.45 25.7825 6.37 25.8475 ;
        RECT  5.45 24.4375 6.37 24.5025 ;
        RECT  5.5175 25.4725 5.5825 25.6075 ;
        RECT  5.7075 25.4725 5.7725 25.6075 ;
        RECT  5.5175 25.4725 5.5825 25.6075 ;
        RECT  5.7075 25.4725 5.7725 25.6075 ;
        RECT  5.7075 25.4725 5.7725 25.6075 ;
        RECT  5.8975 25.4725 5.9625 25.6075 ;
        RECT  5.7075 25.4725 5.7725 25.6075 ;
        RECT  5.8975 25.4725 5.9625 25.6075 ;
        RECT  5.5175 24.6325 5.5825 24.7675 ;
        RECT  5.7075 24.6325 5.7725 24.7675 ;
        RECT  5.5175 24.6325 5.5825 24.7675 ;
        RECT  5.7075 24.6325 5.7725 24.7675 ;
        RECT  5.7075 24.6325 5.7725 24.7675 ;
        RECT  5.8975 24.6325 5.9625 24.7675 ;
        RECT  5.7075 24.6325 5.7725 24.7675 ;
        RECT  5.8975 24.6325 5.9625 24.7675 ;
        RECT  6.0675 24.5875 6.1325 24.7225 ;
        RECT  6.0675 25.5175 6.1325 25.6525 ;
        RECT  5.7675 24.8625 5.9025 24.9275 ;
        RECT  5.51 25.0775 5.645 25.1425 ;
        RECT  5.7075 25.4725 5.7725 25.6075 ;
        RECT  5.8975 24.6325 5.9625 24.7675 ;
        RECT  5.8625 25.0775 5.9975 25.1425 ;
        RECT  6.7975 24.47 6.8625 24.655 ;
        RECT  6.7975 25.585 6.8625 25.815 ;
        RECT  6.4375 24.4375 6.5025 24.5875 ;
        RECT  6.4375 25.4725 6.5025 25.8475 ;
        RECT  6.6275 24.7225 6.6925 25.4725 ;
        RECT  6.495 24.985 6.56 25.12 ;
        RECT  6.66 25.02 6.725 25.085 ;
        RECT  6.37 25.7825 6.93 25.8475 ;
        RECT  6.37 24.4375 6.93 24.5025 ;
        RECT  6.4375 25.4725 6.5025 25.6075 ;
        RECT  6.6275 25.4725 6.6925 25.6075 ;
        RECT  6.4375 25.4725 6.5025 25.6075 ;
        RECT  6.6275 25.4725 6.6925 25.6075 ;
        RECT  6.4375 24.5875 6.5025 24.7225 ;
        RECT  6.6275 24.5875 6.6925 24.7225 ;
        RECT  6.4375 24.5875 6.5025 24.7225 ;
        RECT  6.6275 24.5875 6.6925 24.7225 ;
        RECT  6.7975 24.5875 6.8625 24.7225 ;
        RECT  6.7975 25.5175 6.8625 25.6525 ;
        RECT  6.495 24.985 6.56 25.12 ;
        RECT  4.6325 24.985 4.6975 25.12 ;
        RECT  4.7725 24.7575 4.8375 24.8925 ;
        RECT  5.6325 24.8625 5.7675 24.9275 ;
        RECT  5.3175 26.975 5.3825 27.16 ;
        RECT  5.3175 25.815 5.3825 26.045 ;
        RECT  4.9575 27.0425 5.0225 27.1925 ;
        RECT  4.9575 25.7825 5.0225 26.1575 ;
        RECT  5.1475 26.1575 5.2125 26.9075 ;
        RECT  5.015 26.51 5.08 26.645 ;
        RECT  5.18 26.545 5.245 26.61 ;
        RECT  4.89 25.7825 5.45 25.8475 ;
        RECT  4.89 27.1275 5.45 27.1925 ;
        RECT  4.9575 26.2925 5.0225 26.4275 ;
        RECT  5.1475 26.2925 5.2125 26.4275 ;
        RECT  4.9575 26.2925 5.0225 26.4275 ;
        RECT  5.1475 26.2925 5.2125 26.4275 ;
        RECT  4.9575 26.9975 5.0225 27.1325 ;
        RECT  5.1475 26.9975 5.2125 27.1325 ;
        RECT  4.9575 26.9975 5.0225 27.1325 ;
        RECT  5.1475 26.9975 5.2125 27.1325 ;
        RECT  5.3175 27.0425 5.3825 27.1775 ;
        RECT  5.3175 26.1125 5.3825 26.2475 ;
        RECT  5.015 26.645 5.08 26.78 ;
        RECT  6.0675 26.975 6.1325 27.16 ;
        RECT  6.0675 25.815 6.1325 26.045 ;
        RECT  5.5175 26.9975 5.5825 27.1925 ;
        RECT  5.5175 25.7825 5.5825 26.1575 ;
        RECT  5.8975 25.7825 5.9625 26.1575 ;
        RECT  5.51 26.4875 5.645 26.5525 ;
        RECT  5.8625 26.4875 5.9975 26.5525 ;
        RECT  5.7675 26.7025 5.9025 26.7675 ;
        RECT  5.45 25.7825 6.37 25.8475 ;
        RECT  5.45 27.1275 6.37 27.1925 ;
        RECT  5.5175 26.2925 5.5825 26.4275 ;
        RECT  5.7075 26.2925 5.7725 26.4275 ;
        RECT  5.5175 26.2925 5.5825 26.4275 ;
        RECT  5.7075 26.2925 5.7725 26.4275 ;
        RECT  5.7075 26.2925 5.7725 26.4275 ;
        RECT  5.8975 26.2925 5.9625 26.4275 ;
        RECT  5.7075 26.2925 5.7725 26.4275 ;
        RECT  5.8975 26.2925 5.9625 26.4275 ;
        RECT  5.5175 27.0425 5.5825 27.1775 ;
        RECT  5.7075 27.0425 5.7725 27.1775 ;
        RECT  5.5175 27.0425 5.5825 27.1775 ;
        RECT  5.7075 27.0425 5.7725 27.1775 ;
        RECT  5.7075 27.0425 5.7725 27.1775 ;
        RECT  5.8975 27.0425 5.9625 27.1775 ;
        RECT  5.7075 27.0425 5.7725 27.1775 ;
        RECT  5.8975 27.0425 5.9625 27.1775 ;
        RECT  6.0675 27.0425 6.1325 27.1775 ;
        RECT  6.0675 26.1125 6.1325 26.2475 ;
        RECT  5.7675 26.7775 5.9025 26.8425 ;
        RECT  5.51 26.5625 5.645 26.6275 ;
        RECT  5.7075 26.1575 5.7725 26.2925 ;
        RECT  5.8975 26.9975 5.9625 27.1325 ;
        RECT  5.8625 26.5575 5.9975 26.6225 ;
        RECT  6.7975 26.975 6.8625 27.16 ;
        RECT  6.7975 25.815 6.8625 26.045 ;
        RECT  6.4375 27.0425 6.5025 27.1925 ;
        RECT  6.4375 25.7825 6.5025 26.1575 ;
        RECT  6.6275 26.1575 6.6925 26.9075 ;
        RECT  6.495 26.51 6.56 26.645 ;
        RECT  6.66 26.545 6.725 26.61 ;
        RECT  6.37 25.7825 6.93 25.8475 ;
        RECT  6.37 27.1275 6.93 27.1925 ;
        RECT  6.4375 26.2925 6.5025 26.4275 ;
        RECT  6.6275 26.2925 6.6925 26.4275 ;
        RECT  6.4375 26.2925 6.5025 26.4275 ;
        RECT  6.6275 26.2925 6.6925 26.4275 ;
        RECT  6.4375 26.9975 6.5025 27.1325 ;
        RECT  6.6275 26.9975 6.6925 27.1325 ;
        RECT  6.4375 26.9975 6.5025 27.1325 ;
        RECT  6.6275 26.9975 6.6925 27.1325 ;
        RECT  6.7975 27.0425 6.8625 27.1775 ;
        RECT  6.7975 26.1125 6.8625 26.2475 ;
        RECT  6.495 26.645 6.56 26.78 ;
        RECT  4.6325 26.51 4.6975 26.645 ;
        RECT  4.7725 26.7375 4.8375 26.8725 ;
        RECT  5.6325 26.7025 5.7675 26.7675 ;
        RECT  5.3175 27.16 5.3825 27.345 ;
        RECT  5.3175 28.275 5.3825 28.505 ;
        RECT  4.9575 27.1275 5.0225 27.2775 ;
        RECT  4.9575 28.1625 5.0225 28.5375 ;
        RECT  5.1475 27.4125 5.2125 28.1625 ;
        RECT  5.015 27.675 5.08 27.81 ;
        RECT  5.18 27.71 5.245 27.775 ;
        RECT  4.89 28.4725 5.45 28.5375 ;
        RECT  4.89 27.1275 5.45 27.1925 ;
        RECT  4.9575 28.1625 5.0225 28.2975 ;
        RECT  5.1475 28.1625 5.2125 28.2975 ;
        RECT  4.9575 28.1625 5.0225 28.2975 ;
        RECT  5.1475 28.1625 5.2125 28.2975 ;
        RECT  4.9575 27.2775 5.0225 27.4125 ;
        RECT  5.1475 27.2775 5.2125 27.4125 ;
        RECT  4.9575 27.2775 5.0225 27.4125 ;
        RECT  5.1475 27.2775 5.2125 27.4125 ;
        RECT  5.3175 27.2775 5.3825 27.4125 ;
        RECT  5.3175 28.2075 5.3825 28.3425 ;
        RECT  5.015 27.675 5.08 27.81 ;
        RECT  6.0675 27.16 6.1325 27.345 ;
        RECT  6.0675 28.275 6.1325 28.505 ;
        RECT  5.5175 27.1275 5.5825 27.3225 ;
        RECT  5.5175 28.1625 5.5825 28.5375 ;
        RECT  5.8975 28.1625 5.9625 28.5375 ;
        RECT  5.51 27.7675 5.645 27.8325 ;
        RECT  5.8625 27.7675 5.9975 27.8325 ;
        RECT  5.7675 27.5525 5.9025 27.6175 ;
        RECT  5.45 28.4725 6.37 28.5375 ;
        RECT  5.45 27.1275 6.37 27.1925 ;
        RECT  5.5175 28.1625 5.5825 28.2975 ;
        RECT  5.7075 28.1625 5.7725 28.2975 ;
        RECT  5.5175 28.1625 5.5825 28.2975 ;
        RECT  5.7075 28.1625 5.7725 28.2975 ;
        RECT  5.7075 28.1625 5.7725 28.2975 ;
        RECT  5.8975 28.1625 5.9625 28.2975 ;
        RECT  5.7075 28.1625 5.7725 28.2975 ;
        RECT  5.8975 28.1625 5.9625 28.2975 ;
        RECT  5.5175 27.3225 5.5825 27.4575 ;
        RECT  5.7075 27.3225 5.7725 27.4575 ;
        RECT  5.5175 27.3225 5.5825 27.4575 ;
        RECT  5.7075 27.3225 5.7725 27.4575 ;
        RECT  5.7075 27.3225 5.7725 27.4575 ;
        RECT  5.8975 27.3225 5.9625 27.4575 ;
        RECT  5.7075 27.3225 5.7725 27.4575 ;
        RECT  5.8975 27.3225 5.9625 27.4575 ;
        RECT  6.0675 27.2775 6.1325 27.4125 ;
        RECT  6.0675 28.2075 6.1325 28.3425 ;
        RECT  5.7675 27.5525 5.9025 27.6175 ;
        RECT  5.51 27.7675 5.645 27.8325 ;
        RECT  5.7075 28.1625 5.7725 28.2975 ;
        RECT  5.8975 27.3225 5.9625 27.4575 ;
        RECT  5.8625 27.7675 5.9975 27.8325 ;
        RECT  6.7975 27.16 6.8625 27.345 ;
        RECT  6.7975 28.275 6.8625 28.505 ;
        RECT  6.4375 27.1275 6.5025 27.2775 ;
        RECT  6.4375 28.1625 6.5025 28.5375 ;
        RECT  6.6275 27.4125 6.6925 28.1625 ;
        RECT  6.495 27.675 6.56 27.81 ;
        RECT  6.66 27.71 6.725 27.775 ;
        RECT  6.37 28.4725 6.93 28.5375 ;
        RECT  6.37 27.1275 6.93 27.1925 ;
        RECT  6.4375 28.1625 6.5025 28.2975 ;
        RECT  6.6275 28.1625 6.6925 28.2975 ;
        RECT  6.4375 28.1625 6.5025 28.2975 ;
        RECT  6.6275 28.1625 6.6925 28.2975 ;
        RECT  6.4375 27.2775 6.5025 27.4125 ;
        RECT  6.6275 27.2775 6.6925 27.4125 ;
        RECT  6.4375 27.2775 6.5025 27.4125 ;
        RECT  6.6275 27.2775 6.6925 27.4125 ;
        RECT  6.7975 27.2775 6.8625 27.4125 ;
        RECT  6.7975 28.2075 6.8625 28.3425 ;
        RECT  6.495 27.675 6.56 27.81 ;
        RECT  4.6325 27.675 4.6975 27.81 ;
        RECT  4.7725 27.4475 4.8375 27.5825 ;
        RECT  5.6325 27.5525 5.7675 27.6175 ;
        RECT  5.3175 29.665 5.3825 29.85 ;
        RECT  5.3175 28.505 5.3825 28.735 ;
        RECT  4.9575 29.7325 5.0225 29.8825 ;
        RECT  4.9575 28.4725 5.0225 28.8475 ;
        RECT  5.1475 28.8475 5.2125 29.5975 ;
        RECT  5.015 29.2 5.08 29.335 ;
        RECT  5.18 29.235 5.245 29.3 ;
        RECT  4.89 28.4725 5.45 28.5375 ;
        RECT  4.89 29.8175 5.45 29.8825 ;
        RECT  4.9575 28.9825 5.0225 29.1175 ;
        RECT  5.1475 28.9825 5.2125 29.1175 ;
        RECT  4.9575 28.9825 5.0225 29.1175 ;
        RECT  5.1475 28.9825 5.2125 29.1175 ;
        RECT  4.9575 29.6875 5.0225 29.8225 ;
        RECT  5.1475 29.6875 5.2125 29.8225 ;
        RECT  4.9575 29.6875 5.0225 29.8225 ;
        RECT  5.1475 29.6875 5.2125 29.8225 ;
        RECT  5.3175 29.7325 5.3825 29.8675 ;
        RECT  5.3175 28.8025 5.3825 28.9375 ;
        RECT  5.015 29.335 5.08 29.47 ;
        RECT  6.0675 29.665 6.1325 29.85 ;
        RECT  6.0675 28.505 6.1325 28.735 ;
        RECT  5.5175 29.6875 5.5825 29.8825 ;
        RECT  5.5175 28.4725 5.5825 28.8475 ;
        RECT  5.8975 28.4725 5.9625 28.8475 ;
        RECT  5.51 29.1775 5.645 29.2425 ;
        RECT  5.8625 29.1775 5.9975 29.2425 ;
        RECT  5.7675 29.3925 5.9025 29.4575 ;
        RECT  5.45 28.4725 6.37 28.5375 ;
        RECT  5.45 29.8175 6.37 29.8825 ;
        RECT  5.5175 28.9825 5.5825 29.1175 ;
        RECT  5.7075 28.9825 5.7725 29.1175 ;
        RECT  5.5175 28.9825 5.5825 29.1175 ;
        RECT  5.7075 28.9825 5.7725 29.1175 ;
        RECT  5.7075 28.9825 5.7725 29.1175 ;
        RECT  5.8975 28.9825 5.9625 29.1175 ;
        RECT  5.7075 28.9825 5.7725 29.1175 ;
        RECT  5.8975 28.9825 5.9625 29.1175 ;
        RECT  5.5175 29.7325 5.5825 29.8675 ;
        RECT  5.7075 29.7325 5.7725 29.8675 ;
        RECT  5.5175 29.7325 5.5825 29.8675 ;
        RECT  5.7075 29.7325 5.7725 29.8675 ;
        RECT  5.7075 29.7325 5.7725 29.8675 ;
        RECT  5.8975 29.7325 5.9625 29.8675 ;
        RECT  5.7075 29.7325 5.7725 29.8675 ;
        RECT  5.8975 29.7325 5.9625 29.8675 ;
        RECT  6.0675 29.7325 6.1325 29.8675 ;
        RECT  6.0675 28.8025 6.1325 28.9375 ;
        RECT  5.7675 29.4675 5.9025 29.5325 ;
        RECT  5.51 29.2525 5.645 29.3175 ;
        RECT  5.7075 28.8475 5.7725 28.9825 ;
        RECT  5.8975 29.6875 5.9625 29.8225 ;
        RECT  5.8625 29.2475 5.9975 29.3125 ;
        RECT  6.7975 29.665 6.8625 29.85 ;
        RECT  6.7975 28.505 6.8625 28.735 ;
        RECT  6.4375 29.7325 6.5025 29.8825 ;
        RECT  6.4375 28.4725 6.5025 28.8475 ;
        RECT  6.6275 28.8475 6.6925 29.5975 ;
        RECT  6.495 29.2 6.56 29.335 ;
        RECT  6.66 29.235 6.725 29.3 ;
        RECT  6.37 28.4725 6.93 28.5375 ;
        RECT  6.37 29.8175 6.93 29.8825 ;
        RECT  6.4375 28.9825 6.5025 29.1175 ;
        RECT  6.6275 28.9825 6.6925 29.1175 ;
        RECT  6.4375 28.9825 6.5025 29.1175 ;
        RECT  6.6275 28.9825 6.6925 29.1175 ;
        RECT  6.4375 29.6875 6.5025 29.8225 ;
        RECT  6.6275 29.6875 6.6925 29.8225 ;
        RECT  6.4375 29.6875 6.5025 29.8225 ;
        RECT  6.6275 29.6875 6.6925 29.8225 ;
        RECT  6.7975 29.7325 6.8625 29.8675 ;
        RECT  6.7975 28.8025 6.8625 28.9375 ;
        RECT  6.495 29.335 6.56 29.47 ;
        RECT  4.6325 29.2 4.6975 29.335 ;
        RECT  4.7725 29.4275 4.8375 29.5625 ;
        RECT  5.6325 29.3925 5.7675 29.4575 ;
        RECT  5.3175 29.85 5.3825 30.035 ;
        RECT  5.3175 30.965 5.3825 31.195 ;
        RECT  4.9575 29.8175 5.0225 29.9675 ;
        RECT  4.9575 30.8525 5.0225 31.2275 ;
        RECT  5.1475 30.1025 5.2125 30.8525 ;
        RECT  5.015 30.365 5.08 30.5 ;
        RECT  5.18 30.4 5.245 30.465 ;
        RECT  4.89 31.1625 5.45 31.2275 ;
        RECT  4.89 29.8175 5.45 29.8825 ;
        RECT  4.9575 30.8525 5.0225 30.9875 ;
        RECT  5.1475 30.8525 5.2125 30.9875 ;
        RECT  4.9575 30.8525 5.0225 30.9875 ;
        RECT  5.1475 30.8525 5.2125 30.9875 ;
        RECT  4.9575 29.9675 5.0225 30.1025 ;
        RECT  5.1475 29.9675 5.2125 30.1025 ;
        RECT  4.9575 29.9675 5.0225 30.1025 ;
        RECT  5.1475 29.9675 5.2125 30.1025 ;
        RECT  5.3175 29.9675 5.3825 30.1025 ;
        RECT  5.3175 30.8975 5.3825 31.0325 ;
        RECT  5.015 30.365 5.08 30.5 ;
        RECT  6.0675 29.85 6.1325 30.035 ;
        RECT  6.0675 30.965 6.1325 31.195 ;
        RECT  5.5175 29.8175 5.5825 30.0125 ;
        RECT  5.5175 30.8525 5.5825 31.2275 ;
        RECT  5.8975 30.8525 5.9625 31.2275 ;
        RECT  5.51 30.4575 5.645 30.5225 ;
        RECT  5.8625 30.4575 5.9975 30.5225 ;
        RECT  5.7675 30.2425 5.9025 30.3075 ;
        RECT  5.45 31.1625 6.37 31.2275 ;
        RECT  5.45 29.8175 6.37 29.8825 ;
        RECT  5.5175 30.8525 5.5825 30.9875 ;
        RECT  5.7075 30.8525 5.7725 30.9875 ;
        RECT  5.5175 30.8525 5.5825 30.9875 ;
        RECT  5.7075 30.8525 5.7725 30.9875 ;
        RECT  5.7075 30.8525 5.7725 30.9875 ;
        RECT  5.8975 30.8525 5.9625 30.9875 ;
        RECT  5.7075 30.8525 5.7725 30.9875 ;
        RECT  5.8975 30.8525 5.9625 30.9875 ;
        RECT  5.5175 30.0125 5.5825 30.1475 ;
        RECT  5.7075 30.0125 5.7725 30.1475 ;
        RECT  5.5175 30.0125 5.5825 30.1475 ;
        RECT  5.7075 30.0125 5.7725 30.1475 ;
        RECT  5.7075 30.0125 5.7725 30.1475 ;
        RECT  5.8975 30.0125 5.9625 30.1475 ;
        RECT  5.7075 30.0125 5.7725 30.1475 ;
        RECT  5.8975 30.0125 5.9625 30.1475 ;
        RECT  6.0675 29.9675 6.1325 30.1025 ;
        RECT  6.0675 30.8975 6.1325 31.0325 ;
        RECT  5.7675 30.2425 5.9025 30.3075 ;
        RECT  5.51 30.4575 5.645 30.5225 ;
        RECT  5.7075 30.8525 5.7725 30.9875 ;
        RECT  5.8975 30.0125 5.9625 30.1475 ;
        RECT  5.8625 30.4575 5.9975 30.5225 ;
        RECT  6.7975 29.85 6.8625 30.035 ;
        RECT  6.7975 30.965 6.8625 31.195 ;
        RECT  6.4375 29.8175 6.5025 29.9675 ;
        RECT  6.4375 30.8525 6.5025 31.2275 ;
        RECT  6.6275 30.1025 6.6925 30.8525 ;
        RECT  6.495 30.365 6.56 30.5 ;
        RECT  6.66 30.4 6.725 30.465 ;
        RECT  6.37 31.1625 6.93 31.2275 ;
        RECT  6.37 29.8175 6.93 29.8825 ;
        RECT  6.4375 30.8525 6.5025 30.9875 ;
        RECT  6.6275 30.8525 6.6925 30.9875 ;
        RECT  6.4375 30.8525 6.5025 30.9875 ;
        RECT  6.6275 30.8525 6.6925 30.9875 ;
        RECT  6.4375 29.9675 6.5025 30.1025 ;
        RECT  6.6275 29.9675 6.6925 30.1025 ;
        RECT  6.4375 29.9675 6.5025 30.1025 ;
        RECT  6.6275 29.9675 6.6925 30.1025 ;
        RECT  6.7975 29.9675 6.8625 30.1025 ;
        RECT  6.7975 30.8975 6.8625 31.0325 ;
        RECT  6.495 30.365 6.56 30.5 ;
        RECT  4.6325 30.365 4.6975 30.5 ;
        RECT  4.7725 30.1375 4.8375 30.2725 ;
        RECT  5.6325 30.2425 5.7675 30.3075 ;
        RECT  5.3175 32.355 5.3825 32.54 ;
        RECT  5.3175 31.195 5.3825 31.425 ;
        RECT  4.9575 32.4225 5.0225 32.5725 ;
        RECT  4.9575 31.1625 5.0225 31.5375 ;
        RECT  5.1475 31.5375 5.2125 32.2875 ;
        RECT  5.015 31.89 5.08 32.025 ;
        RECT  5.18 31.925 5.245 31.99 ;
        RECT  4.89 31.1625 5.45 31.2275 ;
        RECT  4.89 32.5075 5.45 32.5725 ;
        RECT  4.9575 31.6725 5.0225 31.8075 ;
        RECT  5.1475 31.6725 5.2125 31.8075 ;
        RECT  4.9575 31.6725 5.0225 31.8075 ;
        RECT  5.1475 31.6725 5.2125 31.8075 ;
        RECT  4.9575 32.3775 5.0225 32.5125 ;
        RECT  5.1475 32.3775 5.2125 32.5125 ;
        RECT  4.9575 32.3775 5.0225 32.5125 ;
        RECT  5.1475 32.3775 5.2125 32.5125 ;
        RECT  5.3175 32.4225 5.3825 32.5575 ;
        RECT  5.3175 31.4925 5.3825 31.6275 ;
        RECT  5.015 32.025 5.08 32.16 ;
        RECT  6.0675 32.355 6.1325 32.54 ;
        RECT  6.0675 31.195 6.1325 31.425 ;
        RECT  5.5175 32.3775 5.5825 32.5725 ;
        RECT  5.5175 31.1625 5.5825 31.5375 ;
        RECT  5.8975 31.1625 5.9625 31.5375 ;
        RECT  5.51 31.8675 5.645 31.9325 ;
        RECT  5.8625 31.8675 5.9975 31.9325 ;
        RECT  5.7675 32.0825 5.9025 32.1475 ;
        RECT  5.45 31.1625 6.37 31.2275 ;
        RECT  5.45 32.5075 6.37 32.5725 ;
        RECT  5.5175 31.6725 5.5825 31.8075 ;
        RECT  5.7075 31.6725 5.7725 31.8075 ;
        RECT  5.5175 31.6725 5.5825 31.8075 ;
        RECT  5.7075 31.6725 5.7725 31.8075 ;
        RECT  5.7075 31.6725 5.7725 31.8075 ;
        RECT  5.8975 31.6725 5.9625 31.8075 ;
        RECT  5.7075 31.6725 5.7725 31.8075 ;
        RECT  5.8975 31.6725 5.9625 31.8075 ;
        RECT  5.5175 32.4225 5.5825 32.5575 ;
        RECT  5.7075 32.4225 5.7725 32.5575 ;
        RECT  5.5175 32.4225 5.5825 32.5575 ;
        RECT  5.7075 32.4225 5.7725 32.5575 ;
        RECT  5.7075 32.4225 5.7725 32.5575 ;
        RECT  5.8975 32.4225 5.9625 32.5575 ;
        RECT  5.7075 32.4225 5.7725 32.5575 ;
        RECT  5.8975 32.4225 5.9625 32.5575 ;
        RECT  6.0675 32.4225 6.1325 32.5575 ;
        RECT  6.0675 31.4925 6.1325 31.6275 ;
        RECT  5.7675 32.1575 5.9025 32.2225 ;
        RECT  5.51 31.9425 5.645 32.0075 ;
        RECT  5.7075 31.5375 5.7725 31.6725 ;
        RECT  5.8975 32.3775 5.9625 32.5125 ;
        RECT  5.8625 31.9375 5.9975 32.0025 ;
        RECT  6.7975 32.355 6.8625 32.54 ;
        RECT  6.7975 31.195 6.8625 31.425 ;
        RECT  6.4375 32.4225 6.5025 32.5725 ;
        RECT  6.4375 31.1625 6.5025 31.5375 ;
        RECT  6.6275 31.5375 6.6925 32.2875 ;
        RECT  6.495 31.89 6.56 32.025 ;
        RECT  6.66 31.925 6.725 31.99 ;
        RECT  6.37 31.1625 6.93 31.2275 ;
        RECT  6.37 32.5075 6.93 32.5725 ;
        RECT  6.4375 31.6725 6.5025 31.8075 ;
        RECT  6.6275 31.6725 6.6925 31.8075 ;
        RECT  6.4375 31.6725 6.5025 31.8075 ;
        RECT  6.6275 31.6725 6.6925 31.8075 ;
        RECT  6.4375 32.3775 6.5025 32.5125 ;
        RECT  6.6275 32.3775 6.6925 32.5125 ;
        RECT  6.4375 32.3775 6.5025 32.5125 ;
        RECT  6.6275 32.3775 6.6925 32.5125 ;
        RECT  6.7975 32.4225 6.8625 32.5575 ;
        RECT  6.7975 31.4925 6.8625 31.6275 ;
        RECT  6.495 32.025 6.56 32.16 ;
        RECT  4.6325 31.89 4.6975 32.025 ;
        RECT  4.7725 32.1175 4.8375 32.2525 ;
        RECT  5.6325 32.0825 5.7675 32.1475 ;
        RECT  5.3175 32.54 5.3825 32.725 ;
        RECT  5.3175 33.655 5.3825 33.885 ;
        RECT  4.9575 32.5075 5.0225 32.6575 ;
        RECT  4.9575 33.5425 5.0225 33.9175 ;
        RECT  5.1475 32.7925 5.2125 33.5425 ;
        RECT  5.015 33.055 5.08 33.19 ;
        RECT  5.18 33.09 5.245 33.155 ;
        RECT  4.89 33.8525 5.45 33.9175 ;
        RECT  4.89 32.5075 5.45 32.5725 ;
        RECT  4.9575 33.5425 5.0225 33.6775 ;
        RECT  5.1475 33.5425 5.2125 33.6775 ;
        RECT  4.9575 33.5425 5.0225 33.6775 ;
        RECT  5.1475 33.5425 5.2125 33.6775 ;
        RECT  4.9575 32.6575 5.0225 32.7925 ;
        RECT  5.1475 32.6575 5.2125 32.7925 ;
        RECT  4.9575 32.6575 5.0225 32.7925 ;
        RECT  5.1475 32.6575 5.2125 32.7925 ;
        RECT  5.3175 32.6575 5.3825 32.7925 ;
        RECT  5.3175 33.5875 5.3825 33.7225 ;
        RECT  5.015 33.055 5.08 33.19 ;
        RECT  6.0675 32.54 6.1325 32.725 ;
        RECT  6.0675 33.655 6.1325 33.885 ;
        RECT  5.5175 32.5075 5.5825 32.7025 ;
        RECT  5.5175 33.5425 5.5825 33.9175 ;
        RECT  5.8975 33.5425 5.9625 33.9175 ;
        RECT  5.51 33.1475 5.645 33.2125 ;
        RECT  5.8625 33.1475 5.9975 33.2125 ;
        RECT  5.7675 32.9325 5.9025 32.9975 ;
        RECT  5.45 33.8525 6.37 33.9175 ;
        RECT  5.45 32.5075 6.37 32.5725 ;
        RECT  5.5175 33.5425 5.5825 33.6775 ;
        RECT  5.7075 33.5425 5.7725 33.6775 ;
        RECT  5.5175 33.5425 5.5825 33.6775 ;
        RECT  5.7075 33.5425 5.7725 33.6775 ;
        RECT  5.7075 33.5425 5.7725 33.6775 ;
        RECT  5.8975 33.5425 5.9625 33.6775 ;
        RECT  5.7075 33.5425 5.7725 33.6775 ;
        RECT  5.8975 33.5425 5.9625 33.6775 ;
        RECT  5.5175 32.7025 5.5825 32.8375 ;
        RECT  5.7075 32.7025 5.7725 32.8375 ;
        RECT  5.5175 32.7025 5.5825 32.8375 ;
        RECT  5.7075 32.7025 5.7725 32.8375 ;
        RECT  5.7075 32.7025 5.7725 32.8375 ;
        RECT  5.8975 32.7025 5.9625 32.8375 ;
        RECT  5.7075 32.7025 5.7725 32.8375 ;
        RECT  5.8975 32.7025 5.9625 32.8375 ;
        RECT  6.0675 32.6575 6.1325 32.7925 ;
        RECT  6.0675 33.5875 6.1325 33.7225 ;
        RECT  5.7675 32.9325 5.9025 32.9975 ;
        RECT  5.51 33.1475 5.645 33.2125 ;
        RECT  5.7075 33.5425 5.7725 33.6775 ;
        RECT  5.8975 32.7025 5.9625 32.8375 ;
        RECT  5.8625 33.1475 5.9975 33.2125 ;
        RECT  6.7975 32.54 6.8625 32.725 ;
        RECT  6.7975 33.655 6.8625 33.885 ;
        RECT  6.4375 32.5075 6.5025 32.6575 ;
        RECT  6.4375 33.5425 6.5025 33.9175 ;
        RECT  6.6275 32.7925 6.6925 33.5425 ;
        RECT  6.495 33.055 6.56 33.19 ;
        RECT  6.66 33.09 6.725 33.155 ;
        RECT  6.37 33.8525 6.93 33.9175 ;
        RECT  6.37 32.5075 6.93 32.5725 ;
        RECT  6.4375 33.5425 6.5025 33.6775 ;
        RECT  6.6275 33.5425 6.6925 33.6775 ;
        RECT  6.4375 33.5425 6.5025 33.6775 ;
        RECT  6.6275 33.5425 6.6925 33.6775 ;
        RECT  6.4375 32.6575 6.5025 32.7925 ;
        RECT  6.6275 32.6575 6.6925 32.7925 ;
        RECT  6.4375 32.6575 6.5025 32.7925 ;
        RECT  6.6275 32.6575 6.6925 32.7925 ;
        RECT  6.7975 32.6575 6.8625 32.7925 ;
        RECT  6.7975 33.5875 6.8625 33.7225 ;
        RECT  6.495 33.055 6.56 33.19 ;
        RECT  4.6325 33.055 4.6975 33.19 ;
        RECT  4.7725 32.8275 4.8375 32.9625 ;
        RECT  5.6325 32.9325 5.7675 32.9975 ;
        RECT  5.3175 35.045 5.3825 35.23 ;
        RECT  5.3175 33.885 5.3825 34.115 ;
        RECT  4.9575 35.1125 5.0225 35.2625 ;
        RECT  4.9575 33.8525 5.0225 34.2275 ;
        RECT  5.1475 34.2275 5.2125 34.9775 ;
        RECT  5.015 34.58 5.08 34.715 ;
        RECT  5.18 34.615 5.245 34.68 ;
        RECT  4.89 33.8525 5.45 33.9175 ;
        RECT  4.89 35.1975 5.45 35.2625 ;
        RECT  4.9575 34.3625 5.0225 34.4975 ;
        RECT  5.1475 34.3625 5.2125 34.4975 ;
        RECT  4.9575 34.3625 5.0225 34.4975 ;
        RECT  5.1475 34.3625 5.2125 34.4975 ;
        RECT  4.9575 35.0675 5.0225 35.2025 ;
        RECT  5.1475 35.0675 5.2125 35.2025 ;
        RECT  4.9575 35.0675 5.0225 35.2025 ;
        RECT  5.1475 35.0675 5.2125 35.2025 ;
        RECT  5.3175 35.1125 5.3825 35.2475 ;
        RECT  5.3175 34.1825 5.3825 34.3175 ;
        RECT  5.015 34.715 5.08 34.85 ;
        RECT  6.0675 35.045 6.1325 35.23 ;
        RECT  6.0675 33.885 6.1325 34.115 ;
        RECT  5.5175 35.0675 5.5825 35.2625 ;
        RECT  5.5175 33.8525 5.5825 34.2275 ;
        RECT  5.8975 33.8525 5.9625 34.2275 ;
        RECT  5.51 34.5575 5.645 34.6225 ;
        RECT  5.8625 34.5575 5.9975 34.6225 ;
        RECT  5.7675 34.7725 5.9025 34.8375 ;
        RECT  5.45 33.8525 6.37 33.9175 ;
        RECT  5.45 35.1975 6.37 35.2625 ;
        RECT  5.5175 34.3625 5.5825 34.4975 ;
        RECT  5.7075 34.3625 5.7725 34.4975 ;
        RECT  5.5175 34.3625 5.5825 34.4975 ;
        RECT  5.7075 34.3625 5.7725 34.4975 ;
        RECT  5.7075 34.3625 5.7725 34.4975 ;
        RECT  5.8975 34.3625 5.9625 34.4975 ;
        RECT  5.7075 34.3625 5.7725 34.4975 ;
        RECT  5.8975 34.3625 5.9625 34.4975 ;
        RECT  5.5175 35.1125 5.5825 35.2475 ;
        RECT  5.7075 35.1125 5.7725 35.2475 ;
        RECT  5.5175 35.1125 5.5825 35.2475 ;
        RECT  5.7075 35.1125 5.7725 35.2475 ;
        RECT  5.7075 35.1125 5.7725 35.2475 ;
        RECT  5.8975 35.1125 5.9625 35.2475 ;
        RECT  5.7075 35.1125 5.7725 35.2475 ;
        RECT  5.8975 35.1125 5.9625 35.2475 ;
        RECT  6.0675 35.1125 6.1325 35.2475 ;
        RECT  6.0675 34.1825 6.1325 34.3175 ;
        RECT  5.7675 34.8475 5.9025 34.9125 ;
        RECT  5.51 34.6325 5.645 34.6975 ;
        RECT  5.7075 34.2275 5.7725 34.3625 ;
        RECT  5.8975 35.0675 5.9625 35.2025 ;
        RECT  5.8625 34.6275 5.9975 34.6925 ;
        RECT  6.7975 35.045 6.8625 35.23 ;
        RECT  6.7975 33.885 6.8625 34.115 ;
        RECT  6.4375 35.1125 6.5025 35.2625 ;
        RECT  6.4375 33.8525 6.5025 34.2275 ;
        RECT  6.6275 34.2275 6.6925 34.9775 ;
        RECT  6.495 34.58 6.56 34.715 ;
        RECT  6.66 34.615 6.725 34.68 ;
        RECT  6.37 33.8525 6.93 33.9175 ;
        RECT  6.37 35.1975 6.93 35.2625 ;
        RECT  6.4375 34.3625 6.5025 34.4975 ;
        RECT  6.6275 34.3625 6.6925 34.4975 ;
        RECT  6.4375 34.3625 6.5025 34.4975 ;
        RECT  6.6275 34.3625 6.6925 34.4975 ;
        RECT  6.4375 35.0675 6.5025 35.2025 ;
        RECT  6.6275 35.0675 6.6925 35.2025 ;
        RECT  6.4375 35.0675 6.5025 35.2025 ;
        RECT  6.6275 35.0675 6.6925 35.2025 ;
        RECT  6.7975 35.1125 6.8625 35.2475 ;
        RECT  6.7975 34.1825 6.8625 34.3175 ;
        RECT  6.495 34.715 6.56 34.85 ;
        RECT  4.6325 34.58 4.6975 34.715 ;
        RECT  4.7725 34.8075 4.8375 34.9425 ;
        RECT  5.6325 34.7725 5.7675 34.8375 ;
        RECT  5.3175 35.23 5.3825 35.415 ;
        RECT  5.3175 36.345 5.3825 36.575 ;
        RECT  4.9575 35.1975 5.0225 35.3475 ;
        RECT  4.9575 36.2325 5.0225 36.6075 ;
        RECT  5.1475 35.4825 5.2125 36.2325 ;
        RECT  5.015 35.745 5.08 35.88 ;
        RECT  5.18 35.78 5.245 35.845 ;
        RECT  4.89 36.5425 5.45 36.6075 ;
        RECT  4.89 35.1975 5.45 35.2625 ;
        RECT  4.9575 36.2325 5.0225 36.3675 ;
        RECT  5.1475 36.2325 5.2125 36.3675 ;
        RECT  4.9575 36.2325 5.0225 36.3675 ;
        RECT  5.1475 36.2325 5.2125 36.3675 ;
        RECT  4.9575 35.3475 5.0225 35.4825 ;
        RECT  5.1475 35.3475 5.2125 35.4825 ;
        RECT  4.9575 35.3475 5.0225 35.4825 ;
        RECT  5.1475 35.3475 5.2125 35.4825 ;
        RECT  5.3175 35.3475 5.3825 35.4825 ;
        RECT  5.3175 36.2775 5.3825 36.4125 ;
        RECT  5.015 35.745 5.08 35.88 ;
        RECT  6.0675 35.23 6.1325 35.415 ;
        RECT  6.0675 36.345 6.1325 36.575 ;
        RECT  5.5175 35.1975 5.5825 35.3925 ;
        RECT  5.5175 36.2325 5.5825 36.6075 ;
        RECT  5.8975 36.2325 5.9625 36.6075 ;
        RECT  5.51 35.8375 5.645 35.9025 ;
        RECT  5.8625 35.8375 5.9975 35.9025 ;
        RECT  5.7675 35.6225 5.9025 35.6875 ;
        RECT  5.45 36.5425 6.37 36.6075 ;
        RECT  5.45 35.1975 6.37 35.2625 ;
        RECT  5.5175 36.2325 5.5825 36.3675 ;
        RECT  5.7075 36.2325 5.7725 36.3675 ;
        RECT  5.5175 36.2325 5.5825 36.3675 ;
        RECT  5.7075 36.2325 5.7725 36.3675 ;
        RECT  5.7075 36.2325 5.7725 36.3675 ;
        RECT  5.8975 36.2325 5.9625 36.3675 ;
        RECT  5.7075 36.2325 5.7725 36.3675 ;
        RECT  5.8975 36.2325 5.9625 36.3675 ;
        RECT  5.5175 35.3925 5.5825 35.5275 ;
        RECT  5.7075 35.3925 5.7725 35.5275 ;
        RECT  5.5175 35.3925 5.5825 35.5275 ;
        RECT  5.7075 35.3925 5.7725 35.5275 ;
        RECT  5.7075 35.3925 5.7725 35.5275 ;
        RECT  5.8975 35.3925 5.9625 35.5275 ;
        RECT  5.7075 35.3925 5.7725 35.5275 ;
        RECT  5.8975 35.3925 5.9625 35.5275 ;
        RECT  6.0675 35.3475 6.1325 35.4825 ;
        RECT  6.0675 36.2775 6.1325 36.4125 ;
        RECT  5.7675 35.6225 5.9025 35.6875 ;
        RECT  5.51 35.8375 5.645 35.9025 ;
        RECT  5.7075 36.2325 5.7725 36.3675 ;
        RECT  5.8975 35.3925 5.9625 35.5275 ;
        RECT  5.8625 35.8375 5.9975 35.9025 ;
        RECT  6.7975 35.23 6.8625 35.415 ;
        RECT  6.7975 36.345 6.8625 36.575 ;
        RECT  6.4375 35.1975 6.5025 35.3475 ;
        RECT  6.4375 36.2325 6.5025 36.6075 ;
        RECT  6.6275 35.4825 6.6925 36.2325 ;
        RECT  6.495 35.745 6.56 35.88 ;
        RECT  6.66 35.78 6.725 35.845 ;
        RECT  6.37 36.5425 6.93 36.6075 ;
        RECT  6.37 35.1975 6.93 35.2625 ;
        RECT  6.4375 36.2325 6.5025 36.3675 ;
        RECT  6.6275 36.2325 6.6925 36.3675 ;
        RECT  6.4375 36.2325 6.5025 36.3675 ;
        RECT  6.6275 36.2325 6.6925 36.3675 ;
        RECT  6.4375 35.3475 6.5025 35.4825 ;
        RECT  6.6275 35.3475 6.6925 35.4825 ;
        RECT  6.4375 35.3475 6.5025 35.4825 ;
        RECT  6.6275 35.3475 6.6925 35.4825 ;
        RECT  6.7975 35.3475 6.8625 35.4825 ;
        RECT  6.7975 36.2775 6.8625 36.4125 ;
        RECT  6.495 35.745 6.56 35.88 ;
        RECT  4.6325 35.745 4.6975 35.88 ;
        RECT  4.7725 35.5175 4.8375 35.6525 ;
        RECT  5.6325 35.6225 5.7675 35.6875 ;
        RECT  5.3175 37.735 5.3825 37.92 ;
        RECT  5.3175 36.575 5.3825 36.805 ;
        RECT  4.9575 37.8025 5.0225 37.9525 ;
        RECT  4.9575 36.5425 5.0225 36.9175 ;
        RECT  5.1475 36.9175 5.2125 37.6675 ;
        RECT  5.015 37.27 5.08 37.405 ;
        RECT  5.18 37.305 5.245 37.37 ;
        RECT  4.89 36.5425 5.45 36.6075 ;
        RECT  4.89 37.8875 5.45 37.9525 ;
        RECT  4.9575 37.0525 5.0225 37.1875 ;
        RECT  5.1475 37.0525 5.2125 37.1875 ;
        RECT  4.9575 37.0525 5.0225 37.1875 ;
        RECT  5.1475 37.0525 5.2125 37.1875 ;
        RECT  4.9575 37.7575 5.0225 37.8925 ;
        RECT  5.1475 37.7575 5.2125 37.8925 ;
        RECT  4.9575 37.7575 5.0225 37.8925 ;
        RECT  5.1475 37.7575 5.2125 37.8925 ;
        RECT  5.3175 37.8025 5.3825 37.9375 ;
        RECT  5.3175 36.8725 5.3825 37.0075 ;
        RECT  5.015 37.405 5.08 37.54 ;
        RECT  6.0675 37.735 6.1325 37.92 ;
        RECT  6.0675 36.575 6.1325 36.805 ;
        RECT  5.5175 37.7575 5.5825 37.9525 ;
        RECT  5.5175 36.5425 5.5825 36.9175 ;
        RECT  5.8975 36.5425 5.9625 36.9175 ;
        RECT  5.51 37.2475 5.645 37.3125 ;
        RECT  5.8625 37.2475 5.9975 37.3125 ;
        RECT  5.7675 37.4625 5.9025 37.5275 ;
        RECT  5.45 36.5425 6.37 36.6075 ;
        RECT  5.45 37.8875 6.37 37.9525 ;
        RECT  5.5175 37.0525 5.5825 37.1875 ;
        RECT  5.7075 37.0525 5.7725 37.1875 ;
        RECT  5.5175 37.0525 5.5825 37.1875 ;
        RECT  5.7075 37.0525 5.7725 37.1875 ;
        RECT  5.7075 37.0525 5.7725 37.1875 ;
        RECT  5.8975 37.0525 5.9625 37.1875 ;
        RECT  5.7075 37.0525 5.7725 37.1875 ;
        RECT  5.8975 37.0525 5.9625 37.1875 ;
        RECT  5.5175 37.8025 5.5825 37.9375 ;
        RECT  5.7075 37.8025 5.7725 37.9375 ;
        RECT  5.5175 37.8025 5.5825 37.9375 ;
        RECT  5.7075 37.8025 5.7725 37.9375 ;
        RECT  5.7075 37.8025 5.7725 37.9375 ;
        RECT  5.8975 37.8025 5.9625 37.9375 ;
        RECT  5.7075 37.8025 5.7725 37.9375 ;
        RECT  5.8975 37.8025 5.9625 37.9375 ;
        RECT  6.0675 37.8025 6.1325 37.9375 ;
        RECT  6.0675 36.8725 6.1325 37.0075 ;
        RECT  5.7675 37.5375 5.9025 37.6025 ;
        RECT  5.51 37.3225 5.645 37.3875 ;
        RECT  5.7075 36.9175 5.7725 37.0525 ;
        RECT  5.8975 37.7575 5.9625 37.8925 ;
        RECT  5.8625 37.3175 5.9975 37.3825 ;
        RECT  6.7975 37.735 6.8625 37.92 ;
        RECT  6.7975 36.575 6.8625 36.805 ;
        RECT  6.4375 37.8025 6.5025 37.9525 ;
        RECT  6.4375 36.5425 6.5025 36.9175 ;
        RECT  6.6275 36.9175 6.6925 37.6675 ;
        RECT  6.495 37.27 6.56 37.405 ;
        RECT  6.66 37.305 6.725 37.37 ;
        RECT  6.37 36.5425 6.93 36.6075 ;
        RECT  6.37 37.8875 6.93 37.9525 ;
        RECT  6.4375 37.0525 6.5025 37.1875 ;
        RECT  6.6275 37.0525 6.6925 37.1875 ;
        RECT  6.4375 37.0525 6.5025 37.1875 ;
        RECT  6.6275 37.0525 6.6925 37.1875 ;
        RECT  6.4375 37.7575 6.5025 37.8925 ;
        RECT  6.6275 37.7575 6.6925 37.8925 ;
        RECT  6.4375 37.7575 6.5025 37.8925 ;
        RECT  6.6275 37.7575 6.6925 37.8925 ;
        RECT  6.7975 37.8025 6.8625 37.9375 ;
        RECT  6.7975 36.8725 6.8625 37.0075 ;
        RECT  6.495 37.405 6.56 37.54 ;
        RECT  4.6325 37.27 4.6975 37.405 ;
        RECT  4.7725 37.4975 4.8375 37.6325 ;
        RECT  5.6325 37.4625 5.7675 37.5275 ;
        RECT  5.3175 37.92 5.3825 38.105 ;
        RECT  5.3175 39.035 5.3825 39.265 ;
        RECT  4.9575 37.8875 5.0225 38.0375 ;
        RECT  4.9575 38.9225 5.0225 39.2975 ;
        RECT  5.1475 38.1725 5.2125 38.9225 ;
        RECT  5.015 38.435 5.08 38.57 ;
        RECT  5.18 38.47 5.245 38.535 ;
        RECT  4.89 39.2325 5.45 39.2975 ;
        RECT  4.89 37.8875 5.45 37.9525 ;
        RECT  4.9575 38.9225 5.0225 39.0575 ;
        RECT  5.1475 38.9225 5.2125 39.0575 ;
        RECT  4.9575 38.9225 5.0225 39.0575 ;
        RECT  5.1475 38.9225 5.2125 39.0575 ;
        RECT  4.9575 38.0375 5.0225 38.1725 ;
        RECT  5.1475 38.0375 5.2125 38.1725 ;
        RECT  4.9575 38.0375 5.0225 38.1725 ;
        RECT  5.1475 38.0375 5.2125 38.1725 ;
        RECT  5.3175 38.0375 5.3825 38.1725 ;
        RECT  5.3175 38.9675 5.3825 39.1025 ;
        RECT  5.015 38.435 5.08 38.57 ;
        RECT  6.0675 37.92 6.1325 38.105 ;
        RECT  6.0675 39.035 6.1325 39.265 ;
        RECT  5.5175 37.8875 5.5825 38.0825 ;
        RECT  5.5175 38.9225 5.5825 39.2975 ;
        RECT  5.8975 38.9225 5.9625 39.2975 ;
        RECT  5.51 38.5275 5.645 38.5925 ;
        RECT  5.8625 38.5275 5.9975 38.5925 ;
        RECT  5.7675 38.3125 5.9025 38.3775 ;
        RECT  5.45 39.2325 6.37 39.2975 ;
        RECT  5.45 37.8875 6.37 37.9525 ;
        RECT  5.5175 38.9225 5.5825 39.0575 ;
        RECT  5.7075 38.9225 5.7725 39.0575 ;
        RECT  5.5175 38.9225 5.5825 39.0575 ;
        RECT  5.7075 38.9225 5.7725 39.0575 ;
        RECT  5.7075 38.9225 5.7725 39.0575 ;
        RECT  5.8975 38.9225 5.9625 39.0575 ;
        RECT  5.7075 38.9225 5.7725 39.0575 ;
        RECT  5.8975 38.9225 5.9625 39.0575 ;
        RECT  5.5175 38.0825 5.5825 38.2175 ;
        RECT  5.7075 38.0825 5.7725 38.2175 ;
        RECT  5.5175 38.0825 5.5825 38.2175 ;
        RECT  5.7075 38.0825 5.7725 38.2175 ;
        RECT  5.7075 38.0825 5.7725 38.2175 ;
        RECT  5.8975 38.0825 5.9625 38.2175 ;
        RECT  5.7075 38.0825 5.7725 38.2175 ;
        RECT  5.8975 38.0825 5.9625 38.2175 ;
        RECT  6.0675 38.0375 6.1325 38.1725 ;
        RECT  6.0675 38.9675 6.1325 39.1025 ;
        RECT  5.7675 38.3125 5.9025 38.3775 ;
        RECT  5.51 38.5275 5.645 38.5925 ;
        RECT  5.7075 38.9225 5.7725 39.0575 ;
        RECT  5.8975 38.0825 5.9625 38.2175 ;
        RECT  5.8625 38.5275 5.9975 38.5925 ;
        RECT  6.7975 37.92 6.8625 38.105 ;
        RECT  6.7975 39.035 6.8625 39.265 ;
        RECT  6.4375 37.8875 6.5025 38.0375 ;
        RECT  6.4375 38.9225 6.5025 39.2975 ;
        RECT  6.6275 38.1725 6.6925 38.9225 ;
        RECT  6.495 38.435 6.56 38.57 ;
        RECT  6.66 38.47 6.725 38.535 ;
        RECT  6.37 39.2325 6.93 39.2975 ;
        RECT  6.37 37.8875 6.93 37.9525 ;
        RECT  6.4375 38.9225 6.5025 39.0575 ;
        RECT  6.6275 38.9225 6.6925 39.0575 ;
        RECT  6.4375 38.9225 6.5025 39.0575 ;
        RECT  6.6275 38.9225 6.6925 39.0575 ;
        RECT  6.4375 38.0375 6.5025 38.1725 ;
        RECT  6.6275 38.0375 6.6925 38.1725 ;
        RECT  6.4375 38.0375 6.5025 38.1725 ;
        RECT  6.6275 38.0375 6.6925 38.1725 ;
        RECT  6.7975 38.0375 6.8625 38.1725 ;
        RECT  6.7975 38.9675 6.8625 39.1025 ;
        RECT  6.495 38.435 6.56 38.57 ;
        RECT  4.6325 38.435 4.6975 38.57 ;
        RECT  4.7725 38.2075 4.8375 38.3425 ;
        RECT  5.6325 38.3125 5.7675 38.3775 ;
        RECT  5.3175 40.425 5.3825 40.61 ;
        RECT  5.3175 39.265 5.3825 39.495 ;
        RECT  4.9575 40.4925 5.0225 40.6425 ;
        RECT  4.9575 39.2325 5.0225 39.6075 ;
        RECT  5.1475 39.6075 5.2125 40.3575 ;
        RECT  5.015 39.96 5.08 40.095 ;
        RECT  5.18 39.995 5.245 40.06 ;
        RECT  4.89 39.2325 5.45 39.2975 ;
        RECT  4.89 40.5775 5.45 40.6425 ;
        RECT  4.9575 39.7425 5.0225 39.8775 ;
        RECT  5.1475 39.7425 5.2125 39.8775 ;
        RECT  4.9575 39.7425 5.0225 39.8775 ;
        RECT  5.1475 39.7425 5.2125 39.8775 ;
        RECT  4.9575 40.4475 5.0225 40.5825 ;
        RECT  5.1475 40.4475 5.2125 40.5825 ;
        RECT  4.9575 40.4475 5.0225 40.5825 ;
        RECT  5.1475 40.4475 5.2125 40.5825 ;
        RECT  5.3175 40.4925 5.3825 40.6275 ;
        RECT  5.3175 39.5625 5.3825 39.6975 ;
        RECT  5.015 40.095 5.08 40.23 ;
        RECT  6.0675 40.425 6.1325 40.61 ;
        RECT  6.0675 39.265 6.1325 39.495 ;
        RECT  5.5175 40.4475 5.5825 40.6425 ;
        RECT  5.5175 39.2325 5.5825 39.6075 ;
        RECT  5.8975 39.2325 5.9625 39.6075 ;
        RECT  5.51 39.9375 5.645 40.0025 ;
        RECT  5.8625 39.9375 5.9975 40.0025 ;
        RECT  5.7675 40.1525 5.9025 40.2175 ;
        RECT  5.45 39.2325 6.37 39.2975 ;
        RECT  5.45 40.5775 6.37 40.6425 ;
        RECT  5.5175 39.7425 5.5825 39.8775 ;
        RECT  5.7075 39.7425 5.7725 39.8775 ;
        RECT  5.5175 39.7425 5.5825 39.8775 ;
        RECT  5.7075 39.7425 5.7725 39.8775 ;
        RECT  5.7075 39.7425 5.7725 39.8775 ;
        RECT  5.8975 39.7425 5.9625 39.8775 ;
        RECT  5.7075 39.7425 5.7725 39.8775 ;
        RECT  5.8975 39.7425 5.9625 39.8775 ;
        RECT  5.5175 40.4925 5.5825 40.6275 ;
        RECT  5.7075 40.4925 5.7725 40.6275 ;
        RECT  5.5175 40.4925 5.5825 40.6275 ;
        RECT  5.7075 40.4925 5.7725 40.6275 ;
        RECT  5.7075 40.4925 5.7725 40.6275 ;
        RECT  5.8975 40.4925 5.9625 40.6275 ;
        RECT  5.7075 40.4925 5.7725 40.6275 ;
        RECT  5.8975 40.4925 5.9625 40.6275 ;
        RECT  6.0675 40.4925 6.1325 40.6275 ;
        RECT  6.0675 39.5625 6.1325 39.6975 ;
        RECT  5.7675 40.2275 5.9025 40.2925 ;
        RECT  5.51 40.0125 5.645 40.0775 ;
        RECT  5.7075 39.6075 5.7725 39.7425 ;
        RECT  5.8975 40.4475 5.9625 40.5825 ;
        RECT  5.8625 40.0075 5.9975 40.0725 ;
        RECT  6.7975 40.425 6.8625 40.61 ;
        RECT  6.7975 39.265 6.8625 39.495 ;
        RECT  6.4375 40.4925 6.5025 40.6425 ;
        RECT  6.4375 39.2325 6.5025 39.6075 ;
        RECT  6.6275 39.6075 6.6925 40.3575 ;
        RECT  6.495 39.96 6.56 40.095 ;
        RECT  6.66 39.995 6.725 40.06 ;
        RECT  6.37 39.2325 6.93 39.2975 ;
        RECT  6.37 40.5775 6.93 40.6425 ;
        RECT  6.4375 39.7425 6.5025 39.8775 ;
        RECT  6.6275 39.7425 6.6925 39.8775 ;
        RECT  6.4375 39.7425 6.5025 39.8775 ;
        RECT  6.6275 39.7425 6.6925 39.8775 ;
        RECT  6.4375 40.4475 6.5025 40.5825 ;
        RECT  6.6275 40.4475 6.6925 40.5825 ;
        RECT  6.4375 40.4475 6.5025 40.5825 ;
        RECT  6.6275 40.4475 6.6925 40.5825 ;
        RECT  6.7975 40.4925 6.8625 40.6275 ;
        RECT  6.7975 39.5625 6.8625 39.6975 ;
        RECT  6.495 40.095 6.56 40.23 ;
        RECT  4.6325 39.96 4.6975 40.095 ;
        RECT  4.7725 40.1875 4.8375 40.3225 ;
        RECT  5.6325 40.1525 5.7675 40.2175 ;
        RECT  0.685 5.1 0.75 7.92 ;
        RECT  0.845 5.1 0.91 7.92 ;
        RECT  3.69 5.1 3.755 7.92 ;
        RECT  6.65 5.1 6.715 7.92 ;
        RECT  1.7 5.1 1.765 7.92 ;
        RECT  4.66 5.1 4.725 7.92 ;
        RECT  3.17 7.315 3.305 7.38 ;
        RECT  3.17 7.5 3.305 7.565 ;
        RECT  1.935 7.315 2.07 7.38 ;
        RECT  1.935 7.5 2.07 7.565 ;
        RECT  3.17 7.505 3.305 7.57 ;
        RECT  3.17 7.69 3.305 7.755 ;
        RECT  6.13 7.505 6.265 7.57 ;
        RECT  6.13 7.69 6.265 7.755 ;
        RECT  1.935 7.505 2.07 7.57 ;
        RECT  1.935 7.69 2.07 7.755 ;
        RECT  6.13 7.315 6.265 7.38 ;
        RECT  6.13 7.5 6.265 7.565 ;
        RECT  1.4 7.505 1.535 7.57 ;
        RECT  1.4 7.69 1.535 7.755 ;
        RECT  4.36 7.365 4.495 7.43 ;
        RECT  4.36 7.55 4.495 7.615 ;
        RECT  4.895 7.315 5.03 7.38 ;
        RECT  4.895 7.5 5.03 7.565 ;
        RECT  4.895 7.505 5.03 7.57 ;
        RECT  4.895 7.69 5.03 7.755 ;
        RECT  5.32 7.315 5.455 7.38 ;
        RECT  5.32 7.5 5.455 7.565 ;
        RECT  2.36 7.315 2.495 7.38 ;
        RECT  2.36 7.5 2.495 7.565 ;
        RECT  5.705 7.315 5.84 7.38 ;
        RECT  5.705 7.5 5.84 7.565 ;
        RECT  5.705 7.505 5.84 7.57 ;
        RECT  5.705 7.69 5.84 7.755 ;
        RECT  2.36 7.505 2.495 7.57 ;
        RECT  2.36 7.69 2.495 7.755 ;
        RECT  5.32 7.505 5.455 7.57 ;
        RECT  5.32 7.69 5.455 7.755 ;
        RECT  2.745 7.505 2.88 7.57 ;
        RECT  2.745 7.69 2.88 7.755 ;
        RECT  2.745 7.315 2.88 7.38 ;
        RECT  2.745 7.5 2.88 7.565 ;
        RECT  0.975 7.505 1.11 7.57 ;
        RECT  0.975 7.69 1.11 7.755 ;
        RECT  3.95 7.43 4.085 7.495 ;
        RECT  3.95 7.615 4.085 7.68 ;
        RECT  0.685 7.5575 0.75 7.6925 ;
        RECT  6.1825 7.69 6.3175 7.755 ;
        RECT  4.3675 7.8 4.5025 7.865 ;
        RECT  3.4675 7.69 3.6025 7.755 ;
        RECT  3.9425 7.2675 4.0775 7.3325 ;
        RECT  6.5475 7.69 6.6825 7.755 ;
        RECT  1.005 7.1825 1.14 7.2475 ;
        RECT  5.0875 7.325 5.2225 7.39 ;
        RECT  3.48 7.3225 3.615 7.3875 ;
        RECT  2.0825 7.3225 2.2175 7.3875 ;
        RECT  0.865 7.8875 1.0 7.9525 ;
        RECT  0.9825 7.3125 1.1175 7.3775 ;
        RECT  2.5925 7.2425 2.6575 7.3775 ;
        RECT  1.5075 7.2725 1.6425 7.3375 ;
        RECT  5.5525 7.2425 5.6175 7.3775 ;
        RECT  6.44 7.365 6.575 7.43 ;
        RECT  2.97 7.445 3.105 7.51 ;
        RECT  5.93 7.455 6.065 7.52 ;
        RECT  4.24 7.6175 4.305 7.7525 ;
        RECT  3.9425 7.1825 4.0775 7.2475 ;
        RECT  1.235 7.7275 1.3 7.8625 ;
        RECT  2.7475 7.6875 2.8825 7.7525 ;
        RECT  6.44 7.3225 6.575 7.3875 ;
        RECT  5.93 7.5 6.065 7.565 ;
        RECT  5.5175 7.1825 5.6525 7.2475 ;
        RECT  0.815 7.1825 0.95 7.2475 ;
        RECT  3.48 7.3225 3.615 7.3875 ;
        RECT  2.5575 7.1825 2.6925 7.2475 ;
        RECT  2.3575 7.6875 2.4925 7.7525 ;
        RECT  2.3575 7.5 2.4925 7.565 ;
        RECT  2.97 7.5 3.105 7.565 ;
        RECT  5.3175 7.69 5.4525 7.755 ;
        RECT  5.3175 7.5 5.4525 7.565 ;
        RECT  0.685 7.18 0.75 7.955 ;
        RECT  3.755 7.82 6.65 7.885 ;
        RECT  6.265 7.315 6.575 7.38 ;
        RECT  5.84 7.69 6.13 7.755 ;
        RECT  5.03 7.69 5.32 7.755 ;
        RECT  6.6525 7.5425 6.715 7.615 ;
        RECT  6.265 7.5 6.65 7.57 ;
        RECT  5.03 7.5 5.32 7.57 ;
        RECT  5.55 7.5 5.7075 7.57 ;
        RECT  5.84 7.315 6.13 7.38 ;
        RECT  5.03 7.315 5.32 7.38 ;
        RECT  5.55 7.185 5.62 7.57 ;
        RECT  6.65 7.18 6.715 7.955 ;
        RECT  4.66 7.18 4.725 7.955 ;
        RECT  1.765 7.82 3.69 7.885 ;
        RECT  3.305 7.315 3.615 7.38 ;
        RECT  2.88 7.69 3.17 7.755 ;
        RECT  4.045 7.615 4.495 7.68 ;
        RECT  3.305 7.5 3.69 7.57 ;
        RECT  2.59 7.5 2.7475 7.57 ;
        RECT  3.6025 7.69 3.69 7.755 ;
        RECT  2.88 7.315 3.17 7.38 ;
        RECT  3.82 7.25 3.885 7.495 ;
        RECT  3.82 7.25 3.9425 7.3325 ;
        RECT  3.9425 7.245 4.0775 7.3125 ;
        RECT  3.69 7.18 3.755 7.955 ;
        RECT  2.07 7.69 2.36 7.755 ;
        RECT  1.5325 7.505 1.7 7.57 ;
        RECT  1.04 7.2475 1.11 7.505 ;
        RECT  0.975 7.69 1.4 7.755 ;
        RECT  2.07 7.5 2.36 7.57 ;
        RECT  1.23 7.69 1.305 7.8625 ;
        RECT  2.07 7.315 2.36 7.38 ;
        RECT  0.91 7.3125 0.9825 7.3775 ;
        RECT  2.59 7.185 2.66 7.57 ;
        RECT  1.62 7.2725 1.735 7.3375 ;
        RECT  0.845 7.18 0.91 7.955 ;
        RECT  1.7 7.18 1.765 7.955 ;
        RECT  0.69 7.75 0.7475 7.815 ;
        RECT  0.93 7.1825 1.0525 7.2475 ;
        RECT  4.4925 7.365 4.66 7.43 ;
        RECT  3.885 7.4275 3.9875 7.495 ;
        RECT  0.685 7.18 0.75 7.955 ;
        RECT  3.69 7.18 3.755 7.955 ;
        RECT  6.65 7.18 6.715 7.955 ;
        RECT  1.7 7.18 1.765 7.955 ;
        RECT  4.66 7.18 4.725 7.955 ;
        RECT  0.845 7.18 0.91 7.955 ;
        RECT  3.17 7.05 3.305 7.115 ;
        RECT  3.17 6.865 3.305 6.93 ;
        RECT  1.935 7.05 2.07 7.115 ;
        RECT  1.935 6.865 2.07 6.93 ;
        RECT  3.17 6.86 3.305 6.925 ;
        RECT  3.17 6.675 3.305 6.74 ;
        RECT  6.13 6.86 6.265 6.925 ;
        RECT  6.13 6.675 6.265 6.74 ;
        RECT  1.935 6.86 2.07 6.925 ;
        RECT  1.935 6.675 2.07 6.74 ;
        RECT  6.13 7.05 6.265 7.115 ;
        RECT  6.13 6.865 6.265 6.93 ;
        RECT  1.4 6.86 1.535 6.925 ;
        RECT  1.4 6.675 1.535 6.74 ;
        RECT  4.36 7.0 4.495 7.065 ;
        RECT  4.36 6.815 4.495 6.88 ;
        RECT  4.895 7.05 5.03 7.115 ;
        RECT  4.895 6.865 5.03 6.93 ;
        RECT  4.895 6.86 5.03 6.925 ;
        RECT  4.895 6.675 5.03 6.74 ;
        RECT  5.32 7.05 5.455 7.115 ;
        RECT  5.32 6.865 5.455 6.93 ;
        RECT  2.36 7.05 2.495 7.115 ;
        RECT  2.36 6.865 2.495 6.93 ;
        RECT  5.705 7.05 5.84 7.115 ;
        RECT  5.705 6.865 5.84 6.93 ;
        RECT  5.705 6.86 5.84 6.925 ;
        RECT  5.705 6.675 5.84 6.74 ;
        RECT  2.36 6.86 2.495 6.925 ;
        RECT  2.36 6.675 2.495 6.74 ;
        RECT  5.32 6.86 5.455 6.925 ;
        RECT  5.32 6.675 5.455 6.74 ;
        RECT  2.745 6.86 2.88 6.925 ;
        RECT  2.745 6.675 2.88 6.74 ;
        RECT  2.745 7.05 2.88 7.115 ;
        RECT  2.745 6.865 2.88 6.93 ;
        RECT  0.975 6.86 1.11 6.925 ;
        RECT  0.975 6.675 1.11 6.74 ;
        RECT  3.95 6.935 4.085 7.0 ;
        RECT  3.95 6.75 4.085 6.815 ;
        RECT  0.685 6.7375 0.75 6.8725 ;
        RECT  6.1825 6.675 6.3175 6.74 ;
        RECT  4.3675 6.565 4.5025 6.63 ;
        RECT  3.4675 6.675 3.6025 6.74 ;
        RECT  3.9425 7.0975 4.0775 7.1625 ;
        RECT  6.5475 6.675 6.6825 6.74 ;
        RECT  1.005 7.1825 1.14 7.2475 ;
        RECT  5.0875 7.04 5.2225 7.105 ;
        RECT  3.48 7.0425 3.615 7.1075 ;
        RECT  2.0825 7.0425 2.2175 7.1075 ;
        RECT  0.865 6.4775 1.0 6.5425 ;
        RECT  0.9825 7.0525 1.1175 7.1175 ;
        RECT  2.5925 7.0525 2.6575 7.1875 ;
        RECT  1.5075 7.0925 1.6425 7.1575 ;
        RECT  5.5525 7.0525 5.6175 7.1875 ;
        RECT  6.44 7.0 6.575 7.065 ;
        RECT  2.97 6.92 3.105 6.985 ;
        RECT  5.93 6.91 6.065 6.975 ;
        RECT  4.24 6.6775 4.305 6.8125 ;
        RECT  3.9425 7.1825 4.0775 7.2475 ;
        RECT  1.235 6.5675 1.3 6.7025 ;
        RECT  2.7475 6.6775 2.8825 6.7425 ;
        RECT  6.44 7.0425 6.575 7.1075 ;
        RECT  5.93 6.865 6.065 6.93 ;
        RECT  5.5175 7.1825 5.6525 7.2475 ;
        RECT  0.815 7.1825 0.95 7.2475 ;
        RECT  3.48 7.0425 3.615 7.1075 ;
        RECT  2.5575 7.1825 2.6925 7.2475 ;
        RECT  2.3575 6.6775 2.4925 6.7425 ;
        RECT  2.3575 6.865 2.4925 6.93 ;
        RECT  2.97 6.865 3.105 6.93 ;
        RECT  5.3175 6.675 5.4525 6.74 ;
        RECT  5.3175 6.865 5.4525 6.93 ;
        RECT  0.685 6.475 0.75 7.25 ;
        RECT  3.755 6.545 6.65 6.61 ;
        RECT  6.265 7.05 6.575 7.115 ;
        RECT  5.84 6.675 6.13 6.74 ;
        RECT  5.03 6.675 5.32 6.74 ;
        RECT  6.6525 6.815 6.715 6.8875 ;
        RECT  6.265 6.86 6.65 6.93 ;
        RECT  5.03 6.86 5.32 6.93 ;
        RECT  5.55 6.86 5.7075 6.93 ;
        RECT  5.84 7.05 6.13 7.115 ;
        RECT  5.03 7.05 5.32 7.115 ;
        RECT  5.55 6.86 5.62 7.245 ;
        RECT  6.65 6.475 6.715 7.25 ;
        RECT  4.66 6.475 4.725 7.25 ;
        RECT  1.765 6.545 3.69 6.61 ;
        RECT  3.305 7.05 3.615 7.115 ;
        RECT  2.88 6.675 3.17 6.74 ;
        RECT  4.045 6.75 4.495 6.815 ;
        RECT  3.305 6.86 3.69 6.93 ;
        RECT  2.59 6.86 2.7475 6.93 ;
        RECT  3.6025 6.675 3.69 6.74 ;
        RECT  2.88 7.05 3.17 7.115 ;
        RECT  3.82 6.935 3.885 7.18 ;
        RECT  3.82 7.0975 3.9425 7.18 ;
        RECT  3.9425 7.1175 4.0775 7.185 ;
        RECT  3.69 6.475 3.755 7.25 ;
        RECT  2.07 6.675 2.36 6.74 ;
        RECT  1.5325 6.86 1.7 6.925 ;
        RECT  1.04 6.925 1.11 7.1825 ;
        RECT  0.975 6.675 1.4 6.74 ;
        RECT  2.07 6.86 2.36 6.93 ;
        RECT  1.23 6.5675 1.305 6.74 ;
        RECT  2.07 7.05 2.36 7.115 ;
        RECT  0.91 7.0525 0.9825 7.1175 ;
        RECT  2.59 6.86 2.66 7.245 ;
        RECT  1.62 7.0925 1.735 7.1575 ;
        RECT  0.845 6.475 0.91 7.25 ;
        RECT  1.7 6.475 1.765 7.25 ;
        RECT  0.69 6.615 0.7475 6.68 ;
        RECT  0.93 7.1825 1.0525 7.2475 ;
        RECT  4.4925 7.0 4.66 7.065 ;
        RECT  3.885 6.935 3.9875 7.0025 ;
        RECT  0.685 6.475 0.75 7.25 ;
        RECT  3.69 6.475 3.755 7.25 ;
        RECT  6.65 6.475 6.715 7.25 ;
        RECT  1.7 6.475 1.765 7.25 ;
        RECT  4.66 6.475 4.725 7.25 ;
        RECT  0.845 6.475 0.91 7.25 ;
        RECT  3.17 5.905 3.305 5.97 ;
        RECT  3.17 6.09 3.305 6.155 ;
        RECT  1.935 5.905 2.07 5.97 ;
        RECT  1.935 6.09 2.07 6.155 ;
        RECT  3.17 6.095 3.305 6.16 ;
        RECT  3.17 6.28 3.305 6.345 ;
        RECT  6.13 6.095 6.265 6.16 ;
        RECT  6.13 6.28 6.265 6.345 ;
        RECT  1.935 6.095 2.07 6.16 ;
        RECT  1.935 6.28 2.07 6.345 ;
        RECT  6.13 5.905 6.265 5.97 ;
        RECT  6.13 6.09 6.265 6.155 ;
        RECT  1.4 6.095 1.535 6.16 ;
        RECT  1.4 6.28 1.535 6.345 ;
        RECT  4.36 5.955 4.495 6.02 ;
        RECT  4.36 6.14 4.495 6.205 ;
        RECT  4.895 5.905 5.03 5.97 ;
        RECT  4.895 6.09 5.03 6.155 ;
        RECT  4.895 6.095 5.03 6.16 ;
        RECT  4.895 6.28 5.03 6.345 ;
        RECT  5.32 5.905 5.455 5.97 ;
        RECT  5.32 6.09 5.455 6.155 ;
        RECT  2.36 5.905 2.495 5.97 ;
        RECT  2.36 6.09 2.495 6.155 ;
        RECT  5.705 5.905 5.84 5.97 ;
        RECT  5.705 6.09 5.84 6.155 ;
        RECT  5.705 6.095 5.84 6.16 ;
        RECT  5.705 6.28 5.84 6.345 ;
        RECT  2.36 6.095 2.495 6.16 ;
        RECT  2.36 6.28 2.495 6.345 ;
        RECT  5.32 6.095 5.455 6.16 ;
        RECT  5.32 6.28 5.455 6.345 ;
        RECT  2.745 6.095 2.88 6.16 ;
        RECT  2.745 6.28 2.88 6.345 ;
        RECT  2.745 5.905 2.88 5.97 ;
        RECT  2.745 6.09 2.88 6.155 ;
        RECT  0.975 6.095 1.11 6.16 ;
        RECT  0.975 6.28 1.11 6.345 ;
        RECT  3.95 6.02 4.085 6.085 ;
        RECT  3.95 6.205 4.085 6.27 ;
        RECT  0.685 6.1475 0.75 6.2825 ;
        RECT  6.1825 6.28 6.3175 6.345 ;
        RECT  4.3675 6.39 4.5025 6.455 ;
        RECT  3.4675 6.28 3.6025 6.345 ;
        RECT  3.9425 5.8575 4.0775 5.9225 ;
        RECT  6.5475 6.28 6.6825 6.345 ;
        RECT  1.005 5.7725 1.14 5.8375 ;
        RECT  5.0875 5.915 5.2225 5.98 ;
        RECT  3.48 5.9125 3.615 5.9775 ;
        RECT  2.0825 5.9125 2.2175 5.9775 ;
        RECT  0.865 6.4775 1.0 6.5425 ;
        RECT  0.9825 5.9025 1.1175 5.9675 ;
        RECT  2.5925 5.8325 2.6575 5.9675 ;
        RECT  1.5075 5.8625 1.6425 5.9275 ;
        RECT  5.5525 5.8325 5.6175 5.9675 ;
        RECT  6.44 5.955 6.575 6.02 ;
        RECT  2.97 6.035 3.105 6.1 ;
        RECT  5.93 6.045 6.065 6.11 ;
        RECT  4.24 6.2075 4.305 6.3425 ;
        RECT  3.9425 5.7725 4.0775 5.8375 ;
        RECT  1.235 6.3175 1.3 6.4525 ;
        RECT  2.7475 6.2775 2.8825 6.3425 ;
        RECT  6.44 5.9125 6.575 5.9775 ;
        RECT  5.93 6.09 6.065 6.155 ;
        RECT  5.5175 5.7725 5.6525 5.8375 ;
        RECT  0.815 5.7725 0.95 5.8375 ;
        RECT  3.48 5.9125 3.615 5.9775 ;
        RECT  2.5575 5.7725 2.6925 5.8375 ;
        RECT  2.3575 6.2775 2.4925 6.3425 ;
        RECT  2.3575 6.09 2.4925 6.155 ;
        RECT  2.97 6.09 3.105 6.155 ;
        RECT  5.3175 6.28 5.4525 6.345 ;
        RECT  5.3175 6.09 5.4525 6.155 ;
        RECT  0.685 5.77 0.75 6.545 ;
        RECT  3.755 6.41 6.65 6.475 ;
        RECT  6.265 5.905 6.575 5.97 ;
        RECT  5.84 6.28 6.13 6.345 ;
        RECT  5.03 6.28 5.32 6.345 ;
        RECT  6.6525 6.1325 6.715 6.205 ;
        RECT  6.265 6.09 6.65 6.16 ;
        RECT  5.03 6.09 5.32 6.16 ;
        RECT  5.55 6.09 5.7075 6.16 ;
        RECT  5.84 5.905 6.13 5.97 ;
        RECT  5.03 5.905 5.32 5.97 ;
        RECT  5.55 5.775 5.62 6.16 ;
        RECT  6.65 5.77 6.715 6.545 ;
        RECT  4.66 5.77 4.725 6.545 ;
        RECT  1.765 6.41 3.69 6.475 ;
        RECT  3.305 5.905 3.615 5.97 ;
        RECT  2.88 6.28 3.17 6.345 ;
        RECT  4.045 6.205 4.495 6.27 ;
        RECT  3.305 6.09 3.69 6.16 ;
        RECT  2.59 6.09 2.7475 6.16 ;
        RECT  3.6025 6.28 3.69 6.345 ;
        RECT  2.88 5.905 3.17 5.97 ;
        RECT  3.82 5.84 3.885 6.085 ;
        RECT  3.82 5.84 3.9425 5.9225 ;
        RECT  3.9425 5.835 4.0775 5.9025 ;
        RECT  3.69 5.77 3.755 6.545 ;
        RECT  2.07 6.28 2.36 6.345 ;
        RECT  1.5325 6.095 1.7 6.16 ;
        RECT  1.04 5.8375 1.11 6.095 ;
        RECT  0.975 6.28 1.4 6.345 ;
        RECT  2.07 6.09 2.36 6.16 ;
        RECT  1.23 6.28 1.305 6.4525 ;
        RECT  2.07 5.905 2.36 5.97 ;
        RECT  0.91 5.9025 0.9825 5.9675 ;
        RECT  2.59 5.775 2.66 6.16 ;
        RECT  1.62 5.8625 1.735 5.9275 ;
        RECT  0.845 5.77 0.91 6.545 ;
        RECT  1.7 5.77 1.765 6.545 ;
        RECT  0.69 6.34 0.7475 6.405 ;
        RECT  0.93 5.7725 1.0525 5.8375 ;
        RECT  4.4925 5.955 4.66 6.02 ;
        RECT  3.885 6.0175 3.9875 6.085 ;
        RECT  0.685 5.77 0.75 6.545 ;
        RECT  3.69 5.77 3.755 6.545 ;
        RECT  6.65 5.77 6.715 6.545 ;
        RECT  1.7 5.77 1.765 6.545 ;
        RECT  4.66 5.77 4.725 6.545 ;
        RECT  0.845 5.77 0.91 6.545 ;
        RECT  3.17 5.64 3.305 5.705 ;
        RECT  3.17 5.455 3.305 5.52 ;
        RECT  1.935 5.64 2.07 5.705 ;
        RECT  1.935 5.455 2.07 5.52 ;
        RECT  3.17 5.45 3.305 5.515 ;
        RECT  3.17 5.265 3.305 5.33 ;
        RECT  6.13 5.45 6.265 5.515 ;
        RECT  6.13 5.265 6.265 5.33 ;
        RECT  1.935 5.45 2.07 5.515 ;
        RECT  1.935 5.265 2.07 5.33 ;
        RECT  6.13 5.64 6.265 5.705 ;
        RECT  6.13 5.455 6.265 5.52 ;
        RECT  1.4 5.45 1.535 5.515 ;
        RECT  1.4 5.265 1.535 5.33 ;
        RECT  4.36 5.59 4.495 5.655 ;
        RECT  4.36 5.405 4.495 5.47 ;
        RECT  4.895 5.64 5.03 5.705 ;
        RECT  4.895 5.455 5.03 5.52 ;
        RECT  4.895 5.45 5.03 5.515 ;
        RECT  4.895 5.265 5.03 5.33 ;
        RECT  5.32 5.64 5.455 5.705 ;
        RECT  5.32 5.455 5.455 5.52 ;
        RECT  2.36 5.64 2.495 5.705 ;
        RECT  2.36 5.455 2.495 5.52 ;
        RECT  5.705 5.64 5.84 5.705 ;
        RECT  5.705 5.455 5.84 5.52 ;
        RECT  5.705 5.45 5.84 5.515 ;
        RECT  5.705 5.265 5.84 5.33 ;
        RECT  2.36 5.45 2.495 5.515 ;
        RECT  2.36 5.265 2.495 5.33 ;
        RECT  5.32 5.45 5.455 5.515 ;
        RECT  5.32 5.265 5.455 5.33 ;
        RECT  2.745 5.45 2.88 5.515 ;
        RECT  2.745 5.265 2.88 5.33 ;
        RECT  2.745 5.64 2.88 5.705 ;
        RECT  2.745 5.455 2.88 5.52 ;
        RECT  0.975 5.45 1.11 5.515 ;
        RECT  0.975 5.265 1.11 5.33 ;
        RECT  3.95 5.525 4.085 5.59 ;
        RECT  3.95 5.34 4.085 5.405 ;
        RECT  0.685 5.3275 0.75 5.4625 ;
        RECT  6.1825 5.265 6.3175 5.33 ;
        RECT  4.3675 5.155 4.5025 5.22 ;
        RECT  3.4675 5.265 3.6025 5.33 ;
        RECT  3.9425 5.6875 4.0775 5.7525 ;
        RECT  6.5475 5.265 6.6825 5.33 ;
        RECT  1.005 5.7725 1.14 5.8375 ;
        RECT  5.0875 5.63 5.2225 5.695 ;
        RECT  3.48 5.6325 3.615 5.6975 ;
        RECT  2.0825 5.6325 2.2175 5.6975 ;
        RECT  0.865 5.0675 1.0 5.1325 ;
        RECT  0.9825 5.6425 1.1175 5.7075 ;
        RECT  2.5925 5.6425 2.6575 5.7775 ;
        RECT  1.5075 5.6825 1.6425 5.7475 ;
        RECT  5.5525 5.6425 5.6175 5.7775 ;
        RECT  6.44 5.59 6.575 5.655 ;
        RECT  2.97 5.51 3.105 5.575 ;
        RECT  5.93 5.5 6.065 5.565 ;
        RECT  4.24 5.2675 4.305 5.4025 ;
        RECT  3.9425 5.7725 4.0775 5.8375 ;
        RECT  1.235 5.1575 1.3 5.2925 ;
        RECT  2.7475 5.2675 2.8825 5.3325 ;
        RECT  6.44 5.6325 6.575 5.6975 ;
        RECT  5.93 5.455 6.065 5.52 ;
        RECT  5.5175 5.7725 5.6525 5.8375 ;
        RECT  0.815 5.7725 0.95 5.8375 ;
        RECT  3.48 5.6325 3.615 5.6975 ;
        RECT  2.5575 5.7725 2.6925 5.8375 ;
        RECT  2.3575 5.2675 2.4925 5.3325 ;
        RECT  2.3575 5.455 2.4925 5.52 ;
        RECT  2.97 5.455 3.105 5.52 ;
        RECT  5.3175 5.265 5.4525 5.33 ;
        RECT  5.3175 5.455 5.4525 5.52 ;
        RECT  0.685 5.065 0.75 5.84 ;
        RECT  3.755 5.135 6.65 5.2 ;
        RECT  6.265 5.64 6.575 5.705 ;
        RECT  5.84 5.265 6.13 5.33 ;
        RECT  5.03 5.265 5.32 5.33 ;
        RECT  6.6525 5.405 6.715 5.4775 ;
        RECT  6.265 5.45 6.65 5.52 ;
        RECT  5.03 5.45 5.32 5.52 ;
        RECT  5.55 5.45 5.7075 5.52 ;
        RECT  5.84 5.64 6.13 5.705 ;
        RECT  5.03 5.64 5.32 5.705 ;
        RECT  5.55 5.45 5.62 5.835 ;
        RECT  6.65 5.065 6.715 5.84 ;
        RECT  4.66 5.065 4.725 5.84 ;
        RECT  1.765 5.135 3.69 5.2 ;
        RECT  3.305 5.64 3.615 5.705 ;
        RECT  2.88 5.265 3.17 5.33 ;
        RECT  4.045 5.34 4.495 5.405 ;
        RECT  3.305 5.45 3.69 5.52 ;
        RECT  2.59 5.45 2.7475 5.52 ;
        RECT  3.6025 5.265 3.69 5.33 ;
        RECT  2.88 5.64 3.17 5.705 ;
        RECT  3.82 5.525 3.885 5.77 ;
        RECT  3.82 5.6875 3.9425 5.77 ;
        RECT  3.9425 5.7075 4.0775 5.775 ;
        RECT  3.69 5.065 3.755 5.84 ;
        RECT  2.07 5.265 2.36 5.33 ;
        RECT  1.5325 5.45 1.7 5.515 ;
        RECT  1.04 5.515 1.11 5.7725 ;
        RECT  0.975 5.265 1.4 5.33 ;
        RECT  2.07 5.45 2.36 5.52 ;
        RECT  1.23 5.1575 1.305 5.33 ;
        RECT  2.07 5.64 2.36 5.705 ;
        RECT  0.91 5.6425 0.9825 5.7075 ;
        RECT  2.59 5.45 2.66 5.835 ;
        RECT  1.62 5.6825 1.735 5.7475 ;
        RECT  0.845 5.065 0.91 5.84 ;
        RECT  1.7 5.065 1.765 5.84 ;
        RECT  0.69 5.205 0.7475 5.27 ;
        RECT  0.93 5.7725 1.0525 5.8375 ;
        RECT  4.4925 5.59 4.66 5.655 ;
        RECT  3.885 5.525 3.9875 5.5925 ;
        RECT  0.685 5.065 0.75 5.84 ;
        RECT  3.69 5.065 3.755 5.84 ;
        RECT  6.65 5.065 6.715 5.84 ;
        RECT  1.7 5.065 1.765 5.84 ;
        RECT  4.66 5.065 4.725 5.84 ;
        RECT  0.845 5.065 0.91 5.84 ;
        RECT  8.2525 19.0575 8.3875 19.1225 ;
        RECT  8.2525 21.7475 8.3875 21.8125 ;
        RECT  8.2525 24.4375 8.3875 24.5025 ;
        RECT  8.2525 27.1275 8.3875 27.1925 ;
        RECT  8.2525 29.8175 8.3875 29.8825 ;
        RECT  8.2525 32.5075 8.3875 32.5725 ;
        RECT  8.2525 35.1975 8.3875 35.2625 ;
        RECT  8.2525 37.8875 8.3875 37.9525 ;
        RECT  8.2525 40.5775 8.3875 40.6425 ;
        RECT  6.785 8.5025 6.92 8.5675 ;
        RECT  7.195 8.5025 7.33 8.5675 ;
        RECT  6.51 9.8475 6.645 9.9125 ;
        RECT  7.4 9.8475 7.535 9.9125 ;
        RECT  6.785 13.8825 6.92 13.9475 ;
        RECT  7.605 13.8825 7.74 13.9475 ;
        RECT  6.51 15.2275 6.645 15.2925 ;
        RECT  7.81 15.2275 7.945 15.2925 ;
        RECT  6.99 8.2975 7.125 8.3625 ;
        RECT  6.99 10.9875 7.125 11.0525 ;
        RECT  6.99 13.6775 7.125 13.7425 ;
        RECT  6.99 16.3675 7.125 16.4325 ;
        RECT  6.8525 7.535 6.9875 7.6 ;
        RECT  7.195 7.535 7.33 7.6 ;
        RECT  6.8525 6.83 6.9875 6.895 ;
        RECT  7.4 6.83 7.535 6.895 ;
        RECT  6.8525 6.125 6.9875 6.19 ;
        RECT  7.605 6.125 7.74 6.19 ;
        RECT  6.8525 5.42 6.9875 5.485 ;
        RECT  7.81 5.42 7.945 5.485 ;
        RECT  6.92 7.8875 7.055 7.9525 ;
        RECT  8.2525 7.8875 8.3875 7.9525 ;
        RECT  6.92 7.1825 7.055 7.2475 ;
        RECT  8.2525 7.1825 8.3875 7.2475 ;
        RECT  6.92 6.4775 7.055 6.5425 ;
        RECT  8.2525 6.4775 8.3875 6.5425 ;
        RECT  6.92 5.7725 7.055 5.8375 ;
        RECT  8.2525 5.7725 8.3875 5.8375 ;
        RECT  6.92 5.0675 7.055 5.1325 ;
        RECT  8.2525 5.0675 8.3875 5.1325 ;
        RECT  9.39 3.795 9.525 3.86 ;
        RECT  8.98 1.61 9.115 1.675 ;
        RECT  9.185 3.1575 9.32 3.2225 ;
        RECT  9.39 41.4775 9.525 41.5425 ;
        RECT  9.595 10.2975 9.73 10.3625 ;
        RECT  9.8 14.3225 9.935 14.3875 ;
        RECT  8.775 8.0925 8.91 8.1575 ;
        RECT  4.5975 40.7825 4.7325 40.8475 ;
        RECT  8.775 40.7825 8.91 40.8475 ;
        RECT  8.4675 3.0275 8.6025 3.0925 ;
        RECT  8.4675 14.4525 8.6025 14.5175 ;
        RECT  8.4675 3.955 8.6025 4.02 ;
        RECT  8.4675 11.23 8.6025 11.295 ;
        RECT  -0.725 19.52 -0.66 19.585 ;
        RECT  -0.7225 19.52 -0.6925 19.585 ;
        RECT  -0.725 19.5525 -0.66 20.1375 ;
        RECT  -0.725 20.6825 -0.66 21.0775 ;
        RECT  -0.725 22.0025 -0.66 22.5875 ;
        RECT  -1.895 22.44 -1.5175 22.505 ;
        RECT  -1.895 25.4 -1.5175 25.465 ;
        RECT  -1.895 20.45 -1.5175 20.515 ;
        RECT  -1.895 23.41 -1.5175 23.475 ;
        RECT  -0.755 19.52 -0.69 19.585 ;
        RECT  -0.725 20.65 -0.66 20.715 ;
        RECT  -2.28 31.335 -2.215 32.1 ;
        RECT  -0.725 24.685 -0.66 26.115 ;
        RECT  -1.895 19.435 -1.69 19.5 ;
        RECT  -2.2775 26.115 -2.2125 28.0525 ;
        RECT  -2.4925 26.525 -2.4275 28.31 ;
        RECT  -0.95 27.55 -0.885 28.12 ;
        RECT  -0.81 27.345 -0.745 28.31 ;
        RECT  -0.67 26.73 -0.605 28.5 ;
        RECT  -0.95 29.06 -0.885 29.125 ;
        RECT  -0.95 28.595 -0.885 29.0925 ;
        RECT  -0.9175 29.06 -0.7225 29.125 ;
        RECT  -0.72 29.225 -0.655 29.29 ;
        RECT  -0.7225 29.225 -0.6875 29.29 ;
        RECT  -0.72 29.2575 -0.655 32.7975 ;
        RECT  -3.64 27.55 -3.575 28.68 ;
        RECT  -3.5 26.73 -3.435 28.87 ;
        RECT  -3.36 26.935 -3.295 29.06 ;
        RECT  -3.64 29.62 -3.575 29.685 ;
        RECT  -3.64 29.155 -3.575 29.6525 ;
        RECT  -3.6075 29.62 -3.4125 29.685 ;
        RECT  -3.445 29.8175 -3.38 30.2125 ;
        RECT  -3.445 30.3775 -3.38 30.7725 ;
        RECT  -2.28 31.3025 -2.215 31.3675 ;
        RECT  -2.28 31.3025 -2.2475 31.3675 ;
        RECT  -2.28 31.21 -2.215 31.335 ;
        RECT  -2.28 30.6175 -2.215 31.0125 ;
        RECT  -2.2775 28.475 -2.2125 28.845 ;
        RECT  -2.2225 29.55 -2.1575 29.99 ;
        RECT  -3.445 30.9375 -3.38 31.175 ;
        RECT  -2.28 30.215 -2.215 30.4525 ;
        RECT  -0.1725 19.23 -0.1075 31.335 ;
        RECT  -0.1725 26.32 -0.1075 27.925 ;
        RECT  -1.5175 19.23 -1.4525 31.335 ;
        RECT  -1.5175 27.14 -1.4525 27.925 ;
        RECT  -2.8625 27.925 -2.7975 31.335 ;
        RECT  -2.8625 26.32 -2.7975 27.925 ;
        RECT  -4.2075 27.925 -4.1425 31.335 ;
        RECT  -4.2075 27.14 -4.1425 27.925 ;
        RECT  -4.2075 31.3025 -4.1425 31.3675 ;
        RECT  -4.2075 31.13 -4.1425 31.335 ;
        RECT  -4.22 31.3025 -4.175 31.3675 ;
        RECT  -0.79 19.355 -0.655 19.42 ;
        RECT  -1.5175 19.23 -1.4525 19.295 ;
        RECT  -0.1725 19.23 -0.1075 19.295 ;
        RECT  -4.01 19.435 -1.895 19.5 ;
        RECT  -4.01 19.595 -1.895 19.66 ;
        RECT  -4.01 22.44 -1.895 22.505 ;
        RECT  -4.01 25.4 -1.895 25.465 ;
        RECT  -4.01 20.45 -1.895 20.515 ;
        RECT  -4.01 23.41 -1.895 23.475 ;
        RECT  -3.47 21.92 -3.405 22.055 ;
        RECT  -3.655 21.92 -3.59 22.055 ;
        RECT  -3.47 20.685 -3.405 20.82 ;
        RECT  -3.655 20.685 -3.59 20.82 ;
        RECT  -3.66 21.92 -3.595 22.055 ;
        RECT  -3.845 21.92 -3.78 22.055 ;
        RECT  -3.66 24.88 -3.595 25.015 ;
        RECT  -3.845 24.88 -3.78 25.015 ;
        RECT  -3.66 20.685 -3.595 20.82 ;
        RECT  -3.845 20.685 -3.78 20.82 ;
        RECT  -3.47 24.88 -3.405 25.015 ;
        RECT  -3.655 24.88 -3.59 25.015 ;
        RECT  -3.66 20.15 -3.595 20.285 ;
        RECT  -3.845 20.15 -3.78 20.285 ;
        RECT  -3.52 23.11 -3.455 23.245 ;
        RECT  -3.705 23.11 -3.64 23.245 ;
        RECT  -3.47 23.645 -3.405 23.78 ;
        RECT  -3.655 23.645 -3.59 23.78 ;
        RECT  -3.66 23.645 -3.595 23.78 ;
        RECT  -3.845 23.645 -3.78 23.78 ;
        RECT  -3.47 24.07 -3.405 24.205 ;
        RECT  -3.655 24.07 -3.59 24.205 ;
        RECT  -3.47 21.11 -3.405 21.245 ;
        RECT  -3.655 21.11 -3.59 21.245 ;
        RECT  -3.47 24.455 -3.405 24.59 ;
        RECT  -3.655 24.455 -3.59 24.59 ;
        RECT  -3.66 24.455 -3.595 24.59 ;
        RECT  -3.845 24.455 -3.78 24.59 ;
        RECT  -3.66 21.11 -3.595 21.245 ;
        RECT  -3.845 21.11 -3.78 21.245 ;
        RECT  -3.66 24.07 -3.595 24.205 ;
        RECT  -3.845 24.07 -3.78 24.205 ;
        RECT  -3.66 21.495 -3.595 21.63 ;
        RECT  -3.845 21.495 -3.78 21.63 ;
        RECT  -3.47 21.495 -3.405 21.63 ;
        RECT  -3.655 21.495 -3.59 21.63 ;
        RECT  -3.66 19.725 -3.595 19.86 ;
        RECT  -3.845 19.725 -3.78 19.86 ;
        RECT  -3.585 22.7 -3.52 22.835 ;
        RECT  -3.77 22.7 -3.705 22.835 ;
        RECT  -3.7825 19.435 -3.6475 19.5 ;
        RECT  -3.845 24.9325 -3.78 25.0675 ;
        RECT  -3.955 23.1175 -3.89 23.2525 ;
        RECT  -3.845 22.2175 -3.78 22.3525 ;
        RECT  -3.4225 22.6925 -3.3575 22.8275 ;
        RECT  -3.845 25.2975 -3.78 25.4325 ;
        RECT  -3.3375 19.755 -3.2725 19.89 ;
        RECT  -3.48 23.8375 -3.415 23.9725 ;
        RECT  -3.4775 22.23 -3.4125 22.365 ;
        RECT  -3.4775 20.8325 -3.4125 20.9675 ;
        RECT  -4.0425 19.615 -3.9775 19.75 ;
        RECT  -3.4675 19.7325 -3.4025 19.8675 ;
        RECT  -3.4675 21.3425 -3.3325 21.4075 ;
        RECT  -3.4275 20.2575 -3.3625 20.3925 ;
        RECT  -3.4675 24.3025 -3.3325 24.3675 ;
        RECT  -3.52 25.19 -3.455 25.325 ;
        RECT  -3.6 21.72 -3.535 21.855 ;
        RECT  -3.61 24.68 -3.545 24.815 ;
        RECT  -3.8425 22.99 -3.7075 23.055 ;
        RECT  -3.3375 22.6925 -3.2725 22.8275 ;
        RECT  -3.9525 19.985 -3.8175 20.05 ;
        RECT  -3.8425 21.4975 -3.7775 21.6325 ;
        RECT  -3.4775 25.19 -3.4125 25.325 ;
        RECT  -3.655 24.68 -3.59 24.815 ;
        RECT  -3.3375 24.2675 -3.2725 24.4025 ;
        RECT  -3.3375 19.565 -3.2725 19.7 ;
        RECT  -3.4775 22.23 -3.4125 22.365 ;
        RECT  -3.3375 21.3075 -3.2725 21.4425 ;
        RECT  -3.8425 21.1075 -3.7775 21.2425 ;
        RECT  -3.655 21.1075 -3.59 21.2425 ;
        RECT  -3.655 21.72 -3.59 21.855 ;
        RECT  -3.845 24.0675 -3.78 24.2025 ;
        RECT  -3.655 24.0675 -3.59 24.2025 ;
        RECT  -4.045 19.435 -3.27 19.5 ;
        RECT  -3.975 22.505 -3.91 25.4 ;
        RECT  -3.47 25.015 -3.405 25.325 ;
        RECT  -3.845 24.59 -3.78 24.88 ;
        RECT  -3.845 23.78 -3.78 24.07 ;
        RECT  -3.705 25.4025 -3.6325 25.465 ;
        RECT  -3.66 25.015 -3.59 25.4 ;
        RECT  -3.66 23.78 -3.59 24.07 ;
        RECT  -3.66 24.3 -3.59 24.4575 ;
        RECT  -3.47 24.59 -3.405 24.88 ;
        RECT  -3.47 23.78 -3.405 24.07 ;
        RECT  -3.66 24.3 -3.275 24.37 ;
        RECT  -4.045 25.4 -3.27 25.465 ;
        RECT  -4.045 23.41 -3.27 23.475 ;
        RECT  -3.975 20.515 -3.91 22.44 ;
        RECT  -3.47 22.055 -3.405 22.365 ;
        RECT  -3.845 21.63 -3.78 21.92 ;
        RECT  -3.77 22.795 -3.705 23.245 ;
        RECT  -3.66 22.055 -3.59 22.44 ;
        RECT  -3.66 21.34 -3.59 21.4975 ;
        RECT  -3.845 22.3525 -3.78 22.44 ;
        RECT  -3.47 21.63 -3.405 21.92 ;
        RECT  -3.585 22.57 -3.34 22.635 ;
        RECT  -3.4225 22.57 -3.34 22.6925 ;
        RECT  -3.4025 22.6925 -3.335 22.8275 ;
        RECT  -4.045 22.44 -3.27 22.505 ;
        RECT  -3.845 20.82 -3.78 21.11 ;
        RECT  -3.66 20.2825 -3.595 20.45 ;
        RECT  -3.595 19.79 -3.3375 19.86 ;
        RECT  -3.845 19.725 -3.78 20.15 ;
        RECT  -3.66 20.82 -3.59 21.11 ;
        RECT  -3.9525 19.98 -3.78 20.055 ;
        RECT  -3.47 20.82 -3.405 21.11 ;
        RECT  -3.4675 19.66 -3.4025 19.7325 ;
        RECT  -3.66 21.34 -3.275 21.41 ;
        RECT  -3.4275 20.37 -3.3625 20.485 ;
        RECT  -4.045 19.595 -3.27 19.66 ;
        RECT  -4.045 20.45 -3.27 20.515 ;
        RECT  -3.905 19.44 -3.84 19.4975 ;
        RECT  -3.3375 19.68 -3.2725 19.8025 ;
        RECT  -3.52 23.2425 -3.455 23.41 ;
        RECT  -3.585 22.635 -3.5175 22.7375 ;
        RECT  -4.045 19.435 -3.27 19.5 ;
        RECT  -4.045 22.44 -3.27 22.505 ;
        RECT  -4.045 25.4 -3.27 25.465 ;
        RECT  -4.045 20.45 -3.27 20.515 ;
        RECT  -4.045 23.41 -3.27 23.475 ;
        RECT  -4.045 19.595 -3.27 19.66 ;
        RECT  -3.205 21.92 -3.14 22.055 ;
        RECT  -3.02 21.92 -2.955 22.055 ;
        RECT  -3.205 20.685 -3.14 20.82 ;
        RECT  -3.02 20.685 -2.955 20.82 ;
        RECT  -3.015 21.92 -2.95 22.055 ;
        RECT  -2.83 21.92 -2.765 22.055 ;
        RECT  -3.015 24.88 -2.95 25.015 ;
        RECT  -2.83 24.88 -2.765 25.015 ;
        RECT  -3.015 20.685 -2.95 20.82 ;
        RECT  -2.83 20.685 -2.765 20.82 ;
        RECT  -3.205 24.88 -3.14 25.015 ;
        RECT  -3.02 24.88 -2.955 25.015 ;
        RECT  -3.015 20.15 -2.95 20.285 ;
        RECT  -2.83 20.15 -2.765 20.285 ;
        RECT  -3.155 23.11 -3.09 23.245 ;
        RECT  -2.97 23.11 -2.905 23.245 ;
        RECT  -3.205 23.645 -3.14 23.78 ;
        RECT  -3.02 23.645 -2.955 23.78 ;
        RECT  -3.015 23.645 -2.95 23.78 ;
        RECT  -2.83 23.645 -2.765 23.78 ;
        RECT  -3.205 24.07 -3.14 24.205 ;
        RECT  -3.02 24.07 -2.955 24.205 ;
        RECT  -3.205 21.11 -3.14 21.245 ;
        RECT  -3.02 21.11 -2.955 21.245 ;
        RECT  -3.205 24.455 -3.14 24.59 ;
        RECT  -3.02 24.455 -2.955 24.59 ;
        RECT  -3.015 24.455 -2.95 24.59 ;
        RECT  -2.83 24.455 -2.765 24.59 ;
        RECT  -3.015 21.11 -2.95 21.245 ;
        RECT  -2.83 21.11 -2.765 21.245 ;
        RECT  -3.015 24.07 -2.95 24.205 ;
        RECT  -2.83 24.07 -2.765 24.205 ;
        RECT  -3.015 21.495 -2.95 21.63 ;
        RECT  -2.83 21.495 -2.765 21.63 ;
        RECT  -3.205 21.495 -3.14 21.63 ;
        RECT  -3.02 21.495 -2.955 21.63 ;
        RECT  -3.015 19.725 -2.95 19.86 ;
        RECT  -2.83 19.725 -2.765 19.86 ;
        RECT  -3.09 22.7 -3.025 22.835 ;
        RECT  -2.905 22.7 -2.84 22.835 ;
        RECT  -2.9625 19.435 -2.8275 19.5 ;
        RECT  -2.83 24.9325 -2.765 25.0675 ;
        RECT  -2.72 23.1175 -2.655 23.2525 ;
        RECT  -2.83 22.2175 -2.765 22.3525 ;
        RECT  -3.2525 22.6925 -3.1875 22.8275 ;
        RECT  -2.83 25.2975 -2.765 25.4325 ;
        RECT  -3.3375 19.755 -3.2725 19.89 ;
        RECT  -3.195 23.8375 -3.13 23.9725 ;
        RECT  -3.1975 22.23 -3.1325 22.365 ;
        RECT  -3.1975 20.8325 -3.1325 20.9675 ;
        RECT  -2.6325 19.615 -2.5675 19.75 ;
        RECT  -3.2075 19.7325 -3.1425 19.8675 ;
        RECT  -3.2775 21.3425 -3.1425 21.4075 ;
        RECT  -3.2475 20.2575 -3.1825 20.3925 ;
        RECT  -3.2775 24.3025 -3.1425 24.3675 ;
        RECT  -3.155 25.19 -3.09 25.325 ;
        RECT  -3.075 21.72 -3.01 21.855 ;
        RECT  -3.065 24.68 -3.0 24.815 ;
        RECT  -2.9025 22.99 -2.7675 23.055 ;
        RECT  -3.3375 22.6925 -3.2725 22.8275 ;
        RECT  -2.7925 19.985 -2.6575 20.05 ;
        RECT  -2.8325 21.4975 -2.7675 21.6325 ;
        RECT  -3.1975 25.19 -3.1325 25.325 ;
        RECT  -3.02 24.68 -2.955 24.815 ;
        RECT  -3.3375 24.2675 -3.2725 24.4025 ;
        RECT  -3.3375 19.565 -3.2725 19.7 ;
        RECT  -3.1975 22.23 -3.1325 22.365 ;
        RECT  -3.3375 21.3075 -3.2725 21.4425 ;
        RECT  -2.8325 21.1075 -2.7675 21.2425 ;
        RECT  -3.02 21.1075 -2.955 21.2425 ;
        RECT  -3.02 21.72 -2.955 21.855 ;
        RECT  -2.83 24.0675 -2.765 24.2025 ;
        RECT  -3.02 24.0675 -2.955 24.2025 ;
        RECT  -3.34 19.435 -2.565 19.5 ;
        RECT  -2.7 22.505 -2.635 25.4 ;
        RECT  -3.205 25.015 -3.14 25.325 ;
        RECT  -2.83 24.59 -2.765 24.88 ;
        RECT  -2.83 23.78 -2.765 24.07 ;
        RECT  -2.9775 25.4025 -2.905 25.465 ;
        RECT  -3.02 25.015 -2.95 25.4 ;
        RECT  -3.02 23.78 -2.95 24.07 ;
        RECT  -3.02 24.3 -2.95 24.4575 ;
        RECT  -3.205 24.59 -3.14 24.88 ;
        RECT  -3.205 23.78 -3.14 24.07 ;
        RECT  -3.335 24.3 -2.95 24.37 ;
        RECT  -3.34 25.4 -2.565 25.465 ;
        RECT  -3.34 23.41 -2.565 23.475 ;
        RECT  -2.7 20.515 -2.635 22.44 ;
        RECT  -3.205 22.055 -3.14 22.365 ;
        RECT  -2.83 21.63 -2.765 21.92 ;
        RECT  -2.905 22.795 -2.84 23.245 ;
        RECT  -3.02 22.055 -2.95 22.44 ;
        RECT  -3.02 21.34 -2.95 21.4975 ;
        RECT  -2.83 22.3525 -2.765 22.44 ;
        RECT  -3.205 21.63 -3.14 21.92 ;
        RECT  -3.27 22.57 -3.025 22.635 ;
        RECT  -3.27 22.57 -3.1875 22.6925 ;
        RECT  -3.275 22.6925 -3.2075 22.8275 ;
        RECT  -3.34 22.44 -2.565 22.505 ;
        RECT  -2.83 20.82 -2.765 21.11 ;
        RECT  -3.015 20.2825 -2.95 20.45 ;
        RECT  -3.2725 19.79 -3.015 19.86 ;
        RECT  -2.83 19.725 -2.765 20.15 ;
        RECT  -3.02 20.82 -2.95 21.11 ;
        RECT  -2.83 19.98 -2.6575 20.055 ;
        RECT  -3.205 20.82 -3.14 21.11 ;
        RECT  -3.2075 19.66 -3.1425 19.7325 ;
        RECT  -3.335 21.34 -2.95 21.41 ;
        RECT  -3.2475 20.37 -3.1825 20.485 ;
        RECT  -3.34 19.595 -2.565 19.66 ;
        RECT  -3.34 20.45 -2.565 20.515 ;
        RECT  -2.77 19.44 -2.705 19.4975 ;
        RECT  -3.3375 19.68 -3.2725 19.8025 ;
        RECT  -3.155 23.2425 -3.09 23.41 ;
        RECT  -3.0925 22.635 -3.025 22.7375 ;
        RECT  -3.34 19.435 -2.565 19.5 ;
        RECT  -3.34 22.44 -2.565 22.505 ;
        RECT  -3.34 25.4 -2.565 25.465 ;
        RECT  -3.34 20.45 -2.565 20.515 ;
        RECT  -3.34 23.41 -2.565 23.475 ;
        RECT  -3.34 19.595 -2.565 19.66 ;
        RECT  -2.06 21.92 -1.995 22.055 ;
        RECT  -2.245 21.92 -2.18 22.055 ;
        RECT  -2.06 20.685 -1.995 20.82 ;
        RECT  -2.245 20.685 -2.18 20.82 ;
        RECT  -2.25 21.92 -2.185 22.055 ;
        RECT  -2.435 21.92 -2.37 22.055 ;
        RECT  -2.25 24.88 -2.185 25.015 ;
        RECT  -2.435 24.88 -2.37 25.015 ;
        RECT  -2.25 20.685 -2.185 20.82 ;
        RECT  -2.435 20.685 -2.37 20.82 ;
        RECT  -2.06 24.88 -1.995 25.015 ;
        RECT  -2.245 24.88 -2.18 25.015 ;
        RECT  -2.25 20.15 -2.185 20.285 ;
        RECT  -2.435 20.15 -2.37 20.285 ;
        RECT  -2.11 23.11 -2.045 23.245 ;
        RECT  -2.295 23.11 -2.23 23.245 ;
        RECT  -2.06 23.645 -1.995 23.78 ;
        RECT  -2.245 23.645 -2.18 23.78 ;
        RECT  -2.25 23.645 -2.185 23.78 ;
        RECT  -2.435 23.645 -2.37 23.78 ;
        RECT  -2.06 24.07 -1.995 24.205 ;
        RECT  -2.245 24.07 -2.18 24.205 ;
        RECT  -2.06 21.11 -1.995 21.245 ;
        RECT  -2.245 21.11 -2.18 21.245 ;
        RECT  -2.06 24.455 -1.995 24.59 ;
        RECT  -2.245 24.455 -2.18 24.59 ;
        RECT  -2.25 24.455 -2.185 24.59 ;
        RECT  -2.435 24.455 -2.37 24.59 ;
        RECT  -2.25 21.11 -2.185 21.245 ;
        RECT  -2.435 21.11 -2.37 21.245 ;
        RECT  -2.25 24.07 -2.185 24.205 ;
        RECT  -2.435 24.07 -2.37 24.205 ;
        RECT  -2.25 21.495 -2.185 21.63 ;
        RECT  -2.435 21.495 -2.37 21.63 ;
        RECT  -2.06 21.495 -1.995 21.63 ;
        RECT  -2.245 21.495 -2.18 21.63 ;
        RECT  -2.25 19.725 -2.185 19.86 ;
        RECT  -2.435 19.725 -2.37 19.86 ;
        RECT  -2.175 22.7 -2.11 22.835 ;
        RECT  -2.36 22.7 -2.295 22.835 ;
        RECT  -2.3725 19.435 -2.2375 19.5 ;
        RECT  -2.435 24.9325 -2.37 25.0675 ;
        RECT  -2.545 23.1175 -2.48 23.2525 ;
        RECT  -2.435 22.2175 -2.37 22.3525 ;
        RECT  -2.0125 22.6925 -1.9475 22.8275 ;
        RECT  -2.435 25.2975 -2.37 25.4325 ;
        RECT  -1.9275 19.755 -1.8625 19.89 ;
        RECT  -2.07 23.8375 -2.005 23.9725 ;
        RECT  -2.0675 22.23 -2.0025 22.365 ;
        RECT  -2.0675 20.8325 -2.0025 20.9675 ;
        RECT  -2.6325 19.615 -2.5675 19.75 ;
        RECT  -2.0575 19.7325 -1.9925 19.8675 ;
        RECT  -2.0575 21.3425 -1.9225 21.4075 ;
        RECT  -2.0175 20.2575 -1.9525 20.3925 ;
        RECT  -2.0575 24.3025 -1.9225 24.3675 ;
        RECT  -2.11 25.19 -2.045 25.325 ;
        RECT  -2.19 21.72 -2.125 21.855 ;
        RECT  -2.2 24.68 -2.135 24.815 ;
        RECT  -2.4325 22.99 -2.2975 23.055 ;
        RECT  -1.9275 22.6925 -1.8625 22.8275 ;
        RECT  -2.5425 19.985 -2.4075 20.05 ;
        RECT  -2.4325 21.4975 -2.3675 21.6325 ;
        RECT  -2.0675 25.19 -2.0025 25.325 ;
        RECT  -2.245 24.68 -2.18 24.815 ;
        RECT  -1.9275 24.2675 -1.8625 24.4025 ;
        RECT  -1.9275 19.565 -1.8625 19.7 ;
        RECT  -2.0675 22.23 -2.0025 22.365 ;
        RECT  -1.9275 21.3075 -1.8625 21.4425 ;
        RECT  -2.4325 21.1075 -2.3675 21.2425 ;
        RECT  -2.245 21.1075 -2.18 21.2425 ;
        RECT  -2.245 21.72 -2.18 21.855 ;
        RECT  -2.435 24.0675 -2.37 24.2025 ;
        RECT  -2.245 24.0675 -2.18 24.2025 ;
        RECT  -2.635 19.435 -1.86 19.5 ;
        RECT  -2.565 22.505 -2.5 25.4 ;
        RECT  -2.06 25.015 -1.995 25.325 ;
        RECT  -2.435 24.59 -2.37 24.88 ;
        RECT  -2.435 23.78 -2.37 24.07 ;
        RECT  -2.295 25.4025 -2.2225 25.465 ;
        RECT  -2.25 25.015 -2.18 25.4 ;
        RECT  -2.25 23.78 -2.18 24.07 ;
        RECT  -2.25 24.3 -2.18 24.4575 ;
        RECT  -2.06 24.59 -1.995 24.88 ;
        RECT  -2.06 23.78 -1.995 24.07 ;
        RECT  -2.25 24.3 -1.865 24.37 ;
        RECT  -2.635 25.4 -1.86 25.465 ;
        RECT  -2.635 23.41 -1.86 23.475 ;
        RECT  -2.565 20.515 -2.5 22.44 ;
        RECT  -2.06 22.055 -1.995 22.365 ;
        RECT  -2.435 21.63 -2.37 21.92 ;
        RECT  -2.36 22.795 -2.295 23.245 ;
        RECT  -2.25 22.055 -2.18 22.44 ;
        RECT  -2.25 21.34 -2.18 21.4975 ;
        RECT  -2.435 22.3525 -2.37 22.44 ;
        RECT  -2.06 21.63 -1.995 21.92 ;
        RECT  -2.175 22.57 -1.93 22.635 ;
        RECT  -2.0125 22.57 -1.93 22.6925 ;
        RECT  -1.9925 22.6925 -1.925 22.8275 ;
        RECT  -2.635 22.44 -1.86 22.505 ;
        RECT  -2.435 20.82 -2.37 21.11 ;
        RECT  -2.25 20.2825 -2.185 20.45 ;
        RECT  -2.185 19.79 -1.9275 19.86 ;
        RECT  -2.435 19.725 -2.37 20.15 ;
        RECT  -2.25 20.82 -2.18 21.11 ;
        RECT  -2.5425 19.98 -2.37 20.055 ;
        RECT  -2.06 20.82 -1.995 21.11 ;
        RECT  -2.0575 19.66 -1.9925 19.7325 ;
        RECT  -2.25 21.34 -1.865 21.41 ;
        RECT  -2.0175 20.37 -1.9525 20.485 ;
        RECT  -2.635 19.595 -1.86 19.66 ;
        RECT  -2.635 20.45 -1.86 20.515 ;
        RECT  -2.495 19.44 -2.43 19.4975 ;
        RECT  -1.9275 19.68 -1.8625 19.8025 ;
        RECT  -2.11 23.2425 -2.045 23.41 ;
        RECT  -2.175 22.635 -2.1075 22.7375 ;
        RECT  -2.635 19.435 -1.86 19.5 ;
        RECT  -2.635 22.44 -1.86 22.505 ;
        RECT  -2.635 25.4 -1.86 25.465 ;
        RECT  -2.635 20.45 -1.86 20.515 ;
        RECT  -2.635 23.41 -1.86 23.475 ;
        RECT  -2.635 19.595 -1.86 19.66 ;
        RECT  -0.325 19.8475 -0.14 19.9125 ;
        RECT  -1.485 19.8475 -1.255 19.9125 ;
        RECT  -1.5175 19.2975 -1.3425 19.7425 ;
        RECT  -1.1425 19.4875 -0.3925 19.5525 ;
        RECT  -0.79 19.355 -0.655 19.42 ;
        RECT  -0.755 19.52 -0.69 19.585 ;
        RECT  -1.5175 19.23 -1.4525 19.98 ;
        RECT  -0.1725 19.23 -0.1075 19.98 ;
        RECT  -1.375 19.2975 -1.21 19.3625 ;
        RECT  -1.375 19.6775 -1.21 19.7425 ;
        RECT  -1.4075 19.2975 -1.3425 19.7425 ;
        RECT  -1.2775 19.4875 -1.1425 19.5525 ;
        RECT  -1.2775 19.2975 -1.1425 19.3625 ;
        RECT  -1.2775 19.6775 -1.1425 19.7425 ;
        RECT  -1.2775 19.4875 -1.1425 19.5525 ;
        RECT  -0.325 19.2975 -0.16 19.3625 ;
        RECT  -0.325 19.6775 -0.16 19.7425 ;
        RECT  -0.1925 19.2975 -0.1275 19.7425 ;
        RECT  -0.3925 19.4875 -0.2575 19.5525 ;
        RECT  -0.3925 19.2975 -0.2575 19.3625 ;
        RECT  -0.3925 19.6775 -0.2575 19.7425 ;
        RECT  -0.3925 19.4875 -0.2575 19.5525 ;
        RECT  -0.3925 19.8475 -0.2575 19.9125 ;
        RECT  -1.3225 19.8475 -1.1875 19.9125 ;
        RECT  -0.79 19.355 -0.655 19.42 ;
        RECT  -0.325 20.7875 -0.14 20.8525 ;
        RECT  -1.485 20.7875 -1.255 20.8525 ;
        RECT  -1.5175 20.0475 -1.2975 20.4925 ;
        RECT  -0.9675 20.6175 -0.5375 20.6825 ;
        RECT  -0.76 20.105 -0.625 20.17 ;
        RECT  -0.725 20.65 -0.66 20.715 ;
        RECT  -1.5175 19.98 -1.4525 20.92 ;
        RECT  -0.1725 19.98 -0.1075 20.92 ;
        RECT  -1.33 20.0475 -1.165 20.1125 ;
        RECT  -1.33 20.4275 -1.165 20.4925 ;
        RECT  -1.165 20.2375 -1.0 20.3025 ;
        RECT  -1.165 20.6175 -1.0 20.6825 ;
        RECT  -1.3625 20.0475 -1.2975 20.4925 ;
        RECT  -1.0325 20.2375 -0.9675 20.6825 ;
        RECT  -1.2325 20.0475 -1.0975 20.1125 ;
        RECT  -1.2325 20.4275 -1.0975 20.4925 ;
        RECT  -1.2325 20.2375 -1.0975 20.3025 ;
        RECT  -1.2325 20.6175 -1.0975 20.6825 ;
        RECT  -0.34 20.0475 -0.175 20.1125 ;
        RECT  -0.34 20.4275 -0.175 20.4925 ;
        RECT  -0.505 20.2375 -0.34 20.3025 ;
        RECT  -0.505 20.6175 -0.34 20.6825 ;
        RECT  -0.2075 20.0475 -0.1425 20.4925 ;
        RECT  -0.5375 20.2375 -0.4725 20.6825 ;
        RECT  -0.4075 20.0475 -0.2725 20.1125 ;
        RECT  -0.4075 20.4275 -0.2725 20.4925 ;
        RECT  -0.4075 20.2375 -0.2725 20.3025 ;
        RECT  -0.4075 20.6175 -0.2725 20.6825 ;
        RECT  -0.3925 20.7875 -0.2575 20.8525 ;
        RECT  -1.3225 20.7875 -1.1875 20.8525 ;
        RECT  -0.76 20.105 -0.625 20.17 ;
        RECT  -0.325 22.2975 -0.14 22.3625 ;
        RECT  -1.485 22.2975 -1.255 22.3625 ;
        RECT  -1.5175 20.9875 -1.2975 22.1925 ;
        RECT  -0.9675 21.9375 -0.5375 22.0025 ;
        RECT  -0.76 21.045 -0.625 21.11 ;
        RECT  -0.725 21.97 -0.66 22.035 ;
        RECT  -1.5175 20.92 -1.4525 22.43 ;
        RECT  -0.1725 20.92 -0.1075 22.43 ;
        RECT  -1.33 20.9875 -1.165 21.0525 ;
        RECT  -1.33 21.3675 -1.165 21.4325 ;
        RECT  -1.33 21.7475 -1.165 21.8125 ;
        RECT  -1.33 22.1275 -1.165 22.1925 ;
        RECT  -1.165 21.1775 -1.0 21.2425 ;
        RECT  -1.165 21.5575 -1.0 21.6225 ;
        RECT  -1.165 21.9375 -1.0 22.0025 ;
        RECT  -1.3625 20.9875 -1.2975 22.1925 ;
        RECT  -1.0325 21.1775 -0.9675 22.0025 ;
        RECT  -1.2325 20.9875 -1.0975 21.0525 ;
        RECT  -1.2325 21.3675 -1.0975 21.4325 ;
        RECT  -1.2325 21.7475 -1.0975 21.8125 ;
        RECT  -1.2325 22.1275 -1.0975 22.1925 ;
        RECT  -1.2325 21.1775 -1.0975 21.2425 ;
        RECT  -1.2325 21.5575 -1.0975 21.6225 ;
        RECT  -1.2325 21.9375 -1.0975 22.0025 ;
        RECT  -0.34 20.9875 -0.175 21.0525 ;
        RECT  -0.34 21.3675 -0.175 21.4325 ;
        RECT  -0.34 21.7475 -0.175 21.8125 ;
        RECT  -0.34 22.1275 -0.175 22.1925 ;
        RECT  -0.505 21.1775 -0.34 21.2425 ;
        RECT  -0.505 21.5575 -0.34 21.6225 ;
        RECT  -0.505 21.9375 -0.34 22.0025 ;
        RECT  -0.2075 20.9875 -0.1425 22.1925 ;
        RECT  -0.5375 21.1775 -0.4725 22.0025 ;
        RECT  -0.4075 20.9875 -0.2725 21.0525 ;
        RECT  -0.4075 21.3675 -0.2725 21.4325 ;
        RECT  -0.4075 21.7475 -0.2725 21.8125 ;
        RECT  -0.4075 22.1275 -0.2725 22.1925 ;
        RECT  -0.4075 21.1775 -0.2725 21.2425 ;
        RECT  -0.4075 21.5575 -0.2725 21.6225 ;
        RECT  -0.4075 21.9375 -0.2725 22.0025 ;
        RECT  -0.3925 22.2975 -0.2575 22.3625 ;
        RECT  -1.3225 22.2975 -1.1875 22.3625 ;
        RECT  -0.76 21.045 -0.625 21.11 ;
        RECT  -0.325 24.9475 -0.14 25.0125 ;
        RECT  -1.485 24.9475 -1.255 25.0125 ;
        RECT  -1.5175 22.4975 -1.2975 24.8425 ;
        RECT  -0.9675 24.5875 -0.5375 24.6525 ;
        RECT  -0.76 22.555 -0.625 22.62 ;
        RECT  -0.725 24.62 -0.66 24.685 ;
        RECT  -1.5175 22.43 -1.4525 25.08 ;
        RECT  -0.1725 22.43 -0.1075 25.08 ;
        RECT  -1.33 22.4975 -1.165 22.5625 ;
        RECT  -1.33 22.8775 -1.165 22.9425 ;
        RECT  -1.33 23.2575 -1.165 23.3225 ;
        RECT  -1.33 23.6375 -1.165 23.7025 ;
        RECT  -1.33 24.0175 -1.165 24.0825 ;
        RECT  -1.33 24.3975 -1.165 24.4625 ;
        RECT  -1.33 24.7775 -1.165 24.8425 ;
        RECT  -1.165 22.6875 -1.0 22.7525 ;
        RECT  -1.165 23.0675 -1.0 23.1325 ;
        RECT  -1.165 23.4475 -1.0 23.5125 ;
        RECT  -1.165 23.8275 -1.0 23.8925 ;
        RECT  -1.165 24.2075 -1.0 24.2725 ;
        RECT  -1.165 24.5875 -1.0 24.6525 ;
        RECT  -1.3625 22.4975 -1.2975 24.8425 ;
        RECT  -1.0325 22.6875 -0.9675 24.6525 ;
        RECT  -1.2325 22.4975 -1.0975 22.5625 ;
        RECT  -1.2325 22.8775 -1.0975 22.9425 ;
        RECT  -1.2325 23.2575 -1.0975 23.3225 ;
        RECT  -1.2325 23.6375 -1.0975 23.7025 ;
        RECT  -1.2325 24.0175 -1.0975 24.0825 ;
        RECT  -1.2325 24.3975 -1.0975 24.4625 ;
        RECT  -1.2325 24.7775 -1.0975 24.8425 ;
        RECT  -1.2325 22.6875 -1.0975 22.7525 ;
        RECT  -1.2325 23.0675 -1.0975 23.1325 ;
        RECT  -1.2325 23.4475 -1.0975 23.5125 ;
        RECT  -1.2325 23.8275 -1.0975 23.8925 ;
        RECT  -1.2325 24.2075 -1.0975 24.2725 ;
        RECT  -1.2325 24.5875 -1.0975 24.6525 ;
        RECT  -0.34 22.4975 -0.175 22.5625 ;
        RECT  -0.34 22.8775 -0.175 22.9425 ;
        RECT  -0.34 23.2575 -0.175 23.3225 ;
        RECT  -0.34 23.6375 -0.175 23.7025 ;
        RECT  -0.34 24.0175 -0.175 24.0825 ;
        RECT  -0.34 24.3975 -0.175 24.4625 ;
        RECT  -0.34 24.7775 -0.175 24.8425 ;
        RECT  -0.505 22.6875 -0.34 22.7525 ;
        RECT  -0.505 23.0675 -0.34 23.1325 ;
        RECT  -0.505 23.4475 -0.34 23.5125 ;
        RECT  -0.505 23.8275 -0.34 23.8925 ;
        RECT  -0.505 24.2075 -0.34 24.2725 ;
        RECT  -0.505 24.5875 -0.34 24.6525 ;
        RECT  -0.2075 22.4975 -0.1425 24.8425 ;
        RECT  -0.5375 22.6875 -0.4725 24.6525 ;
        RECT  -0.4075 22.4975 -0.2725 22.5625 ;
        RECT  -0.4075 22.8775 -0.2725 22.9425 ;
        RECT  -0.4075 23.2575 -0.2725 23.3225 ;
        RECT  -0.4075 23.6375 -0.2725 23.7025 ;
        RECT  -0.4075 24.0175 -0.2725 24.0825 ;
        RECT  -0.4075 24.3975 -0.2725 24.4625 ;
        RECT  -0.4075 24.7775 -0.2725 24.8425 ;
        RECT  -0.4075 22.6875 -0.2725 22.7525 ;
        RECT  -0.4075 23.0675 -0.2725 23.1325 ;
        RECT  -0.4075 23.4475 -0.2725 23.5125 ;
        RECT  -0.4075 23.8275 -0.2725 23.8925 ;
        RECT  -0.4075 24.2075 -0.2725 24.2725 ;
        RECT  -0.4075 24.5875 -0.2725 24.6525 ;
        RECT  -0.3925 24.9475 -0.2575 25.0125 ;
        RECT  -1.3225 24.9475 -1.1875 25.0125 ;
        RECT  -0.76 22.555 -0.625 22.62 ;
        RECT  -0.325 28.7325 -0.14 28.7975 ;
        RECT  -1.485 28.7325 -1.255 28.7975 ;
        RECT  -0.3475 27.9925 -0.1075 28.0575 ;
        RECT  -1.5175 27.9925 -1.1425 28.0575 ;
        RECT  -1.5175 28.3725 -1.1425 28.4375 ;
        RECT  -0.95 28.0525 -0.885 28.1875 ;
        RECT  -0.67 28.4325 -0.605 28.5675 ;
        RECT  -0.81 28.2425 -0.745 28.3775 ;
        RECT  -1.5175 27.925 -1.4525 28.935 ;
        RECT  -0.1725 27.925 -0.1075 28.935 ;
        RECT  -0.985 28.5625 -0.85 28.6275 ;
        RECT  -1.2775 27.9925 -1.1425 28.0575 ;
        RECT  -1.2775 28.1825 -1.1425 28.2475 ;
        RECT  -1.2775 27.9925 -1.1425 28.0575 ;
        RECT  -1.2775 28.1825 -1.1425 28.2475 ;
        RECT  -1.2775 28.1825 -1.1425 28.2475 ;
        RECT  -1.2775 28.3725 -1.1425 28.4375 ;
        RECT  -1.2775 28.1825 -1.1425 28.2475 ;
        RECT  -1.2775 28.3725 -1.1425 28.4375 ;
        RECT  -1.2775 28.3725 -1.1425 28.4375 ;
        RECT  -1.2775 28.5625 -1.1425 28.6275 ;
        RECT  -1.2775 28.3725 -1.1425 28.4375 ;
        RECT  -1.2775 28.5625 -1.1425 28.6275 ;
        RECT  -0.4825 27.9925 -0.3475 28.0575 ;
        RECT  -0.4825 28.1825 -0.3475 28.2475 ;
        RECT  -0.4825 27.9925 -0.3475 28.0575 ;
        RECT  -0.4825 28.1825 -0.3475 28.2475 ;
        RECT  -0.4825 28.1825 -0.3475 28.2475 ;
        RECT  -0.4825 28.3725 -0.3475 28.4375 ;
        RECT  -0.4825 28.1825 -0.3475 28.2475 ;
        RECT  -0.4825 28.3725 -0.3475 28.4375 ;
        RECT  -0.4825 28.3725 -0.3475 28.4375 ;
        RECT  -0.4825 28.5625 -0.3475 28.6275 ;
        RECT  -0.4825 28.3725 -0.3475 28.4375 ;
        RECT  -0.4825 28.5625 -0.3475 28.6275 ;
        RECT  -0.3925 28.7325 -0.2575 28.7975 ;
        RECT  -1.3225 28.7325 -1.1875 28.7975 ;
        RECT  -0.67 28.4325 -0.605 28.5675 ;
        RECT  -0.81 28.2425 -0.745 28.3775 ;
        RECT  -0.95 28.0525 -0.885 28.1875 ;
        RECT  -1.2775 28.1825 -1.1425 28.2475 ;
        RECT  -1.2775 28.5625 -1.1425 28.6275 ;
        RECT  -0.4825 28.5625 -0.3475 28.6275 ;
        RECT  -0.985 28.5625 -0.85 28.6275 ;
        RECT  -0.325 29.3625 -0.14 29.4275 ;
        RECT  -1.485 29.3625 -1.255 29.4275 ;
        RECT  -0.2575 29.0025 -0.1075 29.0675 ;
        RECT  -1.5175 29.0025 -1.1425 29.0675 ;
        RECT  -1.1425 29.1925 -0.3925 29.2575 ;
        RECT  -0.79 29.06 -0.655 29.125 ;
        RECT  -0.755 29.225 -0.69 29.29 ;
        RECT  -1.5175 28.935 -1.4525 29.495 ;
        RECT  -0.1725 28.935 -0.1075 29.495 ;
        RECT  -1.2775 29.0025 -1.1425 29.0675 ;
        RECT  -1.2775 29.1925 -1.1425 29.2575 ;
        RECT  -1.2775 29.0025 -1.1425 29.0675 ;
        RECT  -1.2775 29.1925 -1.1425 29.2575 ;
        RECT  -0.3925 29.0025 -0.2575 29.0675 ;
        RECT  -0.3925 29.1925 -0.2575 29.2575 ;
        RECT  -0.3925 29.0025 -0.2575 29.0675 ;
        RECT  -0.3925 29.1925 -0.2575 29.2575 ;
        RECT  -0.3925 29.3625 -0.2575 29.4275 ;
        RECT  -1.3225 29.3625 -1.1875 29.4275 ;
        RECT  -0.79 29.06 -0.655 29.125 ;
        RECT  -2.83 28.5425 -2.645 28.6075 ;
        RECT  -1.715 28.5425 -1.485 28.6075 ;
        RECT  -2.8625 27.9925 -2.7125 28.0575 ;
        RECT  -2.8625 28.3725 -2.7125 28.4375 ;
        RECT  -1.895 27.9925 -1.4525 28.0575 ;
        RECT  -2.2775 27.985 -2.2125 28.12 ;
        RECT  -2.2775 28.4075 -2.2125 28.5425 ;
        RECT  -2.4925 28.2425 -2.4275 28.3775 ;
        RECT  -1.5175 27.925 -1.4525 28.845 ;
        RECT  -2.8625 27.925 -2.7975 28.845 ;
        RECT  -2.3 27.9925 -2.165 28.0575 ;
        RECT  -2.3 28.1825 -2.165 28.2475 ;
        RECT  -2.3 27.9925 -2.165 28.0575 ;
        RECT  -2.3 28.1825 -2.165 28.2475 ;
        RECT  -2.3 28.1825 -2.165 28.2475 ;
        RECT  -2.3 28.3725 -2.165 28.4375 ;
        RECT  -2.3 28.1825 -2.165 28.2475 ;
        RECT  -2.3 28.3725 -2.165 28.4375 ;
        RECT  -2.8025 27.9925 -2.6675 28.0575 ;
        RECT  -2.8025 28.1825 -2.6675 28.2475 ;
        RECT  -2.8025 27.9925 -2.6675 28.0575 ;
        RECT  -2.8025 28.1825 -2.6675 28.2475 ;
        RECT  -2.8025 28.1825 -2.6675 28.2475 ;
        RECT  -2.8025 28.3725 -2.6675 28.4375 ;
        RECT  -2.8025 28.1825 -2.6675 28.2475 ;
        RECT  -2.8025 28.3725 -2.6675 28.4375 ;
        RECT  -2.8475 28.5425 -2.7125 28.6075 ;
        RECT  -1.9175 28.5425 -1.7825 28.6075 ;
        RECT  -2.5675 28.2425 -2.5025 28.3775 ;
        RECT  -2.3525 27.985 -2.2875 28.12 ;
        RECT  -2.03 28.3725 -1.895 28.4375 ;
        RECT  -2.7475 28.1475 -2.6825 28.2825 ;
        RECT  -2.3475 28.4075 -2.2825 28.5425 ;
        RECT  -2.83 29.6875 -2.645 29.7525 ;
        RECT  -1.715 29.6875 -1.485 29.7525 ;
        RECT  -2.8625 29.1375 -2.6675 29.2025 ;
        RECT  -1.8275 29.1375 -1.4525 29.2025 ;
        RECT  -1.8275 29.5175 -1.4525 29.5825 ;
        RECT  -2.2225 29.13 -2.1575 29.265 ;
        RECT  -2.2225 29.4825 -2.1575 29.6175 ;
        RECT  -2.4375 29.3875 -2.3725 29.5225 ;
        RECT  -1.5175 29.07 -1.4525 29.99 ;
        RECT  -2.8625 29.07 -2.7975 29.99 ;
        RECT  -2.0975 29.1375 -1.9625 29.2025 ;
        RECT  -2.0975 29.3275 -1.9625 29.3925 ;
        RECT  -2.0975 29.1375 -1.9625 29.2025 ;
        RECT  -2.0975 29.3275 -1.9625 29.3925 ;
        RECT  -2.0975 29.3275 -1.9625 29.3925 ;
        RECT  -2.0975 29.5175 -1.9625 29.5825 ;
        RECT  -2.0975 29.3275 -1.9625 29.3925 ;
        RECT  -2.0975 29.5175 -1.9625 29.5825 ;
        RECT  -2.8475 29.1375 -2.7125 29.2025 ;
        RECT  -2.8475 29.3275 -2.7125 29.3925 ;
        RECT  -2.8475 29.1375 -2.7125 29.2025 ;
        RECT  -2.8475 29.3275 -2.7125 29.3925 ;
        RECT  -2.8475 29.3275 -2.7125 29.3925 ;
        RECT  -2.8475 29.5175 -2.7125 29.5825 ;
        RECT  -2.8475 29.3275 -2.7125 29.3925 ;
        RECT  -2.8475 29.5175 -2.7125 29.5825 ;
        RECT  -2.8475 29.6875 -2.7125 29.7525 ;
        RECT  -1.9175 29.6875 -1.7825 29.7525 ;
        RECT  -2.5125 29.3875 -2.4475 29.5225 ;
        RECT  -2.2975 29.13 -2.2325 29.265 ;
        RECT  -1.9625 29.3275 -1.8275 29.3925 ;
        RECT  -2.8025 29.5175 -2.6675 29.5825 ;
        RECT  -2.2925 29.4825 -2.2275 29.6175 ;
        RECT  -2.83 30.2825 -2.645 30.3475 ;
        RECT  -1.715 30.2825 -1.485 30.3475 ;
        RECT  -2.8625 30.6425 -2.7125 30.7075 ;
        RECT  -1.8275 30.6425 -1.4525 30.7075 ;
        RECT  -2.5775 30.4525 -1.8275 30.5175 ;
        RECT  -2.315 30.585 -2.18 30.65 ;
        RECT  -2.28 30.42 -2.215 30.485 ;
        RECT  -1.5175 30.215 -1.4525 30.775 ;
        RECT  -2.8625 30.215 -2.7975 30.775 ;
        RECT  -1.8275 30.6425 -1.6925 30.7075 ;
        RECT  -1.8275 30.4525 -1.6925 30.5175 ;
        RECT  -1.8275 30.6425 -1.6925 30.7075 ;
        RECT  -1.8275 30.4525 -1.6925 30.5175 ;
        RECT  -2.7125 30.6425 -2.5775 30.7075 ;
        RECT  -2.7125 30.4525 -2.5775 30.5175 ;
        RECT  -2.7125 30.6425 -2.5775 30.7075 ;
        RECT  -2.7125 30.4525 -2.5775 30.5175 ;
        RECT  -2.7125 30.2825 -2.5775 30.3475 ;
        RECT  -1.7825 30.2825 -1.6475 30.3475 ;
        RECT  -2.315 30.585 -2.18 30.65 ;
        RECT  -2.83 30.8425 -2.645 30.9075 ;
        RECT  -1.715 30.8425 -1.485 30.9075 ;
        RECT  -2.8625 31.2025 -2.7125 31.2675 ;
        RECT  -1.8275 31.2025 -1.4525 31.2675 ;
        RECT  -2.5775 31.0125 -1.8275 31.0775 ;
        RECT  -2.315 31.145 -2.18 31.21 ;
        RECT  -2.28 30.98 -2.215 31.045 ;
        RECT  -1.5175 30.775 -1.4525 31.335 ;
        RECT  -2.8625 30.775 -2.7975 31.335 ;
        RECT  -1.8275 31.2025 -1.6925 31.2675 ;
        RECT  -1.8275 31.0125 -1.6925 31.0775 ;
        RECT  -1.8275 31.2025 -1.6925 31.2675 ;
        RECT  -1.8275 31.0125 -1.6925 31.0775 ;
        RECT  -2.7125 31.2025 -2.5775 31.2675 ;
        RECT  -2.7125 31.0125 -2.5775 31.0775 ;
        RECT  -2.7125 31.2025 -2.5775 31.2675 ;
        RECT  -2.7125 31.0125 -2.5775 31.0775 ;
        RECT  -2.7125 30.8425 -2.5775 30.9075 ;
        RECT  -1.7825 30.8425 -1.6475 30.9075 ;
        RECT  -2.315 31.145 -2.18 31.21 ;
        RECT  -3.015 29.2925 -2.83 29.3575 ;
        RECT  -4.175 29.2925 -3.945 29.3575 ;
        RECT  -3.0375 28.5525 -2.7975 28.6175 ;
        RECT  -4.2075 28.5525 -3.8325 28.6175 ;
        RECT  -4.2075 28.9325 -3.8325 28.9975 ;
        RECT  -3.64 28.6125 -3.575 28.7475 ;
        RECT  -3.36 28.9925 -3.295 29.1275 ;
        RECT  -3.5 28.8025 -3.435 28.9375 ;
        RECT  -4.2075 28.485 -4.1425 29.495 ;
        RECT  -2.8625 28.485 -2.7975 29.495 ;
        RECT  -3.675 29.1225 -3.54 29.1875 ;
        RECT  -3.9675 28.5525 -3.8325 28.6175 ;
        RECT  -3.9675 28.7425 -3.8325 28.8075 ;
        RECT  -3.9675 28.5525 -3.8325 28.6175 ;
        RECT  -3.9675 28.7425 -3.8325 28.8075 ;
        RECT  -3.9675 28.7425 -3.8325 28.8075 ;
        RECT  -3.9675 28.9325 -3.8325 28.9975 ;
        RECT  -3.9675 28.7425 -3.8325 28.8075 ;
        RECT  -3.9675 28.9325 -3.8325 28.9975 ;
        RECT  -3.9675 28.9325 -3.8325 28.9975 ;
        RECT  -3.9675 29.1225 -3.8325 29.1875 ;
        RECT  -3.9675 28.9325 -3.8325 28.9975 ;
        RECT  -3.9675 29.1225 -3.8325 29.1875 ;
        RECT  -3.1725 28.5525 -3.0375 28.6175 ;
        RECT  -3.1725 28.7425 -3.0375 28.8075 ;
        RECT  -3.1725 28.5525 -3.0375 28.6175 ;
        RECT  -3.1725 28.7425 -3.0375 28.8075 ;
        RECT  -3.1725 28.7425 -3.0375 28.8075 ;
        RECT  -3.1725 28.9325 -3.0375 28.9975 ;
        RECT  -3.1725 28.7425 -3.0375 28.8075 ;
        RECT  -3.1725 28.9325 -3.0375 28.9975 ;
        RECT  -3.1725 28.9325 -3.0375 28.9975 ;
        RECT  -3.1725 29.1225 -3.0375 29.1875 ;
        RECT  -3.1725 28.9325 -3.0375 28.9975 ;
        RECT  -3.1725 29.1225 -3.0375 29.1875 ;
        RECT  -3.0825 29.2925 -2.9475 29.3575 ;
        RECT  -4.0125 29.2925 -3.8775 29.3575 ;
        RECT  -3.36 28.9925 -3.295 29.1275 ;
        RECT  -3.5 28.8025 -3.435 28.9375 ;
        RECT  -3.64 28.6125 -3.575 28.7475 ;
        RECT  -3.9675 28.7425 -3.8325 28.8075 ;
        RECT  -3.9675 29.1225 -3.8325 29.1875 ;
        RECT  -3.1725 29.1225 -3.0375 29.1875 ;
        RECT  -3.675 29.1225 -3.54 29.1875 ;
        RECT  -3.015 29.9225 -2.83 29.9875 ;
        RECT  -4.175 29.9225 -3.945 29.9875 ;
        RECT  -2.9475 29.5625 -2.7975 29.6275 ;
        RECT  -4.2075 29.5625 -3.8325 29.6275 ;
        RECT  -3.8325 29.7525 -3.0825 29.8175 ;
        RECT  -3.48 29.62 -3.345 29.685 ;
        RECT  -3.445 29.785 -3.38 29.85 ;
        RECT  -4.2075 29.495 -4.1425 30.055 ;
        RECT  -2.8625 29.495 -2.7975 30.055 ;
        RECT  -3.9675 29.5625 -3.8325 29.6275 ;
        RECT  -3.9675 29.7525 -3.8325 29.8175 ;
        RECT  -3.9675 29.5625 -3.8325 29.6275 ;
        RECT  -3.9675 29.7525 -3.8325 29.8175 ;
        RECT  -3.0825 29.5625 -2.9475 29.6275 ;
        RECT  -3.0825 29.7525 -2.9475 29.8175 ;
        RECT  -3.0825 29.5625 -2.9475 29.6275 ;
        RECT  -3.0825 29.7525 -2.9475 29.8175 ;
        RECT  -3.0825 29.9225 -2.9475 29.9875 ;
        RECT  -4.0125 29.9225 -3.8775 29.9875 ;
        RECT  -3.48 29.62 -3.345 29.685 ;
        RECT  -3.015 30.4825 -2.83 30.5475 ;
        RECT  -4.175 30.4825 -3.945 30.5475 ;
        RECT  -2.9475 30.1225 -2.7975 30.1875 ;
        RECT  -4.2075 30.1225 -3.8325 30.1875 ;
        RECT  -3.8325 30.3125 -3.0825 30.3775 ;
        RECT  -3.48 30.18 -3.345 30.245 ;
        RECT  -3.445 30.345 -3.38 30.41 ;
        RECT  -4.2075 30.055 -4.1425 30.615 ;
        RECT  -2.8625 30.055 -2.7975 30.615 ;
        RECT  -3.9675 30.1225 -3.8325 30.1875 ;
        RECT  -3.9675 30.3125 -3.8325 30.3775 ;
        RECT  -3.9675 30.1225 -3.8325 30.1875 ;
        RECT  -3.9675 30.3125 -3.8325 30.3775 ;
        RECT  -3.0825 30.1225 -2.9475 30.1875 ;
        RECT  -3.0825 30.3125 -2.9475 30.3775 ;
        RECT  -3.0825 30.1225 -2.9475 30.1875 ;
        RECT  -3.0825 30.3125 -2.9475 30.3775 ;
        RECT  -3.0825 30.4825 -2.9475 30.5475 ;
        RECT  -4.0125 30.4825 -3.8775 30.5475 ;
        RECT  -3.48 30.18 -3.345 30.245 ;
        RECT  -3.015 31.0425 -2.83 31.1075 ;
        RECT  -4.175 31.0425 -3.945 31.1075 ;
        RECT  -2.9475 30.6825 -2.7975 30.7475 ;
        RECT  -4.2075 30.6825 -3.8325 30.7475 ;
        RECT  -3.8325 30.8725 -3.0825 30.9375 ;
        RECT  -3.48 30.74 -3.345 30.805 ;
        RECT  -3.445 30.905 -3.38 30.97 ;
        RECT  -4.2075 30.615 -4.1425 31.175 ;
        RECT  -2.8625 30.615 -2.7975 31.175 ;
        RECT  -3.9675 30.6825 -3.8325 30.7475 ;
        RECT  -3.9675 30.8725 -3.8325 30.9375 ;
        RECT  -3.9675 30.6825 -3.8325 30.7475 ;
        RECT  -3.9675 30.8725 -3.8325 30.9375 ;
        RECT  -3.0825 30.6825 -2.9475 30.7475 ;
        RECT  -3.0825 30.8725 -2.9475 30.9375 ;
        RECT  -3.0825 30.6825 -2.9475 30.7475 ;
        RECT  -3.0825 30.8725 -2.9475 30.9375 ;
        RECT  -3.0825 31.0425 -2.9475 31.1075 ;
        RECT  -4.0125 31.0425 -3.8775 31.1075 ;
        RECT  -3.48 30.74 -3.345 30.805 ;
        RECT  -3.24 33.9075 -2.795 33.9725 ;
        RECT  -3.24 36.3175 -2.795 36.3825 ;
        RECT  -3.24 36.7625 -2.83 36.8275 ;
        RECT  -4.155 35.1125 -3.24 35.1775 ;
        RECT  -4.155 32.4225 -3.24 32.4875 ;
        RECT  -2.28 33.435 -2.215 34.135 ;
        RECT  -2.28 33.6275 -2.215 33.6925 ;
        RECT  -2.28 33.435 -2.215 33.66 ;
        RECT  -3.15 33.6275 -2.2475 33.6925 ;
        RECT  -1.71 33.4975 -1.485 33.5625 ;
        RECT  -1.81 32.6275 -1.745 32.6925 ;
        RECT  -2.28 32.6275 -2.215 32.6925 ;
        RECT  -1.81 32.66 -1.745 33.3075 ;
        RECT  -2.2475 32.6275 -1.7775 32.6925 ;
        RECT  -2.28 32.33 -2.215 32.66 ;
        RECT  -3.0025 32.6275 -2.2475 32.6925 ;
        RECT  -3.425 32.03 -3.0025 32.095 ;
        RECT  -2.315 32.265 -2.18 32.33 ;
        RECT  -2.28 34.135 -2.215 34.34 ;
        RECT  -0.72 31.335 -0.655 34.26 ;
        RECT  -4.22 31.335 -4.155 36.5225 ;
        RECT  -1.5175 31.335 -1.4525 34.135 ;
        RECT  -2.865 31.335 -2.795 32.455 ;
        RECT  -0.1725 31.335 -0.1075 34.135 ;
        RECT  -2.28 31.335 -2.215 32.1 ;
        RECT  -2.83 32.8825 -2.645 32.9475 ;
        RECT  -1.715 32.8825 -1.485 32.9475 ;
        RECT  -2.8625 32.5225 -2.7125 32.5875 ;
        RECT  -1.8275 32.5225 -1.4525 32.5875 ;
        RECT  -2.5775 32.7125 -1.8275 32.7775 ;
        RECT  -2.315 32.58 -2.18 32.645 ;
        RECT  -2.28 32.745 -2.215 32.81 ;
        RECT  -1.5175 32.455 -1.4525 33.015 ;
        RECT  -2.8625 32.455 -2.7975 33.015 ;
        RECT  -2.0975 32.5225 -1.9625 32.5875 ;
        RECT  -2.0975 32.7125 -1.9625 32.7775 ;
        RECT  -2.0975 32.5225 -1.9625 32.5875 ;
        RECT  -2.0975 32.7125 -1.9625 32.7775 ;
        RECT  -2.8025 32.5225 -2.6675 32.5875 ;
        RECT  -2.8025 32.7125 -2.6675 32.7775 ;
        RECT  -2.8025 32.5225 -2.6675 32.5875 ;
        RECT  -2.8025 32.7125 -2.6675 32.7775 ;
        RECT  -2.8475 32.8825 -2.7125 32.9475 ;
        RECT  -1.9175 32.8825 -1.7825 32.9475 ;
        RECT  -2.45 32.58 -2.315 32.645 ;
        RECT  -1.845 33.2175 -1.71 33.2825 ;
        RECT  -1.845 33.0275 -1.71 33.0925 ;
        RECT  -1.845 33.2175 -1.71 33.2825 ;
        RECT  -1.845 33.0275 -1.71 33.0925 ;
        RECT  -2.8625 32.8525 -2.7975 32.9175 ;
        RECT  -0.1725 32.8525 -0.1075 32.9175 ;
        RECT  -2.8625 32.885 -2.7975 33.015 ;
        RECT  -2.83 32.8525 -0.14 32.9175 ;
        RECT  -0.1725 32.885 -0.1075 33.015 ;
        RECT  -2.28 33.93 -2.215 34.135 ;
        RECT  -1.5175 33.015 -1.4525 34.135 ;
        RECT  -2.8625 33.015 -2.7975 34.135 ;
        RECT  -0.1725 33.015 -0.1075 34.135 ;
        RECT  -0.79 33.945 -0.655 34.01 ;
        RECT  -0.325 33.6425 -0.14 33.7075 ;
        RECT  -1.485 33.6425 -1.255 33.7075 ;
        RECT  -0.2575 34.0025 -0.1075 34.0675 ;
        RECT  -1.5175 34.0025 -1.1425 34.0675 ;
        RECT  -1.1425 33.8125 -0.3925 33.8775 ;
        RECT  -0.79 33.945 -0.655 34.01 ;
        RECT  -0.755 33.78 -0.69 33.845 ;
        RECT  -1.5175 33.575 -1.4525 34.135 ;
        RECT  -0.1725 33.575 -0.1075 34.135 ;
        RECT  -1.0075 34.0025 -0.8725 34.0675 ;
        RECT  -1.0075 33.8125 -0.8725 33.8775 ;
        RECT  -1.0075 34.0025 -0.8725 34.0675 ;
        RECT  -1.0075 33.8125 -0.8725 33.8775 ;
        RECT  -0.3025 34.0025 -0.1675 34.0675 ;
        RECT  -0.3025 33.8125 -0.1675 33.8775 ;
        RECT  -0.3025 34.0025 -0.1675 34.0675 ;
        RECT  -0.3025 33.8125 -0.1675 33.8775 ;
        RECT  -0.2575 33.6425 -0.1225 33.7075 ;
        RECT  -1.1875 33.6425 -1.0525 33.7075 ;
        RECT  -0.655 33.945 -0.52 34.01 ;
        RECT  -0.325 33.0825 -0.14 33.1475 ;
        RECT  -1.485 33.0825 -1.255 33.1475 ;
        RECT  -0.2575 33.4425 -0.1075 33.5075 ;
        RECT  -1.5175 33.4425 -1.1425 33.5075 ;
        RECT  -1.1425 33.2525 -0.3925 33.3175 ;
        RECT  -0.79 33.385 -0.655 33.45 ;
        RECT  -0.755 33.22 -0.69 33.285 ;
        RECT  -1.5175 33.015 -1.4525 33.575 ;
        RECT  -0.1725 33.015 -0.1075 33.575 ;
        RECT  -1.0075 33.4425 -0.8725 33.5075 ;
        RECT  -1.0075 33.2525 -0.8725 33.3175 ;
        RECT  -1.0075 33.4425 -0.8725 33.5075 ;
        RECT  -1.0075 33.2525 -0.8725 33.3175 ;
        RECT  -0.3025 33.4425 -0.1675 33.5075 ;
        RECT  -0.3025 33.2525 -0.1675 33.3175 ;
        RECT  -0.3025 33.4425 -0.1675 33.5075 ;
        RECT  -0.3025 33.2525 -0.1675 33.3175 ;
        RECT  -0.2575 33.0825 -0.1225 33.1475 ;
        RECT  -1.1875 33.0825 -1.0525 33.1475 ;
        RECT  -0.655 33.385 -0.52 33.45 ;
        RECT  -0.79 33.385 -0.655 33.45 ;
        RECT  -2.83 33.4425 -2.645 33.5075 ;
        RECT  -1.715 33.4425 -1.485 33.5075 ;
        RECT  -2.8625 33.0825 -2.7125 33.1475 ;
        RECT  -1.8275 33.0825 -1.4525 33.1475 ;
        RECT  -2.5775 33.2725 -1.8275 33.3375 ;
        RECT  -2.315 33.14 -2.18 33.205 ;
        RECT  -2.28 33.305 -2.215 33.37 ;
        RECT  -1.5175 33.015 -1.4525 33.575 ;
        RECT  -2.8625 33.015 -2.7975 33.575 ;
        RECT  -2.0975 33.0825 -1.9625 33.1475 ;
        RECT  -2.0975 33.2725 -1.9625 33.3375 ;
        RECT  -2.0975 33.0825 -1.9625 33.1475 ;
        RECT  -2.0975 33.2725 -1.9625 33.3375 ;
        RECT  -2.8025 33.0825 -2.6675 33.1475 ;
        RECT  -2.8025 33.2725 -2.6675 33.3375 ;
        RECT  -2.8025 33.0825 -2.6675 33.1475 ;
        RECT  -2.8025 33.2725 -2.6675 33.3375 ;
        RECT  -2.8475 33.4425 -2.7125 33.5075 ;
        RECT  -1.9175 33.4425 -1.7825 33.5075 ;
        RECT  -2.45 33.14 -2.315 33.205 ;
        RECT  -2.315 33.14 -2.18 33.205 ;
        RECT  -2.83 34.0025 -2.645 34.0675 ;
        RECT  -1.715 34.0025 -1.485 34.0675 ;
        RECT  -2.8625 33.6425 -2.7125 33.7075 ;
        RECT  -1.8275 33.6425 -1.4525 33.7075 ;
        RECT  -2.5775 33.8325 -1.8275 33.8975 ;
        RECT  -2.315 33.7 -2.18 33.765 ;
        RECT  -2.28 33.865 -2.215 33.93 ;
        RECT  -1.5175 33.575 -1.4525 34.135 ;
        RECT  -2.8625 33.575 -2.7975 34.135 ;
        RECT  -2.0975 33.6425 -1.9625 33.7075 ;
        RECT  -2.0975 33.8325 -1.9625 33.8975 ;
        RECT  -2.0975 33.6425 -1.9625 33.7075 ;
        RECT  -2.0975 33.8325 -1.9625 33.8975 ;
        RECT  -2.8025 33.6425 -2.6675 33.7075 ;
        RECT  -2.8025 33.8325 -2.6675 33.8975 ;
        RECT  -2.8025 33.6425 -2.6675 33.7075 ;
        RECT  -2.8025 33.8325 -2.6675 33.8975 ;
        RECT  -2.8475 34.0025 -2.7125 34.0675 ;
        RECT  -1.9175 34.0025 -1.7825 34.0675 ;
        RECT  -2.45 33.7 -2.315 33.765 ;
        RECT  -2.315 33.7 -2.18 33.765 ;
        RECT  -0.79 33.78 -0.655 33.845 ;
        RECT  -0.79 33.22 -0.655 33.285 ;
        RECT  -2.315 33.305 -2.18 33.37 ;
        RECT  -3.895 34.0575 -3.83 34.1925 ;
        RECT  -3.71 34.0575 -3.645 34.1925 ;
        RECT  -3.54 34.0625 -3.475 34.1975 ;
        RECT  -3.355 34.0625 -3.29 34.1975 ;
        RECT  -3.975 34.4475 -3.91 34.5825 ;
        RECT  -3.79 34.4475 -3.725 34.5825 ;
        RECT  -3.46 34.4475 -3.395 34.5825 ;
        RECT  -3.275 34.4475 -3.21 34.5825 ;
        RECT  -3.975 34.9125 -3.91 35.0475 ;
        RECT  -3.79 34.9125 -3.725 35.0475 ;
        RECT  -3.46 34.9125 -3.395 35.0475 ;
        RECT  -3.275 34.9125 -3.21 35.0475 ;
        RECT  -3.2725 34.0625 -3.2075 34.1975 ;
        RECT  -3.9775 34.5375 -3.9125 34.6725 ;
        RECT  -3.2725 34.5375 -3.2075 34.6725 ;
        RECT  -3.725 34.0575 -3.66 34.1925 ;
        RECT  -3.525 34.0625 -3.46 34.1975 ;
        RECT  -3.7725 34.6525 -3.6375 34.7175 ;
        RECT  -3.5475 34.8025 -3.4125 34.8675 ;
        RECT  -3.65 33.9075 -3.515 33.9725 ;
        RECT  -3.6575 35.1125 -3.5225 35.1775 ;
        RECT  -3.655 33.7675 -3.52 33.8325 ;
        RECT  -4.0125 33.7675 -3.8775 33.8325 ;
        RECT  -3.2925 34.0625 -3.24 34.1975 ;
        RECT  -3.3075 33.7675 -3.1725 33.8325 ;
        RECT  -3.6225 35.1125 -3.5575 35.1775 ;
        RECT  -3.275 33.9075 -3.205 33.9725 ;
        RECT  -3.83 34.2825 -3.725 34.3475 ;
        RECT  -3.79 34.3475 -3.725 34.4475 ;
        RECT  -3.895 34.1925 -3.83 34.3475 ;
        RECT  -3.46 34.2825 -3.355 34.3475 ;
        RECT  -3.46 34.3475 -3.395 34.4475 ;
        RECT  -3.355 34.1975 -3.29 34.3475 ;
        RECT  -3.975 35.0475 -3.91 35.1125 ;
        RECT  -3.275 35.0475 -3.21 35.1125 ;
        RECT  -3.79 34.4475 -3.725 34.9375 ;
        RECT  -3.46 34.4475 -3.395 34.9375 ;
        RECT  -4.035 33.9075 -3.15 33.9725 ;
        RECT  -4.035 35.1125 -3.15 35.1775 ;
        RECT  -4.035 33.7675 -3.15 33.8325 ;
        RECT  -4.035 33.9075 -3.15 33.9725 ;
        RECT  -4.035 35.1125 -3.15 35.1775 ;
        RECT  -4.035 33.6275 -3.15 33.6925 ;
        RECT  -4.035 31.2175 -3.15 31.2825 ;
        RECT  -4.035 32.4225 -3.15 32.4875 ;
        RECT  -4.035 33.7675 -3.15 33.8325 ;
        RECT  -4.035 31.0775 -3.15 31.1425 ;
        RECT  -3.975 32.5525 -3.91 32.6875 ;
        RECT  -3.79 32.5525 -3.725 32.6875 ;
        RECT  -3.275 32.5525 -3.21 32.6875 ;
        RECT  -3.46 32.5525 -3.395 32.6875 ;
        RECT  -3.79 33.0175 -3.725 33.1525 ;
        RECT  -3.975 33.0175 -3.91 33.1525 ;
        RECT  -3.46 33.0175 -3.395 33.1525 ;
        RECT  -3.275 33.0175 -3.21 33.1525 ;
        RECT  -3.895 33.4075 -3.83 33.5425 ;
        RECT  -3.71 33.4075 -3.645 33.5425 ;
        RECT  -3.54 33.4075 -3.475 33.5425 ;
        RECT  -3.355 33.4075 -3.29 33.5425 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.655 32.4225 -3.52 32.4875 ;
        RECT  -3.3075 33.7675 -3.1725 33.8325 ;
        RECT  -4.0125 33.7675 -3.8775 33.8325 ;
        RECT  -3.6425 33.6275 -3.5075 33.6925 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.5475 32.7375 -3.4125 32.8025 ;
        RECT  -3.5475 32.7375 -3.4125 32.8025 ;
        RECT  -3.7725 32.8875 -3.6375 32.9525 ;
        RECT  -3.7725 32.8875 -3.6375 32.9525 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.5275 33.4075 -3.4625 33.5425 ;
        RECT  -3.2725 32.915 -3.2075 33.05 ;
        RECT  -3.2725 32.915 -3.2075 33.05 ;
        RECT  -3.2725 32.915 -3.2075 33.05 ;
        RECT  -3.2725 32.915 -3.2075 33.05 ;
        RECT  -3.2725 32.915 -3.2075 33.05 ;
        RECT  -3.2725 32.915 -3.2075 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.7225 33.4075 -3.6575 33.5425 ;
        RECT  -3.66 33.7675 -3.525 33.8325 ;
        RECT  -3.66 33.7675 -3.525 33.8325 ;
        RECT  -4.0125 33.7675 -3.8775 33.8325 ;
        RECT  -3.655 32.4225 -3.52 32.4875 ;
        RECT  -4.0125 33.7675 -3.8775 33.8325 ;
        RECT  -4.0125 33.7675 -3.8775 33.8325 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.9775 32.915 -3.9125 33.05 ;
        RECT  -3.3075 33.7675 -3.1725 33.8325 ;
        RECT  -3.6325 32.425 -3.5325 32.4875 ;
        RECT  -3.6325 32.4225 -3.5325 32.485 ;
        RECT  -3.9125 33.6275 -3.86 33.69 ;
        RECT  -3.6325 32.425 -3.5325 32.4875 ;
        RECT  -3.98 32.4875 -3.91 32.6875 ;
        RECT  -3.98 33.0175 -3.91 33.1525 ;
        RECT  -3.98 33.0175 -3.91 33.1525 ;
        RECT  -4.035 33.7675 -3.15 33.8325 ;
        RECT  -3.9 33.2525 -3.725 33.3175 ;
        RECT  -3.275 33.0175 -3.205 33.1525 ;
        RECT  -3.46 32.5775 -3.395 33.3175 ;
        RECT  -3.6325 32.4225 -3.5325 32.485 ;
        RECT  -3.2075 33.6275 -3.155 33.69 ;
        RECT  -3.98 33.0175 -3.91 33.1525 ;
        RECT  -4.035 32.4225 -3.15 32.4875 ;
        RECT  -3.79 32.6875 -3.725 33.3175 ;
        RECT  -3.98 33.0175 -3.91 33.1525 ;
        RECT  -3.98 33.0175 -3.91 33.1525 ;
        RECT  -3.36 33.2525 -3.29 33.5425 ;
        RECT  -3.275 33.0175 -3.205 33.1525 ;
        RECT  -4.035 33.6275 -3.15 33.6925 ;
        RECT  -3.98 33.0175 -3.91 33.1525 ;
        RECT  -3.98 32.4875 -3.91 32.6875 ;
        RECT  -3.275 32.4875 -3.205 32.6875 ;
        RECT  -3.9 33.2525 -3.83 33.5425 ;
        RECT  -3.46 33.2525 -3.29 33.3175 ;
        RECT  -4.035 33.6275 -3.15 33.6925 ;
        RECT  -4.035 33.7675 -3.15 33.8325 ;
        RECT  -4.035 32.4225 -3.15 32.4875 ;
        RECT  -3.975 32.2225 -3.91 32.3575 ;
        RECT  -3.79 32.2225 -3.725 32.3575 ;
        RECT  -3.275 32.2225 -3.21 32.3575 ;
        RECT  -3.46 32.2225 -3.395 32.3575 ;
        RECT  -3.79 31.7575 -3.725 31.8925 ;
        RECT  -3.975 31.7575 -3.91 31.8925 ;
        RECT  -3.46 31.7575 -3.395 31.8925 ;
        RECT  -3.275 31.7575 -3.21 31.8925 ;
        RECT  -3.895 31.3675 -3.83 31.5025 ;
        RECT  -3.71 31.3675 -3.645 31.5025 ;
        RECT  -3.54 31.3675 -3.475 31.5025 ;
        RECT  -3.355 31.3675 -3.29 31.5025 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.655 32.4225 -3.52 32.4875 ;
        RECT  -3.3075 31.0775 -3.1725 31.1425 ;
        RECT  -4.0125 31.0775 -3.8775 31.1425 ;
        RECT  -3.6425 31.2175 -3.5075 31.2825 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.5475 32.1075 -3.4125 32.1725 ;
        RECT  -3.5475 32.1075 -3.4125 32.1725 ;
        RECT  -3.7725 31.9575 -3.6375 32.0225 ;
        RECT  -3.7725 31.9575 -3.6375 32.0225 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.5275 31.3675 -3.4625 31.5025 ;
        RECT  -3.2725 31.86 -3.2075 31.995 ;
        RECT  -3.2725 31.86 -3.2075 31.995 ;
        RECT  -3.2725 31.86 -3.2075 31.995 ;
        RECT  -3.2725 31.86 -3.2075 31.995 ;
        RECT  -3.2725 31.86 -3.2075 31.995 ;
        RECT  -3.2725 31.86 -3.2075 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.7225 31.3675 -3.6575 31.5025 ;
        RECT  -3.66 31.0775 -3.525 31.1425 ;
        RECT  -3.66 31.0775 -3.525 31.1425 ;
        RECT  -4.0125 31.0775 -3.8775 31.1425 ;
        RECT  -3.655 32.4225 -3.52 32.4875 ;
        RECT  -4.0125 31.0775 -3.8775 31.1425 ;
        RECT  -4.0125 31.0775 -3.8775 31.1425 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.9775 31.86 -3.9125 31.995 ;
        RECT  -3.3075 31.0775 -3.1725 31.1425 ;
        RECT  -3.6325 32.4225 -3.5325 32.485 ;
        RECT  -3.6325 32.425 -3.5325 32.4875 ;
        RECT  -3.9125 31.22 -3.86 31.2825 ;
        RECT  -3.6325 32.4225 -3.5325 32.485 ;
        RECT  -3.98 32.2225 -3.91 32.4225 ;
        RECT  -3.98 31.7575 -3.91 31.8925 ;
        RECT  -3.98 31.7575 -3.91 31.8925 ;
        RECT  -4.035 31.0775 -3.15 31.1425 ;
        RECT  -3.9 31.5925 -3.725 31.6575 ;
        RECT  -3.275 31.7575 -3.205 31.8925 ;
        RECT  -3.46 31.5925 -3.395 32.3325 ;
        RECT  -3.6325 32.425 -3.5325 32.4875 ;
        RECT  -3.2075 31.22 -3.155 31.2825 ;
        RECT  -3.98 31.7575 -3.91 31.8925 ;
        RECT  -4.035 32.4225 -3.15 32.4875 ;
        RECT  -3.79 31.5925 -3.725 32.2225 ;
        RECT  -3.98 31.7575 -3.91 31.8925 ;
        RECT  -3.98 31.7575 -3.91 31.8925 ;
        RECT  -3.36 31.3675 -3.29 31.6575 ;
        RECT  -3.275 31.7575 -3.205 31.8925 ;
        RECT  -4.035 31.2175 -3.15 31.2825 ;
        RECT  -3.98 31.7575 -3.91 31.8925 ;
        RECT  -3.98 32.2225 -3.91 32.4225 ;
        RECT  -3.275 32.2225 -3.205 32.4225 ;
        RECT  -3.9 31.3675 -3.83 31.6575 ;
        RECT  -3.46 31.5925 -3.29 31.6575 ;
        RECT  -4.035 31.2175 -3.15 31.2825 ;
        RECT  -4.035 31.0775 -3.15 31.1425 ;
        RECT  -4.035 32.4225 -3.15 32.4875 ;
        RECT  -2.8625 33.7725 -2.7975 33.9075 ;
        RECT  -2.8625 36.1825 -2.7975 36.3175 ;
        RECT  -2.8625 34.0 -2.7975 34.135 ;
        RECT  -2.8625 31.625 -2.7975 31.76 ;
        RECT  -2.8975 36.6925 -2.7625 36.7575 ;
        RECT  -3.3075 36.6925 -3.1725 36.7575 ;
        RECT  -2.28 33.2325 -2.215 33.3675 ;
        RECT  -3.07 32.5575 -2.935 32.6225 ;
        RECT  -3.07 31.96 -2.935 32.025 ;
        RECT  -3.4925 31.96 -3.3575 32.025 ;
        RECT  -0.725 26.0475 -0.66 26.1825 ;
        RECT  -0.725 21.9675 -0.66 22.1025 ;
        RECT  -1.7225 19.4 -1.6575 19.535 ;
        RECT  -2.2775 26.0475 -2.2125 26.1825 ;
        RECT  -2.4925 26.4575 -2.4275 26.5925 ;
        RECT  -2.2225 28.995 -2.1575 29.13 ;
        RECT  -2.4375 29.2525 -2.3725 29.3875 ;
        RECT  -0.95 27.4825 -0.885 27.6175 ;
        RECT  -0.81 27.2775 -0.745 27.4125 ;
        RECT  -0.67 26.6625 -0.605 26.7975 ;
        RECT  -3.64 27.4825 -3.575 27.6175 ;
        RECT  -3.5 26.6625 -3.435 26.7975 ;
        RECT  -3.36 26.8675 -3.295 27.0025 ;
        RECT  -2.3125 28.8125 -2.1775 28.8775 ;
        RECT  -2.2575 29.9575 -2.1225 30.0225 ;
        RECT  -3.48 31.1425 -3.345 31.2075 ;
        RECT  -2.315 30.1825 -2.18 30.2475 ;
        RECT  -0.1725 26.2525 -0.1075 26.3875 ;
        RECT  -1.5175 27.0725 -1.4525 27.2075 ;
        RECT  -2.8625 26.2525 -2.7975 26.3875 ;
        RECT  -4.2075 27.0725 -4.1425 27.2075 ;
        RECT  0.1075 27.1075 0.2425 27.1725 ;
        LAYER  via1 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  10.3125 19.0575 10.3775 19.1225 ;
        RECT  11.0175 19.0575 11.0825 19.1225 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  10.5675 19.3825 10.6325 19.4475 ;
        RECT  10.3125 19.875 10.3775 19.94 ;
        RECT  10.3125 19.875 10.3775 19.94 ;
        RECT  10.3125 19.875 10.3775 19.94 ;
        RECT  10.3125 19.875 10.3775 19.94 ;
        RECT  10.3125 19.875 10.3775 19.94 ;
        RECT  10.3125 19.875 10.3775 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  10.7625 19.3825 10.8275 19.4475 ;
        RECT  11.0175 19.0575 11.0825 19.1225 ;
        RECT  11.0175 19.0575 11.0825 19.1225 ;
        RECT  11.0175 19.0575 11.0825 19.1225 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  10.3125 19.0575 10.3775 19.1225 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  10.3125 21.7475 10.3775 21.8125 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  10.5675 21.4225 10.6325 21.4875 ;
        RECT  10.3125 20.93 10.3775 20.995 ;
        RECT  10.3125 20.93 10.3775 20.995 ;
        RECT  10.3125 20.93 10.3775 20.995 ;
        RECT  10.3125 20.93 10.3775 20.995 ;
        RECT  10.3125 20.93 10.3775 20.995 ;
        RECT  10.3125 20.93 10.3775 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  10.7625 21.4225 10.8275 21.4875 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  10.3125 21.7475 10.3775 21.8125 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  10.3125 21.7475 10.3775 21.8125 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  10.5675 22.0725 10.6325 22.1375 ;
        RECT  10.3125 22.565 10.3775 22.63 ;
        RECT  10.3125 22.565 10.3775 22.63 ;
        RECT  10.3125 22.565 10.3775 22.63 ;
        RECT  10.3125 22.565 10.3775 22.63 ;
        RECT  10.3125 22.565 10.3775 22.63 ;
        RECT  10.3125 22.565 10.3775 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  10.7625 22.0725 10.8275 22.1375 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  10.3125 21.7475 10.3775 21.8125 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  10.3125 24.4375 10.3775 24.5025 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  10.5675 24.1125 10.6325 24.1775 ;
        RECT  10.3125 23.62 10.3775 23.685 ;
        RECT  10.3125 23.62 10.3775 23.685 ;
        RECT  10.3125 23.62 10.3775 23.685 ;
        RECT  10.3125 23.62 10.3775 23.685 ;
        RECT  10.3125 23.62 10.3775 23.685 ;
        RECT  10.3125 23.62 10.3775 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  10.7625 24.1125 10.8275 24.1775 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  10.3125 24.4375 10.3775 24.5025 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  10.3125 24.4375 10.3775 24.5025 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  10.5675 24.7625 10.6325 24.8275 ;
        RECT  10.3125 25.255 10.3775 25.32 ;
        RECT  10.3125 25.255 10.3775 25.32 ;
        RECT  10.3125 25.255 10.3775 25.32 ;
        RECT  10.3125 25.255 10.3775 25.32 ;
        RECT  10.3125 25.255 10.3775 25.32 ;
        RECT  10.3125 25.255 10.3775 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  10.7625 24.7625 10.8275 24.8275 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  10.3125 24.4375 10.3775 24.5025 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  10.3125 27.1275 10.3775 27.1925 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  10.5675 26.8025 10.6325 26.8675 ;
        RECT  10.3125 26.31 10.3775 26.375 ;
        RECT  10.3125 26.31 10.3775 26.375 ;
        RECT  10.3125 26.31 10.3775 26.375 ;
        RECT  10.3125 26.31 10.3775 26.375 ;
        RECT  10.3125 26.31 10.3775 26.375 ;
        RECT  10.3125 26.31 10.3775 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  10.7625 26.8025 10.8275 26.8675 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  10.3125 27.1275 10.3775 27.1925 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  10.3125 27.1275 10.3775 27.1925 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  10.5675 27.4525 10.6325 27.5175 ;
        RECT  10.3125 27.945 10.3775 28.01 ;
        RECT  10.3125 27.945 10.3775 28.01 ;
        RECT  10.3125 27.945 10.3775 28.01 ;
        RECT  10.3125 27.945 10.3775 28.01 ;
        RECT  10.3125 27.945 10.3775 28.01 ;
        RECT  10.3125 27.945 10.3775 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  10.7625 27.4525 10.8275 27.5175 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  10.3125 27.1275 10.3775 27.1925 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  10.3125 29.8175 10.3775 29.8825 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  10.5675 29.4925 10.6325 29.5575 ;
        RECT  10.3125 29.0 10.3775 29.065 ;
        RECT  10.3125 29.0 10.3775 29.065 ;
        RECT  10.3125 29.0 10.3775 29.065 ;
        RECT  10.3125 29.0 10.3775 29.065 ;
        RECT  10.3125 29.0 10.3775 29.065 ;
        RECT  10.3125 29.0 10.3775 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  10.7625 29.4925 10.8275 29.5575 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  10.3125 29.8175 10.3775 29.8825 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  10.3125 29.8175 10.3775 29.8825 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  10.5675 30.1425 10.6325 30.2075 ;
        RECT  10.3125 30.635 10.3775 30.7 ;
        RECT  10.3125 30.635 10.3775 30.7 ;
        RECT  10.3125 30.635 10.3775 30.7 ;
        RECT  10.3125 30.635 10.3775 30.7 ;
        RECT  10.3125 30.635 10.3775 30.7 ;
        RECT  10.3125 30.635 10.3775 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  10.7625 30.1425 10.8275 30.2075 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  10.3125 29.8175 10.3775 29.8825 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  10.3125 32.5075 10.3775 32.5725 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  10.5675 32.1825 10.6325 32.2475 ;
        RECT  10.3125 31.69 10.3775 31.755 ;
        RECT  10.3125 31.69 10.3775 31.755 ;
        RECT  10.3125 31.69 10.3775 31.755 ;
        RECT  10.3125 31.69 10.3775 31.755 ;
        RECT  10.3125 31.69 10.3775 31.755 ;
        RECT  10.3125 31.69 10.3775 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  10.7625 32.1825 10.8275 32.2475 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  10.3125 32.5075 10.3775 32.5725 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  10.3125 32.5075 10.3775 32.5725 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  10.5675 32.8325 10.6325 32.8975 ;
        RECT  10.3125 33.325 10.3775 33.39 ;
        RECT  10.3125 33.325 10.3775 33.39 ;
        RECT  10.3125 33.325 10.3775 33.39 ;
        RECT  10.3125 33.325 10.3775 33.39 ;
        RECT  10.3125 33.325 10.3775 33.39 ;
        RECT  10.3125 33.325 10.3775 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  10.7625 32.8325 10.8275 32.8975 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  10.3125 32.5075 10.3775 32.5725 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  10.3125 35.1975 10.3775 35.2625 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  10.5675 34.8725 10.6325 34.9375 ;
        RECT  10.3125 34.38 10.3775 34.445 ;
        RECT  10.3125 34.38 10.3775 34.445 ;
        RECT  10.3125 34.38 10.3775 34.445 ;
        RECT  10.3125 34.38 10.3775 34.445 ;
        RECT  10.3125 34.38 10.3775 34.445 ;
        RECT  10.3125 34.38 10.3775 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  10.7625 34.8725 10.8275 34.9375 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  10.3125 35.1975 10.3775 35.2625 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  10.3125 35.1975 10.3775 35.2625 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  10.5675 35.5225 10.6325 35.5875 ;
        RECT  10.3125 36.015 10.3775 36.08 ;
        RECT  10.3125 36.015 10.3775 36.08 ;
        RECT  10.3125 36.015 10.3775 36.08 ;
        RECT  10.3125 36.015 10.3775 36.08 ;
        RECT  10.3125 36.015 10.3775 36.08 ;
        RECT  10.3125 36.015 10.3775 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  10.7625 35.5225 10.8275 35.5875 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  10.3125 35.1975 10.3775 35.2625 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  10.3125 37.8875 10.3775 37.9525 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  10.5675 37.5625 10.6325 37.6275 ;
        RECT  10.3125 37.07 10.3775 37.135 ;
        RECT  10.3125 37.07 10.3775 37.135 ;
        RECT  10.3125 37.07 10.3775 37.135 ;
        RECT  10.3125 37.07 10.3775 37.135 ;
        RECT  10.3125 37.07 10.3775 37.135 ;
        RECT  10.3125 37.07 10.3775 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  10.7625 37.5625 10.8275 37.6275 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  10.3125 37.8875 10.3775 37.9525 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  10.3125 37.8875 10.3775 37.9525 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  10.5675 38.2125 10.6325 38.2775 ;
        RECT  10.3125 38.705 10.3775 38.77 ;
        RECT  10.3125 38.705 10.3775 38.77 ;
        RECT  10.3125 38.705 10.3775 38.77 ;
        RECT  10.3125 38.705 10.3775 38.77 ;
        RECT  10.3125 38.705 10.3775 38.77 ;
        RECT  10.3125 38.705 10.3775 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  10.7625 38.2125 10.8275 38.2775 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  10.3125 37.8875 10.3775 37.9525 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  10.3125 40.5775 10.3775 40.6425 ;
        RECT  11.0175 40.5775 11.0825 40.6425 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  10.5675 40.2525 10.6325 40.3175 ;
        RECT  10.3125 39.76 10.3775 39.825 ;
        RECT  10.3125 39.76 10.3775 39.825 ;
        RECT  10.3125 39.76 10.3775 39.825 ;
        RECT  10.3125 39.76 10.3775 39.825 ;
        RECT  10.3125 39.76 10.3775 39.825 ;
        RECT  10.3125 39.76 10.3775 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  10.7625 40.2525 10.8275 40.3175 ;
        RECT  11.0175 40.5775 11.0825 40.6425 ;
        RECT  11.0175 40.5775 11.0825 40.6425 ;
        RECT  11.0175 40.5775 11.0825 40.6425 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  10.3125 40.5775 10.3775 40.6425 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.0175 19.0575 11.0825 19.1225 ;
        RECT  11.7225 19.0575 11.7875 19.1225 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.2725 19.3825 11.3375 19.4475 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.4675 19.3825 11.5325 19.4475 ;
        RECT  11.7225 19.0575 11.7875 19.1225 ;
        RECT  11.7225 19.0575 11.7875 19.1225 ;
        RECT  11.7225 19.0575 11.7875 19.1225 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.0175 19.0575 11.0825 19.1225 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.2725 21.4225 11.3375 21.4875 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.4675 21.4225 11.5325 21.4875 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.2725 22.0725 11.3375 22.1375 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.4675 22.0725 11.5325 22.1375 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.2725 24.1125 11.3375 24.1775 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.4675 24.1125 11.5325 24.1775 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.2725 24.7625 11.3375 24.8275 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.4675 24.7625 11.5325 24.8275 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.2725 26.8025 11.3375 26.8675 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.4675 26.8025 11.5325 26.8675 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.2725 27.4525 11.3375 27.5175 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.4675 27.4525 11.5325 27.5175 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.2725 29.4925 11.3375 29.5575 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.4675 29.4925 11.5325 29.5575 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.2725 30.1425 11.3375 30.2075 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.4675 30.1425 11.5325 30.2075 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.2725 32.1825 11.3375 32.2475 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.4675 32.1825 11.5325 32.2475 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.2725 32.8325 11.3375 32.8975 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.4675 32.8325 11.5325 32.8975 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.2725 34.8725 11.3375 34.9375 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.4675 34.8725 11.5325 34.9375 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.2725 35.5225 11.3375 35.5875 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.4675 35.5225 11.5325 35.5875 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.2725 37.5625 11.3375 37.6275 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.4675 37.5625 11.5325 37.6275 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.2725 38.2125 11.3375 38.2775 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.4675 38.2125 11.5325 38.2775 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.0175 40.5775 11.0825 40.6425 ;
        RECT  11.7225 40.5775 11.7875 40.6425 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.2725 40.2525 11.3375 40.3175 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.4675 40.2525 11.5325 40.3175 ;
        RECT  11.7225 40.5775 11.7875 40.6425 ;
        RECT  11.7225 40.5775 11.7875 40.6425 ;
        RECT  11.7225 40.5775 11.7875 40.6425 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.0175 40.5775 11.0825 40.6425 ;
        RECT  10.5075 41.2175 10.5725 41.2825 ;
        RECT  10.6975 41.2175 10.7625 41.2825 ;
        RECT  10.5075 41.8025 10.5725 41.8675 ;
        RECT  10.8875 41.8025 10.9525 41.8675 ;
        RECT  11.2125 41.2175 11.2775 41.2825 ;
        RECT  11.4025 41.2175 11.4675 41.2825 ;
        RECT  11.2125 41.8025 11.2775 41.8675 ;
        RECT  11.5925 41.8025 11.6575 41.8675 ;
        RECT  10.665 16.38 10.73 16.445 ;
        RECT  10.665 18.5225 10.73 18.5875 ;
        RECT  10.4725 17.68 10.5375 17.745 ;
        RECT  10.855 17.27 10.92 17.335 ;
        RECT  10.3125 14.4875 10.3775 14.5525 ;
        RECT  11.0175 14.4875 11.0825 14.5525 ;
        RECT  10.66 18.7275 10.725 18.7925 ;
        RECT  11.37 16.38 11.435 16.445 ;
        RECT  11.37 18.5225 11.435 18.5875 ;
        RECT  11.1775 17.68 11.2425 17.745 ;
        RECT  11.56 17.27 11.625 17.335 ;
        RECT  11.0175 14.4875 11.0825 14.5525 ;
        RECT  11.7225 14.4875 11.7875 14.5525 ;
        RECT  11.365 18.7275 11.43 18.7925 ;
        RECT  10.5875 10.165 10.6525 10.23 ;
        RECT  11.0175 11.8 11.0825 11.865 ;
        RECT  11.0175 11.23 11.0825 11.295 ;
        RECT  10.3125 11.23 10.3775 11.295 ;
        RECT  10.7325 11.435 10.7975 11.5 ;
        RECT  11.0175 13.7275 11.0825 13.7925 ;
        RECT  10.7325 11.025 10.7975 11.09 ;
        RECT  10.5925 11.025 10.6575 11.09 ;
        RECT  11.0175 11.435 11.0825 11.5 ;
        RECT  10.3125 11.435 10.3775 11.5 ;
        RECT  10.485 10.4275 10.55 10.4925 ;
        RECT  10.5925 13.405 10.6575 13.47 ;
        RECT  10.7625 11.8 10.8275 11.865 ;
        RECT  10.4525 12.715 10.5175 12.78 ;
        RECT  10.5925 11.435 10.6575 11.5 ;
        RECT  10.3125 11.8 10.3775 11.865 ;
        RECT  10.7625 12.315 10.8275 12.38 ;
        RECT  10.4975 13.9375 10.5625 14.0025 ;
        RECT  10.3125 13.7275 10.3775 13.7925 ;
        RECT  11.2925 10.165 11.3575 10.23 ;
        RECT  11.7225 11.8 11.7875 11.865 ;
        RECT  11.7225 11.23 11.7875 11.295 ;
        RECT  11.0175 11.23 11.0825 11.295 ;
        RECT  11.4375 11.435 11.5025 11.5 ;
        RECT  11.7225 13.7275 11.7875 13.7925 ;
        RECT  11.4375 11.025 11.5025 11.09 ;
        RECT  11.2975 11.025 11.3625 11.09 ;
        RECT  11.7225 11.435 11.7875 11.5 ;
        RECT  11.0175 11.435 11.0825 11.5 ;
        RECT  11.19 10.4275 11.255 10.4925 ;
        RECT  11.2975 13.405 11.3625 13.47 ;
        RECT  11.4675 11.8 11.5325 11.865 ;
        RECT  11.1575 12.715 11.2225 12.78 ;
        RECT  11.2975 11.435 11.3625 11.5 ;
        RECT  11.0175 11.8 11.0825 11.865 ;
        RECT  11.4675 12.315 11.5325 12.38 ;
        RECT  11.2025 13.9375 11.2675 14.0025 ;
        RECT  11.0175 13.7275 11.0825 13.7925 ;
        RECT  10.51 9.3275 10.575 9.3925 ;
        RECT  11.0175 4.15 11.0825 4.215 ;
        RECT  10.875 8.2325 10.94 8.2975 ;
        RECT  10.8775 6.625 10.9425 6.69 ;
        RECT  10.8775 5.2275 10.9425 5.2925 ;
        RECT  10.3125 4.01 10.3775 4.075 ;
        RECT  11.0175 7.0875 11.0825 7.1525 ;
        RECT  10.5125 5.8925 10.5775 5.9575 ;
        RECT  10.8775 9.585 10.9425 9.65 ;
        RECT  10.7 9.075 10.765 9.14 ;
        RECT  11.0175 8.6625 11.0825 8.7275 ;
        RECT  11.0175 3.96 11.0825 4.025 ;
        RECT  11.0175 5.7025 11.0825 5.7675 ;
        RECT  10.5125 5.5025 10.5775 5.5675 ;
        RECT  10.7 5.5025 10.765 5.5675 ;
        RECT  10.7 6.115 10.765 6.18 ;
        RECT  10.51 8.4625 10.575 8.5275 ;
        RECT  10.7 8.4625 10.765 8.5275 ;
        RECT  11.525 9.3275 11.59 9.3925 ;
        RECT  11.0175 4.15 11.0825 4.215 ;
        RECT  11.16 8.2325 11.225 8.2975 ;
        RECT  11.1575 6.625 11.2225 6.69 ;
        RECT  11.1575 5.2275 11.2225 5.2925 ;
        RECT  11.7225 4.01 11.7875 4.075 ;
        RECT  11.0175 7.0875 11.0825 7.1525 ;
        RECT  11.5225 5.8925 11.5875 5.9575 ;
        RECT  11.1575 9.585 11.2225 9.65 ;
        RECT  11.335 9.075 11.4 9.14 ;
        RECT  11.0175 8.6625 11.0825 8.7275 ;
        RECT  11.0175 3.96 11.0825 4.025 ;
        RECT  11.0175 5.7025 11.0825 5.7675 ;
        RECT  11.5225 5.5025 11.5875 5.5675 ;
        RECT  11.335 5.5025 11.4 5.5675 ;
        RECT  11.335 6.115 11.4 6.18 ;
        RECT  11.525 8.4625 11.59 8.5275 ;
        RECT  11.335 8.4625 11.4 8.5275 ;
        RECT  10.7975 4.5075 10.8625 4.5725 ;
        RECT  10.6975 5.715 10.7625 5.78 ;
        RECT  10.49 5.9925 10.555 6.0575 ;
        RECT  11.0175 6.1825 11.0825 6.2475 ;
        RECT  10.7975 6.015 10.8625 6.08 ;
        RECT  11.0175 4.1225 11.0825 4.1875 ;
        RECT  10.665 5.375 10.73 5.44 ;
        RECT  10.4525 4.275 10.5175 4.34 ;
        RECT  11.5025 4.5075 11.5675 4.5725 ;
        RECT  11.4025 5.715 11.4675 5.78 ;
        RECT  11.195 5.9925 11.26 6.0575 ;
        RECT  11.7225 6.1825 11.7875 6.2475 ;
        RECT  11.5025 6.015 11.5675 6.08 ;
        RECT  11.7225 4.1225 11.7875 4.1875 ;
        RECT  11.37 5.375 11.435 5.44 ;
        RECT  11.1575 4.275 11.2225 4.34 ;
        RECT  4.1125 7.2275 4.1775 7.2925 ;
        RECT  3.9225 8.0675 3.9875 8.1325 ;
        RECT  3.9225 7.6575 3.9875 7.7225 ;
        RECT  4.1125 11.9225 4.1775 11.9875 ;
        RECT  3.9225 11.0825 3.9875 11.1475 ;
        RECT  3.9225 11.5575 3.9875 11.6225 ;
        RECT  4.1125 9.9175 4.1775 9.9825 ;
        RECT  3.9225 10.7575 3.9875 10.8225 ;
        RECT  3.9225 10.3475 3.9875 10.4125 ;
        RECT  4.1125 14.6125 4.1775 14.6775 ;
        RECT  3.9225 13.7725 3.9875 13.8375 ;
        RECT  3.9225 14.2475 3.9875 14.3125 ;
        RECT  5.4675 9.3775 5.5325 9.4425 ;
        RECT  6.8525 8.81 6.9175 8.875 ;
        RECT  5.1925 10.7225 5.2575 10.7875 ;
        RECT  6.5775 10.335 6.6425 10.4 ;
        RECT  6.8525 11.0525 6.9175 11.1175 ;
        RECT  4.9175 11.0525 4.9825 11.1175 ;
        RECT  6.5775 12.3975 6.6425 12.4625 ;
        RECT  4.6425 12.3975 4.7075 12.4625 ;
        RECT  5.4675 8.8675 5.5325 8.9325 ;
        RECT  5.1925 8.6525 5.2575 8.7175 ;
        RECT  4.9175 10.2775 4.9825 10.3425 ;
        RECT  5.1925 10.4925 5.2575 10.5575 ;
        RECT  5.4675 11.5575 5.5325 11.6225 ;
        RECT  4.6425 11.3425 4.7075 11.4075 ;
        RECT  4.9175 12.9675 4.9825 13.0325 ;
        RECT  4.6425 13.1825 4.7075 13.2475 ;
        RECT  4.1125 12.6075 4.1775 12.6725 ;
        RECT  3.9225 13.4475 3.9875 13.5125 ;
        RECT  3.9225 13.0375 3.9875 13.1025 ;
        RECT  4.1125 17.3025 4.1775 17.3675 ;
        RECT  3.9225 16.4625 3.9875 16.5275 ;
        RECT  3.9225 16.9375 3.9875 17.0025 ;
        RECT  4.1125 15.2975 4.1775 15.3625 ;
        RECT  3.9225 16.1375 3.9875 16.2025 ;
        RECT  3.9225 15.7275 3.9875 15.7925 ;
        RECT  4.1125 19.9925 4.1775 20.0575 ;
        RECT  3.9225 19.1525 3.9875 19.2175 ;
        RECT  3.9225 19.6275 3.9875 19.6925 ;
        RECT  5.4675 14.7575 5.5325 14.8225 ;
        RECT  6.8525 14.19 6.9175 14.255 ;
        RECT  5.1925 16.1025 5.2575 16.1675 ;
        RECT  6.5775 15.715 6.6425 15.78 ;
        RECT  6.8525 16.4325 6.9175 16.4975 ;
        RECT  4.9175 16.4325 4.9825 16.4975 ;
        RECT  6.5775 17.7775 6.6425 17.8425 ;
        RECT  4.6425 17.7775 4.7075 17.8425 ;
        RECT  5.4675 14.2475 5.5325 14.3125 ;
        RECT  5.1925 14.0325 5.2575 14.0975 ;
        RECT  4.9175 15.6575 4.9825 15.7225 ;
        RECT  5.1925 15.8725 5.2575 15.9375 ;
        RECT  5.4675 16.9375 5.5325 17.0025 ;
        RECT  4.6425 16.7225 4.7075 16.7875 ;
        RECT  4.9175 18.3475 4.9825 18.4125 ;
        RECT  4.6425 18.5625 4.7075 18.6275 ;
        RECT  3.2125 20.1275 3.2775 20.1925 ;
        RECT  3.4025 19.2875 3.4675 19.3525 ;
        RECT  3.4025 19.6975 3.4675 19.7625 ;
        RECT  3.2125 20.8125 3.2775 20.8775 ;
        RECT  3.4025 21.6525 3.4675 21.7175 ;
        RECT  3.4025 21.1775 3.4675 21.2425 ;
        RECT  3.2125 22.8175 3.2775 22.8825 ;
        RECT  3.4025 21.9775 3.4675 22.0425 ;
        RECT  3.4025 22.3875 3.4675 22.4525 ;
        RECT  3.2125 23.5025 3.2775 23.5675 ;
        RECT  3.4025 24.3425 3.4675 24.4075 ;
        RECT  3.4025 23.8675 3.4675 23.9325 ;
        RECT  3.2125 25.5075 3.2775 25.5725 ;
        RECT  3.4025 24.6675 3.4675 24.7325 ;
        RECT  3.4025 25.0775 3.4675 25.1425 ;
        RECT  3.2125 26.1925 3.2775 26.2575 ;
        RECT  3.4025 27.0325 3.4675 27.0975 ;
        RECT  3.4025 26.5575 3.4675 26.6225 ;
        RECT  3.2125 28.1975 3.2775 28.2625 ;
        RECT  3.4025 27.3575 3.4675 27.4225 ;
        RECT  3.4025 27.7675 3.4675 27.8325 ;
        RECT  3.2125 28.8825 3.2775 28.9475 ;
        RECT  3.4025 29.7225 3.4675 29.7875 ;
        RECT  3.4025 29.2475 3.4675 29.3125 ;
        RECT  3.2125 30.8875 3.2775 30.9525 ;
        RECT  3.4025 30.0475 3.4675 30.1125 ;
        RECT  3.4025 30.4575 3.4675 30.5225 ;
        RECT  3.2125 31.5725 3.2775 31.6375 ;
        RECT  3.4025 32.4125 3.4675 32.4775 ;
        RECT  3.4025 31.9375 3.4675 32.0025 ;
        RECT  3.2125 33.5775 3.2775 33.6425 ;
        RECT  3.4025 32.7375 3.4675 32.8025 ;
        RECT  3.4025 33.1475 3.4675 33.2125 ;
        RECT  3.2125 34.2625 3.2775 34.3275 ;
        RECT  3.4025 35.1025 3.4675 35.1675 ;
        RECT  3.4025 34.6275 3.4675 34.6925 ;
        RECT  3.2125 36.2675 3.2775 36.3325 ;
        RECT  3.4025 35.4275 3.4675 35.4925 ;
        RECT  3.4025 35.8375 3.4675 35.9025 ;
        RECT  3.2125 36.9525 3.2775 37.0175 ;
        RECT  3.4025 37.7925 3.4675 37.8575 ;
        RECT  3.4025 37.3175 3.4675 37.3825 ;
        RECT  3.2125 38.9575 3.2775 39.0225 ;
        RECT  3.4025 38.1175 3.4675 38.1825 ;
        RECT  3.4025 38.5275 3.4675 38.5925 ;
        RECT  3.2125 39.6425 3.2775 39.7075 ;
        RECT  3.4025 40.4825 3.4675 40.5475 ;
        RECT  3.4025 40.0075 3.4675 40.0725 ;
        RECT  1.5575 8.88 1.6225 8.945 ;
        RECT  1.7325 10.405 1.7975 10.47 ;
        RECT  1.9075 11.57 1.9725 11.635 ;
        RECT  2.0825 13.095 2.1475 13.16 ;
        RECT  2.2575 14.26 2.3225 14.325 ;
        RECT  2.4325 15.785 2.4975 15.85 ;
        RECT  2.6075 16.95 2.6725 17.015 ;
        RECT  2.7825 18.475 2.8475 18.54 ;
        RECT  1.5575 19.6975 1.6225 19.7625 ;
        RECT  2.2575 19.4825 2.3225 19.5475 ;
        RECT  1.5575 21.1075 1.6225 21.1725 ;
        RECT  2.4325 21.3225 2.4975 21.3875 ;
        RECT  1.5575 22.3875 1.6225 22.4525 ;
        RECT  2.6075 22.1725 2.6725 22.2375 ;
        RECT  1.5575 23.7975 1.6225 23.8625 ;
        RECT  2.7825 24.0125 2.8475 24.0775 ;
        RECT  1.7325 25.0775 1.7975 25.1425 ;
        RECT  2.2575 24.8625 2.3225 24.9275 ;
        RECT  1.7325 26.4875 1.7975 26.5525 ;
        RECT  2.4325 26.7025 2.4975 26.7675 ;
        RECT  1.7325 27.7675 1.7975 27.8325 ;
        RECT  2.6075 27.5525 2.6725 27.6175 ;
        RECT  1.7325 29.1775 1.7975 29.2425 ;
        RECT  2.7825 29.3925 2.8475 29.4575 ;
        RECT  1.9075 30.4575 1.9725 30.5225 ;
        RECT  2.2575 30.2425 2.3225 30.3075 ;
        RECT  1.9075 31.8675 1.9725 31.9325 ;
        RECT  2.4325 32.0825 2.4975 32.1475 ;
        RECT  1.9075 33.1475 1.9725 33.2125 ;
        RECT  2.6075 32.9325 2.6725 32.9975 ;
        RECT  1.9075 34.5575 1.9725 34.6225 ;
        RECT  2.7825 34.7725 2.8475 34.8375 ;
        RECT  2.0825 35.8375 2.1475 35.9025 ;
        RECT  2.2575 35.6225 2.3225 35.6875 ;
        RECT  2.0825 37.2475 2.1475 37.3125 ;
        RECT  2.4325 37.4625 2.4975 37.5275 ;
        RECT  2.0825 38.5275 2.1475 38.5925 ;
        RECT  2.6075 38.3125 2.6725 38.3775 ;
        RECT  2.0825 39.9375 2.1475 40.0025 ;
        RECT  2.7825 40.1525 2.8475 40.2175 ;
        RECT  5.7075 20.1275 5.7725 20.1925 ;
        RECT  5.8975 19.2875 5.9625 19.3525 ;
        RECT  5.8975 19.6975 5.9625 19.7625 ;
        RECT  4.6325 19.64 4.6975 19.705 ;
        RECT  4.7725 19.4125 4.8375 19.4775 ;
        RECT  5.6675 19.4825 5.7325 19.5475 ;
        RECT  5.7075 20.8125 5.7725 20.8775 ;
        RECT  5.8975 21.6525 5.9625 21.7175 ;
        RECT  5.8975 21.1775 5.9625 21.2425 ;
        RECT  4.6325 21.165 4.6975 21.23 ;
        RECT  4.7725 21.3925 4.8375 21.4575 ;
        RECT  5.6675 21.3225 5.7325 21.3875 ;
        RECT  5.7075 22.8175 5.7725 22.8825 ;
        RECT  5.8975 21.9775 5.9625 22.0425 ;
        RECT  5.8975 22.3875 5.9625 22.4525 ;
        RECT  4.6325 22.33 4.6975 22.395 ;
        RECT  4.7725 22.1025 4.8375 22.1675 ;
        RECT  5.6675 22.1725 5.7325 22.2375 ;
        RECT  5.7075 23.5025 5.7725 23.5675 ;
        RECT  5.8975 24.3425 5.9625 24.4075 ;
        RECT  5.8975 23.8675 5.9625 23.9325 ;
        RECT  4.6325 23.855 4.6975 23.92 ;
        RECT  4.7725 24.0825 4.8375 24.1475 ;
        RECT  5.6675 24.0125 5.7325 24.0775 ;
        RECT  5.7075 25.5075 5.7725 25.5725 ;
        RECT  5.8975 24.6675 5.9625 24.7325 ;
        RECT  5.8975 25.0775 5.9625 25.1425 ;
        RECT  4.6325 25.02 4.6975 25.085 ;
        RECT  4.7725 24.7925 4.8375 24.8575 ;
        RECT  5.6675 24.8625 5.7325 24.9275 ;
        RECT  5.7075 26.1925 5.7725 26.2575 ;
        RECT  5.8975 27.0325 5.9625 27.0975 ;
        RECT  5.8975 26.5575 5.9625 26.6225 ;
        RECT  4.6325 26.545 4.6975 26.61 ;
        RECT  4.7725 26.7725 4.8375 26.8375 ;
        RECT  5.6675 26.7025 5.7325 26.7675 ;
        RECT  5.7075 28.1975 5.7725 28.2625 ;
        RECT  5.8975 27.3575 5.9625 27.4225 ;
        RECT  5.8975 27.7675 5.9625 27.8325 ;
        RECT  4.6325 27.71 4.6975 27.775 ;
        RECT  4.7725 27.4825 4.8375 27.5475 ;
        RECT  5.6675 27.5525 5.7325 27.6175 ;
        RECT  5.7075 28.8825 5.7725 28.9475 ;
        RECT  5.8975 29.7225 5.9625 29.7875 ;
        RECT  5.8975 29.2475 5.9625 29.3125 ;
        RECT  4.6325 29.235 4.6975 29.3 ;
        RECT  4.7725 29.4625 4.8375 29.5275 ;
        RECT  5.6675 29.3925 5.7325 29.4575 ;
        RECT  5.7075 30.8875 5.7725 30.9525 ;
        RECT  5.8975 30.0475 5.9625 30.1125 ;
        RECT  5.8975 30.4575 5.9625 30.5225 ;
        RECT  4.6325 30.4 4.6975 30.465 ;
        RECT  4.7725 30.1725 4.8375 30.2375 ;
        RECT  5.6675 30.2425 5.7325 30.3075 ;
        RECT  5.7075 31.5725 5.7725 31.6375 ;
        RECT  5.8975 32.4125 5.9625 32.4775 ;
        RECT  5.8975 31.9375 5.9625 32.0025 ;
        RECT  4.6325 31.925 4.6975 31.99 ;
        RECT  4.7725 32.1525 4.8375 32.2175 ;
        RECT  5.6675 32.0825 5.7325 32.1475 ;
        RECT  5.7075 33.5775 5.7725 33.6425 ;
        RECT  5.8975 32.7375 5.9625 32.8025 ;
        RECT  5.8975 33.1475 5.9625 33.2125 ;
        RECT  4.6325 33.09 4.6975 33.155 ;
        RECT  4.7725 32.8625 4.8375 32.9275 ;
        RECT  5.6675 32.9325 5.7325 32.9975 ;
        RECT  5.7075 34.2625 5.7725 34.3275 ;
        RECT  5.8975 35.1025 5.9625 35.1675 ;
        RECT  5.8975 34.6275 5.9625 34.6925 ;
        RECT  4.6325 34.615 4.6975 34.68 ;
        RECT  4.7725 34.8425 4.8375 34.9075 ;
        RECT  5.6675 34.7725 5.7325 34.8375 ;
        RECT  5.7075 36.2675 5.7725 36.3325 ;
        RECT  5.8975 35.4275 5.9625 35.4925 ;
        RECT  5.8975 35.8375 5.9625 35.9025 ;
        RECT  4.6325 35.78 4.6975 35.845 ;
        RECT  4.7725 35.5525 4.8375 35.6175 ;
        RECT  5.6675 35.6225 5.7325 35.6875 ;
        RECT  5.7075 36.9525 5.7725 37.0175 ;
        RECT  5.8975 37.7925 5.9625 37.8575 ;
        RECT  5.8975 37.3175 5.9625 37.3825 ;
        RECT  4.6325 37.305 4.6975 37.37 ;
        RECT  4.7725 37.5325 4.8375 37.5975 ;
        RECT  5.6675 37.4625 5.7325 37.5275 ;
        RECT  5.7075 38.9575 5.7725 39.0225 ;
        RECT  5.8975 38.1175 5.9625 38.1825 ;
        RECT  5.8975 38.5275 5.9625 38.5925 ;
        RECT  4.6325 38.47 4.6975 38.535 ;
        RECT  4.7725 38.2425 4.8375 38.3075 ;
        RECT  5.6675 38.3125 5.7325 38.3775 ;
        RECT  5.7075 39.6425 5.7725 39.7075 ;
        RECT  5.8975 40.4825 5.9625 40.5475 ;
        RECT  5.8975 40.0075 5.9625 40.0725 ;
        RECT  4.6325 39.995 4.6975 40.06 ;
        RECT  4.7725 40.2225 4.8375 40.2875 ;
        RECT  5.6675 40.1525 5.7325 40.2175 ;
        RECT  6.2175 7.69 6.2825 7.755 ;
        RECT  1.04 7.1825 1.105 7.2475 ;
        RECT  5.1225 7.325 5.1875 7.39 ;
        RECT  3.515 7.3225 3.58 7.3875 ;
        RECT  2.1175 7.3225 2.1825 7.3875 ;
        RECT  0.9 7.8875 0.965 7.9525 ;
        RECT  3.9775 7.1825 4.0425 7.2475 ;
        RECT  2.7825 7.6875 2.8475 7.7525 ;
        RECT  6.475 7.3225 6.54 7.3875 ;
        RECT  5.965 7.5 6.03 7.565 ;
        RECT  5.5525 7.1825 5.6175 7.2475 ;
        RECT  0.85 7.1825 0.915 7.2475 ;
        RECT  2.5925 7.1825 2.6575 7.2475 ;
        RECT  2.3925 7.6875 2.4575 7.7525 ;
        RECT  2.3925 7.5 2.4575 7.565 ;
        RECT  3.005 7.5 3.07 7.565 ;
        RECT  5.3525 7.69 5.4175 7.755 ;
        RECT  5.3525 7.5 5.4175 7.565 ;
        RECT  6.2175 6.675 6.2825 6.74 ;
        RECT  1.04 7.1825 1.105 7.2475 ;
        RECT  5.1225 7.04 5.1875 7.105 ;
        RECT  3.515 7.0425 3.58 7.1075 ;
        RECT  2.1175 7.0425 2.1825 7.1075 ;
        RECT  0.9 6.4775 0.965 6.5425 ;
        RECT  3.9775 7.1825 4.0425 7.2475 ;
        RECT  2.7825 6.6775 2.8475 6.7425 ;
        RECT  6.475 7.0425 6.54 7.1075 ;
        RECT  5.965 6.865 6.03 6.93 ;
        RECT  5.5525 7.1825 5.6175 7.2475 ;
        RECT  0.85 7.1825 0.915 7.2475 ;
        RECT  2.5925 7.1825 2.6575 7.2475 ;
        RECT  2.3925 6.6775 2.4575 6.7425 ;
        RECT  2.3925 6.865 2.4575 6.93 ;
        RECT  3.005 6.865 3.07 6.93 ;
        RECT  5.3525 6.675 5.4175 6.74 ;
        RECT  5.3525 6.865 5.4175 6.93 ;
        RECT  6.2175 6.28 6.2825 6.345 ;
        RECT  1.04 5.7725 1.105 5.8375 ;
        RECT  5.1225 5.915 5.1875 5.98 ;
        RECT  3.515 5.9125 3.58 5.9775 ;
        RECT  2.1175 5.9125 2.1825 5.9775 ;
        RECT  0.9 6.4775 0.965 6.5425 ;
        RECT  3.9775 5.7725 4.0425 5.8375 ;
        RECT  2.7825 6.2775 2.8475 6.3425 ;
        RECT  6.475 5.9125 6.54 5.9775 ;
        RECT  5.965 6.09 6.03 6.155 ;
        RECT  5.5525 5.7725 5.6175 5.8375 ;
        RECT  0.85 5.7725 0.915 5.8375 ;
        RECT  2.5925 5.7725 2.6575 5.8375 ;
        RECT  2.3925 6.2775 2.4575 6.3425 ;
        RECT  2.3925 6.09 2.4575 6.155 ;
        RECT  3.005 6.09 3.07 6.155 ;
        RECT  5.3525 6.28 5.4175 6.345 ;
        RECT  5.3525 6.09 5.4175 6.155 ;
        RECT  6.2175 5.265 6.2825 5.33 ;
        RECT  1.04 5.7725 1.105 5.8375 ;
        RECT  5.1225 5.63 5.1875 5.695 ;
        RECT  3.515 5.6325 3.58 5.6975 ;
        RECT  2.1175 5.6325 2.1825 5.6975 ;
        RECT  0.9 5.0675 0.965 5.1325 ;
        RECT  3.9775 5.7725 4.0425 5.8375 ;
        RECT  2.7825 5.2675 2.8475 5.3325 ;
        RECT  6.475 5.6325 6.54 5.6975 ;
        RECT  5.965 5.455 6.03 5.52 ;
        RECT  5.5525 5.7725 5.6175 5.8375 ;
        RECT  0.85 5.7725 0.915 5.8375 ;
        RECT  2.5925 5.7725 2.6575 5.8375 ;
        RECT  2.3925 5.2675 2.4575 5.3325 ;
        RECT  2.3925 5.455 2.4575 5.52 ;
        RECT  3.005 5.455 3.07 5.52 ;
        RECT  5.3525 5.265 5.4175 5.33 ;
        RECT  5.3525 5.455 5.4175 5.52 ;
        RECT  8.2875 19.0575 8.3525 19.1225 ;
        RECT  8.2875 21.7475 8.3525 21.8125 ;
        RECT  8.2875 24.4375 8.3525 24.5025 ;
        RECT  8.2875 27.1275 8.3525 27.1925 ;
        RECT  8.2875 29.8175 8.3525 29.8825 ;
        RECT  8.2875 32.5075 8.3525 32.5725 ;
        RECT  8.2875 35.1975 8.3525 35.2625 ;
        RECT  8.2875 37.8875 8.3525 37.9525 ;
        RECT  8.2875 40.5775 8.3525 40.6425 ;
        RECT  6.82 8.5025 6.885 8.5675 ;
        RECT  7.23 8.5025 7.295 8.5675 ;
        RECT  6.545 9.8475 6.61 9.9125 ;
        RECT  7.435 9.8475 7.5 9.9125 ;
        RECT  6.82 13.8825 6.885 13.9475 ;
        RECT  7.64 13.8825 7.705 13.9475 ;
        RECT  6.545 15.2275 6.61 15.2925 ;
        RECT  7.845 15.2275 7.91 15.2925 ;
        RECT  7.025 8.2975 7.09 8.3625 ;
        RECT  7.025 10.9875 7.09 11.0525 ;
        RECT  7.025 13.6775 7.09 13.7425 ;
        RECT  7.025 16.3675 7.09 16.4325 ;
        RECT  6.8875 7.535 6.9525 7.6 ;
        RECT  7.23 7.535 7.295 7.6 ;
        RECT  6.8875 6.83 6.9525 6.895 ;
        RECT  7.435 6.83 7.5 6.895 ;
        RECT  6.8875 6.125 6.9525 6.19 ;
        RECT  7.64 6.125 7.705 6.19 ;
        RECT  6.8875 5.42 6.9525 5.485 ;
        RECT  7.845 5.42 7.91 5.485 ;
        RECT  6.955 7.8875 7.02 7.9525 ;
        RECT  8.2875 7.8875 8.3525 7.9525 ;
        RECT  6.955 7.1825 7.02 7.2475 ;
        RECT  8.2875 7.1825 8.3525 7.2475 ;
        RECT  6.955 6.4775 7.02 6.5425 ;
        RECT  8.2875 6.4775 8.3525 6.5425 ;
        RECT  6.955 5.7725 7.02 5.8375 ;
        RECT  8.2875 5.7725 8.3525 5.8375 ;
        RECT  6.955 5.0675 7.02 5.1325 ;
        RECT  8.2875 5.0675 8.3525 5.1325 ;
        RECT  9.425 3.795 9.49 3.86 ;
        RECT  9.015 1.61 9.08 1.675 ;
        RECT  9.22 3.1575 9.285 3.2225 ;
        RECT  9.425 41.4775 9.49 41.5425 ;
        RECT  9.63 10.2975 9.695 10.3625 ;
        RECT  9.835 14.3225 9.9 14.3875 ;
        RECT  8.81 8.0925 8.875 8.1575 ;
        RECT  4.6325 40.7825 4.6975 40.8475 ;
        RECT  8.81 40.7825 8.875 40.8475 ;
        RECT  8.5025 3.0275 8.5675 3.0925 ;
        RECT  8.5025 14.4525 8.5675 14.5175 ;
        RECT  8.5025 3.955 8.5675 4.02 ;
        RECT  8.5025 11.23 8.5675 11.295 ;
        RECT  -3.845 24.9675 -3.78 25.0325 ;
        RECT  -3.3375 19.79 -3.2725 19.855 ;
        RECT  -3.48 23.8725 -3.415 23.9375 ;
        RECT  -3.4775 22.265 -3.4125 22.33 ;
        RECT  -3.4775 20.8675 -3.4125 20.9325 ;
        RECT  -4.0425 19.65 -3.9775 19.715 ;
        RECT  -3.3375 22.7275 -3.2725 22.7925 ;
        RECT  -3.8425 21.5325 -3.7775 21.5975 ;
        RECT  -3.4775 25.225 -3.4125 25.29 ;
        RECT  -3.655 24.715 -3.59 24.78 ;
        RECT  -3.3375 24.3025 -3.2725 24.3675 ;
        RECT  -3.3375 19.6 -3.2725 19.665 ;
        RECT  -3.3375 21.3425 -3.2725 21.4075 ;
        RECT  -3.8425 21.1425 -3.7775 21.2075 ;
        RECT  -3.655 21.1425 -3.59 21.2075 ;
        RECT  -3.655 21.755 -3.59 21.82 ;
        RECT  -3.845 24.1025 -3.78 24.1675 ;
        RECT  -3.655 24.1025 -3.59 24.1675 ;
        RECT  -2.83 24.9675 -2.765 25.0325 ;
        RECT  -3.3375 19.79 -3.2725 19.855 ;
        RECT  -3.195 23.8725 -3.13 23.9375 ;
        RECT  -3.1975 22.265 -3.1325 22.33 ;
        RECT  -3.1975 20.8675 -3.1325 20.9325 ;
        RECT  -2.6325 19.65 -2.5675 19.715 ;
        RECT  -3.3375 22.7275 -3.2725 22.7925 ;
        RECT  -2.8325 21.5325 -2.7675 21.5975 ;
        RECT  -3.1975 25.225 -3.1325 25.29 ;
        RECT  -3.02 24.715 -2.955 24.78 ;
        RECT  -3.3375 24.3025 -3.2725 24.3675 ;
        RECT  -3.3375 19.6 -3.2725 19.665 ;
        RECT  -3.3375 21.3425 -3.2725 21.4075 ;
        RECT  -2.8325 21.1425 -2.7675 21.2075 ;
        RECT  -3.02 21.1425 -2.955 21.2075 ;
        RECT  -3.02 21.755 -2.955 21.82 ;
        RECT  -2.83 24.1025 -2.765 24.1675 ;
        RECT  -3.02 24.1025 -2.955 24.1675 ;
        RECT  -2.435 24.9675 -2.37 25.0325 ;
        RECT  -1.9275 19.79 -1.8625 19.855 ;
        RECT  -2.07 23.8725 -2.005 23.9375 ;
        RECT  -2.0675 22.265 -2.0025 22.33 ;
        RECT  -2.0675 20.8675 -2.0025 20.9325 ;
        RECT  -2.6325 19.65 -2.5675 19.715 ;
        RECT  -1.9275 22.7275 -1.8625 22.7925 ;
        RECT  -2.4325 21.5325 -2.3675 21.5975 ;
        RECT  -2.0675 25.225 -2.0025 25.29 ;
        RECT  -2.245 24.715 -2.18 24.78 ;
        RECT  -1.9275 24.3025 -1.8625 24.3675 ;
        RECT  -1.9275 19.6 -1.8625 19.665 ;
        RECT  -1.9275 21.3425 -1.8625 21.4075 ;
        RECT  -2.4325 21.1425 -2.3675 21.2075 ;
        RECT  -2.245 21.1425 -2.18 21.2075 ;
        RECT  -2.245 21.755 -2.18 21.82 ;
        RECT  -2.435 24.1025 -2.37 24.1675 ;
        RECT  -2.245 24.1025 -2.18 24.1675 ;
        RECT  -1.2425 28.1825 -1.1775 28.2475 ;
        RECT  -1.2425 28.5625 -1.1775 28.6275 ;
        RECT  -0.4475 28.5625 -0.3825 28.6275 ;
        RECT  -0.95 28.5625 -0.885 28.6275 ;
        RECT  -1.995 28.3725 -1.93 28.4375 ;
        RECT  -2.7475 28.1825 -2.6825 28.2475 ;
        RECT  -2.3475 28.4425 -2.2825 28.5075 ;
        RECT  -1.9275 29.3275 -1.8625 29.3925 ;
        RECT  -2.7675 29.5175 -2.7025 29.5825 ;
        RECT  -2.2925 29.5175 -2.2275 29.5825 ;
        RECT  -3.9325 28.7425 -3.8675 28.8075 ;
        RECT  -3.9325 29.1225 -3.8675 29.1875 ;
        RECT  -3.1375 29.1225 -3.0725 29.1875 ;
        RECT  -3.64 29.1225 -3.575 29.1875 ;
        RECT  -0.755 33.385 -0.69 33.45 ;
        RECT  -2.28 33.14 -2.215 33.205 ;
        RECT  -2.28 33.7 -2.215 33.765 ;
        RECT  -0.755 33.78 -0.69 33.845 ;
        RECT  -0.755 33.22 -0.69 33.285 ;
        RECT  -2.28 33.305 -2.215 33.37 ;
        RECT  -3.2725 34.0975 -3.2075 34.1625 ;
        RECT  -3.9775 34.5725 -3.9125 34.6375 ;
        RECT  -3.2725 34.5725 -3.2075 34.6375 ;
        RECT  -3.725 34.0925 -3.66 34.1575 ;
        RECT  -3.525 34.0975 -3.46 34.1625 ;
        RECT  -3.9775 33.7675 -3.9125 33.8325 ;
        RECT  -3.2725 33.7675 -3.2075 33.8325 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.2725 33.7675 -3.2075 33.8325 ;
        RECT  -3.9775 33.7675 -3.9125 33.8325 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.5275 33.4425 -3.4625 33.5075 ;
        RECT  -3.2725 32.95 -3.2075 33.015 ;
        RECT  -3.2725 32.95 -3.2075 33.015 ;
        RECT  -3.2725 32.95 -3.2075 33.015 ;
        RECT  -3.2725 32.95 -3.2075 33.015 ;
        RECT  -3.2725 32.95 -3.2075 33.015 ;
        RECT  -3.2725 32.95 -3.2075 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.7225 33.4425 -3.6575 33.5075 ;
        RECT  -3.9775 33.7675 -3.9125 33.8325 ;
        RECT  -3.9775 33.7675 -3.9125 33.8325 ;
        RECT  -3.9775 33.7675 -3.9125 33.8325 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.9775 32.95 -3.9125 33.015 ;
        RECT  -3.2725 33.7675 -3.2075 33.8325 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.2725 31.0775 -3.2075 31.1425 ;
        RECT  -3.9775 31.0775 -3.9125 31.1425 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.5275 31.4025 -3.4625 31.4675 ;
        RECT  -3.2725 31.895 -3.2075 31.96 ;
        RECT  -3.2725 31.895 -3.2075 31.96 ;
        RECT  -3.2725 31.895 -3.2075 31.96 ;
        RECT  -3.2725 31.895 -3.2075 31.96 ;
        RECT  -3.2725 31.895 -3.2075 31.96 ;
        RECT  -3.2725 31.895 -3.2075 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.7225 31.4025 -3.6575 31.4675 ;
        RECT  -3.9775 31.0775 -3.9125 31.1425 ;
        RECT  -3.9775 31.0775 -3.9125 31.1425 ;
        RECT  -3.9775 31.0775 -3.9125 31.1425 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.9775 31.895 -3.9125 31.96 ;
        RECT  -3.2725 31.0775 -3.2075 31.1425 ;
        RECT  -2.8625 33.8075 -2.7975 33.8725 ;
        RECT  -2.8625 36.2175 -2.7975 36.2825 ;
        RECT  -2.8625 34.035 -2.7975 34.1 ;
        RECT  -2.8625 31.66 -2.7975 31.725 ;
        RECT  -2.8625 36.6925 -2.7975 36.7575 ;
        RECT  -3.2725 36.6925 -3.2075 36.7575 ;
        RECT  -3.035 32.5575 -2.97 32.6225 ;
        RECT  -3.035 31.96 -2.97 32.025 ;
        RECT  -3.4575 31.96 -3.3925 32.025 ;
        RECT  -0.725 26.0825 -0.66 26.1475 ;
        RECT  -0.725 22.0025 -0.66 22.0675 ;
        RECT  -1.7225 19.435 -1.6575 19.5 ;
        RECT  -2.2775 26.0825 -2.2125 26.1475 ;
        RECT  -2.4925 26.4925 -2.4275 26.5575 ;
        RECT  -2.2225 29.03 -2.1575 29.095 ;
        RECT  -2.4375 29.2875 -2.3725 29.3525 ;
        RECT  -0.95 27.5175 -0.885 27.5825 ;
        RECT  -0.81 27.3125 -0.745 27.3775 ;
        RECT  -0.67 26.6975 -0.605 26.7625 ;
        RECT  -3.64 27.5175 -3.575 27.5825 ;
        RECT  -3.5 26.6975 -3.435 26.7625 ;
        RECT  -3.36 26.9025 -3.295 26.9675 ;
        RECT  -2.2775 28.8125 -2.2125 28.8775 ;
        RECT  -2.2225 29.9575 -2.1575 30.0225 ;
        RECT  -3.445 31.1425 -3.38 31.2075 ;
        RECT  -2.28 30.1825 -2.215 30.2475 ;
        RECT  -0.1725 26.2875 -0.1075 26.3525 ;
        RECT  -1.5175 27.1075 -1.4525 27.1725 ;
        RECT  -2.8625 26.2875 -2.7975 26.3525 ;
        RECT  -4.2075 27.1075 -4.1425 27.1725 ;
        RECT  0.1425 27.1075 0.2075 27.1725 ;
        LAYER  metal2 ;
        RECT  9.8325 30.01 9.9025 30.215 ;
        RECT  9.6275 30.97 9.6975 31.175 ;
        RECT  9.2175 28.64 9.2875 28.845 ;
        RECT  9.0125 29.785 9.0825 29.99 ;
        RECT  9.4225 27.345 9.4925 27.55 ;
        RECT  8.8075 25.91 8.8775 26.115 ;
        RECT  -0.14 27.105 0.175 27.175 ;
        RECT  8.3925 26.115 8.4625 26.32 ;
        RECT  10.6625 0.0 10.7325 0.14 ;
        RECT  11.3675 0.0 11.4375 0.14 ;
        RECT  8.2525 0.0 8.6025 42.27 ;
        RECT  8.8075 0.0 8.8775 42.27 ;
        RECT  9.0125 0.0 9.0825 42.27 ;
        RECT  9.2175 0.0 9.2875 42.27 ;
        RECT  9.4225 0.0 9.4925 42.27 ;
        RECT  9.6275 0.0 9.6975 42.27 ;
        RECT  9.8325 0.0 9.9025 42.27 ;
        RECT  7.2275 4.69 7.2975 19.09 ;
        RECT  7.4325 4.69 7.5025 19.09 ;
        RECT  7.6375 4.69 7.7075 19.09 ;
        RECT  7.8425 4.69 7.9125 19.09 ;
        RECT  10.495 40.71 10.565 41.06 ;
        RECT  10.83 40.71 10.9 41.06 ;
        RECT  11.2 40.71 11.27 41.06 ;
        RECT  11.535 40.71 11.605 41.06 ;
        RECT  10.6625 0.44 10.7325 0.51 ;
        RECT  10.4875 0.44 10.6975 0.51 ;
        RECT  10.6625 0.475 10.7325 0.615 ;
        RECT  11.3675 0.44 11.4375 0.51 ;
        RECT  11.1925 0.44 11.4025 0.51 ;
        RECT  11.3675 0.475 11.4375 0.615 ;
        RECT  4.63 40.61 4.7 40.815 ;
        RECT  10.6625 0.0 10.7325 0.14 ;
        RECT  11.3675 0.0 11.4375 0.14 ;
        RECT  9.6275 0.0 9.6975 42.27 ;
        RECT  9.4225 0.0 9.4925 42.27 ;
        RECT  8.8075 0.0 8.8775 42.27 ;
        RECT  9.8325 0.0 9.9025 42.27 ;
        RECT  9.0125 0.0 9.0825 42.27 ;
        RECT  8.2525 0.0 8.6025 42.27 ;
        RECT  9.2175 0.0 9.2875 42.27 ;
        RECT  10.83 18.99 10.9 40.71 ;
        RECT  11.2 18.99 11.27 40.71 ;
        RECT  11.535 18.99 11.605 40.71 ;
        RECT  10.495 18.99 10.565 40.71 ;
        RECT  10.31 18.99 10.38 40.71 ;
        RECT  11.015 18.99 11.085 40.71 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  10.2775 19.055 10.4125 19.125 ;
        RECT  10.9825 19.055 11.1175 19.125 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  10.565 19.3475 10.635 19.4825 ;
        RECT  10.31 19.84 10.38 19.975 ;
        RECT  10.31 19.84 10.38 19.975 ;
        RECT  10.31 19.84 10.38 19.975 ;
        RECT  10.31 19.84 10.38 19.975 ;
        RECT  10.31 19.84 10.38 19.975 ;
        RECT  10.31 19.84 10.38 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  10.76 19.3475 10.83 19.4825 ;
        RECT  10.9825 19.055 11.1175 19.125 ;
        RECT  10.9825 19.055 11.1175 19.125 ;
        RECT  10.9825 19.055 11.1175 19.125 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  10.2775 19.055 10.4125 19.125 ;
        RECT  11.015 19.0575 11.085 20.4675 ;
        RECT  10.315 19.06 10.375 19.1175 ;
        RECT  10.5025 19.065 10.5575 19.1175 ;
        RECT  10.8375 19.0575 10.895 19.1175 ;
        RECT  11.02 19.065 11.08 19.1225 ;
        RECT  10.83 18.99 10.9 20.535 ;
        RECT  10.495 18.99 10.565 20.535 ;
        RECT  10.31 18.99 10.38 20.535 ;
        RECT  11.015 18.99 11.085 20.535 ;
        RECT  10.495 18.99 10.565 20.535 ;
        RECT  10.31 18.99 10.38 20.535 ;
        RECT  11.015 18.99 11.085 20.535 ;
        RECT  10.83 18.99 10.9 20.535 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  10.2775 21.745 10.4125 21.815 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  10.565 21.3875 10.635 21.5225 ;
        RECT  10.31 20.895 10.38 21.03 ;
        RECT  10.31 20.895 10.38 21.03 ;
        RECT  10.31 20.895 10.38 21.03 ;
        RECT  10.31 20.895 10.38 21.03 ;
        RECT  10.31 20.895 10.38 21.03 ;
        RECT  10.31 20.895 10.38 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  10.76 21.3875 10.83 21.5225 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  10.2775 21.745 10.4125 21.815 ;
        RECT  11.015 20.4025 11.085 21.8125 ;
        RECT  10.315 21.7525 10.375 21.81 ;
        RECT  10.5025 21.7525 10.5575 21.805 ;
        RECT  10.8375 21.7525 10.895 21.8125 ;
        RECT  11.02 21.7475 11.08 21.805 ;
        RECT  10.83 20.335 10.9 21.88 ;
        RECT  10.495 20.335 10.565 21.88 ;
        RECT  10.31 20.335 10.38 21.88 ;
        RECT  11.015 20.335 11.085 21.88 ;
        RECT  10.495 20.335 10.565 21.88 ;
        RECT  10.31 20.335 10.38 21.88 ;
        RECT  11.015 20.335 11.085 21.88 ;
        RECT  10.83 20.335 10.9 21.88 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  10.2775 21.745 10.4125 21.815 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  10.565 22.0375 10.635 22.1725 ;
        RECT  10.31 22.53 10.38 22.665 ;
        RECT  10.31 22.53 10.38 22.665 ;
        RECT  10.31 22.53 10.38 22.665 ;
        RECT  10.31 22.53 10.38 22.665 ;
        RECT  10.31 22.53 10.38 22.665 ;
        RECT  10.31 22.53 10.38 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  10.76 22.0375 10.83 22.1725 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  10.2775 21.745 10.4125 21.815 ;
        RECT  11.015 21.7475 11.085 23.1575 ;
        RECT  10.315 21.75 10.375 21.8075 ;
        RECT  10.5025 21.755 10.5575 21.8075 ;
        RECT  10.8375 21.7475 10.895 21.8075 ;
        RECT  11.02 21.755 11.08 21.8125 ;
        RECT  10.83 21.68 10.9 23.225 ;
        RECT  10.495 21.68 10.565 23.225 ;
        RECT  10.31 21.68 10.38 23.225 ;
        RECT  11.015 21.68 11.085 23.225 ;
        RECT  10.495 21.68 10.565 23.225 ;
        RECT  10.31 21.68 10.38 23.225 ;
        RECT  11.015 21.68 11.085 23.225 ;
        RECT  10.83 21.68 10.9 23.225 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  10.2775 24.435 10.4125 24.505 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  10.565 24.0775 10.635 24.2125 ;
        RECT  10.31 23.585 10.38 23.72 ;
        RECT  10.31 23.585 10.38 23.72 ;
        RECT  10.31 23.585 10.38 23.72 ;
        RECT  10.31 23.585 10.38 23.72 ;
        RECT  10.31 23.585 10.38 23.72 ;
        RECT  10.31 23.585 10.38 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  10.76 24.0775 10.83 24.2125 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  10.2775 24.435 10.4125 24.505 ;
        RECT  11.015 23.0925 11.085 24.5025 ;
        RECT  10.315 24.4425 10.375 24.5 ;
        RECT  10.5025 24.4425 10.5575 24.495 ;
        RECT  10.8375 24.4425 10.895 24.5025 ;
        RECT  11.02 24.4375 11.08 24.495 ;
        RECT  10.83 23.025 10.9 24.57 ;
        RECT  10.495 23.025 10.565 24.57 ;
        RECT  10.31 23.025 10.38 24.57 ;
        RECT  11.015 23.025 11.085 24.57 ;
        RECT  10.495 23.025 10.565 24.57 ;
        RECT  10.31 23.025 10.38 24.57 ;
        RECT  11.015 23.025 11.085 24.57 ;
        RECT  10.83 23.025 10.9 24.57 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  10.2775 24.435 10.4125 24.505 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  10.565 24.7275 10.635 24.8625 ;
        RECT  10.31 25.22 10.38 25.355 ;
        RECT  10.31 25.22 10.38 25.355 ;
        RECT  10.31 25.22 10.38 25.355 ;
        RECT  10.31 25.22 10.38 25.355 ;
        RECT  10.31 25.22 10.38 25.355 ;
        RECT  10.31 25.22 10.38 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  10.76 24.7275 10.83 24.8625 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  10.2775 24.435 10.4125 24.505 ;
        RECT  11.015 24.4375 11.085 25.8475 ;
        RECT  10.315 24.44 10.375 24.4975 ;
        RECT  10.5025 24.445 10.5575 24.4975 ;
        RECT  10.8375 24.4375 10.895 24.4975 ;
        RECT  11.02 24.445 11.08 24.5025 ;
        RECT  10.83 24.37 10.9 25.915 ;
        RECT  10.495 24.37 10.565 25.915 ;
        RECT  10.31 24.37 10.38 25.915 ;
        RECT  11.015 24.37 11.085 25.915 ;
        RECT  10.495 24.37 10.565 25.915 ;
        RECT  10.31 24.37 10.38 25.915 ;
        RECT  11.015 24.37 11.085 25.915 ;
        RECT  10.83 24.37 10.9 25.915 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  10.2775 27.125 10.4125 27.195 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  10.565 26.7675 10.635 26.9025 ;
        RECT  10.31 26.275 10.38 26.41 ;
        RECT  10.31 26.275 10.38 26.41 ;
        RECT  10.31 26.275 10.38 26.41 ;
        RECT  10.31 26.275 10.38 26.41 ;
        RECT  10.31 26.275 10.38 26.41 ;
        RECT  10.31 26.275 10.38 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  10.76 26.7675 10.83 26.9025 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  10.2775 27.125 10.4125 27.195 ;
        RECT  11.015 25.7825 11.085 27.1925 ;
        RECT  10.315 27.1325 10.375 27.19 ;
        RECT  10.5025 27.1325 10.5575 27.185 ;
        RECT  10.8375 27.1325 10.895 27.1925 ;
        RECT  11.02 27.1275 11.08 27.185 ;
        RECT  10.83 25.715 10.9 27.26 ;
        RECT  10.495 25.715 10.565 27.26 ;
        RECT  10.31 25.715 10.38 27.26 ;
        RECT  11.015 25.715 11.085 27.26 ;
        RECT  10.495 25.715 10.565 27.26 ;
        RECT  10.31 25.715 10.38 27.26 ;
        RECT  11.015 25.715 11.085 27.26 ;
        RECT  10.83 25.715 10.9 27.26 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  10.2775 27.125 10.4125 27.195 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  10.565 27.4175 10.635 27.5525 ;
        RECT  10.31 27.91 10.38 28.045 ;
        RECT  10.31 27.91 10.38 28.045 ;
        RECT  10.31 27.91 10.38 28.045 ;
        RECT  10.31 27.91 10.38 28.045 ;
        RECT  10.31 27.91 10.38 28.045 ;
        RECT  10.31 27.91 10.38 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  10.76 27.4175 10.83 27.5525 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  10.2775 27.125 10.4125 27.195 ;
        RECT  11.015 27.1275 11.085 28.5375 ;
        RECT  10.315 27.13 10.375 27.1875 ;
        RECT  10.5025 27.135 10.5575 27.1875 ;
        RECT  10.8375 27.1275 10.895 27.1875 ;
        RECT  11.02 27.135 11.08 27.1925 ;
        RECT  10.83 27.06 10.9 28.605 ;
        RECT  10.495 27.06 10.565 28.605 ;
        RECT  10.31 27.06 10.38 28.605 ;
        RECT  11.015 27.06 11.085 28.605 ;
        RECT  10.495 27.06 10.565 28.605 ;
        RECT  10.31 27.06 10.38 28.605 ;
        RECT  11.015 27.06 11.085 28.605 ;
        RECT  10.83 27.06 10.9 28.605 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  10.2775 29.815 10.4125 29.885 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  10.565 29.4575 10.635 29.5925 ;
        RECT  10.31 28.965 10.38 29.1 ;
        RECT  10.31 28.965 10.38 29.1 ;
        RECT  10.31 28.965 10.38 29.1 ;
        RECT  10.31 28.965 10.38 29.1 ;
        RECT  10.31 28.965 10.38 29.1 ;
        RECT  10.31 28.965 10.38 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  10.76 29.4575 10.83 29.5925 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  10.2775 29.815 10.4125 29.885 ;
        RECT  11.015 28.4725 11.085 29.8825 ;
        RECT  10.315 29.8225 10.375 29.88 ;
        RECT  10.5025 29.8225 10.5575 29.875 ;
        RECT  10.8375 29.8225 10.895 29.8825 ;
        RECT  11.02 29.8175 11.08 29.875 ;
        RECT  10.83 28.405 10.9 29.95 ;
        RECT  10.495 28.405 10.565 29.95 ;
        RECT  10.31 28.405 10.38 29.95 ;
        RECT  11.015 28.405 11.085 29.95 ;
        RECT  10.495 28.405 10.565 29.95 ;
        RECT  10.31 28.405 10.38 29.95 ;
        RECT  11.015 28.405 11.085 29.95 ;
        RECT  10.83 28.405 10.9 29.95 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  10.2775 29.815 10.4125 29.885 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  10.565 30.1075 10.635 30.2425 ;
        RECT  10.31 30.6 10.38 30.735 ;
        RECT  10.31 30.6 10.38 30.735 ;
        RECT  10.31 30.6 10.38 30.735 ;
        RECT  10.31 30.6 10.38 30.735 ;
        RECT  10.31 30.6 10.38 30.735 ;
        RECT  10.31 30.6 10.38 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  10.76 30.1075 10.83 30.2425 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  10.2775 29.815 10.4125 29.885 ;
        RECT  11.015 29.8175 11.085 31.2275 ;
        RECT  10.315 29.82 10.375 29.8775 ;
        RECT  10.5025 29.825 10.5575 29.8775 ;
        RECT  10.8375 29.8175 10.895 29.8775 ;
        RECT  11.02 29.825 11.08 29.8825 ;
        RECT  10.83 29.75 10.9 31.295 ;
        RECT  10.495 29.75 10.565 31.295 ;
        RECT  10.31 29.75 10.38 31.295 ;
        RECT  11.015 29.75 11.085 31.295 ;
        RECT  10.495 29.75 10.565 31.295 ;
        RECT  10.31 29.75 10.38 31.295 ;
        RECT  11.015 29.75 11.085 31.295 ;
        RECT  10.83 29.75 10.9 31.295 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  10.2775 32.505 10.4125 32.575 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  10.565 32.1475 10.635 32.2825 ;
        RECT  10.31 31.655 10.38 31.79 ;
        RECT  10.31 31.655 10.38 31.79 ;
        RECT  10.31 31.655 10.38 31.79 ;
        RECT  10.31 31.655 10.38 31.79 ;
        RECT  10.31 31.655 10.38 31.79 ;
        RECT  10.31 31.655 10.38 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  10.76 32.1475 10.83 32.2825 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  10.2775 32.505 10.4125 32.575 ;
        RECT  11.015 31.1625 11.085 32.5725 ;
        RECT  10.315 32.5125 10.375 32.57 ;
        RECT  10.5025 32.5125 10.5575 32.565 ;
        RECT  10.8375 32.5125 10.895 32.5725 ;
        RECT  11.02 32.5075 11.08 32.565 ;
        RECT  10.83 31.095 10.9 32.64 ;
        RECT  10.495 31.095 10.565 32.64 ;
        RECT  10.31 31.095 10.38 32.64 ;
        RECT  11.015 31.095 11.085 32.64 ;
        RECT  10.495 31.095 10.565 32.64 ;
        RECT  10.31 31.095 10.38 32.64 ;
        RECT  11.015 31.095 11.085 32.64 ;
        RECT  10.83 31.095 10.9 32.64 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  10.2775 32.505 10.4125 32.575 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  10.565 32.7975 10.635 32.9325 ;
        RECT  10.31 33.29 10.38 33.425 ;
        RECT  10.31 33.29 10.38 33.425 ;
        RECT  10.31 33.29 10.38 33.425 ;
        RECT  10.31 33.29 10.38 33.425 ;
        RECT  10.31 33.29 10.38 33.425 ;
        RECT  10.31 33.29 10.38 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  10.76 32.7975 10.83 32.9325 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  10.2775 32.505 10.4125 32.575 ;
        RECT  11.015 32.5075 11.085 33.9175 ;
        RECT  10.315 32.51 10.375 32.5675 ;
        RECT  10.5025 32.515 10.5575 32.5675 ;
        RECT  10.8375 32.5075 10.895 32.5675 ;
        RECT  11.02 32.515 11.08 32.5725 ;
        RECT  10.83 32.44 10.9 33.985 ;
        RECT  10.495 32.44 10.565 33.985 ;
        RECT  10.31 32.44 10.38 33.985 ;
        RECT  11.015 32.44 11.085 33.985 ;
        RECT  10.495 32.44 10.565 33.985 ;
        RECT  10.31 32.44 10.38 33.985 ;
        RECT  11.015 32.44 11.085 33.985 ;
        RECT  10.83 32.44 10.9 33.985 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  10.2775 35.195 10.4125 35.265 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  10.565 34.8375 10.635 34.9725 ;
        RECT  10.31 34.345 10.38 34.48 ;
        RECT  10.31 34.345 10.38 34.48 ;
        RECT  10.31 34.345 10.38 34.48 ;
        RECT  10.31 34.345 10.38 34.48 ;
        RECT  10.31 34.345 10.38 34.48 ;
        RECT  10.31 34.345 10.38 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  10.76 34.8375 10.83 34.9725 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  10.2775 35.195 10.4125 35.265 ;
        RECT  11.015 33.8525 11.085 35.2625 ;
        RECT  10.315 35.2025 10.375 35.26 ;
        RECT  10.5025 35.2025 10.5575 35.255 ;
        RECT  10.8375 35.2025 10.895 35.2625 ;
        RECT  11.02 35.1975 11.08 35.255 ;
        RECT  10.83 33.785 10.9 35.33 ;
        RECT  10.495 33.785 10.565 35.33 ;
        RECT  10.31 33.785 10.38 35.33 ;
        RECT  11.015 33.785 11.085 35.33 ;
        RECT  10.495 33.785 10.565 35.33 ;
        RECT  10.31 33.785 10.38 35.33 ;
        RECT  11.015 33.785 11.085 35.33 ;
        RECT  10.83 33.785 10.9 35.33 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  10.2775 35.195 10.4125 35.265 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  10.565 35.4875 10.635 35.6225 ;
        RECT  10.31 35.98 10.38 36.115 ;
        RECT  10.31 35.98 10.38 36.115 ;
        RECT  10.31 35.98 10.38 36.115 ;
        RECT  10.31 35.98 10.38 36.115 ;
        RECT  10.31 35.98 10.38 36.115 ;
        RECT  10.31 35.98 10.38 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  10.76 35.4875 10.83 35.6225 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  10.2775 35.195 10.4125 35.265 ;
        RECT  11.015 35.1975 11.085 36.6075 ;
        RECT  10.315 35.2 10.375 35.2575 ;
        RECT  10.5025 35.205 10.5575 35.2575 ;
        RECT  10.8375 35.1975 10.895 35.2575 ;
        RECT  11.02 35.205 11.08 35.2625 ;
        RECT  10.83 35.13 10.9 36.675 ;
        RECT  10.495 35.13 10.565 36.675 ;
        RECT  10.31 35.13 10.38 36.675 ;
        RECT  11.015 35.13 11.085 36.675 ;
        RECT  10.495 35.13 10.565 36.675 ;
        RECT  10.31 35.13 10.38 36.675 ;
        RECT  11.015 35.13 11.085 36.675 ;
        RECT  10.83 35.13 10.9 36.675 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  10.2775 37.885 10.4125 37.955 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  10.565 37.5275 10.635 37.6625 ;
        RECT  10.31 37.035 10.38 37.17 ;
        RECT  10.31 37.035 10.38 37.17 ;
        RECT  10.31 37.035 10.38 37.17 ;
        RECT  10.31 37.035 10.38 37.17 ;
        RECT  10.31 37.035 10.38 37.17 ;
        RECT  10.31 37.035 10.38 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  10.76 37.5275 10.83 37.6625 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  10.2775 37.885 10.4125 37.955 ;
        RECT  11.015 36.5425 11.085 37.9525 ;
        RECT  10.315 37.8925 10.375 37.95 ;
        RECT  10.5025 37.8925 10.5575 37.945 ;
        RECT  10.8375 37.8925 10.895 37.9525 ;
        RECT  11.02 37.8875 11.08 37.945 ;
        RECT  10.83 36.475 10.9 38.02 ;
        RECT  10.495 36.475 10.565 38.02 ;
        RECT  10.31 36.475 10.38 38.02 ;
        RECT  11.015 36.475 11.085 38.02 ;
        RECT  10.495 36.475 10.565 38.02 ;
        RECT  10.31 36.475 10.38 38.02 ;
        RECT  11.015 36.475 11.085 38.02 ;
        RECT  10.83 36.475 10.9 38.02 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  10.2775 37.885 10.4125 37.955 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  10.565 38.1775 10.635 38.3125 ;
        RECT  10.31 38.67 10.38 38.805 ;
        RECT  10.31 38.67 10.38 38.805 ;
        RECT  10.31 38.67 10.38 38.805 ;
        RECT  10.31 38.67 10.38 38.805 ;
        RECT  10.31 38.67 10.38 38.805 ;
        RECT  10.31 38.67 10.38 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  10.76 38.1775 10.83 38.3125 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  10.2775 37.885 10.4125 37.955 ;
        RECT  11.015 37.8875 11.085 39.2975 ;
        RECT  10.315 37.89 10.375 37.9475 ;
        RECT  10.5025 37.895 10.5575 37.9475 ;
        RECT  10.8375 37.8875 10.895 37.9475 ;
        RECT  11.02 37.895 11.08 37.9525 ;
        RECT  10.83 37.82 10.9 39.365 ;
        RECT  10.495 37.82 10.565 39.365 ;
        RECT  10.31 37.82 10.38 39.365 ;
        RECT  11.015 37.82 11.085 39.365 ;
        RECT  10.495 37.82 10.565 39.365 ;
        RECT  10.31 37.82 10.38 39.365 ;
        RECT  11.015 37.82 11.085 39.365 ;
        RECT  10.83 37.82 10.9 39.365 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  10.2775 40.575 10.4125 40.645 ;
        RECT  10.9825 40.575 11.1175 40.645 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  10.565 40.2175 10.635 40.3525 ;
        RECT  10.31 39.725 10.38 39.86 ;
        RECT  10.31 39.725 10.38 39.86 ;
        RECT  10.31 39.725 10.38 39.86 ;
        RECT  10.31 39.725 10.38 39.86 ;
        RECT  10.31 39.725 10.38 39.86 ;
        RECT  10.31 39.725 10.38 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  10.76 40.2175 10.83 40.3525 ;
        RECT  10.9825 40.575 11.1175 40.645 ;
        RECT  10.9825 40.575 11.1175 40.645 ;
        RECT  10.9825 40.575 11.1175 40.645 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  10.2775 40.575 10.4125 40.645 ;
        RECT  11.015 39.2325 11.085 40.6425 ;
        RECT  10.315 40.5825 10.375 40.64 ;
        RECT  10.5025 40.5825 10.5575 40.635 ;
        RECT  10.8375 40.5825 10.895 40.6425 ;
        RECT  11.02 40.5775 11.08 40.635 ;
        RECT  10.83 39.165 10.9 40.71 ;
        RECT  10.495 39.165 10.565 40.71 ;
        RECT  10.31 39.165 10.38 40.71 ;
        RECT  11.015 39.165 11.085 40.71 ;
        RECT  10.495 39.165 10.565 40.71 ;
        RECT  10.31 39.165 10.38 40.71 ;
        RECT  11.015 39.165 11.085 40.71 ;
        RECT  10.83 39.165 10.9 40.71 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  10.9825 19.055 11.1175 19.125 ;
        RECT  11.6875 19.055 11.8225 19.125 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.27 19.3475 11.34 19.4825 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.465 19.3475 11.535 19.4825 ;
        RECT  11.6875 19.055 11.8225 19.125 ;
        RECT  11.6875 19.055 11.8225 19.125 ;
        RECT  11.6875 19.055 11.8225 19.125 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  10.9825 19.055 11.1175 19.125 ;
        RECT  11.72 19.0575 11.79 20.4675 ;
        RECT  11.02 19.06 11.08 19.1175 ;
        RECT  11.2075 19.065 11.2625 19.1175 ;
        RECT  11.5425 19.0575 11.6 19.1175 ;
        RECT  11.725 19.065 11.785 19.1225 ;
        RECT  11.535 18.99 11.605 20.535 ;
        RECT  11.2 18.99 11.27 20.535 ;
        RECT  11.015 18.99 11.085 20.535 ;
        RECT  11.72 18.99 11.79 20.535 ;
        RECT  11.2 18.99 11.27 20.535 ;
        RECT  11.015 18.99 11.085 20.535 ;
        RECT  11.72 18.99 11.79 20.535 ;
        RECT  11.535 18.99 11.605 20.535 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.27 21.3875 11.34 21.5225 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.465 21.3875 11.535 21.5225 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.72 20.4025 11.79 21.8125 ;
        RECT  11.02 21.7525 11.08 21.81 ;
        RECT  11.2075 21.7525 11.2625 21.805 ;
        RECT  11.5425 21.7525 11.6 21.8125 ;
        RECT  11.725 21.7475 11.785 21.805 ;
        RECT  11.535 20.335 11.605 21.88 ;
        RECT  11.2 20.335 11.27 21.88 ;
        RECT  11.015 20.335 11.085 21.88 ;
        RECT  11.72 20.335 11.79 21.88 ;
        RECT  11.2 20.335 11.27 21.88 ;
        RECT  11.015 20.335 11.085 21.88 ;
        RECT  11.72 20.335 11.79 21.88 ;
        RECT  11.535 20.335 11.605 21.88 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.27 22.0375 11.34 22.1725 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.465 22.0375 11.535 22.1725 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.72 21.7475 11.79 23.1575 ;
        RECT  11.02 21.75 11.08 21.8075 ;
        RECT  11.2075 21.755 11.2625 21.8075 ;
        RECT  11.5425 21.7475 11.6 21.8075 ;
        RECT  11.725 21.755 11.785 21.8125 ;
        RECT  11.535 21.68 11.605 23.225 ;
        RECT  11.2 21.68 11.27 23.225 ;
        RECT  11.015 21.68 11.085 23.225 ;
        RECT  11.72 21.68 11.79 23.225 ;
        RECT  11.2 21.68 11.27 23.225 ;
        RECT  11.015 21.68 11.085 23.225 ;
        RECT  11.72 21.68 11.79 23.225 ;
        RECT  11.535 21.68 11.605 23.225 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.27 24.0775 11.34 24.2125 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.465 24.0775 11.535 24.2125 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.72 23.0925 11.79 24.5025 ;
        RECT  11.02 24.4425 11.08 24.5 ;
        RECT  11.2075 24.4425 11.2625 24.495 ;
        RECT  11.5425 24.4425 11.6 24.5025 ;
        RECT  11.725 24.4375 11.785 24.495 ;
        RECT  11.535 23.025 11.605 24.57 ;
        RECT  11.2 23.025 11.27 24.57 ;
        RECT  11.015 23.025 11.085 24.57 ;
        RECT  11.72 23.025 11.79 24.57 ;
        RECT  11.2 23.025 11.27 24.57 ;
        RECT  11.015 23.025 11.085 24.57 ;
        RECT  11.72 23.025 11.79 24.57 ;
        RECT  11.535 23.025 11.605 24.57 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.27 24.7275 11.34 24.8625 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.465 24.7275 11.535 24.8625 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.72 24.4375 11.79 25.8475 ;
        RECT  11.02 24.44 11.08 24.4975 ;
        RECT  11.2075 24.445 11.2625 24.4975 ;
        RECT  11.5425 24.4375 11.6 24.4975 ;
        RECT  11.725 24.445 11.785 24.5025 ;
        RECT  11.535 24.37 11.605 25.915 ;
        RECT  11.2 24.37 11.27 25.915 ;
        RECT  11.015 24.37 11.085 25.915 ;
        RECT  11.72 24.37 11.79 25.915 ;
        RECT  11.2 24.37 11.27 25.915 ;
        RECT  11.015 24.37 11.085 25.915 ;
        RECT  11.72 24.37 11.79 25.915 ;
        RECT  11.535 24.37 11.605 25.915 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.27 26.7675 11.34 26.9025 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.465 26.7675 11.535 26.9025 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.72 25.7825 11.79 27.1925 ;
        RECT  11.02 27.1325 11.08 27.19 ;
        RECT  11.2075 27.1325 11.2625 27.185 ;
        RECT  11.5425 27.1325 11.6 27.1925 ;
        RECT  11.725 27.1275 11.785 27.185 ;
        RECT  11.535 25.715 11.605 27.26 ;
        RECT  11.2 25.715 11.27 27.26 ;
        RECT  11.015 25.715 11.085 27.26 ;
        RECT  11.72 25.715 11.79 27.26 ;
        RECT  11.2 25.715 11.27 27.26 ;
        RECT  11.015 25.715 11.085 27.26 ;
        RECT  11.72 25.715 11.79 27.26 ;
        RECT  11.535 25.715 11.605 27.26 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.27 27.4175 11.34 27.5525 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.465 27.4175 11.535 27.5525 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.72 27.1275 11.79 28.5375 ;
        RECT  11.02 27.13 11.08 27.1875 ;
        RECT  11.2075 27.135 11.2625 27.1875 ;
        RECT  11.5425 27.1275 11.6 27.1875 ;
        RECT  11.725 27.135 11.785 27.1925 ;
        RECT  11.535 27.06 11.605 28.605 ;
        RECT  11.2 27.06 11.27 28.605 ;
        RECT  11.015 27.06 11.085 28.605 ;
        RECT  11.72 27.06 11.79 28.605 ;
        RECT  11.2 27.06 11.27 28.605 ;
        RECT  11.015 27.06 11.085 28.605 ;
        RECT  11.72 27.06 11.79 28.605 ;
        RECT  11.535 27.06 11.605 28.605 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.27 29.4575 11.34 29.5925 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.465 29.4575 11.535 29.5925 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.72 28.4725 11.79 29.8825 ;
        RECT  11.02 29.8225 11.08 29.88 ;
        RECT  11.2075 29.8225 11.2625 29.875 ;
        RECT  11.5425 29.8225 11.6 29.8825 ;
        RECT  11.725 29.8175 11.785 29.875 ;
        RECT  11.535 28.405 11.605 29.95 ;
        RECT  11.2 28.405 11.27 29.95 ;
        RECT  11.015 28.405 11.085 29.95 ;
        RECT  11.72 28.405 11.79 29.95 ;
        RECT  11.2 28.405 11.27 29.95 ;
        RECT  11.015 28.405 11.085 29.95 ;
        RECT  11.72 28.405 11.79 29.95 ;
        RECT  11.535 28.405 11.605 29.95 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.27 30.1075 11.34 30.2425 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.465 30.1075 11.535 30.2425 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.72 29.8175 11.79 31.2275 ;
        RECT  11.02 29.82 11.08 29.8775 ;
        RECT  11.2075 29.825 11.2625 29.8775 ;
        RECT  11.5425 29.8175 11.6 29.8775 ;
        RECT  11.725 29.825 11.785 29.8825 ;
        RECT  11.535 29.75 11.605 31.295 ;
        RECT  11.2 29.75 11.27 31.295 ;
        RECT  11.015 29.75 11.085 31.295 ;
        RECT  11.72 29.75 11.79 31.295 ;
        RECT  11.2 29.75 11.27 31.295 ;
        RECT  11.015 29.75 11.085 31.295 ;
        RECT  11.72 29.75 11.79 31.295 ;
        RECT  11.535 29.75 11.605 31.295 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.27 32.1475 11.34 32.2825 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.465 32.1475 11.535 32.2825 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.72 31.1625 11.79 32.5725 ;
        RECT  11.02 32.5125 11.08 32.57 ;
        RECT  11.2075 32.5125 11.2625 32.565 ;
        RECT  11.5425 32.5125 11.6 32.5725 ;
        RECT  11.725 32.5075 11.785 32.565 ;
        RECT  11.535 31.095 11.605 32.64 ;
        RECT  11.2 31.095 11.27 32.64 ;
        RECT  11.015 31.095 11.085 32.64 ;
        RECT  11.72 31.095 11.79 32.64 ;
        RECT  11.2 31.095 11.27 32.64 ;
        RECT  11.015 31.095 11.085 32.64 ;
        RECT  11.72 31.095 11.79 32.64 ;
        RECT  11.535 31.095 11.605 32.64 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.27 32.7975 11.34 32.9325 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.465 32.7975 11.535 32.9325 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.72 32.5075 11.79 33.9175 ;
        RECT  11.02 32.51 11.08 32.5675 ;
        RECT  11.2075 32.515 11.2625 32.5675 ;
        RECT  11.5425 32.5075 11.6 32.5675 ;
        RECT  11.725 32.515 11.785 32.5725 ;
        RECT  11.535 32.44 11.605 33.985 ;
        RECT  11.2 32.44 11.27 33.985 ;
        RECT  11.015 32.44 11.085 33.985 ;
        RECT  11.72 32.44 11.79 33.985 ;
        RECT  11.2 32.44 11.27 33.985 ;
        RECT  11.015 32.44 11.085 33.985 ;
        RECT  11.72 32.44 11.79 33.985 ;
        RECT  11.535 32.44 11.605 33.985 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.27 34.8375 11.34 34.9725 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.465 34.8375 11.535 34.9725 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.72 33.8525 11.79 35.2625 ;
        RECT  11.02 35.2025 11.08 35.26 ;
        RECT  11.2075 35.2025 11.2625 35.255 ;
        RECT  11.5425 35.2025 11.6 35.2625 ;
        RECT  11.725 35.1975 11.785 35.255 ;
        RECT  11.535 33.785 11.605 35.33 ;
        RECT  11.2 33.785 11.27 35.33 ;
        RECT  11.015 33.785 11.085 35.33 ;
        RECT  11.72 33.785 11.79 35.33 ;
        RECT  11.2 33.785 11.27 35.33 ;
        RECT  11.015 33.785 11.085 35.33 ;
        RECT  11.72 33.785 11.79 35.33 ;
        RECT  11.535 33.785 11.605 35.33 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.27 35.4875 11.34 35.6225 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.465 35.4875 11.535 35.6225 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.72 35.1975 11.79 36.6075 ;
        RECT  11.02 35.2 11.08 35.2575 ;
        RECT  11.2075 35.205 11.2625 35.2575 ;
        RECT  11.5425 35.1975 11.6 35.2575 ;
        RECT  11.725 35.205 11.785 35.2625 ;
        RECT  11.535 35.13 11.605 36.675 ;
        RECT  11.2 35.13 11.27 36.675 ;
        RECT  11.015 35.13 11.085 36.675 ;
        RECT  11.72 35.13 11.79 36.675 ;
        RECT  11.2 35.13 11.27 36.675 ;
        RECT  11.015 35.13 11.085 36.675 ;
        RECT  11.72 35.13 11.79 36.675 ;
        RECT  11.535 35.13 11.605 36.675 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.27 37.5275 11.34 37.6625 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.465 37.5275 11.535 37.6625 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.72 36.5425 11.79 37.9525 ;
        RECT  11.02 37.8925 11.08 37.95 ;
        RECT  11.2075 37.8925 11.2625 37.945 ;
        RECT  11.5425 37.8925 11.6 37.9525 ;
        RECT  11.725 37.8875 11.785 37.945 ;
        RECT  11.535 36.475 11.605 38.02 ;
        RECT  11.2 36.475 11.27 38.02 ;
        RECT  11.015 36.475 11.085 38.02 ;
        RECT  11.72 36.475 11.79 38.02 ;
        RECT  11.2 36.475 11.27 38.02 ;
        RECT  11.015 36.475 11.085 38.02 ;
        RECT  11.72 36.475 11.79 38.02 ;
        RECT  11.535 36.475 11.605 38.02 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.27 38.1775 11.34 38.3125 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.465 38.1775 11.535 38.3125 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.72 37.8875 11.79 39.2975 ;
        RECT  11.02 37.89 11.08 37.9475 ;
        RECT  11.2075 37.895 11.2625 37.9475 ;
        RECT  11.5425 37.8875 11.6 37.9475 ;
        RECT  11.725 37.895 11.785 37.9525 ;
        RECT  11.535 37.82 11.605 39.365 ;
        RECT  11.2 37.82 11.27 39.365 ;
        RECT  11.015 37.82 11.085 39.365 ;
        RECT  11.72 37.82 11.79 39.365 ;
        RECT  11.2 37.82 11.27 39.365 ;
        RECT  11.015 37.82 11.085 39.365 ;
        RECT  11.72 37.82 11.79 39.365 ;
        RECT  11.535 37.82 11.605 39.365 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  10.9825 40.575 11.1175 40.645 ;
        RECT  11.6875 40.575 11.8225 40.645 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.27 40.2175 11.34 40.3525 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.465 40.2175 11.535 40.3525 ;
        RECT  11.6875 40.575 11.8225 40.645 ;
        RECT  11.6875 40.575 11.8225 40.645 ;
        RECT  11.6875 40.575 11.8225 40.645 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  10.9825 40.575 11.1175 40.645 ;
        RECT  11.72 39.2325 11.79 40.6425 ;
        RECT  11.02 40.5825 11.08 40.64 ;
        RECT  11.2075 40.5825 11.2625 40.635 ;
        RECT  11.5425 40.5825 11.6 40.6425 ;
        RECT  11.725 40.5775 11.785 40.635 ;
        RECT  11.535 39.165 11.605 40.71 ;
        RECT  11.2 39.165 11.27 40.71 ;
        RECT  11.015 39.165 11.085 40.71 ;
        RECT  11.72 39.165 11.79 40.71 ;
        RECT  11.2 39.165 11.27 40.71 ;
        RECT  11.015 39.165 11.085 40.71 ;
        RECT  11.72 39.165 11.79 40.71 ;
        RECT  11.535 39.165 11.605 40.71 ;
        RECT  11.2 41.06 11.27 42.27 ;
        RECT  10.495 41.06 10.565 42.27 ;
        RECT  11.535 41.06 11.605 42.27 ;
        RECT  10.83 41.06 10.9 42.27 ;
        RECT  10.495 41.1825 10.5725 41.3175 ;
        RECT  10.6975 41.1825 10.9 41.3175 ;
        RECT  10.495 41.7675 10.5725 41.9025 ;
        RECT  10.83 41.7675 10.9525 41.9025 ;
        RECT  10.495 41.06 10.565 42.27 ;
        RECT  10.83 41.06 10.9 42.27 ;
        RECT  10.505 41.1825 10.575 41.3175 ;
        RECT  10.695 41.1825 10.765 41.3175 ;
        RECT  10.505 41.7675 10.575 41.9025 ;
        RECT  10.885 41.7675 10.955 41.9025 ;
        RECT  11.2 41.1825 11.2775 41.3175 ;
        RECT  11.4025 41.1825 11.605 41.3175 ;
        RECT  11.2 41.7675 11.2775 41.9025 ;
        RECT  11.535 41.7675 11.6575 41.9025 ;
        RECT  11.2 41.06 11.27 42.27 ;
        RECT  11.535 41.06 11.605 42.27 ;
        RECT  11.21 41.1825 11.28 41.3175 ;
        RECT  11.4 41.1825 11.47 41.3175 ;
        RECT  11.21 41.7675 11.28 41.9025 ;
        RECT  11.59 41.7675 11.66 41.9025 ;
        RECT  11.2 14.205 11.27 19.09 ;
        RECT  10.495 14.205 10.565 19.09 ;
        RECT  11.535 14.205 11.605 18.29 ;
        RECT  10.83 14.205 10.9 18.29 ;
        RECT  10.31 14.205 10.38 19.09 ;
        RECT  10.495 14.205 10.565 19.09 ;
        RECT  10.83 14.205 10.9 17.75 ;
        RECT  10.6625 16.48 10.7325 18.49 ;
        RECT  10.83 15.005 10.9 19.09 ;
        RECT  11.015 14.205 11.085 19.09 ;
        RECT  10.835 19.04 10.895 19.09 ;
        RECT  10.495 19.03 10.565 19.09 ;
        RECT  10.6575 19.035 10.7275 19.09 ;
        RECT  10.6575 18.6925 10.7275 19.09 ;
        RECT  10.6625 16.345 10.7325 16.48 ;
        RECT  10.6625 18.4875 10.7325 18.6225 ;
        RECT  10.47 17.645 10.54 17.78 ;
        RECT  10.8525 17.235 10.9225 17.37 ;
        RECT  10.31 14.4525 10.38 14.5875 ;
        RECT  11.015 14.4525 11.085 14.5875 ;
        RECT  10.6575 18.6925 10.7275 18.8275 ;
        RECT  10.6575 18.95 10.7275 19.09 ;
        RECT  10.83 15.005 10.9 19.09 ;
        RECT  10.495 14.205 10.565 19.09 ;
        RECT  11.015 14.205 11.085 19.09 ;
        RECT  11.2 14.205 11.27 19.09 ;
        RECT  11.535 14.205 11.605 17.75 ;
        RECT  11.3675 16.48 11.4375 18.49 ;
        RECT  11.535 15.005 11.605 19.09 ;
        RECT  11.72 14.205 11.79 19.09 ;
        RECT  11.54 19.04 11.6 19.09 ;
        RECT  11.2 19.03 11.27 19.09 ;
        RECT  11.3625 19.035 11.4325 19.09 ;
        RECT  11.3625 18.6925 11.4325 19.09 ;
        RECT  11.3675 16.345 11.4375 16.48 ;
        RECT  11.3675 18.4875 11.4375 18.6225 ;
        RECT  11.175 17.645 11.245 17.78 ;
        RECT  11.5575 17.235 11.6275 17.37 ;
        RECT  11.015 14.4525 11.085 14.5875 ;
        RECT  11.72 14.4525 11.79 14.5875 ;
        RECT  11.3625 18.6925 11.4325 18.8275 ;
        RECT  11.3625 18.95 11.4325 19.09 ;
        RECT  11.535 15.005 11.605 19.09 ;
        RECT  11.2 14.205 11.27 19.09 ;
        RECT  10.6625 10.03 10.7325 10.17 ;
        RECT  11.3675 10.03 11.4375 10.17 ;
        RECT  10.495 13.905 10.565 14.205 ;
        RECT  11.2 13.905 11.27 14.205 ;
        RECT  11.535 11.765 11.605 14.205 ;
        RECT  10.83 11.765 10.9 14.205 ;
        RECT  10.5525 10.1625 10.6875 10.2325 ;
        RECT  11.015 11.765 11.085 11.9 ;
        RECT  11.015 11.195 11.085 11.33 ;
        RECT  10.31 11.195 10.38 11.33 ;
        RECT  10.73 11.4 10.8 11.535 ;
        RECT  11.015 13.6925 11.085 13.8275 ;
        RECT  10.73 10.99 10.8 11.125 ;
        RECT  10.59 10.99 10.66 11.125 ;
        RECT  11.015 11.4 11.085 11.535 ;
        RECT  10.31 11.4 10.38 11.535 ;
        RECT  10.45 10.425 10.585 10.495 ;
        RECT  10.59 13.37 10.66 13.505 ;
        RECT  10.76 11.765 10.83 11.9 ;
        RECT  10.45 12.68 10.52 12.815 ;
        RECT  10.59 11.4 10.66 11.535 ;
        RECT  10.31 11.765 10.38 11.9 ;
        RECT  10.76 12.28 10.83 12.415 ;
        RECT  10.495 13.9025 10.565 14.0375 ;
        RECT  10.31 13.6925 10.38 13.8275 ;
        RECT  10.495 13.905 10.565 14.205 ;
        RECT  10.495 14.14 10.565 14.205 ;
        RECT  10.8325 14.145 10.8975 14.205 ;
        RECT  10.665 10.035 10.73 10.0975 ;
        RECT  11.015 10.03 11.085 14.205 ;
        RECT  10.31 10.03 10.38 14.205 ;
        RECT  10.83 11.765 10.9 14.205 ;
        RECT  10.54 10.1625 10.7325 10.2325 ;
        RECT  10.73 11.125 10.8 11.4 ;
        RECT  10.45 10.495 10.52 12.815 ;
        RECT  10.59 11.125 10.66 11.4 ;
        RECT  10.59 11.4 10.66 13.4975 ;
        RECT  10.6625 10.03 10.7325 10.17 ;
        RECT  10.6625 10.03 10.7325 10.17 ;
        RECT  10.83 11.765 10.9 14.205 ;
        RECT  10.495 13.905 10.565 14.205 ;
        RECT  11.2575 10.1625 11.3925 10.2325 ;
        RECT  11.72 11.765 11.79 11.9 ;
        RECT  11.72 11.195 11.79 11.33 ;
        RECT  11.015 11.195 11.085 11.33 ;
        RECT  11.435 11.4 11.505 11.535 ;
        RECT  11.72 13.6925 11.79 13.8275 ;
        RECT  11.435 10.99 11.505 11.125 ;
        RECT  11.295 10.99 11.365 11.125 ;
        RECT  11.72 11.4 11.79 11.535 ;
        RECT  11.015 11.4 11.085 11.535 ;
        RECT  11.155 10.425 11.29 10.495 ;
        RECT  11.295 13.37 11.365 13.505 ;
        RECT  11.465 11.765 11.535 11.9 ;
        RECT  11.155 12.68 11.225 12.815 ;
        RECT  11.295 11.4 11.365 11.535 ;
        RECT  11.015 11.765 11.085 11.9 ;
        RECT  11.465 12.28 11.535 12.415 ;
        RECT  11.2 13.9025 11.27 14.0375 ;
        RECT  11.015 13.6925 11.085 13.8275 ;
        RECT  11.2 13.905 11.27 14.205 ;
        RECT  11.2 14.14 11.27 14.205 ;
        RECT  11.5375 14.145 11.6025 14.205 ;
        RECT  11.37 10.035 11.435 10.0975 ;
        RECT  11.72 10.03 11.79 14.205 ;
        RECT  11.015 10.03 11.085 14.205 ;
        RECT  11.535 11.765 11.605 14.205 ;
        RECT  11.245 10.1625 11.4375 10.2325 ;
        RECT  11.435 11.125 11.505 11.4 ;
        RECT  11.155 10.495 11.225 12.815 ;
        RECT  11.295 11.125 11.365 11.4 ;
        RECT  11.295 11.4 11.365 13.4975 ;
        RECT  11.3675 10.03 11.4375 10.17 ;
        RECT  11.3675 10.03 11.4375 10.17 ;
        RECT  11.535 11.765 11.605 14.205 ;
        RECT  11.2 13.905 11.27 14.205 ;
        RECT  11.5225 9.3425 11.5925 10.03 ;
        RECT  11.3675 3.59 11.4375 3.735 ;
        RECT  10.6625 3.59 10.7325 3.735 ;
        RECT  10.31 3.59 10.38 10.03 ;
        RECT  11.015 3.59 11.085 10.03 ;
        RECT  11.72 3.59 11.79 10.03 ;
        RECT  10.5075 9.3425 10.5775 10.03 ;
        RECT  10.6625 9.76 10.7325 10.03 ;
        RECT  11.3675 9.76 11.4375 10.03 ;
        RECT  10.5075 9.2925 10.5775 9.4275 ;
        RECT  11.015 4.115 11.085 4.25 ;
        RECT  10.8725 8.1975 10.9425 8.3325 ;
        RECT  10.875 6.59 10.945 6.725 ;
        RECT  10.875 5.1925 10.945 5.3275 ;
        RECT  10.31 3.975 10.38 4.11 ;
        RECT  10.6625 3.59 10.7325 3.73 ;
        RECT  11.015 7.0525 11.085 7.1875 ;
        RECT  10.51 5.8575 10.58 5.9925 ;
        RECT  10.875 9.55 10.945 9.685 ;
        RECT  10.6975 9.04 10.7675 9.175 ;
        RECT  11.015 8.6275 11.085 8.7625 ;
        RECT  11.015 3.925 11.085 4.06 ;
        RECT  11.015 5.6675 11.085 5.8025 ;
        RECT  10.51 5.4675 10.58 5.6025 ;
        RECT  10.6975 5.4675 10.7675 5.6025 ;
        RECT  10.6975 6.08 10.7675 6.215 ;
        RECT  10.5075 8.4275 10.5775 8.5625 ;
        RECT  10.6975 8.4275 10.7675 8.5625 ;
        RECT  10.7325 9.76 10.875 9.83 ;
        RECT  10.6625 3.59 10.7325 3.735 ;
        RECT  10.7275 3.665 10.875 3.735 ;
        RECT  10.6625 9.76 10.7325 10.03 ;
        RECT  10.3125 9.5525 10.375 9.6125 ;
        RECT  10.31 3.59 10.38 10.03 ;
        RECT  10.665 9.965 10.73 10.025 ;
        RECT  10.875 9.55 10.945 9.83 ;
        RECT  10.875 3.665 10.945 5.3275 ;
        RECT  10.5075 9.3425 10.5775 10.03 ;
        RECT  10.875 6.725 10.945 8.3325 ;
        RECT  10.6975 8.4275 10.7675 9.145 ;
        RECT  10.51 5.4675 10.58 5.9925 ;
        RECT  10.5125 9.8925 10.575 9.9525 ;
        RECT  10.5075 8.4275 10.5775 9.3675 ;
        RECT  10.6625 3.595 10.73 3.66 ;
        RECT  11.015 3.59 11.085 10.03 ;
        RECT  10.6975 5.4675 10.7675 6.185 ;
        RECT  10.6625 3.59 10.7325 3.735 ;
        RECT  10.6625 9.76 10.7325 10.03 ;
        RECT  10.5075 9.3425 10.5775 10.03 ;
        RECT  10.31 3.59 10.38 10.03 ;
        RECT  11.015 3.59 11.085 10.03 ;
        RECT  11.5225 9.2925 11.5925 9.4275 ;
        RECT  11.015 4.115 11.085 4.25 ;
        RECT  11.1575 8.1975 11.2275 8.3325 ;
        RECT  11.155 6.59 11.225 6.725 ;
        RECT  11.155 5.1925 11.225 5.3275 ;
        RECT  11.72 3.975 11.79 4.11 ;
        RECT  11.3675 3.59 11.4375 3.73 ;
        RECT  11.015 7.0525 11.085 7.1875 ;
        RECT  11.52 5.8575 11.59 5.9925 ;
        RECT  11.155 9.55 11.225 9.685 ;
        RECT  11.3325 9.04 11.4025 9.175 ;
        RECT  11.015 8.6275 11.085 8.7625 ;
        RECT  11.015 3.925 11.085 4.06 ;
        RECT  11.015 5.6675 11.085 5.8025 ;
        RECT  11.52 5.4675 11.59 5.6025 ;
        RECT  11.3325 5.4675 11.4025 5.6025 ;
        RECT  11.3325 6.08 11.4025 6.215 ;
        RECT  11.5225 8.4275 11.5925 8.5625 ;
        RECT  11.3325 8.4275 11.4025 8.5625 ;
        RECT  11.225 9.76 11.3675 9.83 ;
        RECT  11.3675 3.59 11.4375 3.735 ;
        RECT  11.225 3.665 11.3725 3.735 ;
        RECT  11.3675 9.76 11.4375 10.03 ;
        RECT  11.725 9.5525 11.7875 9.6125 ;
        RECT  11.72 3.59 11.79 10.03 ;
        RECT  11.37 9.965 11.435 10.025 ;
        RECT  11.155 9.55 11.225 9.83 ;
        RECT  11.155 3.665 11.225 5.3275 ;
        RECT  11.5225 9.3425 11.5925 10.03 ;
        RECT  11.155 6.725 11.225 8.3325 ;
        RECT  11.3325 8.4275 11.4025 9.145 ;
        RECT  11.52 5.4675 11.59 5.9925 ;
        RECT  11.525 9.8925 11.5875 9.9525 ;
        RECT  11.5225 8.4275 11.5925 9.3675 ;
        RECT  11.37 3.595 11.4375 3.66 ;
        RECT  11.015 3.59 11.085 10.03 ;
        RECT  11.3325 5.4675 11.4025 6.185 ;
        RECT  11.3675 3.59 11.4375 3.735 ;
        RECT  11.3675 9.76 11.4375 10.03 ;
        RECT  11.5225 9.3425 11.5925 10.03 ;
        RECT  11.72 3.59 11.79 10.03 ;
        RECT  11.015 3.59 11.085 10.03 ;
        RECT  10.6625 0.615 10.7325 0.855 ;
        RECT  10.6625 3.24 10.7325 3.59 ;
        RECT  11.3675 3.24 11.4375 3.59 ;
        RECT  11.3675 0.615 11.4375 0.855 ;
        RECT  10.45 3.87 10.52 4.24 ;
        RECT  10.5225 4.505 10.7625 4.575 ;
        RECT  10.7625 4.505 10.8975 4.575 ;
        RECT  11.015 4.1625 11.085 4.22 ;
        RECT  11.015 3.59 11.085 6.565 ;
        RECT  10.695 5.4425 10.765 5.68 ;
        RECT  10.835 6.0125 10.905 6.395 ;
        RECT  10.4525 4.505 10.5225 6.0925 ;
        RECT  10.6625 3.745 10.7325 3.8075 ;
        RECT  10.6625 6.5075 10.7325 6.56 ;
        RECT  10.6625 6.325 10.7325 6.565 ;
        RECT  10.7325 6.325 10.835 6.395 ;
        RECT  10.6625 3.59 10.7325 3.94 ;
        RECT  10.45 3.87 10.6625 3.94 ;
        RECT  10.695 5.68 10.765 5.815 ;
        RECT  10.4875 5.9575 10.5575 6.0925 ;
        RECT  11.015 6.1475 11.085 6.2825 ;
        RECT  10.7625 6.0125 10.8975 6.0825 ;
        RECT  10.6625 3.7425 10.7325 3.8825 ;
        RECT  11.015 4.0875 11.085 4.2225 ;
        RECT  10.63 5.3725 10.765 5.4425 ;
        RECT  11.015 3.59 11.085 6.565 ;
        RECT  10.6625 6.325 10.7325 6.565 ;
        RECT  10.6625 3.59 10.7325 3.94 ;
        RECT  10.45 4.24 10.52 4.375 ;
        RECT  11.155 3.87 11.225 4.24 ;
        RECT  11.2275 4.505 11.4675 4.575 ;
        RECT  11.4675 4.505 11.6025 4.575 ;
        RECT  11.72 4.1625 11.79 4.22 ;
        RECT  11.72 3.59 11.79 6.565 ;
        RECT  11.4 5.4425 11.47 5.68 ;
        RECT  11.54 6.0125 11.61 6.395 ;
        RECT  11.1575 4.505 11.2275 6.0925 ;
        RECT  11.3675 3.745 11.4375 3.8075 ;
        RECT  11.3675 6.5075 11.4375 6.56 ;
        RECT  11.3675 6.325 11.4375 6.565 ;
        RECT  11.4375 6.325 11.54 6.395 ;
        RECT  11.3675 3.59 11.4375 3.94 ;
        RECT  11.155 3.87 11.3675 3.94 ;
        RECT  11.4 5.68 11.47 5.815 ;
        RECT  11.1925 5.9575 11.2625 6.0925 ;
        RECT  11.72 6.1475 11.79 6.2825 ;
        RECT  11.4675 6.0125 11.6025 6.0825 ;
        RECT  11.3675 3.7425 11.4375 3.8825 ;
        RECT  11.72 4.0875 11.79 4.2225 ;
        RECT  11.335 5.3725 11.47 5.4425 ;
        RECT  11.72 3.59 11.79 6.565 ;
        RECT  11.3675 6.325 11.4375 6.565 ;
        RECT  11.3675 3.59 11.4375 3.94 ;
        RECT  11.155 4.24 11.225 4.375 ;
        RECT  1.555 8.33 1.625 40.61 ;
        RECT  1.73 8.33 1.8 40.61 ;
        RECT  1.905 8.33 1.975 40.61 ;
        RECT  2.08 8.33 2.15 40.61 ;
        RECT  2.255 8.33 2.325 40.61 ;
        RECT  2.43 8.33 2.5 40.61 ;
        RECT  2.605 8.33 2.675 40.61 ;
        RECT  2.78 8.33 2.85 40.61 ;
        RECT  6.575 13.71 6.645 18.95 ;
        RECT  6.575 8.33 6.645 13.57 ;
        RECT  6.85 8.33 6.92 13.57 ;
        RECT  6.85 13.71 6.92 18.95 ;
        RECT  4.915 8.33 4.985 13.57 ;
        RECT  4.64 8.33 4.71 13.57 ;
        RECT  5.465 8.33 5.535 13.57 ;
        RECT  5.19 8.33 5.26 13.57 ;
        RECT  6.85 8.33 6.92 13.57 ;
        RECT  6.575 8.33 6.645 13.57 ;
        RECT  4.11 7.655 4.18 7.725 ;
        RECT  3.92 7.655 3.99 7.725 ;
        RECT  4.11 7.3275 4.18 7.69 ;
        RECT  3.955 7.655 4.145 7.725 ;
        RECT  3.92 7.69 3.99 8.0325 ;
        RECT  4.11 7.1925 4.18 7.3275 ;
        RECT  3.92 8.0325 3.99 8.1675 ;
        RECT  3.8875 7.655 4.0225 7.725 ;
        RECT  4.11 11.625 4.18 11.695 ;
        RECT  3.92 11.625 3.99 11.695 ;
        RECT  4.11 11.66 4.18 12.0225 ;
        RECT  3.955 11.625 4.145 11.695 ;
        RECT  3.92 11.3175 3.99 11.66 ;
        RECT  4.11 11.8875 4.18 12.0225 ;
        RECT  3.92 11.0475 3.99 11.1825 ;
        RECT  3.8875 11.555 4.0225 11.625 ;
        RECT  4.11 10.345 4.18 10.415 ;
        RECT  3.92 10.345 3.99 10.415 ;
        RECT  4.11 10.0175 4.18 10.38 ;
        RECT  3.955 10.345 4.145 10.415 ;
        RECT  3.92 10.38 3.99 10.7225 ;
        RECT  4.11 9.8825 4.18 10.0175 ;
        RECT  3.92 10.7225 3.99 10.8575 ;
        RECT  3.8875 10.345 4.0225 10.415 ;
        RECT  4.11 14.315 4.18 14.385 ;
        RECT  3.92 14.315 3.99 14.385 ;
        RECT  4.11 14.35 4.18 14.7125 ;
        RECT  3.955 14.315 4.145 14.385 ;
        RECT  3.92 14.0075 3.99 14.35 ;
        RECT  4.11 14.5775 4.18 14.7125 ;
        RECT  3.92 13.7375 3.99 13.8725 ;
        RECT  3.8875 14.245 4.0225 14.315 ;
        RECT  5.4325 9.375 5.5675 9.445 ;
        RECT  6.8175 8.8075 6.9525 8.8775 ;
        RECT  5.1575 10.72 5.2925 10.79 ;
        RECT  6.5425 10.3325 6.6775 10.4025 ;
        RECT  6.8175 11.05 6.9525 11.12 ;
        RECT  4.8825 11.05 5.0175 11.12 ;
        RECT  6.5425 12.395 6.6775 12.465 ;
        RECT  4.6075 12.395 4.7425 12.465 ;
        RECT  5.4325 8.865 5.5675 8.935 ;
        RECT  5.1575 8.65 5.2925 8.72 ;
        RECT  4.8825 10.275 5.0175 10.345 ;
        RECT  5.1575 10.49 5.2925 10.56 ;
        RECT  5.4325 11.555 5.5675 11.625 ;
        RECT  4.6075 11.34 4.7425 11.41 ;
        RECT  4.8825 12.965 5.0175 13.035 ;
        RECT  4.6075 13.18 4.7425 13.25 ;
        RECT  4.915 13.71 4.985 18.95 ;
        RECT  4.64 13.71 4.71 18.95 ;
        RECT  5.465 13.71 5.535 18.95 ;
        RECT  5.19 13.71 5.26 18.95 ;
        RECT  6.85 13.71 6.92 18.95 ;
        RECT  6.575 13.71 6.645 18.95 ;
        RECT  4.11 13.035 4.18 13.105 ;
        RECT  3.92 13.035 3.99 13.105 ;
        RECT  4.11 12.7075 4.18 13.07 ;
        RECT  3.955 13.035 4.145 13.105 ;
        RECT  3.92 13.07 3.99 13.4125 ;
        RECT  4.11 12.5725 4.18 12.7075 ;
        RECT  3.92 13.4125 3.99 13.5475 ;
        RECT  3.8875 13.035 4.0225 13.105 ;
        RECT  4.11 17.005 4.18 17.075 ;
        RECT  3.92 17.005 3.99 17.075 ;
        RECT  4.11 17.04 4.18 17.4025 ;
        RECT  3.955 17.005 4.145 17.075 ;
        RECT  3.92 16.6975 3.99 17.04 ;
        RECT  4.11 17.2675 4.18 17.4025 ;
        RECT  3.92 16.4275 3.99 16.5625 ;
        RECT  3.8875 16.935 4.0225 17.005 ;
        RECT  4.11 15.725 4.18 15.795 ;
        RECT  3.92 15.725 3.99 15.795 ;
        RECT  4.11 15.3975 4.18 15.76 ;
        RECT  3.955 15.725 4.145 15.795 ;
        RECT  3.92 15.76 3.99 16.1025 ;
        RECT  4.11 15.2625 4.18 15.3975 ;
        RECT  3.92 16.1025 3.99 16.2375 ;
        RECT  3.8875 15.725 4.0225 15.795 ;
        RECT  4.11 19.695 4.18 19.765 ;
        RECT  3.92 19.695 3.99 19.765 ;
        RECT  4.11 19.73 4.18 20.0925 ;
        RECT  3.955 19.695 4.145 19.765 ;
        RECT  3.92 19.3875 3.99 19.73 ;
        RECT  4.11 19.9575 4.18 20.0925 ;
        RECT  3.92 19.1175 3.99 19.2525 ;
        RECT  3.8875 19.625 4.0225 19.695 ;
        RECT  5.4325 14.755 5.5675 14.825 ;
        RECT  6.8175 14.1875 6.9525 14.2575 ;
        RECT  5.1575 16.1 5.2925 16.17 ;
        RECT  6.5425 15.7125 6.6775 15.7825 ;
        RECT  6.8175 16.43 6.9525 16.5 ;
        RECT  4.8825 16.43 5.0175 16.5 ;
        RECT  6.5425 17.775 6.6775 17.845 ;
        RECT  4.6075 17.775 4.7425 17.845 ;
        RECT  5.4325 14.245 5.5675 14.315 ;
        RECT  5.1575 14.03 5.2925 14.1 ;
        RECT  4.8825 15.655 5.0175 15.725 ;
        RECT  5.1575 15.87 5.2925 15.94 ;
        RECT  5.4325 16.935 5.5675 17.005 ;
        RECT  4.6075 16.72 4.7425 16.79 ;
        RECT  4.8825 18.345 5.0175 18.415 ;
        RECT  4.6075 18.56 4.7425 18.63 ;
        RECT  3.21 19.695 3.28 19.765 ;
        RECT  3.4 19.695 3.47 19.765 ;
        RECT  3.21 19.73 3.28 20.0925 ;
        RECT  3.245 19.695 3.435 19.765 ;
        RECT  3.4 19.3875 3.47 19.73 ;
        RECT  3.21 20.0925 3.28 20.2275 ;
        RECT  3.4 19.2525 3.47 19.3875 ;
        RECT  3.3675 19.695 3.5025 19.765 ;
        RECT  3.21 21.105 3.28 21.175 ;
        RECT  3.4 21.105 3.47 21.175 ;
        RECT  3.21 20.7775 3.28 21.14 ;
        RECT  3.245 21.105 3.435 21.175 ;
        RECT  3.4 21.14 3.47 21.4825 ;
        RECT  3.21 20.7775 3.28 20.9125 ;
        RECT  3.4 21.6175 3.47 21.7525 ;
        RECT  3.3675 21.175 3.5025 21.245 ;
        RECT  3.21 22.385 3.28 22.455 ;
        RECT  3.4 22.385 3.47 22.455 ;
        RECT  3.21 22.42 3.28 22.7825 ;
        RECT  3.245 22.385 3.435 22.455 ;
        RECT  3.4 22.0775 3.47 22.42 ;
        RECT  3.21 22.7825 3.28 22.9175 ;
        RECT  3.4 21.9425 3.47 22.0775 ;
        RECT  3.3675 22.385 3.5025 22.455 ;
        RECT  3.21 23.795 3.28 23.865 ;
        RECT  3.4 23.795 3.47 23.865 ;
        RECT  3.21 23.4675 3.28 23.83 ;
        RECT  3.245 23.795 3.435 23.865 ;
        RECT  3.4 23.83 3.47 24.1725 ;
        RECT  3.21 23.4675 3.28 23.6025 ;
        RECT  3.4 24.3075 3.47 24.4425 ;
        RECT  3.3675 23.865 3.5025 23.935 ;
        RECT  3.21 25.075 3.28 25.145 ;
        RECT  3.4 25.075 3.47 25.145 ;
        RECT  3.21 25.11 3.28 25.4725 ;
        RECT  3.245 25.075 3.435 25.145 ;
        RECT  3.4 24.7675 3.47 25.11 ;
        RECT  3.21 25.4725 3.28 25.6075 ;
        RECT  3.4 24.6325 3.47 24.7675 ;
        RECT  3.3675 25.075 3.5025 25.145 ;
        RECT  3.21 26.485 3.28 26.555 ;
        RECT  3.4 26.485 3.47 26.555 ;
        RECT  3.21 26.1575 3.28 26.52 ;
        RECT  3.245 26.485 3.435 26.555 ;
        RECT  3.4 26.52 3.47 26.8625 ;
        RECT  3.21 26.1575 3.28 26.2925 ;
        RECT  3.4 26.9975 3.47 27.1325 ;
        RECT  3.3675 26.555 3.5025 26.625 ;
        RECT  3.21 27.765 3.28 27.835 ;
        RECT  3.4 27.765 3.47 27.835 ;
        RECT  3.21 27.8 3.28 28.1625 ;
        RECT  3.245 27.765 3.435 27.835 ;
        RECT  3.4 27.4575 3.47 27.8 ;
        RECT  3.21 28.1625 3.28 28.2975 ;
        RECT  3.4 27.3225 3.47 27.4575 ;
        RECT  3.3675 27.765 3.5025 27.835 ;
        RECT  3.21 29.175 3.28 29.245 ;
        RECT  3.4 29.175 3.47 29.245 ;
        RECT  3.21 28.8475 3.28 29.21 ;
        RECT  3.245 29.175 3.435 29.245 ;
        RECT  3.4 29.21 3.47 29.5525 ;
        RECT  3.21 28.8475 3.28 28.9825 ;
        RECT  3.4 29.6875 3.47 29.8225 ;
        RECT  3.3675 29.245 3.5025 29.315 ;
        RECT  3.21 30.455 3.28 30.525 ;
        RECT  3.4 30.455 3.47 30.525 ;
        RECT  3.21 30.49 3.28 30.8525 ;
        RECT  3.245 30.455 3.435 30.525 ;
        RECT  3.4 30.1475 3.47 30.49 ;
        RECT  3.21 30.8525 3.28 30.9875 ;
        RECT  3.4 30.0125 3.47 30.1475 ;
        RECT  3.3675 30.455 3.5025 30.525 ;
        RECT  3.21 31.865 3.28 31.935 ;
        RECT  3.4 31.865 3.47 31.935 ;
        RECT  3.21 31.5375 3.28 31.9 ;
        RECT  3.245 31.865 3.435 31.935 ;
        RECT  3.4 31.9 3.47 32.2425 ;
        RECT  3.21 31.5375 3.28 31.6725 ;
        RECT  3.4 32.3775 3.47 32.5125 ;
        RECT  3.3675 31.935 3.5025 32.005 ;
        RECT  3.21 33.145 3.28 33.215 ;
        RECT  3.4 33.145 3.47 33.215 ;
        RECT  3.21 33.18 3.28 33.5425 ;
        RECT  3.245 33.145 3.435 33.215 ;
        RECT  3.4 32.8375 3.47 33.18 ;
        RECT  3.21 33.5425 3.28 33.6775 ;
        RECT  3.4 32.7025 3.47 32.8375 ;
        RECT  3.3675 33.145 3.5025 33.215 ;
        RECT  3.21 34.555 3.28 34.625 ;
        RECT  3.4 34.555 3.47 34.625 ;
        RECT  3.21 34.2275 3.28 34.59 ;
        RECT  3.245 34.555 3.435 34.625 ;
        RECT  3.4 34.59 3.47 34.9325 ;
        RECT  3.21 34.2275 3.28 34.3625 ;
        RECT  3.4 35.0675 3.47 35.2025 ;
        RECT  3.3675 34.625 3.5025 34.695 ;
        RECT  3.21 35.835 3.28 35.905 ;
        RECT  3.4 35.835 3.47 35.905 ;
        RECT  3.21 35.87 3.28 36.2325 ;
        RECT  3.245 35.835 3.435 35.905 ;
        RECT  3.4 35.5275 3.47 35.87 ;
        RECT  3.21 36.2325 3.28 36.3675 ;
        RECT  3.4 35.3925 3.47 35.5275 ;
        RECT  3.3675 35.835 3.5025 35.905 ;
        RECT  3.21 37.245 3.28 37.315 ;
        RECT  3.4 37.245 3.47 37.315 ;
        RECT  3.21 36.9175 3.28 37.28 ;
        RECT  3.245 37.245 3.435 37.315 ;
        RECT  3.4 37.28 3.47 37.6225 ;
        RECT  3.21 36.9175 3.28 37.0525 ;
        RECT  3.4 37.7575 3.47 37.8925 ;
        RECT  3.3675 37.315 3.5025 37.385 ;
        RECT  3.21 38.525 3.28 38.595 ;
        RECT  3.4 38.525 3.47 38.595 ;
        RECT  3.21 38.56 3.28 38.9225 ;
        RECT  3.245 38.525 3.435 38.595 ;
        RECT  3.4 38.2175 3.47 38.56 ;
        RECT  3.21 38.9225 3.28 39.0575 ;
        RECT  3.4 38.0825 3.47 38.2175 ;
        RECT  3.3675 38.525 3.5025 38.595 ;
        RECT  3.21 39.935 3.28 40.005 ;
        RECT  3.4 39.935 3.47 40.005 ;
        RECT  3.21 39.6075 3.28 39.97 ;
        RECT  3.245 39.935 3.435 40.005 ;
        RECT  3.4 39.97 3.47 40.3125 ;
        RECT  3.21 39.6075 3.28 39.7425 ;
        RECT  3.4 40.4475 3.47 40.5825 ;
        RECT  3.3675 40.005 3.5025 40.075 ;
        RECT  1.5225 8.8775 1.6575 8.9475 ;
        RECT  1.6975 10.4025 1.8325 10.4725 ;
        RECT  1.8725 11.5675 2.0075 11.6375 ;
        RECT  2.0475 13.0925 2.1825 13.1625 ;
        RECT  2.2225 14.2575 2.3575 14.3275 ;
        RECT  2.3975 15.7825 2.5325 15.8525 ;
        RECT  2.5725 16.9475 2.7075 17.0175 ;
        RECT  2.7475 18.4725 2.8825 18.5425 ;
        RECT  1.5225 19.695 1.6575 19.765 ;
        RECT  2.2225 19.48 2.3575 19.55 ;
        RECT  1.5225 21.105 1.6575 21.175 ;
        RECT  2.3975 21.32 2.5325 21.39 ;
        RECT  1.5225 22.385 1.6575 22.455 ;
        RECT  2.5725 22.17 2.7075 22.24 ;
        RECT  1.5225 23.795 1.6575 23.865 ;
        RECT  2.7475 24.01 2.8825 24.08 ;
        RECT  1.6975 25.075 1.8325 25.145 ;
        RECT  2.2225 24.86 2.3575 24.93 ;
        RECT  1.6975 26.485 1.8325 26.555 ;
        RECT  2.3975 26.7 2.5325 26.77 ;
        RECT  1.6975 27.765 1.8325 27.835 ;
        RECT  2.5725 27.55 2.7075 27.62 ;
        RECT  1.6975 29.175 1.8325 29.245 ;
        RECT  2.7475 29.39 2.8825 29.46 ;
        RECT  1.8725 30.455 2.0075 30.525 ;
        RECT  2.2225 30.24 2.3575 30.31 ;
        RECT  1.8725 31.865 2.0075 31.935 ;
        RECT  2.3975 32.08 2.5325 32.15 ;
        RECT  1.8725 33.145 2.0075 33.215 ;
        RECT  2.5725 32.93 2.7075 33.0 ;
        RECT  1.8725 34.555 2.0075 34.625 ;
        RECT  2.7475 34.77 2.8825 34.84 ;
        RECT  2.0475 35.835 2.1825 35.905 ;
        RECT  2.2225 35.62 2.3575 35.69 ;
        RECT  2.0475 37.245 2.1825 37.315 ;
        RECT  2.3975 37.46 2.5325 37.53 ;
        RECT  2.0475 38.525 2.1825 38.595 ;
        RECT  2.5725 38.31 2.7075 38.38 ;
        RECT  2.0475 39.935 2.1825 40.005 ;
        RECT  2.7475 40.15 2.8825 40.22 ;
        RECT  4.77 19.48 4.84 19.55 ;
        RECT  4.77 19.445 4.84 19.515 ;
        RECT  4.805 19.48 5.7675 19.55 ;
        RECT  4.77 21.32 4.84 21.39 ;
        RECT  4.77 21.355 4.84 21.425 ;
        RECT  4.805 21.32 5.7675 21.39 ;
        RECT  4.77 22.17 4.84 22.24 ;
        RECT  4.77 22.135 4.84 22.205 ;
        RECT  4.805 22.17 5.7675 22.24 ;
        RECT  4.77 24.01 4.84 24.08 ;
        RECT  4.77 24.045 4.84 24.115 ;
        RECT  4.805 24.01 5.7675 24.08 ;
        RECT  4.77 24.86 4.84 24.93 ;
        RECT  4.77 24.825 4.84 24.895 ;
        RECT  4.805 24.86 5.7675 24.93 ;
        RECT  4.77 26.7 4.84 26.77 ;
        RECT  4.77 26.735 4.84 26.805 ;
        RECT  4.805 26.7 5.7675 26.77 ;
        RECT  4.77 27.55 4.84 27.62 ;
        RECT  4.77 27.515 4.84 27.585 ;
        RECT  4.805 27.55 5.7675 27.62 ;
        RECT  4.77 29.39 4.84 29.46 ;
        RECT  4.77 29.425 4.84 29.495 ;
        RECT  4.805 29.39 5.7675 29.46 ;
        RECT  4.77 30.24 4.84 30.31 ;
        RECT  4.77 30.205 4.84 30.275 ;
        RECT  4.805 30.24 5.7675 30.31 ;
        RECT  4.77 32.08 4.84 32.15 ;
        RECT  4.77 32.115 4.84 32.185 ;
        RECT  4.805 32.08 5.7675 32.15 ;
        RECT  4.77 32.93 4.84 33.0 ;
        RECT  4.77 32.895 4.84 32.965 ;
        RECT  4.805 32.93 5.7675 33.0 ;
        RECT  4.77 34.77 4.84 34.84 ;
        RECT  4.77 34.805 4.84 34.875 ;
        RECT  4.805 34.77 5.7675 34.84 ;
        RECT  4.77 35.62 4.84 35.69 ;
        RECT  4.77 35.585 4.84 35.655 ;
        RECT  4.805 35.62 5.7675 35.69 ;
        RECT  4.77 37.46 4.84 37.53 ;
        RECT  4.77 37.495 4.84 37.565 ;
        RECT  4.805 37.46 5.7675 37.53 ;
        RECT  4.77 38.31 4.84 38.38 ;
        RECT  4.77 38.275 4.84 38.345 ;
        RECT  4.805 38.31 5.7675 38.38 ;
        RECT  4.77 40.15 4.84 40.22 ;
        RECT  4.77 40.185 4.84 40.255 ;
        RECT  4.805 40.15 5.7675 40.22 ;
        RECT  4.63 19.09 4.7 40.61 ;
        RECT  5.705 19.695 5.775 19.765 ;
        RECT  5.895 19.695 5.965 19.765 ;
        RECT  5.705 19.73 5.775 20.0925 ;
        RECT  5.74 19.695 5.93 19.765 ;
        RECT  5.895 19.3875 5.965 19.73 ;
        RECT  5.705 20.0925 5.775 20.2275 ;
        RECT  5.895 19.2525 5.965 19.3875 ;
        RECT  5.8625 19.695 5.9975 19.765 ;
        RECT  4.63 19.605 4.7 19.74 ;
        RECT  4.77 19.3775 4.84 19.5125 ;
        RECT  5.6325 19.48 5.7675 19.55 ;
        RECT  5.705 21.105 5.775 21.175 ;
        RECT  5.895 21.105 5.965 21.175 ;
        RECT  5.705 20.7775 5.775 21.14 ;
        RECT  5.74 21.105 5.93 21.175 ;
        RECT  5.895 21.14 5.965 21.4825 ;
        RECT  5.705 20.7775 5.775 20.9125 ;
        RECT  5.895 21.6175 5.965 21.7525 ;
        RECT  5.8625 21.175 5.9975 21.245 ;
        RECT  4.63 21.13 4.7 21.265 ;
        RECT  4.77 21.3575 4.84 21.4925 ;
        RECT  5.6325 21.32 5.7675 21.39 ;
        RECT  5.705 22.385 5.775 22.455 ;
        RECT  5.895 22.385 5.965 22.455 ;
        RECT  5.705 22.42 5.775 22.7825 ;
        RECT  5.74 22.385 5.93 22.455 ;
        RECT  5.895 22.0775 5.965 22.42 ;
        RECT  5.705 22.7825 5.775 22.9175 ;
        RECT  5.895 21.9425 5.965 22.0775 ;
        RECT  5.8625 22.385 5.9975 22.455 ;
        RECT  4.63 22.295 4.7 22.43 ;
        RECT  4.77 22.0675 4.84 22.2025 ;
        RECT  5.6325 22.17 5.7675 22.24 ;
        RECT  5.705 23.795 5.775 23.865 ;
        RECT  5.895 23.795 5.965 23.865 ;
        RECT  5.705 23.4675 5.775 23.83 ;
        RECT  5.74 23.795 5.93 23.865 ;
        RECT  5.895 23.83 5.965 24.1725 ;
        RECT  5.705 23.4675 5.775 23.6025 ;
        RECT  5.895 24.3075 5.965 24.4425 ;
        RECT  5.8625 23.865 5.9975 23.935 ;
        RECT  4.63 23.82 4.7 23.955 ;
        RECT  4.77 24.0475 4.84 24.1825 ;
        RECT  5.6325 24.01 5.7675 24.08 ;
        RECT  5.705 25.075 5.775 25.145 ;
        RECT  5.895 25.075 5.965 25.145 ;
        RECT  5.705 25.11 5.775 25.4725 ;
        RECT  5.74 25.075 5.93 25.145 ;
        RECT  5.895 24.7675 5.965 25.11 ;
        RECT  5.705 25.4725 5.775 25.6075 ;
        RECT  5.895 24.6325 5.965 24.7675 ;
        RECT  5.8625 25.075 5.9975 25.145 ;
        RECT  4.63 24.985 4.7 25.12 ;
        RECT  4.77 24.7575 4.84 24.8925 ;
        RECT  5.6325 24.86 5.7675 24.93 ;
        RECT  5.705 26.485 5.775 26.555 ;
        RECT  5.895 26.485 5.965 26.555 ;
        RECT  5.705 26.1575 5.775 26.52 ;
        RECT  5.74 26.485 5.93 26.555 ;
        RECT  5.895 26.52 5.965 26.8625 ;
        RECT  5.705 26.1575 5.775 26.2925 ;
        RECT  5.895 26.9975 5.965 27.1325 ;
        RECT  5.8625 26.555 5.9975 26.625 ;
        RECT  4.63 26.51 4.7 26.645 ;
        RECT  4.77 26.7375 4.84 26.8725 ;
        RECT  5.6325 26.7 5.7675 26.77 ;
        RECT  5.705 27.765 5.775 27.835 ;
        RECT  5.895 27.765 5.965 27.835 ;
        RECT  5.705 27.8 5.775 28.1625 ;
        RECT  5.74 27.765 5.93 27.835 ;
        RECT  5.895 27.4575 5.965 27.8 ;
        RECT  5.705 28.1625 5.775 28.2975 ;
        RECT  5.895 27.3225 5.965 27.4575 ;
        RECT  5.8625 27.765 5.9975 27.835 ;
        RECT  4.63 27.675 4.7 27.81 ;
        RECT  4.77 27.4475 4.84 27.5825 ;
        RECT  5.6325 27.55 5.7675 27.62 ;
        RECT  5.705 29.175 5.775 29.245 ;
        RECT  5.895 29.175 5.965 29.245 ;
        RECT  5.705 28.8475 5.775 29.21 ;
        RECT  5.74 29.175 5.93 29.245 ;
        RECT  5.895 29.21 5.965 29.5525 ;
        RECT  5.705 28.8475 5.775 28.9825 ;
        RECT  5.895 29.6875 5.965 29.8225 ;
        RECT  5.8625 29.245 5.9975 29.315 ;
        RECT  4.63 29.2 4.7 29.335 ;
        RECT  4.77 29.4275 4.84 29.5625 ;
        RECT  5.6325 29.39 5.7675 29.46 ;
        RECT  5.705 30.455 5.775 30.525 ;
        RECT  5.895 30.455 5.965 30.525 ;
        RECT  5.705 30.49 5.775 30.8525 ;
        RECT  5.74 30.455 5.93 30.525 ;
        RECT  5.895 30.1475 5.965 30.49 ;
        RECT  5.705 30.8525 5.775 30.9875 ;
        RECT  5.895 30.0125 5.965 30.1475 ;
        RECT  5.8625 30.455 5.9975 30.525 ;
        RECT  4.63 30.365 4.7 30.5 ;
        RECT  4.77 30.1375 4.84 30.2725 ;
        RECT  5.6325 30.24 5.7675 30.31 ;
        RECT  5.705 31.865 5.775 31.935 ;
        RECT  5.895 31.865 5.965 31.935 ;
        RECT  5.705 31.5375 5.775 31.9 ;
        RECT  5.74 31.865 5.93 31.935 ;
        RECT  5.895 31.9 5.965 32.2425 ;
        RECT  5.705 31.5375 5.775 31.6725 ;
        RECT  5.895 32.3775 5.965 32.5125 ;
        RECT  5.8625 31.935 5.9975 32.005 ;
        RECT  4.63 31.89 4.7 32.025 ;
        RECT  4.77 32.1175 4.84 32.2525 ;
        RECT  5.6325 32.08 5.7675 32.15 ;
        RECT  5.705 33.145 5.775 33.215 ;
        RECT  5.895 33.145 5.965 33.215 ;
        RECT  5.705 33.18 5.775 33.5425 ;
        RECT  5.74 33.145 5.93 33.215 ;
        RECT  5.895 32.8375 5.965 33.18 ;
        RECT  5.705 33.5425 5.775 33.6775 ;
        RECT  5.895 32.7025 5.965 32.8375 ;
        RECT  5.8625 33.145 5.9975 33.215 ;
        RECT  4.63 33.055 4.7 33.19 ;
        RECT  4.77 32.8275 4.84 32.9625 ;
        RECT  5.6325 32.93 5.7675 33.0 ;
        RECT  5.705 34.555 5.775 34.625 ;
        RECT  5.895 34.555 5.965 34.625 ;
        RECT  5.705 34.2275 5.775 34.59 ;
        RECT  5.74 34.555 5.93 34.625 ;
        RECT  5.895 34.59 5.965 34.9325 ;
        RECT  5.705 34.2275 5.775 34.3625 ;
        RECT  5.895 35.0675 5.965 35.2025 ;
        RECT  5.8625 34.625 5.9975 34.695 ;
        RECT  4.63 34.58 4.7 34.715 ;
        RECT  4.77 34.8075 4.84 34.9425 ;
        RECT  5.6325 34.77 5.7675 34.84 ;
        RECT  5.705 35.835 5.775 35.905 ;
        RECT  5.895 35.835 5.965 35.905 ;
        RECT  5.705 35.87 5.775 36.2325 ;
        RECT  5.74 35.835 5.93 35.905 ;
        RECT  5.895 35.5275 5.965 35.87 ;
        RECT  5.705 36.2325 5.775 36.3675 ;
        RECT  5.895 35.3925 5.965 35.5275 ;
        RECT  5.8625 35.835 5.9975 35.905 ;
        RECT  4.63 35.745 4.7 35.88 ;
        RECT  4.77 35.5175 4.84 35.6525 ;
        RECT  5.6325 35.62 5.7675 35.69 ;
        RECT  5.705 37.245 5.775 37.315 ;
        RECT  5.895 37.245 5.965 37.315 ;
        RECT  5.705 36.9175 5.775 37.28 ;
        RECT  5.74 37.245 5.93 37.315 ;
        RECT  5.895 37.28 5.965 37.6225 ;
        RECT  5.705 36.9175 5.775 37.0525 ;
        RECT  5.895 37.7575 5.965 37.8925 ;
        RECT  5.8625 37.315 5.9975 37.385 ;
        RECT  4.63 37.27 4.7 37.405 ;
        RECT  4.77 37.4975 4.84 37.6325 ;
        RECT  5.6325 37.46 5.7675 37.53 ;
        RECT  5.705 38.525 5.775 38.595 ;
        RECT  5.895 38.525 5.965 38.595 ;
        RECT  5.705 38.56 5.775 38.9225 ;
        RECT  5.74 38.525 5.93 38.595 ;
        RECT  5.895 38.2175 5.965 38.56 ;
        RECT  5.705 38.9225 5.775 39.0575 ;
        RECT  5.895 38.0825 5.965 38.2175 ;
        RECT  5.8625 38.525 5.9975 38.595 ;
        RECT  4.63 38.435 4.7 38.57 ;
        RECT  4.77 38.2075 4.84 38.3425 ;
        RECT  5.6325 38.31 5.7675 38.38 ;
        RECT  5.705 39.935 5.775 40.005 ;
        RECT  5.895 39.935 5.965 40.005 ;
        RECT  5.705 39.6075 5.775 39.97 ;
        RECT  5.74 39.935 5.93 40.005 ;
        RECT  5.895 39.97 5.965 40.3125 ;
        RECT  5.705 39.6075 5.775 39.7425 ;
        RECT  5.895 40.4475 5.965 40.5825 ;
        RECT  5.8625 40.005 5.9975 40.075 ;
        RECT  4.63 39.96 4.7 40.095 ;
        RECT  4.77 40.1875 4.84 40.3225 ;
        RECT  5.6325 40.15 5.7675 40.22 ;
        RECT  6.2325 6.6725 6.92 6.7425 ;
        RECT  0.48 5.4175 0.625 5.4875 ;
        RECT  6.2325 6.2775 6.92 6.3475 ;
        RECT  6.2325 5.2625 6.92 5.3325 ;
        RECT  0.48 6.8275 0.625 6.8975 ;
        RECT  0.48 7.5325 0.625 7.6025 ;
        RECT  0.48 6.1225 0.625 6.1925 ;
        RECT  0.48 7.885 6.92 7.955 ;
        RECT  0.48 7.18 6.92 7.25 ;
        RECT  0.48 6.475 6.92 6.545 ;
        RECT  0.48 5.77 6.92 5.84 ;
        RECT  0.48 5.065 6.92 5.135 ;
        RECT  6.2325 7.6875 6.92 7.7575 ;
        RECT  6.65 7.5325 6.92 7.6025 ;
        RECT  6.65 6.8275 6.92 6.8975 ;
        RECT  6.65 5.4175 6.92 5.4875 ;
        RECT  6.65 6.1225 6.92 6.1925 ;
        RECT  6.1825 7.6875 6.3175 7.7575 ;
        RECT  1.005 7.18 1.14 7.25 ;
        RECT  5.0875 7.3225 5.2225 7.3925 ;
        RECT  3.48 7.32 3.615 7.39 ;
        RECT  2.0825 7.32 2.2175 7.39 ;
        RECT  0.865 7.885 1.0 7.955 ;
        RECT  0.48 7.5325 0.62 7.6025 ;
        RECT  3.9425 7.18 4.0775 7.25 ;
        RECT  2.7475 7.685 2.8825 7.755 ;
        RECT  6.44 7.32 6.575 7.39 ;
        RECT  5.93 7.4975 6.065 7.5675 ;
        RECT  5.5175 7.18 5.6525 7.25 ;
        RECT  0.815 7.18 0.95 7.25 ;
        RECT  2.5575 7.18 2.6925 7.25 ;
        RECT  2.3575 7.685 2.4925 7.755 ;
        RECT  2.3575 7.4975 2.4925 7.5675 ;
        RECT  2.97 7.4975 3.105 7.5675 ;
        RECT  5.3175 7.6875 5.4525 7.7575 ;
        RECT  5.3175 7.4975 5.4525 7.5675 ;
        RECT  6.65 7.39 6.72 7.5325 ;
        RECT  0.48 7.5325 0.625 7.6025 ;
        RECT  0.555 7.39 0.625 7.5375 ;
        RECT  6.65 7.5325 6.92 7.6025 ;
        RECT  6.4425 7.89 6.5025 7.9525 ;
        RECT  0.48 7.885 6.92 7.955 ;
        RECT  6.855 7.535 6.915 7.6 ;
        RECT  6.44 7.32 6.72 7.39 ;
        RECT  0.555 7.32 2.2175 7.39 ;
        RECT  6.2325 7.6875 6.92 7.7575 ;
        RECT  3.615 7.32 5.2225 7.39 ;
        RECT  5.3175 7.4975 6.035 7.5675 ;
        RECT  2.3575 7.685 2.8825 7.755 ;
        RECT  6.7825 7.69 6.8425 7.7525 ;
        RECT  5.3175 7.6875 6.2575 7.7575 ;
        RECT  0.485 7.535 0.55 7.6025 ;
        RECT  0.48 7.18 6.92 7.25 ;
        RECT  2.3575 7.4975 3.075 7.5675 ;
        RECT  0.48 7.5325 0.625 7.6025 ;
        RECT  6.65 7.5325 6.92 7.6025 ;
        RECT  6.2325 7.6875 6.92 7.7575 ;
        RECT  0.48 7.885 6.92 7.955 ;
        RECT  0.48 7.18 6.92 7.25 ;
        RECT  6.1825 6.6725 6.3175 6.7425 ;
        RECT  1.005 7.18 1.14 7.25 ;
        RECT  5.0875 7.0375 5.2225 7.1075 ;
        RECT  3.48 7.04 3.615 7.11 ;
        RECT  2.0825 7.04 2.2175 7.11 ;
        RECT  0.865 6.475 1.0 6.545 ;
        RECT  0.48 6.8275 0.62 6.8975 ;
        RECT  3.9425 7.18 4.0775 7.25 ;
        RECT  2.7475 6.675 2.8825 6.745 ;
        RECT  6.44 7.04 6.575 7.11 ;
        RECT  5.93 6.8625 6.065 6.9325 ;
        RECT  5.5175 7.18 5.6525 7.25 ;
        RECT  0.815 7.18 0.95 7.25 ;
        RECT  2.5575 7.18 2.6925 7.25 ;
        RECT  2.3575 6.675 2.4925 6.745 ;
        RECT  2.3575 6.8625 2.4925 6.9325 ;
        RECT  2.97 6.8625 3.105 6.9325 ;
        RECT  5.3175 6.6725 5.4525 6.7425 ;
        RECT  5.3175 6.8625 5.4525 6.9325 ;
        RECT  6.65 6.8975 6.72 7.04 ;
        RECT  0.48 6.8275 0.625 6.8975 ;
        RECT  0.555 6.8925 0.625 7.04 ;
        RECT  6.65 6.8275 6.92 6.8975 ;
        RECT  6.4425 6.4775 6.5025 6.54 ;
        RECT  0.48 6.475 6.92 6.545 ;
        RECT  6.855 6.83 6.915 6.895 ;
        RECT  6.44 7.04 6.72 7.11 ;
        RECT  0.555 7.04 2.2175 7.11 ;
        RECT  6.2325 6.6725 6.92 6.7425 ;
        RECT  3.615 7.04 5.2225 7.11 ;
        RECT  5.3175 6.8625 6.035 6.9325 ;
        RECT  2.3575 6.675 2.8825 6.745 ;
        RECT  6.7825 6.6775 6.8425 6.74 ;
        RECT  5.3175 6.6725 6.2575 6.7425 ;
        RECT  0.485 6.8275 0.55 6.895 ;
        RECT  0.48 7.18 6.92 7.25 ;
        RECT  2.3575 6.8625 3.075 6.9325 ;
        RECT  0.48 6.8275 0.625 6.8975 ;
        RECT  6.65 6.8275 6.92 6.8975 ;
        RECT  6.2325 6.6725 6.92 6.7425 ;
        RECT  0.48 6.475 6.92 6.545 ;
        RECT  0.48 7.18 6.92 7.25 ;
        RECT  6.1825 6.2775 6.3175 6.3475 ;
        RECT  1.005 5.77 1.14 5.84 ;
        RECT  5.0875 5.9125 5.2225 5.9825 ;
        RECT  3.48 5.91 3.615 5.98 ;
        RECT  2.0825 5.91 2.2175 5.98 ;
        RECT  0.865 6.475 1.0 6.545 ;
        RECT  0.48 6.1225 0.62 6.1925 ;
        RECT  3.9425 5.77 4.0775 5.84 ;
        RECT  2.7475 6.275 2.8825 6.345 ;
        RECT  6.44 5.91 6.575 5.98 ;
        RECT  5.93 6.0875 6.065 6.1575 ;
        RECT  5.5175 5.77 5.6525 5.84 ;
        RECT  0.815 5.77 0.95 5.84 ;
        RECT  2.5575 5.77 2.6925 5.84 ;
        RECT  2.3575 6.275 2.4925 6.345 ;
        RECT  2.3575 6.0875 2.4925 6.1575 ;
        RECT  2.97 6.0875 3.105 6.1575 ;
        RECT  5.3175 6.2775 5.4525 6.3475 ;
        RECT  5.3175 6.0875 5.4525 6.1575 ;
        RECT  6.65 5.98 6.72 6.1225 ;
        RECT  0.48 6.1225 0.625 6.1925 ;
        RECT  0.555 5.98 0.625 6.1275 ;
        RECT  6.65 6.1225 6.92 6.1925 ;
        RECT  6.4425 6.48 6.5025 6.5425 ;
        RECT  0.48 6.475 6.92 6.545 ;
        RECT  6.855 6.125 6.915 6.19 ;
        RECT  6.44 5.91 6.72 5.98 ;
        RECT  0.555 5.91 2.2175 5.98 ;
        RECT  6.2325 6.2775 6.92 6.3475 ;
        RECT  3.615 5.91 5.2225 5.98 ;
        RECT  5.3175 6.0875 6.035 6.1575 ;
        RECT  2.3575 6.275 2.8825 6.345 ;
        RECT  6.7825 6.28 6.8425 6.3425 ;
        RECT  5.3175 6.2775 6.2575 6.3475 ;
        RECT  0.485 6.125 0.55 6.1925 ;
        RECT  0.48 5.77 6.92 5.84 ;
        RECT  2.3575 6.0875 3.075 6.1575 ;
        RECT  0.48 6.1225 0.625 6.1925 ;
        RECT  6.65 6.1225 6.92 6.1925 ;
        RECT  6.2325 6.2775 6.92 6.3475 ;
        RECT  0.48 6.475 6.92 6.545 ;
        RECT  0.48 5.77 6.92 5.84 ;
        RECT  6.1825 5.2625 6.3175 5.3325 ;
        RECT  1.005 5.77 1.14 5.84 ;
        RECT  5.0875 5.6275 5.2225 5.6975 ;
        RECT  3.48 5.63 3.615 5.7 ;
        RECT  2.0825 5.63 2.2175 5.7 ;
        RECT  0.865 5.065 1.0 5.135 ;
        RECT  0.48 5.4175 0.62 5.4875 ;
        RECT  3.9425 5.77 4.0775 5.84 ;
        RECT  2.7475 5.265 2.8825 5.335 ;
        RECT  6.44 5.63 6.575 5.7 ;
        RECT  5.93 5.4525 6.065 5.5225 ;
        RECT  5.5175 5.77 5.6525 5.84 ;
        RECT  0.815 5.77 0.95 5.84 ;
        RECT  2.5575 5.77 2.6925 5.84 ;
        RECT  2.3575 5.265 2.4925 5.335 ;
        RECT  2.3575 5.4525 2.4925 5.5225 ;
        RECT  2.97 5.4525 3.105 5.5225 ;
        RECT  5.3175 5.2625 5.4525 5.3325 ;
        RECT  5.3175 5.4525 5.4525 5.5225 ;
        RECT  6.65 5.4875 6.72 5.63 ;
        RECT  0.48 5.4175 0.625 5.4875 ;
        RECT  0.555 5.4825 0.625 5.63 ;
        RECT  6.65 5.4175 6.92 5.4875 ;
        RECT  6.4425 5.0675 6.5025 5.13 ;
        RECT  0.48 5.065 6.92 5.135 ;
        RECT  6.855 5.42 6.915 5.485 ;
        RECT  6.44 5.63 6.72 5.7 ;
        RECT  0.555 5.63 2.2175 5.7 ;
        RECT  6.2325 5.2625 6.92 5.3325 ;
        RECT  3.615 5.63 5.2225 5.7 ;
        RECT  5.3175 5.4525 6.035 5.5225 ;
        RECT  2.3575 5.265 2.8825 5.335 ;
        RECT  6.7825 5.2675 6.8425 5.33 ;
        RECT  5.3175 5.2625 6.2575 5.3325 ;
        RECT  0.485 5.4175 0.55 5.485 ;
        RECT  0.48 5.77 6.92 5.84 ;
        RECT  2.3575 5.4525 3.075 5.5225 ;
        RECT  0.48 5.4175 0.625 5.4875 ;
        RECT  6.65 5.4175 6.92 5.4875 ;
        RECT  6.2325 5.2625 6.92 5.3325 ;
        RECT  0.48 5.065 6.92 5.135 ;
        RECT  0.48 5.77 6.92 5.84 ;
        RECT  10.4525 0.44 10.5225 0.575 ;
        RECT  11.1575 0.44 11.2275 0.575 ;
        RECT  10.6625 0.0 10.7325 0.135 ;
        RECT  11.3675 0.0 11.4375 0.135 ;
        RECT  8.2525 19.055 8.3875 19.125 ;
        RECT  8.2525 21.745 8.3875 21.815 ;
        RECT  8.2525 24.435 8.3875 24.505 ;
        RECT  8.2525 27.125 8.3875 27.195 ;
        RECT  8.2525 29.815 8.3875 29.885 ;
        RECT  8.2525 32.505 8.3875 32.575 ;
        RECT  8.2525 35.195 8.3875 35.265 ;
        RECT  8.2525 37.885 8.3875 37.955 ;
        RECT  8.2525 40.575 8.3875 40.645 ;
        RECT  6.785 8.5 6.92 8.57 ;
        RECT  7.195 8.5 7.33 8.57 ;
        RECT  6.51 9.845 6.645 9.915 ;
        RECT  7.4 9.845 7.535 9.915 ;
        RECT  6.785 13.88 6.92 13.95 ;
        RECT  7.605 13.88 7.74 13.95 ;
        RECT  6.51 15.225 6.645 15.295 ;
        RECT  7.81 15.225 7.945 15.295 ;
        RECT  6.99 8.295 7.125 8.365 ;
        RECT  6.99 8.295 7.125 8.365 ;
        RECT  8.185 8.295 8.32 8.365 ;
        RECT  6.99 10.985 7.125 11.055 ;
        RECT  6.99 10.985 7.125 11.055 ;
        RECT  8.185 10.985 8.32 11.055 ;
        RECT  6.99 13.675 7.125 13.745 ;
        RECT  6.99 13.675 7.125 13.745 ;
        RECT  8.185 13.675 8.32 13.745 ;
        RECT  6.99 16.365 7.125 16.435 ;
        RECT  6.99 16.365 7.125 16.435 ;
        RECT  8.185 16.365 8.32 16.435 ;
        RECT  6.8525 7.5325 6.9875 7.6025 ;
        RECT  7.195 7.5325 7.33 7.6025 ;
        RECT  6.8525 6.8275 6.9875 6.8975 ;
        RECT  7.4 6.8275 7.535 6.8975 ;
        RECT  6.8525 6.1225 6.9875 6.1925 ;
        RECT  7.605 6.1225 7.74 6.1925 ;
        RECT  6.8525 5.4175 6.9875 5.4875 ;
        RECT  7.81 5.4175 7.945 5.4875 ;
        RECT  6.92 7.885 7.055 7.955 ;
        RECT  8.2525 7.885 8.3875 7.955 ;
        RECT  6.92 7.18 7.055 7.25 ;
        RECT  8.2525 7.18 8.3875 7.25 ;
        RECT  6.92 6.475 7.055 6.545 ;
        RECT  8.2525 6.475 8.3875 6.545 ;
        RECT  6.92 5.77 7.055 5.84 ;
        RECT  8.2525 5.77 8.3875 5.84 ;
        RECT  6.92 5.065 7.055 5.135 ;
        RECT  8.2525 5.065 8.3875 5.135 ;
        RECT  9.39 3.7925 9.525 3.8625 ;
        RECT  8.98 1.6075 9.115 1.6775 ;
        RECT  9.185 3.155 9.32 3.225 ;
        RECT  9.39 41.475 9.525 41.545 ;
        RECT  9.595 10.295 9.73 10.365 ;
        RECT  9.8 14.32 9.935 14.39 ;
        RECT  8.775 8.09 8.91 8.16 ;
        RECT  4.5975 40.78 4.7325 40.85 ;
        RECT  8.775 40.78 8.91 40.85 ;
        RECT  8.4675 3.025 8.6025 3.095 ;
        RECT  8.4675 14.45 8.6025 14.52 ;
        RECT  8.4675 3.9525 8.6025 4.0225 ;
        RECT  8.4675 11.2275 8.6025 11.2975 ;
        RECT  -4.175 26.49 -0.14 26.56 ;
        RECT  -4.175 26.695 -0.14 26.765 ;
        RECT  -4.175 26.9 -0.14 26.97 ;
        RECT  -4.175 27.31 -0.14 27.38 ;
        RECT  -1.725 19.4675 -1.655 26.115 ;
        RECT  -0.345 26.285 -0.14 26.355 ;
        RECT  -1.485 27.105 -1.28 27.175 ;
        RECT  -2.83 26.285 -2.625 26.355 ;
        RECT  -4.175 27.105 -3.97 27.175 ;
        RECT  -4.175 27.515 -0.14 27.585 ;
        RECT  -3.4125 31.14 -0.14 31.21 ;
        RECT  -4.175 26.08 -0.14 26.15 ;
        RECT  -2.19 29.955 -0.14 30.025 ;
        RECT  -4.175 27.105 -0.14 27.175 ;
        RECT  -4.175 26.285 -0.14 26.355 ;
        RECT  -2.2475 30.18 -0.14 30.25 ;
        RECT  -2.245 28.81 -0.14 28.88 ;
        RECT  -2.8325 24.9825 -2.7625 25.67 ;
        RECT  -2.4375 24.9825 -2.3675 25.67 ;
        RECT  -2.9875 19.23 -2.9175 19.375 ;
        RECT  -3.6925 19.23 -3.6225 19.375 ;
        RECT  -2.2825 19.23 -2.2125 19.375 ;
        RECT  -4.045 19.23 -3.975 25.67 ;
        RECT  -3.34 19.23 -3.27 25.67 ;
        RECT  -2.635 19.23 -2.565 25.67 ;
        RECT  -1.93 19.23 -1.86 25.67 ;
        RECT  -3.8475 24.9825 -3.7775 25.67 ;
        RECT  -3.6925 25.4 -3.6225 25.67 ;
        RECT  -2.9875 25.4 -2.9175 25.67 ;
        RECT  -2.2825 25.4 -2.2125 25.67 ;
        RECT  -3.8475 24.9325 -3.7775 25.0675 ;
        RECT  -3.34 19.755 -3.27 19.89 ;
        RECT  -3.4825 23.8375 -3.4125 23.9725 ;
        RECT  -3.48 22.23 -3.41 22.365 ;
        RECT  -3.48 20.8325 -3.41 20.9675 ;
        RECT  -4.045 19.615 -3.975 19.75 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -3.34 22.6925 -3.27 22.8275 ;
        RECT  -3.845 21.4975 -3.775 21.6325 ;
        RECT  -3.48 25.19 -3.41 25.325 ;
        RECT  -3.6575 24.68 -3.5875 24.815 ;
        RECT  -3.34 24.2675 -3.27 24.4025 ;
        RECT  -3.34 19.565 -3.27 19.7 ;
        RECT  -3.34 21.3075 -3.27 21.4425 ;
        RECT  -3.845 21.1075 -3.775 21.2425 ;
        RECT  -3.6575 21.1075 -3.5875 21.2425 ;
        RECT  -3.6575 21.72 -3.5875 21.855 ;
        RECT  -3.8475 24.0675 -3.7775 24.2025 ;
        RECT  -3.6575 24.0675 -3.5875 24.2025 ;
        RECT  -3.6225 25.4 -3.48 25.47 ;
        RECT  -3.6925 19.23 -3.6225 19.375 ;
        RECT  -3.6275 19.305 -3.48 19.375 ;
        RECT  -3.6925 25.4 -3.6225 25.67 ;
        RECT  -4.0425 25.1925 -3.98 25.2525 ;
        RECT  -4.045 19.23 -3.975 25.67 ;
        RECT  -3.69 25.605 -3.625 25.665 ;
        RECT  -3.48 25.19 -3.41 25.47 ;
        RECT  -3.48 19.305 -3.41 20.9675 ;
        RECT  -3.8475 24.9825 -3.7775 25.67 ;
        RECT  -3.48 22.365 -3.41 23.9725 ;
        RECT  -3.6575 24.0675 -3.5875 24.785 ;
        RECT  -3.845 21.1075 -3.775 21.6325 ;
        RECT  -3.8425 25.5325 -3.78 25.5925 ;
        RECT  -3.8475 24.0675 -3.7775 25.0075 ;
        RECT  -3.6925 19.235 -3.625 19.3 ;
        RECT  -3.34 19.23 -3.27 25.67 ;
        RECT  -3.6575 21.1075 -3.5875 21.825 ;
        RECT  -3.6925 19.23 -3.6225 19.375 ;
        RECT  -3.6925 25.4 -3.6225 25.67 ;
        RECT  -3.8475 24.9825 -3.7775 25.67 ;
        RECT  -4.045 19.23 -3.975 25.67 ;
        RECT  -3.34 19.23 -3.27 25.67 ;
        RECT  -2.8325 24.9325 -2.7625 25.0675 ;
        RECT  -3.34 19.755 -3.27 19.89 ;
        RECT  -3.1975 23.8375 -3.1275 23.9725 ;
        RECT  -3.2 22.23 -3.13 22.365 ;
        RECT  -3.2 20.8325 -3.13 20.9675 ;
        RECT  -2.635 19.615 -2.565 19.75 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -3.34 22.6925 -3.27 22.8275 ;
        RECT  -2.835 21.4975 -2.765 21.6325 ;
        RECT  -3.2 25.19 -3.13 25.325 ;
        RECT  -3.0225 24.68 -2.9525 24.815 ;
        RECT  -3.34 24.2675 -3.27 24.4025 ;
        RECT  -3.34 19.565 -3.27 19.7 ;
        RECT  -3.34 21.3075 -3.27 21.4425 ;
        RECT  -2.835 21.1075 -2.765 21.2425 ;
        RECT  -3.0225 21.1075 -2.9525 21.2425 ;
        RECT  -3.0225 21.72 -2.9525 21.855 ;
        RECT  -2.8325 24.0675 -2.7625 24.2025 ;
        RECT  -3.0225 24.0675 -2.9525 24.2025 ;
        RECT  -3.13 25.4 -2.9875 25.47 ;
        RECT  -2.9875 19.23 -2.9175 19.375 ;
        RECT  -3.13 19.305 -2.9825 19.375 ;
        RECT  -2.9875 25.4 -2.9175 25.67 ;
        RECT  -2.63 25.1925 -2.5675 25.2525 ;
        RECT  -2.635 19.23 -2.565 25.67 ;
        RECT  -2.985 25.605 -2.92 25.665 ;
        RECT  -3.2 25.19 -3.13 25.47 ;
        RECT  -3.2 19.305 -3.13 20.9675 ;
        RECT  -2.8325 24.9825 -2.7625 25.67 ;
        RECT  -3.2 22.365 -3.13 23.9725 ;
        RECT  -3.0225 24.0675 -2.9525 24.785 ;
        RECT  -2.835 21.1075 -2.765 21.6325 ;
        RECT  -2.83 25.5325 -2.7675 25.5925 ;
        RECT  -2.8325 24.0675 -2.7625 25.0075 ;
        RECT  -2.985 19.235 -2.9175 19.3 ;
        RECT  -3.34 19.23 -3.27 25.67 ;
        RECT  -3.0225 21.1075 -2.9525 21.825 ;
        RECT  -2.9875 19.23 -2.9175 19.375 ;
        RECT  -2.9875 25.4 -2.9175 25.67 ;
        RECT  -2.8325 24.9825 -2.7625 25.67 ;
        RECT  -2.635 19.23 -2.565 25.67 ;
        RECT  -3.34 19.23 -3.27 25.67 ;
        RECT  -2.4375 24.9325 -2.3675 25.0675 ;
        RECT  -1.93 19.755 -1.86 19.89 ;
        RECT  -2.0725 23.8375 -2.0025 23.9725 ;
        RECT  -2.07 22.23 -2.0 22.365 ;
        RECT  -2.07 20.8325 -2.0 20.9675 ;
        RECT  -2.635 19.615 -2.565 19.75 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -1.93 22.6925 -1.86 22.8275 ;
        RECT  -2.435 21.4975 -2.365 21.6325 ;
        RECT  -2.07 25.19 -2.0 25.325 ;
        RECT  -2.2475 24.68 -2.1775 24.815 ;
        RECT  -1.93 24.2675 -1.86 24.4025 ;
        RECT  -1.93 19.565 -1.86 19.7 ;
        RECT  -1.93 21.3075 -1.86 21.4425 ;
        RECT  -2.435 21.1075 -2.365 21.2425 ;
        RECT  -2.2475 21.1075 -2.1775 21.2425 ;
        RECT  -2.2475 21.72 -2.1775 21.855 ;
        RECT  -2.4375 24.0675 -2.3675 24.2025 ;
        RECT  -2.2475 24.0675 -2.1775 24.2025 ;
        RECT  -2.2125 25.4 -2.07 25.47 ;
        RECT  -2.2825 19.23 -2.2125 19.375 ;
        RECT  -2.2175 19.305 -2.07 19.375 ;
        RECT  -2.2825 25.4 -2.2125 25.67 ;
        RECT  -2.6325 25.1925 -2.57 25.2525 ;
        RECT  -2.635 19.23 -2.565 25.67 ;
        RECT  -2.28 25.605 -2.215 25.665 ;
        RECT  -2.07 25.19 -2.0 25.47 ;
        RECT  -2.07 19.305 -2.0 20.9675 ;
        RECT  -2.4375 24.9825 -2.3675 25.67 ;
        RECT  -2.07 22.365 -2.0 23.9725 ;
        RECT  -2.2475 24.0675 -2.1775 24.785 ;
        RECT  -2.435 21.1075 -2.365 21.6325 ;
        RECT  -2.4325 25.5325 -2.37 25.5925 ;
        RECT  -2.4375 24.0675 -2.3675 25.0075 ;
        RECT  -2.2825 19.235 -2.215 19.3 ;
        RECT  -1.93 19.23 -1.86 25.67 ;
        RECT  -2.2475 21.1075 -2.1775 21.825 ;
        RECT  -2.2825 19.23 -2.2125 19.375 ;
        RECT  -2.2825 25.4 -2.2125 25.67 ;
        RECT  -2.4375 24.9825 -2.3675 25.67 ;
        RECT  -2.635 19.23 -2.565 25.67 ;
        RECT  -1.93 19.23 -1.86 25.67 ;
        RECT  -1.1425 28.56 -0.4825 28.63 ;
        RECT  -0.9525 28.18 -0.8825 28.25 ;
        RECT  -0.9525 28.56 -0.8825 28.63 ;
        RECT  -1.1425 28.18 -0.9175 28.25 ;
        RECT  -0.9525 28.215 -0.8825 28.595 ;
        RECT  -0.9175 28.56 -0.4825 28.63 ;
        RECT  -1.2775 28.18 -1.1425 28.25 ;
        RECT  -1.2775 28.56 -1.1425 28.63 ;
        RECT  -0.4825 28.56 -0.3475 28.63 ;
        RECT  -0.985 28.56 -0.85 28.63 ;
        RECT  -2.28 28.37 -2.21 28.44 ;
        RECT  -2.245 28.37 -1.895 28.44 ;
        RECT  -2.28 28.405 -2.21 28.475 ;
        RECT  -2.68 28.37 -2.61 28.44 ;
        RECT  -2.68 28.2475 -2.61 28.405 ;
        RECT  -2.645 28.37 -2.245 28.44 ;
        RECT  -2.03 28.37 -1.895 28.44 ;
        RECT  -2.75 28.1475 -2.68 28.2825 ;
        RECT  -2.35 28.4075 -2.28 28.5425 ;
        RECT  -2.225 29.325 -2.155 29.395 ;
        RECT  -2.225 29.515 -2.155 29.585 ;
        RECT  -2.19 29.325 -1.8275 29.395 ;
        RECT  -2.225 29.36 -2.155 29.55 ;
        RECT  -2.5325 29.515 -2.19 29.585 ;
        RECT  -1.9625 29.325 -1.8275 29.395 ;
        RECT  -2.8025 29.515 -2.6675 29.585 ;
        RECT  -2.295 29.4825 -2.225 29.6175 ;
        RECT  -3.8325 29.12 -3.1725 29.19 ;
        RECT  -3.6425 28.74 -3.5725 28.81 ;
        RECT  -3.6425 29.12 -3.5725 29.19 ;
        RECT  -3.8325 28.74 -3.6075 28.81 ;
        RECT  -3.6425 28.775 -3.5725 29.155 ;
        RECT  -3.6075 29.12 -3.1725 29.19 ;
        RECT  -3.9675 28.74 -3.8325 28.81 ;
        RECT  -3.9675 29.12 -3.8325 29.19 ;
        RECT  -3.1725 29.12 -3.0375 29.19 ;
        RECT  -3.675 29.12 -3.54 29.19 ;
        RECT  -3.8475 25.6025 -3.7775 25.7375 ;
        RECT  -3.8475 27.2775 -3.7775 27.4125 ;
        RECT  -3.6925 25.6025 -3.6225 25.7375 ;
        RECT  -3.6925 26.4575 -3.6225 26.5925 ;
        RECT  -2.8325 25.6025 -2.7625 25.7375 ;
        RECT  -2.8325 26.6625 -2.7625 26.7975 ;
        RECT  -2.4375 25.6025 -2.3675 25.7375 ;
        RECT  -2.4375 26.8675 -2.3675 27.0025 ;
        RECT  -4.045 25.6025 -3.975 25.7375 ;
        RECT  -4.045 26.2525 -3.975 26.3875 ;
        RECT  -3.34 25.6025 -3.27 25.7375 ;
        RECT  -3.34 26.2525 -3.27 26.3875 ;
        RECT  -2.635 25.6025 -2.565 25.7375 ;
        RECT  -2.635 26.2525 -2.565 26.3875 ;
        RECT  -1.93 25.6025 -1.86 25.7375 ;
        RECT  -1.93 26.2525 -1.86 26.3875 ;
        RECT  -2.865 31.895 -2.795 36.695 ;
        RECT  -2.865 32.455 -2.795 32.66 ;
        RECT  -2.865 32.66 -2.795 36.795 ;
        RECT  -3.275 36.59 -3.205 36.795 ;
        RECT  -3.0375 32.0625 -2.9675 32.66 ;
        RECT  -3.46 32.0625 -3.39 32.3425 ;
        RECT  -0.7575 33.4175 -0.6875 33.8125 ;
        RECT  -1.52 33.2175 -1.45 33.2875 ;
        RECT  -1.52 33.1375 -1.45 33.2075 ;
        RECT  -1.485 33.2175 -0.7225 33.2875 ;
        RECT  -1.52 33.1725 -1.45 33.2525 ;
        RECT  -2.2475 33.1375 -1.485 33.2075 ;
        RECT  -2.2825 33.3375 -2.2125 33.7325 ;
        RECT  -0.79 33.3825 -0.655 33.4525 ;
        RECT  -2.315 33.1375 -2.18 33.2075 ;
        RECT  -2.315 33.6975 -2.18 33.7675 ;
        RECT  -0.79 33.7775 -0.655 33.8475 ;
        RECT  -0.79 33.2175 -0.655 33.2875 ;
        RECT  -2.315 33.3025 -2.18 33.3725 ;
        RECT  -3.275 34.0625 -3.205 34.1975 ;
        RECT  -3.98 34.5375 -3.91 34.6725 ;
        RECT  -3.275 34.5375 -3.205 34.6725 ;
        RECT  -3.7275 34.0575 -3.6575 34.1925 ;
        RECT  -3.5275 34.0625 -3.4575 34.1975 ;
        RECT  -4.0125 33.765 -3.8775 33.835 ;
        RECT  -3.3075 33.765 -3.1725 33.835 ;
        RECT  -3.795 33.7675 -3.725 33.8325 ;
        RECT  -3.46 33.7675 -3.39 33.8325 ;
        RECT  -3.275 33.765 -3.205 33.835 ;
        RECT  -3.46 33.7 -3.39 35.2575 ;
        RECT  -3.795 33.7 -3.725 35.265 ;
        RECT  -3.98 33.7 -3.91 35.2675 ;
        RECT  -3.275 33.7 -3.205 35.245 ;
        RECT  -3.46 33.7 -3.39 35.2575 ;
        RECT  -3.275 33.7 -3.205 35.245 ;
        RECT  -3.795 33.7 -3.725 35.265 ;
        RECT  -3.46 31.01 -3.39 33.9 ;
        RECT  -3.275 31.01 -3.205 33.9 ;
        RECT  -3.98 31.01 -3.91 33.9 ;
        RECT  -3.795 31.01 -3.725 33.9 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.3075 33.765 -3.1725 33.835 ;
        RECT  -4.0125 33.765 -3.8775 33.835 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.53 33.4075 -3.46 33.5425 ;
        RECT  -3.275 32.915 -3.205 33.05 ;
        RECT  -3.275 32.915 -3.205 33.05 ;
        RECT  -3.275 32.915 -3.205 33.05 ;
        RECT  -3.275 32.915 -3.205 33.05 ;
        RECT  -3.275 32.915 -3.205 33.05 ;
        RECT  -3.275 32.915 -3.205 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.725 33.4075 -3.655 33.5425 ;
        RECT  -4.0125 33.765 -3.8775 33.835 ;
        RECT  -4.0125 33.765 -3.8775 33.835 ;
        RECT  -4.0125 33.765 -3.8775 33.835 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.98 32.915 -3.91 33.05 ;
        RECT  -3.3075 33.765 -3.1725 33.835 ;
        RECT  -3.98 32.4225 -3.91 33.8325 ;
        RECT  -3.27 33.7725 -3.21 33.83 ;
        RECT  -3.4525 33.7725 -3.3975 33.825 ;
        RECT  -3.79 33.7725 -3.7325 33.8325 ;
        RECT  -3.975 33.7675 -3.915 33.825 ;
        RECT  -3.795 32.355 -3.725 33.9 ;
        RECT  -3.46 32.355 -3.39 33.9 ;
        RECT  -3.275 32.355 -3.205 33.9 ;
        RECT  -3.98 32.355 -3.91 33.9 ;
        RECT  -3.46 32.355 -3.39 33.9 ;
        RECT  -3.275 32.355 -3.205 33.9 ;
        RECT  -3.98 32.355 -3.91 33.9 ;
        RECT  -3.795 32.355 -3.725 33.9 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.3075 31.075 -3.1725 31.145 ;
        RECT  -4.0125 31.075 -3.8775 31.145 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.53 31.3675 -3.46 31.5025 ;
        RECT  -3.275 31.86 -3.205 31.995 ;
        RECT  -3.275 31.86 -3.205 31.995 ;
        RECT  -3.275 31.86 -3.205 31.995 ;
        RECT  -3.275 31.86 -3.205 31.995 ;
        RECT  -3.275 31.86 -3.205 31.995 ;
        RECT  -3.275 31.86 -3.205 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.725 31.3675 -3.655 31.5025 ;
        RECT  -4.0125 31.075 -3.8775 31.145 ;
        RECT  -4.0125 31.075 -3.8775 31.145 ;
        RECT  -4.0125 31.075 -3.8775 31.145 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.98 31.86 -3.91 31.995 ;
        RECT  -3.3075 31.075 -3.1725 31.145 ;
        RECT  -3.98 31.0775 -3.91 32.4875 ;
        RECT  -3.27 31.08 -3.21 31.1375 ;
        RECT  -3.4525 31.085 -3.3975 31.1375 ;
        RECT  -3.79 31.0775 -3.7325 31.1375 ;
        RECT  -3.975 31.085 -3.915 31.1425 ;
        RECT  -3.795 31.01 -3.725 32.555 ;
        RECT  -3.46 31.01 -3.39 32.555 ;
        RECT  -3.275 31.01 -3.205 32.555 ;
        RECT  -3.98 31.01 -3.91 32.555 ;
        RECT  -3.46 31.01 -3.39 32.555 ;
        RECT  -3.275 31.01 -3.205 32.555 ;
        RECT  -3.98 31.01 -3.91 32.555 ;
        RECT  -3.795 31.01 -3.725 32.555 ;
        RECT  -2.865 33.7725 -2.795 33.9075 ;
        RECT  -2.865 36.1825 -2.795 36.3175 ;
        RECT  -2.865 34.0 -2.795 34.135 ;
        RECT  -2.865 31.625 -2.795 31.76 ;
        RECT  -2.8975 36.69 -2.7625 36.76 ;
        RECT  -3.3075 36.69 -3.1725 36.76 ;
        RECT  -3.07 32.555 -2.935 32.625 ;
        RECT  -3.07 31.9575 -2.935 32.0275 ;
        RECT  -3.4925 31.9575 -3.3575 32.0275 ;
        RECT  -0.7275 26.0475 -0.6575 26.1825 ;
        RECT  -0.7275 21.9675 -0.6575 22.1025 ;
        RECT  -0.7275 27.4825 -0.6575 27.6175 ;
        RECT  -0.7275 21.9675 -0.6575 22.1025 ;
        RECT  -1.725 19.4 -1.655 19.535 ;
        RECT  -2.28 26.0475 -2.21 26.1825 ;
        RECT  -2.495 26.4575 -2.425 26.5925 ;
        RECT  -2.225 28.995 -2.155 29.13 ;
        RECT  -2.225 28.995 -2.155 29.13 ;
        RECT  -2.225 27.4825 -2.155 27.6175 ;
        RECT  -2.44 29.2525 -2.37 29.3875 ;
        RECT  -2.44 29.2525 -2.37 29.3875 ;
        RECT  -2.44 27.2775 -2.37 27.4125 ;
        RECT  -0.9525 27.4825 -0.8825 27.6175 ;
        RECT  -0.8125 27.2775 -0.7425 27.4125 ;
        RECT  -0.6725 26.6625 -0.6025 26.7975 ;
        RECT  -3.6425 27.4825 -3.5725 27.6175 ;
        RECT  -3.5025 26.6625 -3.4325 26.7975 ;
        RECT  -3.3625 26.8675 -3.2925 27.0025 ;
        RECT  -2.3125 28.81 -2.1775 28.88 ;
        RECT  -2.2575 29.955 -2.1225 30.025 ;
        RECT  -3.48 31.14 -3.345 31.21 ;
        RECT  -2.315 30.18 -2.18 30.25 ;
        RECT  -0.175 26.2525 -0.105 26.3875 ;
        RECT  -1.52 27.0725 -1.45 27.2075 ;
        RECT  -2.865 26.2525 -2.795 26.3875 ;
        RECT  -4.21 27.0725 -4.14 27.2075 ;
        RECT  9.8 30.18 9.935 30.25 ;
        RECT  -0.275 30.18 -0.14 30.25 ;
        RECT  9.595 31.14 9.73 31.21 ;
        RECT  -0.275 31.14 -0.14 31.21 ;
        RECT  9.185 28.81 9.32 28.88 ;
        RECT  -0.275 28.81 -0.14 28.88 ;
        RECT  8.98 29.955 9.115 30.025 ;
        RECT  -0.275 29.955 -0.14 30.025 ;
        RECT  9.39 27.515 9.525 27.585 ;
        RECT  -0.275 27.515 -0.14 27.585 ;
        RECT  8.775 26.08 8.91 26.15 ;
        RECT  -0.275 26.08 -0.14 26.15 ;
        RECT  0.1075 27.105 0.2425 27.175 ;
        RECT  8.36 26.285 8.495 26.355 ;
        RECT  -0.275 26.285 -0.14 26.355 ;
        LAYER  via2 ;
        RECT  10.6575 18.985 10.7275 19.055 ;
        RECT  11.3625 18.985 11.4325 19.055 ;
        RECT  10.6625 3.625 10.7325 3.695 ;
        RECT  11.3675 3.625 11.4375 3.695 ;
        RECT  10.6625 3.7775 10.7325 3.8475 ;
        RECT  11.3675 3.7775 11.4375 3.8475 ;
        RECT  0.515 7.5325 0.585 7.6025 ;
        RECT  0.515 6.8275 0.585 6.8975 ;
        RECT  0.515 6.1225 0.585 6.1925 ;
        RECT  0.515 5.4175 0.585 5.4875 ;
        RECT  10.455 0.475 10.52 0.54 ;
        RECT  11.16 0.475 11.225 0.54 ;
        RECT  10.665 0.035 10.73 0.1 ;
        RECT  11.37 0.035 11.435 0.1 ;
        RECT  7.025 8.2975 7.09 8.3625 ;
        RECT  8.22 8.2975 8.285 8.3625 ;
        RECT  7.025 10.9875 7.09 11.0525 ;
        RECT  8.22 10.9875 8.285 11.0525 ;
        RECT  7.025 13.6775 7.09 13.7425 ;
        RECT  8.22 13.6775 8.285 13.7425 ;
        RECT  7.025 16.3675 7.09 16.4325 ;
        RECT  8.22 16.3675 8.285 16.4325 ;
        RECT  -3.6925 19.265 -3.6225 19.335 ;
        RECT  -2.9875 19.265 -2.9175 19.335 ;
        RECT  -2.2825 19.265 -2.2125 19.335 ;
        RECT  -3.845 25.6375 -3.78 25.7025 ;
        RECT  -3.845 27.3125 -3.78 27.3775 ;
        RECT  -3.69 25.6375 -3.625 25.7025 ;
        RECT  -3.69 26.4925 -3.625 26.5575 ;
        RECT  -2.83 25.6375 -2.765 25.7025 ;
        RECT  -2.83 26.6975 -2.765 26.7625 ;
        RECT  -2.435 25.6375 -2.37 25.7025 ;
        RECT  -2.435 26.9025 -2.37 26.9675 ;
        RECT  -4.0425 25.6375 -3.9775 25.7025 ;
        RECT  -4.0425 26.2875 -3.9775 26.3525 ;
        RECT  -3.3375 25.6375 -3.2725 25.7025 ;
        RECT  -3.3375 26.2875 -3.2725 26.3525 ;
        RECT  -2.6325 25.6375 -2.5675 25.7025 ;
        RECT  -2.6325 26.2875 -2.5675 26.3525 ;
        RECT  -1.9275 25.6375 -1.8625 25.7025 ;
        RECT  -1.9275 26.2875 -1.8625 26.3525 ;
        RECT  -0.725 22.0025 -0.66 22.0675 ;
        RECT  -0.725 27.5175 -0.66 27.5825 ;
        RECT  -2.2225 29.03 -2.1575 29.095 ;
        RECT  -2.2225 27.5175 -2.1575 27.5825 ;
        RECT  -2.4375 29.2875 -2.3725 29.3525 ;
        RECT  -2.4375 27.3125 -2.3725 27.3775 ;
        RECT  9.835 30.1825 9.9 30.2475 ;
        RECT  -0.24 30.1825 -0.175 30.2475 ;
        RECT  9.63 31.1425 9.695 31.2075 ;
        RECT  -0.24 31.1425 -0.175 31.2075 ;
        RECT  9.22 28.8125 9.285 28.8775 ;
        RECT  -0.24 28.8125 -0.175 28.8775 ;
        RECT  9.015 29.9575 9.08 30.0225 ;
        RECT  -0.24 29.9575 -0.175 30.0225 ;
        RECT  9.425 27.5175 9.49 27.5825 ;
        RECT  -0.24 27.5175 -0.175 27.5825 ;
        RECT  8.81 26.0825 8.875 26.1475 ;
        RECT  -0.24 26.0825 -0.175 26.1475 ;
        RECT  8.395 26.2875 8.46 26.3525 ;
        RECT  -0.24 26.2875 -0.175 26.3525 ;
        LAYER  metal3 ;
        RECT  -0.14 30.18 9.8675 30.25 ;
        RECT  -0.14 31.14 9.6625 31.21 ;
        RECT  -0.14 28.81 9.2525 28.88 ;
        RECT  -0.14 29.955 9.0475 30.025 ;
        RECT  -0.14 27.515 9.4575 27.585 ;
        RECT  -0.14 26.08 8.8425 26.15 ;
        RECT  -0.14 26.285 8.4275 26.355 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  0.0 5.4175 0.48 5.4875 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  0.0 6.8275 0.48 6.8975 ;
        RECT  0.0 7.5325 0.48 7.6025 ;
        RECT  0.0 6.1225 0.48 6.1925 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  10.4525 18.985 10.5225 19.055 ;
        RECT  10.4525 0.475 10.5225 19.02 ;
        RECT  10.4875 18.985 10.6575 19.055 ;
        RECT  11.1575 18.985 11.2275 19.055 ;
        RECT  11.1575 0.475 11.2275 19.02 ;
        RECT  11.1925 18.985 11.3625 19.055 ;
        RECT  10.6625 0.0 10.7325 3.59 ;
        RECT  11.3675 0.0 11.4375 3.59 ;
        RECT  7.0575 8.295 8.2525 8.365 ;
        RECT  7.0575 10.985 8.2525 11.055 ;
        RECT  7.0575 13.675 8.2525 13.745 ;
        RECT  7.0575 16.365 8.2525 16.435 ;
        RECT  0.0 5.4175 0.48 5.4875 ;
        RECT  0.0 6.8275 0.48 6.8975 ;
        RECT  0.0 7.5325 0.48 7.6025 ;
        RECT  0.0 6.1225 0.48 6.1925 ;
        RECT  10.6575 18.95 10.7275 19.09 ;
        RECT  11.3625 18.95 11.4325 19.09 ;
        RECT  10.6575 18.95 10.7275 19.09 ;
        RECT  10.6575 18.95 10.7275 19.09 ;
        RECT  11.3625 18.95 11.4325 19.09 ;
        RECT  11.3625 18.95 11.4325 19.09 ;
        RECT  11.3675 3.59 11.4375 3.73 ;
        RECT  10.6625 3.59 10.7325 3.73 ;
        RECT  10.6625 3.59 10.7325 3.73 ;
        RECT  10.6625 3.59 10.7325 3.73 ;
        RECT  11.3675 3.59 11.4375 3.73 ;
        RECT  11.3675 3.59 11.4375 3.73 ;
        RECT  10.6625 3.7425 10.7325 3.8825 ;
        RECT  11.3675 3.7425 11.4375 3.8825 ;
        RECT  0.48 5.4175 0.62 5.4875 ;
        RECT  0.48 6.8275 0.62 6.8975 ;
        RECT  0.48 7.5325 0.62 7.6025 ;
        RECT  0.48 6.1225 0.62 6.1925 ;
        RECT  0.48 7.5325 0.62 7.6025 ;
        RECT  0.48 7.5325 0.62 7.6025 ;
        RECT  0.48 6.8275 0.62 6.8975 ;
        RECT  0.48 6.8275 0.62 6.8975 ;
        RECT  0.48 6.1225 0.62 6.1925 ;
        RECT  0.48 6.1225 0.62 6.1925 ;
        RECT  0.48 5.4175 0.62 5.4875 ;
        RECT  0.48 5.4175 0.62 5.4875 ;
        RECT  10.4525 0.44 10.5225 0.575 ;
        RECT  11.1575 0.44 11.2275 0.575 ;
        RECT  10.6625 0.0 10.7325 0.135 ;
        RECT  11.3675 0.0 11.4375 0.135 ;
        RECT  6.99 8.295 7.125 8.365 ;
        RECT  8.185 8.295 8.32 8.365 ;
        RECT  6.99 10.985 7.125 11.055 ;
        RECT  8.185 10.985 8.32 11.055 ;
        RECT  6.99 13.675 7.125 13.745 ;
        RECT  8.185 13.675 8.32 13.745 ;
        RECT  6.99 16.365 7.125 16.435 ;
        RECT  8.185 16.365 8.32 16.435 ;
        RECT  -3.8475 25.67 -3.7775 27.345 ;
        RECT  -3.6925 25.67 -3.6225 26.525 ;
        RECT  -2.8325 25.67 -2.7625 26.73 ;
        RECT  -2.4375 25.67 -2.3675 26.935 ;
        RECT  -4.045 25.67 -3.975 26.32 ;
        RECT  -3.34 25.67 -3.27 26.32 ;
        RECT  -2.635 25.67 -2.565 26.32 ;
        RECT  -1.93 25.67 -1.86 26.32 ;
        RECT  -0.7275 22.035 -0.6575 27.55 ;
        RECT  -2.225 27.55 -2.155 29.0625 ;
        RECT  -2.44 27.345 -2.37 29.32 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -3.8475 25.6025 -3.7775 25.7375 ;
        RECT  -3.8475 27.2775 -3.7775 27.4125 ;
        RECT  -3.6925 25.6025 -3.6225 25.7375 ;
        RECT  -3.6925 26.4575 -3.6225 26.5925 ;
        RECT  -2.8325 25.6025 -2.7625 25.7375 ;
        RECT  -2.8325 26.6625 -2.7625 26.7975 ;
        RECT  -2.4375 25.6025 -2.3675 25.7375 ;
        RECT  -2.4375 26.8675 -2.3675 27.0025 ;
        RECT  -4.045 25.6025 -3.975 25.7375 ;
        RECT  -4.045 26.2525 -3.975 26.3875 ;
        RECT  -3.34 25.6025 -3.27 25.7375 ;
        RECT  -3.34 26.2525 -3.27 26.3875 ;
        RECT  -2.635 25.6025 -2.565 25.7375 ;
        RECT  -2.635 26.2525 -2.565 26.3875 ;
        RECT  -1.93 25.6025 -1.86 25.7375 ;
        RECT  -1.93 26.2525 -1.86 26.3875 ;
        RECT  -0.7275 21.9675 -0.6575 22.1025 ;
        RECT  -0.7275 27.4825 -0.6575 27.6175 ;
        RECT  -2.225 28.995 -2.155 29.13 ;
        RECT  -2.225 27.4825 -2.155 27.6175 ;
        RECT  -2.44 29.2525 -2.37 29.3875 ;
        RECT  -2.44 27.2775 -2.37 27.4125 ;
        RECT  9.8 30.18 9.935 30.25 ;
        RECT  -0.275 30.18 -0.14 30.25 ;
        RECT  9.595 31.14 9.73 31.21 ;
        RECT  -0.275 31.14 -0.14 31.21 ;
        RECT  9.185 28.81 9.32 28.88 ;
        RECT  -0.275 28.81 -0.14 28.88 ;
        RECT  8.98 29.955 9.115 30.025 ;
        RECT  -0.275 29.955 -0.14 30.025 ;
        RECT  9.39 27.515 9.525 27.585 ;
        RECT  -0.275 27.515 -0.14 27.585 ;
        RECT  8.775 26.08 8.91 26.15 ;
        RECT  -0.275 26.08 -0.14 26.15 ;
        RECT  8.36 26.285 8.495 26.355 ;
        RECT  -0.275 26.285 -0.14 26.355 ;
    END
END    sram_2_16_1_freepdk45
END    LIBRARY
