magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1296 -1277 2768 2731
<< nwell >>
rect -36 679 1508 1471
<< locali >>
rect 0 1397 1472 1431
rect 64 636 98 702
rect 196 652 449 686
rect 547 664 707 698
rect 809 690 1073 724
rect 1281 690 1315 724
rect 809 681 843 690
rect 0 -17 1472 17
use pinv_5  pinv_5_0
timestamp 1595931502
transform 1 0 992 0 1 0
box -36 -17 516 1471
use pinv_3  pinv_3_0
timestamp 1595931502
transform 1 0 626 0 1 0
box -36 -17 402 1471
use pinv_7  pinv_7_0
timestamp 1595931502
transform 1 0 368 0 1 0
box -36 -17 294 1471
use pinv_4  pinv_4_0
timestamp 1595931502
transform 1 0 0 0 1 0
box -36 -17 404 1471
<< labels >>
rlabel corelocali s 736 0 736 0 4 gnd
rlabel corelocali s 1298 707 1298 707 4 Z
rlabel corelocali s 736 1414 736 1414 4 vdd
rlabel corelocali s 81 669 81 669 4 A
<< properties >>
string FIXED_BBOX 0 0 1472 1414
<< end >>
