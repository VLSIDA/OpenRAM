magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1296 -1277 1776 2731
<< nwell >>
rect -36 679 516 1471
<< poly >>
rect 114 740 144 907
rect 81 674 144 740
rect 114 507 144 674
<< locali >>
rect 0 1397 480 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 64 674 98 740
rect 272 724 306 1096
rect 272 690 323 724
rect 272 318 306 690
rect 62 17 96 218
rect 274 17 308 218
rect 0 -17 480 17
use pmos_m3_w2_000_sli_dli_da_p  pmos_m3_w2_000_sli_dli_da_p_0
timestamp 1595931502
transform 1 0 54 0 1 963
box -59 -56 425 454
use contact_12  contact_12_0
timestamp 1595931502
transform 1 0 48 0 1 674
box 0 0 66 66
use nmos_m3_w2_000_sli_dli_da_p  nmos_m3_w2_000_sli_dli_da_p_0
timestamp 1595931502
transform 1 0 54 0 1 51
box 0 -26 366 456
<< labels >>
rlabel corelocali s 240 0 240 0 4 gnd
rlabel corelocali s 306 707 306 707 4 Z
rlabel corelocali s 240 1414 240 1414 4 vdd
rlabel corelocali s 81 707 81 707 4 A
<< properties >>
string FIXED_BBOX 0 0 480 1414
<< end >>
