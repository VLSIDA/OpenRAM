*********************************************
* Transistor Models
* Note: These models are approximate 
*       and should be substituted with actual
*       models from MOSIS or SCN3ME
*********************************************

.MODEL p PMOS (LEVEL=4 VTO=-0.921340 KP=366.0244-6
+ NSUB=6E16 U0=212 VFB=0.395 GAMMA=0.2370 TOX=13.9n
+ TNOM=27)

