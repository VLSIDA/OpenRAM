*********************************************
* Transistor Models
* Note: These models are approximate 
*       and should be substituted with actual
*       models from MOSIS or SCN3ME
*********************************************

.MODEL n NMOS (LEVEL=49 VTHO=0.669845 KP=113.7771E-6
+ NSUB=6E16 U0=460 K1=0.5705 TOX=13.9n VERSION=3.3.0)

