magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1190 -1316 3224 1750
<< locali >>
rect 70 282 136 316
rect 549 314 970 348
rect 70 174 136 208
rect 936 197 970 314
rect 1079 130 1946 164
<< metal1 >>
rect 246 -30 294 402
rect 670 -32 720 402
rect 1098 0 1126 395
rect 1596 0 1624 395
use pinv_dec_0  pinv_dec_0_0
timestamp 1595931502
transform 1 0 876 0 1 0
box 44 0 1088 490
use nand2_dec  nand2_dec_0
timestamp 1595931502
transform 1 0 0 0 1 0
box 70 -56 888 476
<< labels >>
rlabel metal1 s 270 186 270 186 4 gnd
rlabel metal1 s 1112 197 1112 197 4 gnd
rlabel corelocali s 103 191 103 191 4 B
rlabel corelocali s 1512 147 1512 147 4 Z
rlabel metal1 s 1610 197 1610 197 4 vdd
rlabel metal1 s 695 185 695 185 4 vdd
rlabel corelocali s 103 299 103 299 4 A
<< properties >>
string FIXED_BBOX 0 0 1946 395
<< end >>
