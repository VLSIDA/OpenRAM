magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1296 -1277 1774 2731
<< nwell >>
rect -36 679 514 1471
<< poly >>
rect 114 303 144 1113
rect 96 237 144 303
rect 114 225 144 237
rect 214 225 244 1113
rect 314 551 344 1113
rect 314 485 362 551
rect 314 225 344 485
<< locali >>
rect 0 1397 478 1431
rect 62 1218 96 1397
rect 162 1184 196 1251
rect 262 1218 296 1397
rect 362 1184 396 1251
rect 162 1150 464 1184
rect 345 485 379 551
rect 212 361 246 427
rect 79 237 113 303
rect 430 158 464 1150
rect 379 92 464 158
rect 62 17 96 92
rect 0 -17 478 17
use nmos_m1_w0_740_sactive_dli  nmos_m1_w0_740_sactive_dli_0
timestamp 1595931502
transform 1 0 254 0 1 51
box 0 -26 150 174
use pmos_m1_w1_120_sli_dli  pmos_m1_w1_120_sli_dli_2
timestamp 1595931502
transform 1 0 54 0 1 1139
box -59 -54 209 278
use pmos_m1_w1_120_sli_dli  pmos_m1_w1_120_sli_dli_1
timestamp 1595931502
transform 1 0 154 0 1 1139
box -59 -54 209 278
use pmos_m1_w1_120_sli_dli  pmos_m1_w1_120_sli_dli_0
timestamp 1595931502
transform 1 0 254 0 1 1139
box -59 -54 209 278
use contact_12  contact_12_2
timestamp 1595931502
transform 1 0 63 0 1 237
box 0 0 66 66
use contact_12  contact_12_1
timestamp 1595931502
transform 1 0 196 0 1 361
box 0 0 66 66
use contact_12  contact_12_0
timestamp 1595931502
transform 1 0 329 0 1 485
box 0 0 66 66
use nmos_m1_w0_740_sli_dactive  nmos_m1_w0_740_sli_dactive_0
timestamp 1595931502
transform 1 0 54 0 1 51
box 0 -26 150 174
use nmos_m1_w0_740_sactive_dactive  nmos_m1_w0_740_sactive_dactive_0
timestamp 1595931502
transform 1 0 154 0 1 51
box 0 -26 150 174
<< labels >>
rlabel corelocali s 239 0 239 0 4 gnd
rlabel corelocali s 229 394 229 394 4 B
rlabel corelocali s 96 270 96 270 4 A
rlabel corelocali s 447 1167 447 1167 4 Z
rlabel corelocali s 362 518 362 518 4 C
rlabel corelocali s 239 1414 239 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 478 1414
<< end >>
