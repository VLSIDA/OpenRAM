magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1302 -1260 5046 9160
<< ndiffc >>
rect 1652 7488 1686 7490
rect 2058 7488 2092 7490
rect 1844 7331 1847 7363
rect 1897 7331 1900 7363
rect 1290 7204 1324 7206
rect 2420 7204 2454 7206
rect 1290 7172 1324 7174
rect 2420 7172 2454 7174
rect 1290 7046 1324 7048
rect 2420 7046 2454 7048
rect 1290 7014 1324 7016
rect 2420 7014 2454 7016
rect 1262 6857 1265 6889
rect 1711 6857 1714 6889
rect 1844 6857 1847 6889
rect 1897 6857 1900 6889
rect 2030 6857 2033 6889
rect 2479 6857 2482 6889
rect 1290 6698 1324 6732
rect 1652 6698 1686 6732
rect 2058 6698 2092 6732
rect 2420 6698 2454 6732
rect 1262 6541 1265 6573
rect 1711 6541 1714 6573
rect 1844 6541 1847 6573
rect 1897 6541 1900 6573
rect 2030 6541 2033 6573
rect 2479 6541 2482 6573
rect 1290 6414 1324 6416
rect 2420 6414 2454 6416
rect 1290 6382 1324 6384
rect 2420 6382 2454 6384
rect 1290 6256 1324 6258
rect 2420 6256 2454 6258
rect 1290 6224 1324 6226
rect 2420 6224 2454 6226
rect 1262 6067 1265 6099
rect 1711 6067 1714 6099
rect 1844 6067 1847 6099
rect 1897 6067 1900 6099
rect 2030 6067 2033 6099
rect 2479 6067 2482 6099
rect 1290 5908 1324 5942
rect 1652 5908 1686 5942
rect 2058 5908 2092 5942
rect 2420 5908 2454 5942
rect 1262 5751 1265 5783
rect 1711 5751 1714 5783
rect 1844 5751 1847 5783
rect 1897 5751 1900 5783
rect 2030 5751 2033 5783
rect 2479 5751 2482 5783
rect 1290 5624 1324 5626
rect 2420 5624 2454 5626
rect 1290 5592 1324 5594
rect 2420 5592 2454 5594
rect 1290 5466 1324 5468
rect 2420 5466 2454 5468
rect 1290 5434 1324 5436
rect 2420 5434 2454 5436
rect 1262 5277 1265 5309
rect 1711 5277 1714 5309
rect 1844 5277 1847 5309
rect 1897 5277 1900 5309
rect 2030 5277 2033 5309
rect 2479 5277 2482 5309
rect 1290 5118 1324 5152
rect 1652 5118 1686 5152
rect 2058 5118 2092 5152
rect 2420 5118 2454 5152
rect 1262 4961 1265 4993
rect 1711 4961 1714 4993
rect 1844 4961 1847 4993
rect 1897 4961 1900 4993
rect 2030 4961 2033 4993
rect 2479 4961 2482 4993
rect 1290 4834 1324 4836
rect 2420 4834 2454 4836
rect 1290 4802 1324 4804
rect 2420 4802 2454 4804
rect 1290 4676 1324 4678
rect 2420 4676 2454 4678
rect 1290 4644 1324 4646
rect 2420 4644 2454 4646
rect 1262 4487 1265 4519
rect 1711 4487 1714 4519
rect 1844 4487 1847 4519
rect 1897 4487 1900 4519
rect 2030 4487 2033 4519
rect 2479 4487 2482 4519
rect 1290 4328 1324 4362
rect 1652 4328 1686 4362
rect 2058 4328 2092 4362
rect 2420 4328 2454 4362
rect 1262 4171 1265 4203
rect 1711 4171 1714 4203
rect 1844 4171 1847 4203
rect 1897 4171 1900 4203
rect 2030 4171 2033 4203
rect 2479 4171 2482 4203
rect 1290 4044 1324 4046
rect 2420 4044 2454 4046
rect 1290 4012 1324 4014
rect 2420 4012 2454 4014
rect 1290 3886 1324 3888
rect 2420 3886 2454 3888
rect 1290 3854 1324 3856
rect 2420 3854 2454 3856
rect 1262 3697 1265 3729
rect 1711 3697 1714 3729
rect 1844 3697 1847 3729
rect 1897 3697 1900 3729
rect 2030 3697 2033 3729
rect 2479 3697 2482 3729
rect 1290 3538 1324 3572
rect 1652 3538 1686 3572
rect 2058 3538 2092 3572
rect 2420 3538 2454 3572
rect 1262 3381 1265 3413
rect 1711 3381 1714 3413
rect 1844 3381 1847 3413
rect 1897 3381 1900 3413
rect 2030 3381 2033 3413
rect 2479 3381 2482 3413
rect 1290 3254 1324 3256
rect 2420 3254 2454 3256
rect 1290 3222 1324 3224
rect 2420 3222 2454 3224
rect 1290 3096 1324 3098
rect 2420 3096 2454 3098
rect 1290 3064 1324 3066
rect 2420 3064 2454 3066
rect 1262 2907 1265 2939
rect 1711 2907 1714 2939
rect 1844 2907 1847 2939
rect 1897 2907 1900 2939
rect 2030 2907 2033 2939
rect 2479 2907 2482 2939
rect 1290 2748 1324 2782
rect 1652 2748 1686 2782
rect 2058 2748 2092 2782
rect 2420 2748 2454 2782
rect 1262 2591 1265 2623
rect 1711 2591 1714 2623
rect 1844 2591 1847 2623
rect 1897 2591 1900 2623
rect 2030 2591 2033 2623
rect 2479 2591 2482 2623
rect 1290 2464 1324 2466
rect 2420 2464 2454 2466
rect 1290 2432 1324 2434
rect 2420 2432 2454 2434
rect 1290 2306 1324 2308
rect 2420 2306 2454 2308
rect 1290 2274 1324 2276
rect 2420 2274 2454 2276
rect 1262 2117 1265 2149
rect 1711 2117 1714 2149
rect 1844 2117 1847 2149
rect 1897 2117 1900 2149
rect 2030 2117 2033 2149
rect 2479 2117 2482 2149
rect 1290 1958 1324 1992
rect 1652 1958 1686 1992
rect 2058 1958 2092 1992
rect 2420 1958 2454 1992
rect 1262 1801 1265 1833
rect 1711 1801 1714 1833
rect 1844 1801 1847 1833
rect 1897 1801 1900 1833
rect 2030 1801 2033 1833
rect 2479 1801 2482 1833
rect 1290 1674 1324 1676
rect 2420 1674 2454 1676
rect 1290 1642 1324 1644
rect 2420 1642 2454 1644
rect 1290 1516 1324 1518
rect 2420 1516 2454 1518
rect 1290 1484 1324 1486
rect 2420 1484 2454 1486
rect 1262 1327 1265 1359
rect 1711 1327 1714 1359
rect 1844 1327 1847 1359
rect 1897 1327 1900 1359
rect 2030 1327 2033 1359
rect 2479 1327 2482 1359
rect 1290 1168 1324 1202
rect 1652 1168 1686 1202
rect 2058 1168 2092 1202
rect 2420 1168 2454 1202
rect 1262 1011 1265 1043
rect 1711 1011 1714 1043
rect 1844 1011 1847 1043
rect 1897 1011 1900 1043
rect 2030 1011 2033 1043
rect 2479 1011 2482 1043
rect 1290 884 1324 886
rect 2420 884 2454 886
rect 1290 852 1324 854
rect 2420 852 2454 854
rect 1290 726 1324 728
rect 2420 726 2454 728
rect 1290 694 1324 696
rect 2420 694 2454 696
rect 1844 537 1847 569
rect 1897 537 1900 569
rect 1652 410 1686 412
rect 2058 410 2092 412
<< locali >>
rect 1290 7505 1324 7522
rect 1652 7505 1686 7520
rect 2058 7505 2092 7520
rect 2420 7505 2454 7522
rect 1234 7363 1265 7364
rect 1234 7331 1248 7363
rect 1234 7330 1265 7331
rect 1355 7323 1357 7351
rect 1387 7317 1389 7351
rect 1587 7343 1589 7377
rect 1619 7343 1621 7371
rect 1711 7363 1745 7364
rect 1813 7363 1844 7364
rect 1900 7363 1931 7364
rect 1999 7363 2033 7364
rect 2123 7343 2125 7371
rect 2155 7343 2157 7377
rect 2479 7363 2510 7364
rect 1711 7330 1745 7331
rect 1813 7330 1844 7331
rect 1900 7330 1931 7331
rect 1999 7330 2033 7331
rect 2355 7317 2357 7351
rect 2387 7323 2389 7351
rect 2496 7331 2510 7363
rect 2479 7330 2510 7331
rect 1441 6937 1444 6971
rect 1472 6937 1475 6971
rect 2269 6937 2272 6971
rect 2300 6937 2303 6971
rect 1234 6889 1262 6890
rect 1234 6857 1248 6889
rect 1355 6869 1357 6897
rect 1387 6869 1389 6903
rect 1234 6856 1262 6857
rect 1441 6856 1444 6890
rect 1472 6856 1475 6890
rect 1714 6889 1745 6890
rect 1813 6889 1844 6890
rect 1900 6889 1931 6890
rect 1999 6889 2030 6890
rect 1519 6852 1526 6886
rect 1587 6843 1589 6877
rect 1619 6849 1621 6877
rect 1714 6856 1745 6857
rect 1813 6856 1844 6857
rect 1900 6856 1931 6857
rect 1999 6856 2030 6857
rect 2123 6849 2125 6877
rect 2155 6843 2157 6877
rect 2218 6852 2225 6886
rect 2269 6856 2272 6890
rect 2300 6856 2303 6890
rect 2355 6869 2357 6903
rect 2387 6869 2389 6897
rect 2482 6889 2510 6890
rect 2496 6857 2510 6889
rect 2482 6856 2510 6857
rect 1441 6775 1444 6809
rect 1472 6775 1475 6809
rect 2269 6775 2272 6809
rect 2300 6775 2303 6809
rect 1441 6621 1444 6655
rect 1472 6621 1475 6655
rect 2269 6621 2272 6655
rect 2300 6621 2303 6655
rect 1234 6573 1262 6574
rect 1234 6541 1248 6573
rect 1234 6540 1262 6541
rect 1355 6533 1357 6561
rect 1387 6527 1389 6561
rect 1441 6540 1444 6574
rect 1472 6540 1475 6574
rect 1519 6544 1526 6578
rect 1587 6553 1589 6587
rect 1619 6553 1621 6581
rect 1714 6573 1745 6574
rect 1813 6573 1844 6574
rect 1900 6573 1931 6574
rect 1999 6573 2030 6574
rect 2123 6553 2125 6581
rect 2155 6553 2157 6587
rect 2218 6544 2225 6578
rect 1714 6540 1745 6541
rect 1813 6540 1844 6541
rect 1900 6540 1931 6541
rect 1999 6540 2030 6541
rect 2269 6540 2272 6574
rect 2300 6540 2303 6574
rect 2482 6573 2510 6574
rect 2355 6527 2357 6561
rect 2387 6533 2389 6561
rect 2496 6541 2510 6573
rect 2482 6540 2510 6541
rect 1441 6459 1444 6493
rect 1472 6459 1475 6493
rect 2269 6459 2272 6493
rect 2300 6459 2303 6493
rect 1441 6147 1444 6181
rect 1472 6147 1475 6181
rect 2269 6147 2272 6181
rect 2300 6147 2303 6181
rect 1234 6099 1262 6100
rect 1234 6067 1248 6099
rect 1355 6079 1357 6107
rect 1387 6079 1389 6113
rect 1234 6066 1262 6067
rect 1441 6066 1444 6100
rect 1472 6066 1475 6100
rect 1714 6099 1745 6100
rect 1813 6099 1844 6100
rect 1900 6099 1931 6100
rect 1999 6099 2030 6100
rect 1519 6062 1526 6096
rect 1587 6053 1589 6087
rect 1619 6059 1621 6087
rect 1714 6066 1745 6067
rect 1813 6066 1844 6067
rect 1900 6066 1931 6067
rect 1999 6066 2030 6067
rect 2123 6059 2125 6087
rect 2155 6053 2157 6087
rect 2218 6062 2225 6096
rect 2269 6066 2272 6100
rect 2300 6066 2303 6100
rect 2355 6079 2357 6113
rect 2387 6079 2389 6107
rect 2482 6099 2510 6100
rect 2496 6067 2510 6099
rect 2482 6066 2510 6067
rect 1441 5985 1444 6019
rect 1472 5985 1475 6019
rect 2269 5985 2272 6019
rect 2300 5985 2303 6019
rect 1441 5831 1444 5865
rect 1472 5831 1475 5865
rect 2269 5831 2272 5865
rect 2300 5831 2303 5865
rect 1234 5783 1262 5784
rect 1234 5751 1248 5783
rect 1234 5750 1262 5751
rect 1355 5743 1357 5771
rect 1387 5737 1389 5771
rect 1441 5750 1444 5784
rect 1472 5750 1475 5784
rect 1519 5754 1526 5788
rect 1587 5763 1589 5797
rect 1619 5763 1621 5791
rect 1714 5783 1745 5784
rect 1813 5783 1844 5784
rect 1900 5783 1931 5784
rect 1999 5783 2030 5784
rect 2123 5763 2125 5791
rect 2155 5763 2157 5797
rect 2218 5754 2225 5788
rect 1714 5750 1745 5751
rect 1813 5750 1844 5751
rect 1900 5750 1931 5751
rect 1999 5750 2030 5751
rect 2269 5750 2272 5784
rect 2300 5750 2303 5784
rect 2482 5783 2510 5784
rect 2355 5737 2357 5771
rect 2387 5743 2389 5771
rect 2496 5751 2510 5783
rect 2482 5750 2510 5751
rect 1441 5669 1444 5703
rect 1472 5669 1475 5703
rect 2269 5669 2272 5703
rect 2300 5669 2303 5703
rect 1441 5357 1444 5391
rect 1472 5357 1475 5391
rect 2269 5357 2272 5391
rect 2300 5357 2303 5391
rect 1234 5309 1262 5310
rect 1234 5277 1248 5309
rect 1355 5289 1357 5317
rect 1387 5289 1389 5323
rect 1234 5276 1262 5277
rect 1441 5276 1444 5310
rect 1472 5276 1475 5310
rect 1714 5309 1745 5310
rect 1813 5309 1844 5310
rect 1900 5309 1931 5310
rect 1999 5309 2030 5310
rect 1519 5272 1526 5306
rect 1587 5263 1589 5297
rect 1619 5269 1621 5297
rect 1714 5276 1745 5277
rect 1813 5276 1844 5277
rect 1900 5276 1931 5277
rect 1999 5276 2030 5277
rect 2123 5269 2125 5297
rect 2155 5263 2157 5297
rect 2218 5272 2225 5306
rect 2269 5276 2272 5310
rect 2300 5276 2303 5310
rect 2355 5289 2357 5323
rect 2387 5289 2389 5317
rect 2482 5309 2510 5310
rect 2496 5277 2510 5309
rect 2482 5276 2510 5277
rect 1441 5195 1444 5229
rect 1472 5195 1475 5229
rect 2269 5195 2272 5229
rect 2300 5195 2303 5229
rect 1441 5041 1444 5075
rect 1472 5041 1475 5075
rect 2269 5041 2272 5075
rect 2300 5041 2303 5075
rect 1234 4993 1262 4994
rect 1234 4961 1248 4993
rect 1234 4960 1262 4961
rect 1355 4953 1357 4981
rect 1387 4947 1389 4981
rect 1441 4960 1444 4994
rect 1472 4960 1475 4994
rect 1519 4964 1526 4998
rect 1587 4973 1589 5007
rect 1619 4973 1621 5001
rect 1714 4993 1745 4994
rect 1813 4993 1844 4994
rect 1900 4993 1931 4994
rect 1999 4993 2030 4994
rect 2123 4973 2125 5001
rect 2155 4973 2157 5007
rect 2218 4964 2225 4998
rect 1714 4960 1745 4961
rect 1813 4960 1844 4961
rect 1900 4960 1931 4961
rect 1999 4960 2030 4961
rect 2269 4960 2272 4994
rect 2300 4960 2303 4994
rect 2482 4993 2510 4994
rect 2355 4947 2357 4981
rect 2387 4953 2389 4981
rect 2496 4961 2510 4993
rect 2482 4960 2510 4961
rect 1441 4879 1444 4913
rect 1472 4879 1475 4913
rect 2269 4879 2272 4913
rect 2300 4879 2303 4913
rect 1441 4567 1444 4601
rect 1472 4567 1475 4601
rect 2269 4567 2272 4601
rect 2300 4567 2303 4601
rect 1234 4519 1262 4520
rect 1234 4487 1248 4519
rect 1355 4499 1357 4527
rect 1387 4499 1389 4533
rect 1234 4486 1262 4487
rect 1441 4486 1444 4520
rect 1472 4486 1475 4520
rect 1714 4519 1745 4520
rect 1813 4519 1844 4520
rect 1900 4519 1931 4520
rect 1999 4519 2030 4520
rect 1519 4482 1526 4516
rect 1587 4473 1589 4507
rect 1619 4479 1621 4507
rect 1714 4486 1745 4487
rect 1813 4486 1844 4487
rect 1900 4486 1931 4487
rect 1999 4486 2030 4487
rect 2123 4479 2125 4507
rect 2155 4473 2157 4507
rect 2218 4482 2225 4516
rect 2269 4486 2272 4520
rect 2300 4486 2303 4520
rect 2355 4499 2357 4533
rect 2387 4499 2389 4527
rect 2482 4519 2510 4520
rect 2496 4487 2510 4519
rect 2482 4486 2510 4487
rect 1441 4405 1444 4439
rect 1472 4405 1475 4439
rect 2269 4405 2272 4439
rect 2300 4405 2303 4439
rect 1441 4251 1444 4285
rect 1472 4251 1475 4285
rect 2269 4251 2272 4285
rect 2300 4251 2303 4285
rect 1234 4203 1262 4204
rect 1234 4171 1248 4203
rect 1234 4170 1262 4171
rect 1355 4163 1357 4191
rect 1387 4157 1389 4191
rect 1441 4170 1444 4204
rect 1472 4170 1475 4204
rect 1519 4174 1526 4208
rect 1587 4183 1589 4217
rect 1619 4183 1621 4211
rect 1714 4203 1745 4204
rect 1813 4203 1844 4204
rect 1900 4203 1931 4204
rect 1999 4203 2030 4204
rect 2123 4183 2125 4211
rect 2155 4183 2157 4217
rect 2218 4174 2225 4208
rect 1714 4170 1745 4171
rect 1813 4170 1844 4171
rect 1900 4170 1931 4171
rect 1999 4170 2030 4171
rect 2269 4170 2272 4204
rect 2300 4170 2303 4204
rect 2482 4203 2510 4204
rect 2355 4157 2357 4191
rect 2387 4163 2389 4191
rect 2496 4171 2510 4203
rect 2482 4170 2510 4171
rect 1441 4089 1444 4123
rect 1472 4089 1475 4123
rect 2269 4089 2272 4123
rect 2300 4089 2303 4123
rect 1441 3777 1444 3811
rect 1472 3777 1475 3811
rect 2269 3777 2272 3811
rect 2300 3777 2303 3811
rect 1234 3729 1262 3730
rect 1234 3697 1248 3729
rect 1355 3709 1357 3737
rect 1387 3709 1389 3743
rect 1234 3696 1262 3697
rect 1441 3696 1444 3730
rect 1472 3696 1475 3730
rect 1714 3729 1745 3730
rect 1813 3729 1844 3730
rect 1900 3729 1931 3730
rect 1999 3729 2030 3730
rect 1519 3692 1526 3726
rect 1587 3683 1589 3717
rect 1619 3689 1621 3717
rect 1714 3696 1745 3697
rect 1813 3696 1844 3697
rect 1900 3696 1931 3697
rect 1999 3696 2030 3697
rect 2123 3689 2125 3717
rect 2155 3683 2157 3717
rect 2218 3692 2225 3726
rect 2269 3696 2272 3730
rect 2300 3696 2303 3730
rect 2355 3709 2357 3743
rect 2387 3709 2389 3737
rect 2482 3729 2510 3730
rect 2496 3697 2510 3729
rect 2482 3696 2510 3697
rect 1441 3615 1444 3649
rect 1472 3615 1475 3649
rect 2269 3615 2272 3649
rect 2300 3615 2303 3649
rect 1441 3461 1444 3495
rect 1472 3461 1475 3495
rect 2269 3461 2272 3495
rect 2300 3461 2303 3495
rect 1234 3413 1262 3414
rect 1234 3381 1248 3413
rect 1234 3380 1262 3381
rect 1355 3373 1357 3401
rect 1387 3367 1389 3401
rect 1441 3380 1444 3414
rect 1472 3380 1475 3414
rect 1519 3384 1526 3418
rect 1587 3393 1589 3427
rect 1619 3393 1621 3421
rect 1714 3413 1745 3414
rect 1813 3413 1844 3414
rect 1900 3413 1931 3414
rect 1999 3413 2030 3414
rect 2123 3393 2125 3421
rect 2155 3393 2157 3427
rect 2218 3384 2225 3418
rect 1714 3380 1745 3381
rect 1813 3380 1844 3381
rect 1900 3380 1931 3381
rect 1999 3380 2030 3381
rect 2269 3380 2272 3414
rect 2300 3380 2303 3414
rect 2482 3413 2510 3414
rect 2355 3367 2357 3401
rect 2387 3373 2389 3401
rect 2496 3381 2510 3413
rect 2482 3380 2510 3381
rect 1441 3299 1444 3333
rect 1472 3299 1475 3333
rect 2269 3299 2272 3333
rect 2300 3299 2303 3333
rect 1441 2987 1444 3021
rect 1472 2987 1475 3021
rect 2269 2987 2272 3021
rect 2300 2987 2303 3021
rect 1234 2939 1262 2940
rect 1234 2907 1248 2939
rect 1355 2919 1357 2947
rect 1387 2919 1389 2953
rect 1234 2906 1262 2907
rect 1441 2906 1444 2940
rect 1472 2906 1475 2940
rect 1714 2939 1745 2940
rect 1813 2939 1844 2940
rect 1900 2939 1931 2940
rect 1999 2939 2030 2940
rect 1519 2902 1526 2936
rect 1587 2893 1589 2927
rect 1619 2899 1621 2927
rect 1714 2906 1745 2907
rect 1813 2906 1844 2907
rect 1900 2906 1931 2907
rect 1999 2906 2030 2907
rect 2123 2899 2125 2927
rect 2155 2893 2157 2927
rect 2218 2902 2225 2936
rect 2269 2906 2272 2940
rect 2300 2906 2303 2940
rect 2355 2919 2357 2953
rect 2387 2919 2389 2947
rect 2482 2939 2510 2940
rect 2496 2907 2510 2939
rect 2482 2906 2510 2907
rect 1441 2825 1444 2859
rect 1472 2825 1475 2859
rect 2269 2825 2272 2859
rect 2300 2825 2303 2859
rect 1441 2671 1444 2705
rect 1472 2671 1475 2705
rect 2269 2671 2272 2705
rect 2300 2671 2303 2705
rect 1234 2623 1262 2624
rect 1234 2591 1248 2623
rect 1234 2590 1262 2591
rect 1355 2583 1357 2611
rect 1387 2577 1389 2611
rect 1441 2590 1444 2624
rect 1472 2590 1475 2624
rect 1519 2594 1526 2628
rect 1587 2603 1589 2637
rect 1619 2603 1621 2631
rect 1714 2623 1745 2624
rect 1813 2623 1844 2624
rect 1900 2623 1931 2624
rect 1999 2623 2030 2624
rect 2123 2603 2125 2631
rect 2155 2603 2157 2637
rect 2218 2594 2225 2628
rect 1714 2590 1745 2591
rect 1813 2590 1844 2591
rect 1900 2590 1931 2591
rect 1999 2590 2030 2591
rect 2269 2590 2272 2624
rect 2300 2590 2303 2624
rect 2482 2623 2510 2624
rect 2355 2577 2357 2611
rect 2387 2583 2389 2611
rect 2496 2591 2510 2623
rect 2482 2590 2510 2591
rect 1441 2509 1444 2543
rect 1472 2509 1475 2543
rect 2269 2509 2272 2543
rect 2300 2509 2303 2543
rect 1441 2197 1444 2231
rect 1472 2197 1475 2231
rect 2269 2197 2272 2231
rect 2300 2197 2303 2231
rect 1234 2149 1262 2150
rect 1234 2117 1248 2149
rect 1355 2129 1357 2157
rect 1387 2129 1389 2163
rect 1234 2116 1262 2117
rect 1441 2116 1444 2150
rect 1472 2116 1475 2150
rect 1714 2149 1745 2150
rect 1813 2149 1844 2150
rect 1900 2149 1931 2150
rect 1999 2149 2030 2150
rect 1519 2112 1526 2146
rect 1587 2103 1589 2137
rect 1619 2109 1621 2137
rect 1714 2116 1745 2117
rect 1813 2116 1844 2117
rect 1900 2116 1931 2117
rect 1999 2116 2030 2117
rect 2123 2109 2125 2137
rect 2155 2103 2157 2137
rect 2218 2112 2225 2146
rect 2269 2116 2272 2150
rect 2300 2116 2303 2150
rect 2355 2129 2357 2163
rect 2387 2129 2389 2157
rect 2482 2149 2510 2150
rect 2496 2117 2510 2149
rect 2482 2116 2510 2117
rect 1441 2035 1444 2069
rect 1472 2035 1475 2069
rect 2269 2035 2272 2069
rect 2300 2035 2303 2069
rect 1441 1881 1444 1915
rect 1472 1881 1475 1915
rect 2269 1881 2272 1915
rect 2300 1881 2303 1915
rect 1234 1833 1262 1834
rect 1234 1801 1248 1833
rect 1234 1800 1262 1801
rect 1355 1793 1357 1821
rect 1387 1787 1389 1821
rect 1441 1800 1444 1834
rect 1472 1800 1475 1834
rect 1519 1804 1526 1838
rect 1587 1813 1589 1847
rect 1619 1813 1621 1841
rect 1714 1833 1745 1834
rect 1813 1833 1844 1834
rect 1900 1833 1931 1834
rect 1999 1833 2030 1834
rect 2123 1813 2125 1841
rect 2155 1813 2157 1847
rect 2218 1804 2225 1838
rect 1714 1800 1745 1801
rect 1813 1800 1844 1801
rect 1900 1800 1931 1801
rect 1999 1800 2030 1801
rect 2269 1800 2272 1834
rect 2300 1800 2303 1834
rect 2482 1833 2510 1834
rect 2355 1787 2357 1821
rect 2387 1793 2389 1821
rect 2496 1801 2510 1833
rect 2482 1800 2510 1801
rect 1441 1719 1444 1753
rect 1472 1719 1475 1753
rect 2269 1719 2272 1753
rect 2300 1719 2303 1753
rect 1441 1407 1444 1441
rect 1472 1407 1475 1441
rect 2269 1407 2272 1441
rect 2300 1407 2303 1441
rect 1234 1359 1262 1360
rect 1234 1327 1248 1359
rect 1355 1339 1357 1367
rect 1387 1339 1389 1373
rect 1234 1326 1262 1327
rect 1441 1326 1444 1360
rect 1472 1326 1475 1360
rect 1714 1359 1745 1360
rect 1813 1359 1844 1360
rect 1900 1359 1931 1360
rect 1999 1359 2030 1360
rect 1519 1322 1526 1356
rect 1587 1313 1589 1347
rect 1619 1319 1621 1347
rect 1714 1326 1745 1327
rect 1813 1326 1844 1327
rect 1900 1326 1931 1327
rect 1999 1326 2030 1327
rect 2123 1319 2125 1347
rect 2155 1313 2157 1347
rect 2218 1322 2225 1356
rect 2269 1326 2272 1360
rect 2300 1326 2303 1360
rect 2355 1339 2357 1373
rect 2387 1339 2389 1367
rect 2482 1359 2510 1360
rect 2496 1327 2510 1359
rect 2482 1326 2510 1327
rect 1441 1245 1444 1279
rect 1472 1245 1475 1279
rect 2269 1245 2272 1279
rect 2300 1245 2303 1279
rect 1441 1091 1444 1125
rect 1472 1091 1475 1125
rect 2269 1091 2272 1125
rect 2300 1091 2303 1125
rect 1234 1043 1262 1044
rect 1234 1011 1248 1043
rect 1234 1010 1262 1011
rect 1355 1003 1357 1031
rect 1387 997 1389 1031
rect 1441 1010 1444 1044
rect 1472 1010 1475 1044
rect 1519 1014 1526 1048
rect 1587 1023 1589 1057
rect 1619 1023 1621 1051
rect 1714 1043 1745 1044
rect 1813 1043 1844 1044
rect 1900 1043 1931 1044
rect 1999 1043 2030 1044
rect 2123 1023 2125 1051
rect 2155 1023 2157 1057
rect 2218 1014 2225 1048
rect 1714 1010 1745 1011
rect 1813 1010 1844 1011
rect 1900 1010 1931 1011
rect 1999 1010 2030 1011
rect 2269 1010 2272 1044
rect 2300 1010 2303 1044
rect 2482 1043 2510 1044
rect 2355 997 2357 1031
rect 2387 1003 2389 1031
rect 2496 1011 2510 1043
rect 2482 1010 2510 1011
rect 1441 929 1444 963
rect 1472 929 1475 963
rect 2269 929 2272 963
rect 2300 929 2303 963
rect 1234 569 1265 570
rect 1234 537 1248 569
rect 1355 549 1357 577
rect 1387 549 1389 583
rect 1711 569 1745 570
rect 1813 569 1844 570
rect 1900 569 1931 570
rect 1999 569 2033 570
rect 1234 536 1265 537
rect 1587 523 1589 557
rect 1619 529 1621 557
rect 1711 536 1745 537
rect 1813 536 1844 537
rect 1900 536 1931 537
rect 1999 536 2033 537
rect 2123 529 2125 557
rect 2155 523 2157 557
rect 2355 549 2357 583
rect 2387 549 2389 577
rect 2479 569 2510 570
rect 2496 537 2510 569
rect 2479 536 2510 537
rect 1290 378 1324 395
rect 1652 380 1686 395
rect 2058 380 2092 395
rect 2420 378 2454 395
<< metal1 >>
rect 846 0 882 7900
rect 918 0 954 7900
rect 990 7189 1026 7530
rect 990 6399 1026 7031
rect 990 5609 1026 6241
rect 990 4819 1026 5451
rect 990 4029 1026 4661
rect 990 3239 1026 3871
rect 990 2449 1026 3081
rect 990 1659 1026 2291
rect 990 869 1026 1501
rect 990 370 1026 711
rect 1062 0 1098 7900
rect 1134 0 1170 7900
rect 1326 0 1362 7900
rect 1398 0 1434 7900
rect 1542 0 1578 7900
rect 1614 0 1650 7900
rect 2094 0 2130 7900
rect 2166 0 2202 7900
rect 2310 0 2346 7900
rect 2382 0 2418 7900
rect 2574 0 2610 7900
rect 2646 0 2682 7900
rect 2718 7189 2754 7530
rect 2718 6399 2754 7031
rect 2718 5609 2754 6241
rect 2718 4819 2754 5451
rect 2718 4029 2754 4661
rect 2718 3239 2754 3871
rect 2718 2449 2754 3081
rect 2718 1659 2754 2291
rect 2718 869 2754 1501
rect 2718 370 2754 711
rect 2790 0 2826 7900
rect 2862 0 2898 7900
<< metal2 >>
rect 954 7309 1062 7385
rect 2682 7309 2790 7385
rect 0 7213 3744 7261
rect 954 7055 1062 7165
rect 2682 7055 2790 7165
rect 0 6959 3744 7007
rect 954 6835 1062 6911
rect 2682 6835 2790 6911
rect 0 6739 3744 6787
rect 0 6643 3744 6691
rect 954 6519 1062 6595
rect 2682 6519 2790 6595
rect 0 6423 3744 6471
rect 954 6265 1062 6375
rect 2682 6265 2790 6375
rect 0 6169 3744 6217
rect 954 6045 1062 6121
rect 2682 6045 2790 6121
rect 0 5949 3744 5997
rect 0 5853 3744 5901
rect 954 5729 1062 5805
rect 2682 5729 2790 5805
rect 0 5633 3744 5681
rect 954 5475 1062 5585
rect 2682 5475 2790 5585
rect 0 5379 3744 5427
rect 954 5255 1062 5331
rect 2682 5255 2790 5331
rect 0 5159 3744 5207
rect 0 5063 3744 5111
rect 954 4939 1062 5015
rect 2682 4939 2790 5015
rect 0 4843 3744 4891
rect 954 4685 1062 4795
rect 2682 4685 2790 4795
rect 0 4589 3744 4637
rect 954 4465 1062 4541
rect 2682 4465 2790 4541
rect 0 4369 3744 4417
rect 0 4273 3744 4321
rect 954 4149 1062 4225
rect 2682 4149 2790 4225
rect 0 4053 3744 4101
rect 954 3895 1062 4005
rect 2682 3895 2790 4005
rect 0 3799 3744 3847
rect 954 3675 1062 3751
rect 2682 3675 2790 3751
rect 0 3579 3744 3627
rect 0 3483 3744 3531
rect 954 3359 1062 3435
rect 2682 3359 2790 3435
rect 0 3263 3744 3311
rect 954 3105 1062 3215
rect 2682 3105 2790 3215
rect 0 3009 3744 3057
rect 954 2885 1062 2961
rect 2682 2885 2790 2961
rect 0 2789 3744 2837
rect 0 2693 3744 2741
rect 954 2569 1062 2645
rect 2682 2569 2790 2645
rect 0 2473 3744 2521
rect 954 2315 1062 2425
rect 2682 2315 2790 2425
rect 0 2219 3744 2267
rect 954 2095 1062 2171
rect 2682 2095 2790 2171
rect 0 1999 3744 2047
rect 0 1903 3744 1951
rect 954 1779 1062 1855
rect 2682 1779 2790 1855
rect 0 1683 3744 1731
rect 954 1525 1062 1635
rect 2682 1525 2790 1635
rect 0 1429 3744 1477
rect 954 1305 1062 1381
rect 2682 1305 2790 1381
rect 0 1209 3744 1257
rect 0 1113 3744 1161
rect 954 989 1062 1065
rect 2682 989 2790 1065
rect 0 893 3744 941
rect 954 735 1062 845
rect 2682 735 2790 845
rect 954 515 1062 591
rect 2682 515 2790 591
rect 0 419 3744 467
<< metal3 >>
rect 887 7622 985 7720
rect 1530 7641 1590 7701
rect 2154 7641 2214 7701
rect 2759 7622 2857 7720
rect 210 7317 270 7377
rect 3474 7317 3534 7377
rect 210 7080 270 7140
rect 3474 7080 3534 7140
rect 210 6843 270 6903
rect 3474 6843 3534 6903
rect 210 6527 270 6587
rect 3474 6527 3534 6587
rect 210 6290 270 6350
rect 3474 6290 3534 6350
rect 210 6053 270 6113
rect 3474 6053 3534 6113
rect 210 5737 270 5797
rect 3474 5737 3534 5797
rect 210 5500 270 5560
rect 3474 5500 3534 5560
rect 210 5263 270 5323
rect 3474 5263 3534 5323
rect 210 4947 270 5007
rect 3474 4947 3534 5007
rect 210 4710 270 4770
rect 3474 4710 3534 4770
rect 210 4473 270 4533
rect 3474 4473 3534 4533
rect 210 4157 270 4217
rect 3474 4157 3534 4217
rect 210 3920 270 3980
rect 3474 3920 3534 3980
rect 210 3683 270 3743
rect 3474 3683 3534 3743
rect 210 3367 270 3427
rect 3474 3367 3534 3427
rect 210 3130 270 3190
rect 3474 3130 3534 3190
rect 210 2893 270 2953
rect 3474 2893 3534 2953
rect 210 2577 270 2637
rect 3474 2577 3534 2637
rect 210 2340 270 2400
rect 3474 2340 3534 2400
rect 210 2103 270 2163
rect 3474 2103 3534 2163
rect 210 1787 270 1847
rect 3474 1787 3534 1847
rect 210 1550 270 1610
rect 3474 1550 3534 1610
rect 210 1313 270 1373
rect 3474 1313 3534 1373
rect 210 997 270 1057
rect 3474 997 3534 1057
rect 210 760 270 820
rect 3474 760 3534 820
rect 210 523 270 583
rect 3474 523 3534 583
rect 887 180 985 278
rect 1530 199 1590 259
rect 2154 199 2214 259
rect 2759 180 2857 278
use replica_column_0  replica_column_0_0
timestamp 1595931502
transform 1 0 2496 0 1 0
box -42 0 624 7900
use row_cap_array_0  row_cap_array_0_0
timestamp 1595931502
transform 1 0 3120 0 1 0
box 0 419 666 7481
use row_cap_array  row_cap_array_0
timestamp 1595931502
transform 1 0 0 0 1 0
box -42 419 624 7481
use col_cap_array  col_cap_array_0
timestamp 1595931502
transform 1 0 1248 0 -1 7900
box 0 0 1248 474
use col_cap_array  col_cap_array_1
timestamp 1595931502
transform 1 0 1248 0 1 0
box 0 0 1248 474
use dummy_array  dummy_array_0
timestamp 1595931502
transform 1 0 1248 0 1 7110
box -42 -104 1290 420
use dummy_array  dummy_array_1
timestamp 1595931502
transform 1 0 1248 0 -1 790
box -42 -104 1290 420
use replica_column  replica_column_0
timestamp 1595931502
transform 1 0 624 0 1 0
box 0 0 666 7900
use bitcell_array  bitcell_array_0
timestamp 1595931502
transform 1 0 1248 0 1 790
box -42 -104 1290 6424
<< labels >>
rlabel metal1 s 1416 3950 1416 3950 4 br0_0
rlabel metal2 s 1872 7237 1872 7237 4 rbl_wl1_1
rlabel metal2 s 1872 6983 1872 6983 4 wl1_15
rlabel metal2 s 1872 2717 1872 2717 4 wl0_4
rlabel metal2 s 1872 1707 1872 1707 4 wl1_2
rlabel metal1 s 2184 3950 2184 3950 4 bl1_1
rlabel metal2 s 1872 1453 1872 1453 4 wl1_1
rlabel metal1 s 2880 3950 2880 3950 4 rbl_br1_1
rlabel metal2 s 1872 1137 1872 1137 4 wl0_0
rlabel metal2 s 1872 5183 1872 5183 4 wl0_11
rlabel metal2 s 1872 2497 1872 2497 4 wl1_4
rlabel metal3 s 240 6320 240 6320 4 gnd
rlabel metal2 s 2736 6873 2736 6873 4 gnd
rlabel metal3 s 3504 1343 3504 1343 4 gnd
rlabel metal2 s 1008 7110 1008 7110 4 gnd
rlabel metal2 s 2736 4503 2736 4503 4 gnd
rlabel metal2 s 2736 4740 2736 4740 4 gnd
rlabel metal2 s 1008 5767 1008 5767 4 gnd
rlabel metal3 s 240 5767 240 5767 4 gnd
rlabel metal2 s 2736 2133 2736 2133 4 gnd
rlabel metal3 s 3504 2370 3504 2370 4 gnd
rlabel metal2 s 1008 1027 1008 1027 4 gnd
rlabel metal2 s 1008 5530 1008 5530 4 gnd
rlabel metal2 s 2736 3950 2736 3950 4 gnd
rlabel metal2 s 2736 1027 2736 1027 4 gnd
rlabel metal3 s 3504 2133 3504 2133 4 gnd
rlabel metal2 s 2736 4187 2736 4187 4 gnd
rlabel metal3 s 3504 1817 3504 1817 4 gnd
rlabel metal3 s 240 7110 240 7110 4 gnd
rlabel metal3 s 240 2607 240 2607 4 gnd
rlabel metal2 s 2736 1343 2736 1343 4 gnd
rlabel metal2 s 2736 3160 2736 3160 4 gnd
rlabel metal3 s 3504 5293 3504 5293 4 gnd
rlabel metal2 s 1008 5293 1008 5293 4 gnd
rlabel metal3 s 240 2370 240 2370 4 gnd
rlabel metal3 s 3504 4740 3504 4740 4 gnd
rlabel metal2 s 2736 553 2736 553 4 gnd
rlabel metal2 s 1008 2370 1008 2370 4 gnd
rlabel metal3 s 3504 7110 3504 7110 4 gnd
rlabel metal2 s 1008 4503 1008 4503 4 gnd
rlabel metal3 s 3504 6557 3504 6557 4 gnd
rlabel metal3 s 3504 3950 3504 3950 4 gnd
rlabel metal2 s 2736 6320 2736 6320 4 gnd
rlabel metal3 s 3504 2923 3504 2923 4 gnd
rlabel metal2 s 1008 3713 1008 3713 4 gnd
rlabel metal3 s 240 1580 240 1580 4 gnd
rlabel metal3 s 3504 4503 3504 4503 4 gnd
rlabel metal3 s 240 790 240 790 4 gnd
rlabel metal2 s 1008 7347 1008 7347 4 gnd
rlabel metal2 s 2736 2923 2736 2923 4 gnd
rlabel metal2 s 2736 7347 2736 7347 4 gnd
rlabel metal3 s 240 3397 240 3397 4 gnd
rlabel metal3 s 240 5293 240 5293 4 gnd
rlabel metal3 s 240 3713 240 3713 4 gnd
rlabel metal3 s 240 2133 240 2133 4 gnd
rlabel metal3 s 240 1343 240 1343 4 gnd
rlabel metal3 s 3504 3160 3504 3160 4 gnd
rlabel metal2 s 1008 1817 1008 1817 4 gnd
rlabel metal2 s 2736 4977 2736 4977 4 gnd
rlabel metal3 s 240 3950 240 3950 4 gnd
rlabel metal3 s 240 4977 240 4977 4 gnd
rlabel metal2 s 2736 6083 2736 6083 4 gnd
rlabel metal2 s 1008 4977 1008 4977 4 gnd
rlabel metal3 s 3504 790 3504 790 4 gnd
rlabel metal3 s 3504 1580 3504 1580 4 gnd
rlabel metal2 s 1008 553 1008 553 4 gnd
rlabel metal3 s 3504 6873 3504 6873 4 gnd
rlabel metal2 s 1008 2607 1008 2607 4 gnd
rlabel metal3 s 240 7347 240 7347 4 gnd
rlabel metal3 s 3504 2607 3504 2607 4 gnd
rlabel metal2 s 1008 6557 1008 6557 4 gnd
rlabel metal3 s 240 6083 240 6083 4 gnd
rlabel metal2 s 2736 7110 2736 7110 4 gnd
rlabel metal3 s 240 4187 240 4187 4 gnd
rlabel metal2 s 2736 5530 2736 5530 4 gnd
rlabel metal2 s 1008 4740 1008 4740 4 gnd
rlabel metal3 s 240 6873 240 6873 4 gnd
rlabel metal2 s 2736 5293 2736 5293 4 gnd
rlabel metal2 s 1008 1580 1008 1580 4 gnd
rlabel metal2 s 2736 3713 2736 3713 4 gnd
rlabel metal2 s 2736 5767 2736 5767 4 gnd
rlabel metal2 s 1008 6320 1008 6320 4 gnd
rlabel metal3 s 240 3160 240 3160 4 gnd
rlabel metal3 s 3504 6083 3504 6083 4 gnd
rlabel metal3 s 240 4740 240 4740 4 gnd
rlabel metal2 s 2736 1580 2736 1580 4 gnd
rlabel metal3 s 3504 6320 3504 6320 4 gnd
rlabel metal2 s 1008 2133 1008 2133 4 gnd
rlabel metal2 s 1008 4187 1008 4187 4 gnd
rlabel metal2 s 1008 790 1008 790 4 gnd
rlabel metal2 s 2736 6557 2736 6557 4 gnd
rlabel metal3 s 3504 4187 3504 4187 4 gnd
rlabel metal3 s 3504 7347 3504 7347 4 gnd
rlabel metal3 s 240 2923 240 2923 4 gnd
rlabel metal3 s 240 6557 240 6557 4 gnd
rlabel metal2 s 1008 6083 1008 6083 4 gnd
rlabel metal2 s 1008 6873 1008 6873 4 gnd
rlabel metal3 s 3504 3397 3504 3397 4 gnd
rlabel metal3 s 3504 553 3504 553 4 gnd
rlabel metal2 s 2736 790 2736 790 4 gnd
rlabel metal3 s 3504 3713 3504 3713 4 gnd
rlabel metal3 s 240 5530 240 5530 4 gnd
rlabel metal3 s 3504 5767 3504 5767 4 gnd
rlabel metal2 s 2736 2370 2736 2370 4 gnd
rlabel metal2 s 1008 3950 1008 3950 4 gnd
rlabel metal2 s 1008 3397 1008 3397 4 gnd
rlabel metal2 s 1008 1343 1008 1343 4 gnd
rlabel metal3 s 3504 4977 3504 4977 4 gnd
rlabel metal3 s 240 1817 240 1817 4 gnd
rlabel metal3 s 3504 5530 3504 5530 4 gnd
rlabel metal2 s 2736 3397 2736 3397 4 gnd
rlabel metal2 s 1008 2923 1008 2923 4 gnd
rlabel metal3 s 240 1027 240 1027 4 gnd
rlabel metal2 s 2736 2607 2736 2607 4 gnd
rlabel metal3 s 3504 1027 3504 1027 4 gnd
rlabel metal2 s 1008 3160 1008 3160 4 gnd
rlabel metal3 s 240 4503 240 4503 4 gnd
rlabel metal2 s 2736 1817 2736 1817 4 gnd
rlabel metal3 s 240 553 240 553 4 gnd
rlabel metal2 s 1872 917 1872 917 4 wl1_0
rlabel metal1 s 2736 2120 2736 2120 4 vdd
rlabel metal1 s 2736 1039 2736 1039 4 vdd
rlabel metal1 s 1008 2120 1008 2120 4 vdd
rlabel metal1 s 2736 6860 2736 6860 4 vdd
rlabel metal1 s 2736 1829 2736 1829 4 vdd
rlabel metal3 s 936 229 936 229 4 vdd
rlabel metal1 s 1008 3409 1008 3409 4 vdd
rlabel metal3 s 1560 7671 1560 7671 4 vdd
rlabel metal1 s 1008 5280 1008 5280 4 vdd
rlabel metal1 s 1008 4989 1008 4989 4 vdd
rlabel metal1 s 2736 6070 2736 6070 4 vdd
rlabel metal1 s 1008 1039 1008 1039 4 vdd
rlabel metal1 s 2736 4490 2736 4490 4 vdd
rlabel metal1 s 2736 540 2736 540 4 vdd
rlabel metal1 s 2736 1330 2736 1330 4 vdd
rlabel metal3 s 2808 229 2808 229 4 vdd
rlabel metal1 s 2736 2619 2736 2619 4 vdd
rlabel metal1 s 1008 5779 1008 5779 4 vdd
rlabel metal1 s 2736 7359 2736 7359 4 vdd
rlabel metal1 s 2736 4989 2736 4989 4 vdd
rlabel metal3 s 936 7671 936 7671 4 vdd
rlabel metal1 s 1008 3700 1008 3700 4 vdd
rlabel metal1 s 2736 3409 2736 3409 4 vdd
rlabel metal1 s 1008 6569 1008 6569 4 vdd
rlabel metal1 s 2736 2910 2736 2910 4 vdd
rlabel metal1 s 1008 1330 1008 1330 4 vdd
rlabel metal1 s 1008 6860 1008 6860 4 vdd
rlabel metal1 s 1008 2910 1008 2910 4 vdd
rlabel metal1 s 1008 2619 1008 2619 4 vdd
rlabel metal1 s 2736 5779 2736 5779 4 vdd
rlabel metal1 s 2736 5280 2736 5280 4 vdd
rlabel metal3 s 2184 229 2184 229 4 vdd
rlabel metal3 s 2184 7671 2184 7671 4 vdd
rlabel metal1 s 2736 4199 2736 4199 4 vdd
rlabel metal1 s 1008 7359 1008 7359 4 vdd
rlabel metal3 s 2808 7671 2808 7671 4 vdd
rlabel metal1 s 1008 1829 1008 1829 4 vdd
rlabel metal3 s 1560 229 1560 229 4 vdd
rlabel metal1 s 1008 6070 1008 6070 4 vdd
rlabel metal1 s 2736 6569 2736 6569 4 vdd
rlabel metal1 s 2736 3700 2736 3700 4 vdd
rlabel metal1 s 1008 540 1008 540 4 vdd
rlabel metal1 s 1008 4490 1008 4490 4 vdd
rlabel metal1 s 1008 4199 1008 4199 4 vdd
rlabel metal2 s 1872 443 1872 443 4 rbl_wl0_0
rlabel metal1 s 1152 3950 1152 3950 4 rbl_bl0_0
rlabel metal2 s 1872 6667 1872 6667 4 wl0_14
rlabel metal1 s 1344 3950 1344 3950 4 bl0_0
rlabel metal2 s 1872 2813 1872 2813 4 wl0_5
rlabel metal2 s 1872 5973 1872 5973 4 wl0_13
rlabel metal2 s 1872 2243 1872 2243 4 wl1_3
rlabel metal1 s 2592 3950 2592 3950 4 rbl_bl0_1
rlabel metal1 s 1560 3950 1560 3950 4 bl1_0
rlabel metal2 s 1872 5403 1872 5403 4 wl1_11
rlabel metal1 s 2328 3950 2328 3950 4 br0_1
rlabel metal1 s 1632 3950 1632 3950 4 br1_0
rlabel metal1 s 1080 3950 1080 3950 4 rbl_br0_0
rlabel metal1 s 2664 3950 2664 3950 4 rbl_br0_1
rlabel metal2 s 1872 6193 1872 6193 4 wl1_13
rlabel metal2 s 1872 4613 1872 4613 4 wl1_9
rlabel metal2 s 1872 1927 1872 1927 4 wl0_2
rlabel metal2 s 1872 3823 1872 3823 4 wl1_7
rlabel metal2 s 1872 6447 1872 6447 4 wl1_14
rlabel metal1 s 2808 3950 2808 3950 4 rbl_bl1_1
rlabel metal1 s 2112 3950 2112 3950 4 br1_1
rlabel metal2 s 1872 4867 1872 4867 4 wl1_10
rlabel metal2 s 1872 2023 1872 2023 4 wl0_3
rlabel metal2 s 1872 3287 1872 3287 4 wl1_6
rlabel metal2 s 1872 3507 1872 3507 4 wl0_6
rlabel metal2 s 1872 4393 1872 4393 4 wl0_9
rlabel metal2 s 1872 3603 1872 3603 4 wl0_7
rlabel metal1 s 936 3950 936 3950 4 rbl_bl1_0
rlabel metal2 s 1872 6763 1872 6763 4 wl0_15
rlabel metal2 s 1872 4077 1872 4077 4 wl1_8
rlabel metal2 s 1872 5877 1872 5877 4 wl0_12
rlabel metal2 s 1872 5657 1872 5657 4 wl1_12
rlabel metal2 s 1872 3033 1872 3033 4 wl1_5
rlabel metal1 s 864 3950 864 3950 4 rbl_br1_0
rlabel metal2 s 1872 1233 1872 1233 4 wl0_1
rlabel metal1 s 2400 3950 2400 3950 4 bl0_1
rlabel metal2 s 1872 5087 1872 5087 4 wl0_10
rlabel metal2 s 1872 4297 1872 4297 4 wl0_8
<< properties >>
string FIXED_BBOX 0 0 3744 7900
<< end >>
