magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1260 -1286 1626 1652
<< scnmos >>
rect 60 0 90 336
rect 168 0 198 336
rect 276 0 306 336
<< ndiff >>
rect 0 0 60 336
rect 90 0 168 336
rect 198 0 276 336
rect 306 0 366 336
<< poly >>
rect 60 362 306 392
rect 60 336 90 362
rect 168 336 198 362
rect 276 336 306 362
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
<< locali >>
rect 112 235 358 269
rect 8 135 42 201
rect 112 168 146 235
rect 220 135 254 201
rect 324 168 358 235
use contact_17  contact_17_3
timestamp 1595931502
transform 1 0 0 0 1 135
box 0 0 50 66
use contact_17  contact_17_2
timestamp 1595931502
transform 1 0 104 0 1 135
box 0 0 50 66
use contact_17  contact_17_1
timestamp 1595931502
transform 1 0 212 0 1 135
box 0 0 50 66
use contact_17  contact_17_0
timestamp 1595931502
transform 1 0 316 0 1 135
box 0 0 50 66
<< labels >>
rlabel poly s 183 377 183 377 4 G
rlabel corelocali s 237 168 237 168 4 S
rlabel corelocali s 25 168 25 168 4 S
rlabel corelocali s 235 252 235 252 4 D
<< properties >>
string FIXED_BBOX -25 -26 391 362
<< end >>
