MACRO sram_2_16_1_scn3me_subm
    CLASS RING ;
    ORIGIN 53.7 0.0 ;
    FOREIGN  sram 0.0 0.0 ;
    SIZE 203.4 BY 444.6 ;
    SYMMETRY X Y R90 ;
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  145.8 0.0 150.3 444.6 ;
        RECT  145.8 0.0 150.3 444.6 ;
        RECT  0.0 0.0 4.5 444.6 ;
        RECT  0.0 0.0 4.5 444.6 ;
        END
    END vdd
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal2 ;
        RECT  95.25 0.0 99.75 444.6 ;
        RECT  95.25 0.0 99.75 444.6 ;
        END
    END gnd
    PIN DATA[0]
        DIRECTION INOUT ;
        PORT
        LAYER metal2 ;
        RECT  127.2 0.0 128.1 1.8 ;
        RECT  127.2 0.0 128.1 1.8 ;
        END
    END DATA[0]
    PIN DATA[1]
        DIRECTION INOUT ;
        PORT
        LAYER metal2 ;
        RECT  137.4 0.0 138.3 1.8 ;
        RECT  137.4 0.0 138.3 1.8 ;
        END
    END DATA[1]
    PIN ADDR[0]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 75.0 7.2 76.5 ;
        RECT  0.0 75.0 7.2 76.5 ;
        END
    END ADDR[0]
    PIN ADDR[1]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 64.8 7.2 66.3 ;
        RECT  0.0 64.8 7.2 66.3 ;
        END
    END ADDR[1]
    PIN ADDR[2]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 54.6 7.2 56.1 ;
        RECT  0.0 54.6 7.2 56.1 ;
        END
    END ADDR[2]
    PIN ADDR[3]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 44.4 7.2 45.9 ;
        RECT  0.0 44.4 7.2 45.9 ;
        END
    END ADDR[3]
    PIN CSb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        END
    END CSb
    PIN OEb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        END
    END OEb
    PIN WEb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        END
    END WEb
    PIN clk
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -10.05 204.6 -8.85 205.8 ;
        RECT  -10.05 204.6 -8.85 205.8 ;
        RECT  -10.05 204.6 -8.85 205.8 ;
        RECT  -10.05 204.6 -8.85 205.8 ;
        END
    END clk
    OBS
        LAYER  metal1 ;
        RECT  1.8 295.65 2.7 298.35 ;
        RECT  -10.05 204.6 -8.85 205.8 ;
        RECT  145.8 0.0 150.3 444.6 ;
        RECT  0.0 0.0 4.5 444.6 ;
        RECT  44.7 205.2 45.6 206.1 ;
        RECT  44.7 202.95 45.6 203.85 ;
        RECT  43.35 205.2 45.15 206.1 ;
        RECT  44.7 203.4 45.6 205.65 ;
        RECT  45.15 202.95 47.1 203.85 ;
        RECT  102.15 205.2 103.05 206.1 ;
        RECT  102.15 201.45 103.05 202.35 ;
        RECT  83.25 205.2 102.6 206.1 ;
        RECT  102.15 201.9 103.05 205.65 ;
        RECT  102.6 201.45 122.1 202.35 ;
        RECT  44.7 220.5 45.6 221.4 ;
        RECT  44.7 222.75 45.6 223.65 ;
        RECT  43.35 220.5 45.15 221.4 ;
        RECT  44.7 220.95 45.6 223.2 ;
        RECT  45.15 222.75 47.1 223.65 ;
        RECT  102.15 220.5 103.05 221.4 ;
        RECT  102.15 224.25 103.05 225.15 ;
        RECT  83.25 220.5 102.6 221.4 ;
        RECT  102.15 220.95 103.05 224.7 ;
        RECT  102.6 224.25 122.1 225.15 ;
        RECT  44.7 233.4 45.6 234.3 ;
        RECT  44.7 231.15 45.6 232.05 ;
        RECT  43.35 233.4 45.15 234.3 ;
        RECT  44.7 231.6 45.6 233.85 ;
        RECT  45.15 231.15 47.1 232.05 ;
        RECT  102.15 233.4 103.05 234.3 ;
        RECT  102.15 229.65 103.05 230.55 ;
        RECT  83.25 233.4 102.6 234.3 ;
        RECT  102.15 230.1 103.05 233.85 ;
        RECT  102.6 229.65 122.1 230.55 ;
        RECT  44.7 248.7 45.6 249.6 ;
        RECT  44.7 250.95 45.6 251.85 ;
        RECT  43.35 248.7 45.15 249.6 ;
        RECT  44.7 249.15 45.6 251.4 ;
        RECT  45.15 250.95 47.1 251.85 ;
        RECT  102.15 248.7 103.05 249.6 ;
        RECT  102.15 252.45 103.05 253.35 ;
        RECT  83.25 248.7 102.6 249.6 ;
        RECT  102.15 249.15 103.05 252.9 ;
        RECT  102.6 252.45 122.1 253.35 ;
        RECT  44.7 261.6 45.6 262.5 ;
        RECT  44.7 259.35 45.6 260.25 ;
        RECT  43.35 261.6 45.15 262.5 ;
        RECT  44.7 259.8 45.6 262.05 ;
        RECT  45.15 259.35 47.1 260.25 ;
        RECT  102.15 261.6 103.05 262.5 ;
        RECT  102.15 257.85 103.05 258.75 ;
        RECT  83.25 261.6 102.6 262.5 ;
        RECT  102.15 258.3 103.05 262.05 ;
        RECT  102.6 257.85 122.1 258.75 ;
        RECT  44.7 276.9 45.6 277.8 ;
        RECT  44.7 279.15 45.6 280.05 ;
        RECT  43.35 276.9 45.15 277.8 ;
        RECT  44.7 277.35 45.6 279.6 ;
        RECT  45.15 279.15 47.1 280.05 ;
        RECT  102.15 276.9 103.05 277.8 ;
        RECT  102.15 280.65 103.05 281.55 ;
        RECT  83.25 276.9 102.6 277.8 ;
        RECT  102.15 277.35 103.05 281.1 ;
        RECT  102.6 280.65 122.1 281.55 ;
        RECT  44.7 289.8 45.6 290.7 ;
        RECT  44.7 287.55 45.6 288.45 ;
        RECT  43.35 289.8 45.15 290.7 ;
        RECT  44.7 288.0 45.6 290.25 ;
        RECT  45.15 287.55 47.1 288.45 ;
        RECT  102.15 289.8 103.05 290.7 ;
        RECT  102.15 286.05 103.05 286.95 ;
        RECT  83.25 289.8 102.6 290.7 ;
        RECT  102.15 286.5 103.05 290.25 ;
        RECT  102.6 286.05 122.1 286.95 ;
        RECT  44.7 305.1 45.6 306.0 ;
        RECT  44.7 307.35 45.6 308.25 ;
        RECT  43.35 305.1 45.15 306.0 ;
        RECT  44.7 305.55 45.6 307.8 ;
        RECT  45.15 307.35 47.1 308.25 ;
        RECT  102.15 305.1 103.05 306.0 ;
        RECT  102.15 308.85 103.05 309.75 ;
        RECT  83.25 305.1 102.6 306.0 ;
        RECT  102.15 305.55 103.05 309.3 ;
        RECT  102.6 308.85 122.1 309.75 ;
        RECT  44.7 318.0 45.6 318.9 ;
        RECT  44.7 315.75 45.6 316.65 ;
        RECT  43.35 318.0 45.15 318.9 ;
        RECT  44.7 316.2 45.6 318.45 ;
        RECT  45.15 315.75 47.1 316.65 ;
        RECT  102.15 318.0 103.05 318.9 ;
        RECT  102.15 314.25 103.05 315.15 ;
        RECT  83.25 318.0 102.6 318.9 ;
        RECT  102.15 314.7 103.05 318.45 ;
        RECT  102.6 314.25 122.1 315.15 ;
        RECT  44.7 333.3 45.6 334.2 ;
        RECT  44.7 335.55 45.6 336.45 ;
        RECT  43.35 333.3 45.15 334.2 ;
        RECT  44.7 333.75 45.6 336.0 ;
        RECT  45.15 335.55 47.1 336.45 ;
        RECT  102.15 333.3 103.05 334.2 ;
        RECT  102.15 337.05 103.05 337.95 ;
        RECT  83.25 333.3 102.6 334.2 ;
        RECT  102.15 333.75 103.05 337.5 ;
        RECT  102.6 337.05 122.1 337.95 ;
        RECT  44.7 346.2 45.6 347.1 ;
        RECT  44.7 343.95 45.6 344.85 ;
        RECT  43.35 346.2 45.15 347.1 ;
        RECT  44.7 344.4 45.6 346.65 ;
        RECT  45.15 343.95 47.1 344.85 ;
        RECT  102.15 346.2 103.05 347.1 ;
        RECT  102.15 342.45 103.05 343.35 ;
        RECT  83.25 346.2 102.6 347.1 ;
        RECT  102.15 342.9 103.05 346.65 ;
        RECT  102.6 342.45 122.1 343.35 ;
        RECT  44.7 361.5 45.6 362.4 ;
        RECT  44.7 363.75 45.6 364.65 ;
        RECT  43.35 361.5 45.15 362.4 ;
        RECT  44.7 361.95 45.6 364.2 ;
        RECT  45.15 363.75 47.1 364.65 ;
        RECT  102.15 361.5 103.05 362.4 ;
        RECT  102.15 365.25 103.05 366.15 ;
        RECT  83.25 361.5 102.6 362.4 ;
        RECT  102.15 361.95 103.05 365.7 ;
        RECT  102.6 365.25 122.1 366.15 ;
        RECT  44.7 374.4 45.6 375.3 ;
        RECT  44.7 372.15 45.6 373.05 ;
        RECT  43.35 374.4 45.15 375.3 ;
        RECT  44.7 372.6 45.6 374.85 ;
        RECT  45.15 372.15 47.1 373.05 ;
        RECT  102.15 374.4 103.05 375.3 ;
        RECT  102.15 370.65 103.05 371.55 ;
        RECT  83.25 374.4 102.6 375.3 ;
        RECT  102.15 371.1 103.05 374.85 ;
        RECT  102.6 370.65 122.1 371.55 ;
        RECT  44.7 389.7 45.6 390.6 ;
        RECT  44.7 391.95 45.6 392.85 ;
        RECT  43.35 389.7 45.15 390.6 ;
        RECT  44.7 390.15 45.6 392.4 ;
        RECT  45.15 391.95 47.1 392.85 ;
        RECT  102.15 389.7 103.05 390.6 ;
        RECT  102.15 393.45 103.05 394.35 ;
        RECT  83.25 389.7 102.6 390.6 ;
        RECT  102.15 390.15 103.05 393.9 ;
        RECT  102.6 393.45 122.1 394.35 ;
        RECT  44.7 402.6 45.6 403.5 ;
        RECT  44.7 400.35 45.6 401.25 ;
        RECT  43.35 402.6 45.15 403.5 ;
        RECT  44.7 400.8 45.6 403.05 ;
        RECT  45.15 400.35 47.1 401.25 ;
        RECT  102.15 402.6 103.05 403.5 ;
        RECT  102.15 398.85 103.05 399.75 ;
        RECT  83.25 402.6 102.6 403.5 ;
        RECT  102.15 399.3 103.05 403.05 ;
        RECT  102.6 398.85 122.1 399.75 ;
        RECT  44.7 417.9 45.6 418.8 ;
        RECT  44.7 420.15 45.6 421.05 ;
        RECT  43.35 417.9 45.15 418.8 ;
        RECT  44.7 418.35 45.6 420.6 ;
        RECT  45.15 420.15 47.1 421.05 ;
        RECT  102.15 417.9 103.05 418.8 ;
        RECT  102.15 421.65 103.05 422.55 ;
        RECT  83.25 417.9 102.6 418.8 ;
        RECT  102.15 418.35 103.05 422.1 ;
        RECT  102.6 421.65 122.1 422.55 ;
        RECT  53.4 198.75 122.7 199.65 ;
        RECT  53.4 226.95 122.7 227.85 ;
        RECT  53.4 255.15 122.7 256.05 ;
        RECT  53.4 283.35 122.7 284.25 ;
        RECT  53.4 311.55 122.7 312.45 ;
        RECT  53.4 339.75 122.7 340.65 ;
        RECT  53.4 367.95 122.7 368.85 ;
        RECT  53.4 396.15 122.7 397.05 ;
        RECT  53.4 424.35 122.7 425.25 ;
        RECT  0.0 212.85 150.3 213.75 ;
        RECT  0.0 241.05 150.3 241.95 ;
        RECT  0.0 269.25 150.3 270.15 ;
        RECT  0.0 297.45 150.3 298.35 ;
        RECT  0.0 325.65 150.3 326.55 ;
        RECT  0.0 353.85 150.3 354.75 ;
        RECT  0.0 382.05 150.3 382.95 ;
        RECT  0.0 410.25 150.3 411.15 ;
        RECT  77.7 88.65 82.2 89.55 ;
        RECT  74.7 102.75 84.9 103.65 ;
        RECT  77.7 145.05 87.6 145.95 ;
        RECT  74.7 159.15 90.3 160.05 ;
        RECT  77.7 85.95 79.2 86.85 ;
        RECT  77.7 114.15 79.2 115.05 ;
        RECT  77.7 142.35 79.2 143.25 ;
        RECT  77.7 170.55 79.2 171.45 ;
        RECT  0.0 100.05 77.7 100.95 ;
        RECT  0.0 128.25 77.7 129.15 ;
        RECT  0.0 156.45 77.7 157.35 ;
        RECT  0.0 184.65 77.7 185.55 ;
        RECT  66.3 75.45 82.2 76.35 ;
        RECT  66.3 65.25 84.9 66.15 ;
        RECT  66.3 55.05 87.6 55.95 ;
        RECT  66.3 44.85 90.3 45.75 ;
        RECT  66.3 70.35 96.45 71.25 ;
        RECT  66.3 49.95 96.45 50.85 ;
        RECT  62.7 37.65 63.6 38.55 ;
        RECT  62.7 38.1 63.6 40.2 ;
        RECT  0.0 37.65 63.15 38.55 ;
        RECT  111.0 32.4 122.7 33.3 ;
        RECT  105.6 27.9 122.7 28.8 ;
        RECT  108.3 25.5 122.7 26.4 ;
        RECT  111.0 429.6 122.7 430.5 ;
        RECT  113.7 96.9 122.7 97.8 ;
        RECT  116.4 195.0 122.7 195.9 ;
        RECT  8.7 82.65 9.6 83.55 ;
        RECT  8.7 81.0 9.6 83.1 ;
        RECT  9.15 82.65 102.9 83.55 ;
        RECT  50.25 426.45 103.8 427.35 ;
        RECT  122.7 443.7 145.8 444.6 ;
        RECT  122.7 167.7 145.8 168.6 ;
        RECT  122.7 99.0 145.8 99.9 ;
        RECT  122.7 86.4 145.8 87.3 ;
        RECT  122.7 9.6 145.8 10.5 ;
        RECT  99.75 23.4 122.7 24.3 ;
        RECT  99.75 192.9 122.7 193.8 ;
        RECT  99.75 94.8 122.7 95.7 ;
        RECT  145.8 0.0 150.3 444.6 ;
        RECT  0.0 0.0 4.5 444.6 ;
        RECT  122.1 257.7 143.7 258.9 ;
        RECT  122.1 201.3 143.7 202.5 ;
        RECT  122.1 229.5 143.7 230.7 ;
        RECT  122.1 421.5 143.7 422.7 ;
        RECT  122.1 314.1 143.7 315.3 ;
        RECT  122.1 285.9 143.7 287.1 ;
        RECT  122.1 393.3 143.7 394.5 ;
        RECT  122.1 365.1 143.7 366.3 ;
        RECT  122.1 252.3 143.7 253.5 ;
        RECT  122.1 280.5 143.7 281.7 ;
        RECT  122.1 224.1 143.7 225.3 ;
        RECT  122.1 398.7 143.7 399.9 ;
        RECT  122.1 342.3 143.7 343.5 ;
        RECT  122.1 336.9 143.7 338.1 ;
        RECT  122.1 212.7 143.7 213.6 ;
        RECT  122.1 240.9 143.7 241.8 ;
        RECT  122.1 269.1 143.7 270.0 ;
        RECT  122.1 297.3 143.7 298.2 ;
        RECT  122.1 325.5 143.7 326.4 ;
        RECT  122.1 353.7 143.7 354.6 ;
        RECT  122.1 381.9 143.7 382.8 ;
        RECT  122.1 410.1 143.7 411.0 ;
        RECT  122.1 370.5 143.7 371.7 ;
        RECT  122.1 308.7 143.7 309.9 ;
        RECT  128.4 199.2 131.1 200.4 ;
        RECT  124.2 199.2 126.9 200.4 ;
        RECT  122.1 201.3 133.5 202.5 ;
        RECT  127.8 202.5 129.0 202.8 ;
        RECT  132.3 204.0 133.5 209.7 ;
        RECT  129.9 204.0 131.1 205.2 ;
        RECT  125.7 204.0 126.9 205.2 ;
        RECT  129.6 205.2 130.8 205.8 ;
        RECT  129.0 205.8 130.8 207.0 ;
        RECT  129.6 207.0 130.8 210.6 ;
        RECT  126.0 205.2 127.2 208.5 ;
        RECT  126.0 208.5 128.4 209.7 ;
        RECT  123.3 204.0 124.5 209.7 ;
        RECT  126.0 209.7 127.2 210.6 ;
        RECT  132.3 210.6 133.5 212.7 ;
        RECT  129.3 210.6 130.5 211.8 ;
        RECT  126.3 210.6 127.5 211.8 ;
        RECT  123.3 210.6 124.5 212.7 ;
        RECT  122.1 212.7 133.5 213.9 ;
        RECT  122.1 201.3 133.5 202.5 ;
        RECT  122.1 212.7 133.5 213.9 ;
        RECT  128.4 226.2 131.1 227.4 ;
        RECT  124.2 226.2 126.9 227.4 ;
        RECT  122.1 224.1 133.5 225.3 ;
        RECT  127.8 223.8 129.0 224.1 ;
        RECT  132.3 216.9 133.5 222.6 ;
        RECT  129.9 221.4 131.1 222.6 ;
        RECT  125.7 221.4 126.9 222.6 ;
        RECT  129.6 220.8 130.8 221.4 ;
        RECT  129.0 219.6 130.8 220.8 ;
        RECT  129.6 216.0 130.8 219.6 ;
        RECT  126.0 218.1 127.2 221.4 ;
        RECT  126.0 216.9 128.4 218.1 ;
        RECT  123.3 216.9 124.5 222.6 ;
        RECT  126.0 216.0 127.2 216.9 ;
        RECT  132.3 213.9 133.5 216.0 ;
        RECT  129.3 214.8 130.5 216.0 ;
        RECT  126.3 214.8 127.5 216.0 ;
        RECT  123.3 213.9 124.5 216.0 ;
        RECT  122.1 212.7 133.5 213.9 ;
        RECT  122.1 224.1 133.5 225.3 ;
        RECT  122.1 212.7 133.5 213.9 ;
        RECT  128.4 227.4 131.1 228.6 ;
        RECT  124.2 227.4 126.9 228.6 ;
        RECT  122.1 229.5 133.5 230.7 ;
        RECT  127.8 230.7 129.0 231.0 ;
        RECT  132.3 232.2 133.5 237.9 ;
        RECT  129.9 232.2 131.1 233.4 ;
        RECT  125.7 232.2 126.9 233.4 ;
        RECT  129.6 233.4 130.8 234.0 ;
        RECT  129.0 234.0 130.8 235.2 ;
        RECT  129.6 235.2 130.8 238.8 ;
        RECT  126.0 233.4 127.2 236.7 ;
        RECT  126.0 236.7 128.4 237.9 ;
        RECT  123.3 232.2 124.5 237.9 ;
        RECT  126.0 237.9 127.2 238.8 ;
        RECT  132.3 238.8 133.5 240.9 ;
        RECT  129.3 238.8 130.5 240.0 ;
        RECT  126.3 238.8 127.5 240.0 ;
        RECT  123.3 238.8 124.5 240.9 ;
        RECT  122.1 240.9 133.5 242.1 ;
        RECT  122.1 229.5 133.5 230.7 ;
        RECT  122.1 240.9 133.5 242.1 ;
        RECT  128.4 254.4 131.1 255.6 ;
        RECT  124.2 254.4 126.9 255.6 ;
        RECT  122.1 252.3 133.5 253.5 ;
        RECT  127.8 252.0 129.0 252.3 ;
        RECT  132.3 245.1 133.5 250.8 ;
        RECT  129.9 249.6 131.1 250.8 ;
        RECT  125.7 249.6 126.9 250.8 ;
        RECT  129.6 249.0 130.8 249.6 ;
        RECT  129.0 247.8 130.8 249.0 ;
        RECT  129.6 244.2 130.8 247.8 ;
        RECT  126.0 246.3 127.2 249.6 ;
        RECT  126.0 245.1 128.4 246.3 ;
        RECT  123.3 245.1 124.5 250.8 ;
        RECT  126.0 244.2 127.2 245.1 ;
        RECT  132.3 242.1 133.5 244.2 ;
        RECT  129.3 243.0 130.5 244.2 ;
        RECT  126.3 243.0 127.5 244.2 ;
        RECT  123.3 242.1 124.5 244.2 ;
        RECT  122.1 240.9 133.5 242.1 ;
        RECT  122.1 252.3 133.5 253.5 ;
        RECT  122.1 240.9 133.5 242.1 ;
        RECT  128.4 255.6 131.1 256.8 ;
        RECT  124.2 255.6 126.9 256.8 ;
        RECT  122.1 257.7 133.5 258.9 ;
        RECT  127.8 258.9 129.0 259.2 ;
        RECT  132.3 260.4 133.5 266.1 ;
        RECT  129.9 260.4 131.1 261.6 ;
        RECT  125.7 260.4 126.9 261.6 ;
        RECT  129.6 261.6 130.8 262.2 ;
        RECT  129.0 262.2 130.8 263.4 ;
        RECT  129.6 263.4 130.8 267.0 ;
        RECT  126.0 261.6 127.2 264.9 ;
        RECT  126.0 264.9 128.4 266.1 ;
        RECT  123.3 260.4 124.5 266.1 ;
        RECT  126.0 266.1 127.2 267.0 ;
        RECT  132.3 267.0 133.5 269.1 ;
        RECT  129.3 267.0 130.5 268.2 ;
        RECT  126.3 267.0 127.5 268.2 ;
        RECT  123.3 267.0 124.5 269.1 ;
        RECT  122.1 269.1 133.5 270.3 ;
        RECT  122.1 257.7 133.5 258.9 ;
        RECT  122.1 269.1 133.5 270.3 ;
        RECT  128.4 282.6 131.1 283.8 ;
        RECT  124.2 282.6 126.9 283.8 ;
        RECT  122.1 280.5 133.5 281.7 ;
        RECT  127.8 280.2 129.0 280.5 ;
        RECT  132.3 273.3 133.5 279.0 ;
        RECT  129.9 277.8 131.1 279.0 ;
        RECT  125.7 277.8 126.9 279.0 ;
        RECT  129.6 277.2 130.8 277.8 ;
        RECT  129.0 276.0 130.8 277.2 ;
        RECT  129.6 272.4 130.8 276.0 ;
        RECT  126.0 274.5 127.2 277.8 ;
        RECT  126.0 273.3 128.4 274.5 ;
        RECT  123.3 273.3 124.5 279.0 ;
        RECT  126.0 272.4 127.2 273.3 ;
        RECT  132.3 270.3 133.5 272.4 ;
        RECT  129.3 271.2 130.5 272.4 ;
        RECT  126.3 271.2 127.5 272.4 ;
        RECT  123.3 270.3 124.5 272.4 ;
        RECT  122.1 269.1 133.5 270.3 ;
        RECT  122.1 280.5 133.5 281.7 ;
        RECT  122.1 269.1 133.5 270.3 ;
        RECT  128.4 283.8 131.1 285.0 ;
        RECT  124.2 283.8 126.9 285.0 ;
        RECT  122.1 285.9 133.5 287.1 ;
        RECT  127.8 287.1 129.0 287.4 ;
        RECT  132.3 288.6 133.5 294.3 ;
        RECT  129.9 288.6 131.1 289.8 ;
        RECT  125.7 288.6 126.9 289.8 ;
        RECT  129.6 289.8 130.8 290.4 ;
        RECT  129.0 290.4 130.8 291.6 ;
        RECT  129.6 291.6 130.8 295.2 ;
        RECT  126.0 289.8 127.2 293.1 ;
        RECT  126.0 293.1 128.4 294.3 ;
        RECT  123.3 288.6 124.5 294.3 ;
        RECT  126.0 294.3 127.2 295.2 ;
        RECT  132.3 295.2 133.5 297.3 ;
        RECT  129.3 295.2 130.5 296.4 ;
        RECT  126.3 295.2 127.5 296.4 ;
        RECT  123.3 295.2 124.5 297.3 ;
        RECT  122.1 297.3 133.5 298.5 ;
        RECT  122.1 285.9 133.5 287.1 ;
        RECT  122.1 297.3 133.5 298.5 ;
        RECT  128.4 310.8 131.1 312.0 ;
        RECT  124.2 310.8 126.9 312.0 ;
        RECT  122.1 308.7 133.5 309.9 ;
        RECT  127.8 308.4 129.0 308.7 ;
        RECT  132.3 301.5 133.5 307.2 ;
        RECT  129.9 306.0 131.1 307.2 ;
        RECT  125.7 306.0 126.9 307.2 ;
        RECT  129.6 305.4 130.8 306.0 ;
        RECT  129.0 304.2 130.8 305.4 ;
        RECT  129.6 300.6 130.8 304.2 ;
        RECT  126.0 302.7 127.2 306.0 ;
        RECT  126.0 301.5 128.4 302.7 ;
        RECT  123.3 301.5 124.5 307.2 ;
        RECT  126.0 300.6 127.2 301.5 ;
        RECT  132.3 298.5 133.5 300.6 ;
        RECT  129.3 299.4 130.5 300.6 ;
        RECT  126.3 299.4 127.5 300.6 ;
        RECT  123.3 298.5 124.5 300.6 ;
        RECT  122.1 297.3 133.5 298.5 ;
        RECT  122.1 308.7 133.5 309.9 ;
        RECT  122.1 297.3 133.5 298.5 ;
        RECT  128.4 312.0 131.1 313.2 ;
        RECT  124.2 312.0 126.9 313.2 ;
        RECT  122.1 314.1 133.5 315.3 ;
        RECT  127.8 315.3 129.0 315.6 ;
        RECT  132.3 316.8 133.5 322.5 ;
        RECT  129.9 316.8 131.1 318.0 ;
        RECT  125.7 316.8 126.9 318.0 ;
        RECT  129.6 318.0 130.8 318.6 ;
        RECT  129.0 318.6 130.8 319.8 ;
        RECT  129.6 319.8 130.8 323.4 ;
        RECT  126.0 318.0 127.2 321.3 ;
        RECT  126.0 321.3 128.4 322.5 ;
        RECT  123.3 316.8 124.5 322.5 ;
        RECT  126.0 322.5 127.2 323.4 ;
        RECT  132.3 323.4 133.5 325.5 ;
        RECT  129.3 323.4 130.5 324.6 ;
        RECT  126.3 323.4 127.5 324.6 ;
        RECT  123.3 323.4 124.5 325.5 ;
        RECT  122.1 325.5 133.5 326.7 ;
        RECT  122.1 314.1 133.5 315.3 ;
        RECT  122.1 325.5 133.5 326.7 ;
        RECT  128.4 339.0 131.1 340.2 ;
        RECT  124.2 339.0 126.9 340.2 ;
        RECT  122.1 336.9 133.5 338.1 ;
        RECT  127.8 336.6 129.0 336.9 ;
        RECT  132.3 329.7 133.5 335.4 ;
        RECT  129.9 334.2 131.1 335.4 ;
        RECT  125.7 334.2 126.9 335.4 ;
        RECT  129.6 333.6 130.8 334.2 ;
        RECT  129.0 332.4 130.8 333.6 ;
        RECT  129.6 328.8 130.8 332.4 ;
        RECT  126.0 330.9 127.2 334.2 ;
        RECT  126.0 329.7 128.4 330.9 ;
        RECT  123.3 329.7 124.5 335.4 ;
        RECT  126.0 328.8 127.2 329.7 ;
        RECT  132.3 326.7 133.5 328.8 ;
        RECT  129.3 327.6 130.5 328.8 ;
        RECT  126.3 327.6 127.5 328.8 ;
        RECT  123.3 326.7 124.5 328.8 ;
        RECT  122.1 325.5 133.5 326.7 ;
        RECT  122.1 336.9 133.5 338.1 ;
        RECT  122.1 325.5 133.5 326.7 ;
        RECT  128.4 340.2 131.1 341.4 ;
        RECT  124.2 340.2 126.9 341.4 ;
        RECT  122.1 342.3 133.5 343.5 ;
        RECT  127.8 343.5 129.0 343.8 ;
        RECT  132.3 345.0 133.5 350.7 ;
        RECT  129.9 345.0 131.1 346.2 ;
        RECT  125.7 345.0 126.9 346.2 ;
        RECT  129.6 346.2 130.8 346.8 ;
        RECT  129.0 346.8 130.8 348.0 ;
        RECT  129.6 348.0 130.8 351.6 ;
        RECT  126.0 346.2 127.2 349.5 ;
        RECT  126.0 349.5 128.4 350.7 ;
        RECT  123.3 345.0 124.5 350.7 ;
        RECT  126.0 350.7 127.2 351.6 ;
        RECT  132.3 351.6 133.5 353.7 ;
        RECT  129.3 351.6 130.5 352.8 ;
        RECT  126.3 351.6 127.5 352.8 ;
        RECT  123.3 351.6 124.5 353.7 ;
        RECT  122.1 353.7 133.5 354.9 ;
        RECT  122.1 342.3 133.5 343.5 ;
        RECT  122.1 353.7 133.5 354.9 ;
        RECT  128.4 367.2 131.1 368.4 ;
        RECT  124.2 367.2 126.9 368.4 ;
        RECT  122.1 365.1 133.5 366.3 ;
        RECT  127.8 364.8 129.0 365.1 ;
        RECT  132.3 357.9 133.5 363.6 ;
        RECT  129.9 362.4 131.1 363.6 ;
        RECT  125.7 362.4 126.9 363.6 ;
        RECT  129.6 361.8 130.8 362.4 ;
        RECT  129.0 360.6 130.8 361.8 ;
        RECT  129.6 357.0 130.8 360.6 ;
        RECT  126.0 359.1 127.2 362.4 ;
        RECT  126.0 357.9 128.4 359.1 ;
        RECT  123.3 357.9 124.5 363.6 ;
        RECT  126.0 357.0 127.2 357.9 ;
        RECT  132.3 354.9 133.5 357.0 ;
        RECT  129.3 355.8 130.5 357.0 ;
        RECT  126.3 355.8 127.5 357.0 ;
        RECT  123.3 354.9 124.5 357.0 ;
        RECT  122.1 353.7 133.5 354.9 ;
        RECT  122.1 365.1 133.5 366.3 ;
        RECT  122.1 353.7 133.5 354.9 ;
        RECT  128.4 368.4 131.1 369.6 ;
        RECT  124.2 368.4 126.9 369.6 ;
        RECT  122.1 370.5 133.5 371.7 ;
        RECT  127.8 371.7 129.0 372.0 ;
        RECT  132.3 373.2 133.5 378.9 ;
        RECT  129.9 373.2 131.1 374.4 ;
        RECT  125.7 373.2 126.9 374.4 ;
        RECT  129.6 374.4 130.8 375.0 ;
        RECT  129.0 375.0 130.8 376.2 ;
        RECT  129.6 376.2 130.8 379.8 ;
        RECT  126.0 374.4 127.2 377.7 ;
        RECT  126.0 377.7 128.4 378.9 ;
        RECT  123.3 373.2 124.5 378.9 ;
        RECT  126.0 378.9 127.2 379.8 ;
        RECT  132.3 379.8 133.5 381.9 ;
        RECT  129.3 379.8 130.5 381.0 ;
        RECT  126.3 379.8 127.5 381.0 ;
        RECT  123.3 379.8 124.5 381.9 ;
        RECT  122.1 381.9 133.5 383.1 ;
        RECT  122.1 370.5 133.5 371.7 ;
        RECT  122.1 381.9 133.5 383.1 ;
        RECT  128.4 395.4 131.1 396.6 ;
        RECT  124.2 395.4 126.9 396.6 ;
        RECT  122.1 393.3 133.5 394.5 ;
        RECT  127.8 393.0 129.0 393.3 ;
        RECT  132.3 386.1 133.5 391.8 ;
        RECT  129.9 390.6 131.1 391.8 ;
        RECT  125.7 390.6 126.9 391.8 ;
        RECT  129.6 390.0 130.8 390.6 ;
        RECT  129.0 388.8 130.8 390.0 ;
        RECT  129.6 385.2 130.8 388.8 ;
        RECT  126.0 387.3 127.2 390.6 ;
        RECT  126.0 386.1 128.4 387.3 ;
        RECT  123.3 386.1 124.5 391.8 ;
        RECT  126.0 385.2 127.2 386.1 ;
        RECT  132.3 383.1 133.5 385.2 ;
        RECT  129.3 384.0 130.5 385.2 ;
        RECT  126.3 384.0 127.5 385.2 ;
        RECT  123.3 383.1 124.5 385.2 ;
        RECT  122.1 381.9 133.5 383.1 ;
        RECT  122.1 393.3 133.5 394.5 ;
        RECT  122.1 381.9 133.5 383.1 ;
        RECT  128.4 396.6 131.1 397.8 ;
        RECT  124.2 396.6 126.9 397.8 ;
        RECT  122.1 398.7 133.5 399.9 ;
        RECT  127.8 399.9 129.0 400.2 ;
        RECT  132.3 401.4 133.5 407.1 ;
        RECT  129.9 401.4 131.1 402.6 ;
        RECT  125.7 401.4 126.9 402.6 ;
        RECT  129.6 402.6 130.8 403.2 ;
        RECT  129.0 403.2 130.8 404.4 ;
        RECT  129.6 404.4 130.8 408.0 ;
        RECT  126.0 402.6 127.2 405.9 ;
        RECT  126.0 405.9 128.4 407.1 ;
        RECT  123.3 401.4 124.5 407.1 ;
        RECT  126.0 407.1 127.2 408.0 ;
        RECT  132.3 408.0 133.5 410.1 ;
        RECT  129.3 408.0 130.5 409.2 ;
        RECT  126.3 408.0 127.5 409.2 ;
        RECT  123.3 408.0 124.5 410.1 ;
        RECT  122.1 410.1 133.5 411.3 ;
        RECT  122.1 398.7 133.5 399.9 ;
        RECT  122.1 410.1 133.5 411.3 ;
        RECT  128.4 423.6 131.1 424.8 ;
        RECT  124.2 423.6 126.9 424.8 ;
        RECT  122.1 421.5 133.5 422.7 ;
        RECT  127.8 421.2 129.0 421.5 ;
        RECT  132.3 414.3 133.5 420.0 ;
        RECT  129.9 418.8 131.1 420.0 ;
        RECT  125.7 418.8 126.9 420.0 ;
        RECT  129.6 418.2 130.8 418.8 ;
        RECT  129.0 417.0 130.8 418.2 ;
        RECT  129.6 413.4 130.8 417.0 ;
        RECT  126.0 415.5 127.2 418.8 ;
        RECT  126.0 414.3 128.4 415.5 ;
        RECT  123.3 414.3 124.5 420.0 ;
        RECT  126.0 413.4 127.2 414.3 ;
        RECT  132.3 411.3 133.5 413.4 ;
        RECT  129.3 412.2 130.5 413.4 ;
        RECT  126.3 412.2 127.5 413.4 ;
        RECT  123.3 411.3 124.5 413.4 ;
        RECT  122.1 410.1 133.5 411.3 ;
        RECT  122.1 421.5 133.5 422.7 ;
        RECT  122.1 410.1 133.5 411.3 ;
        RECT  138.6 199.2 141.3 200.4 ;
        RECT  134.4 199.2 137.1 200.4 ;
        RECT  132.3 201.3 143.7 202.5 ;
        RECT  138.0 202.5 139.2 202.8 ;
        RECT  142.5 204.0 143.7 209.7 ;
        RECT  140.1 204.0 141.3 205.2 ;
        RECT  135.9 204.0 137.1 205.2 ;
        RECT  139.8 205.2 141.0 205.8 ;
        RECT  139.2 205.8 141.0 207.0 ;
        RECT  139.8 207.0 141.0 210.6 ;
        RECT  136.2 205.2 137.4 208.5 ;
        RECT  136.2 208.5 138.6 209.7 ;
        RECT  133.5 204.0 134.7 209.7 ;
        RECT  136.2 209.7 137.4 210.6 ;
        RECT  142.5 210.6 143.7 212.7 ;
        RECT  139.5 210.6 140.7 211.8 ;
        RECT  136.5 210.6 137.7 211.8 ;
        RECT  133.5 210.6 134.7 212.7 ;
        RECT  132.3 212.7 143.7 213.9 ;
        RECT  132.3 201.3 143.7 202.5 ;
        RECT  132.3 212.7 143.7 213.9 ;
        RECT  138.6 226.2 141.3 227.4 ;
        RECT  134.4 226.2 137.1 227.4 ;
        RECT  132.3 224.1 143.7 225.3 ;
        RECT  138.0 223.8 139.2 224.1 ;
        RECT  142.5 216.9 143.7 222.6 ;
        RECT  140.1 221.4 141.3 222.6 ;
        RECT  135.9 221.4 137.1 222.6 ;
        RECT  139.8 220.8 141.0 221.4 ;
        RECT  139.2 219.6 141.0 220.8 ;
        RECT  139.8 216.0 141.0 219.6 ;
        RECT  136.2 218.1 137.4 221.4 ;
        RECT  136.2 216.9 138.6 218.1 ;
        RECT  133.5 216.9 134.7 222.6 ;
        RECT  136.2 216.0 137.4 216.9 ;
        RECT  142.5 213.9 143.7 216.0 ;
        RECT  139.5 214.8 140.7 216.0 ;
        RECT  136.5 214.8 137.7 216.0 ;
        RECT  133.5 213.9 134.7 216.0 ;
        RECT  132.3 212.7 143.7 213.9 ;
        RECT  132.3 224.1 143.7 225.3 ;
        RECT  132.3 212.7 143.7 213.9 ;
        RECT  138.6 227.4 141.3 228.6 ;
        RECT  134.4 227.4 137.1 228.6 ;
        RECT  132.3 229.5 143.7 230.7 ;
        RECT  138.0 230.7 139.2 231.0 ;
        RECT  142.5 232.2 143.7 237.9 ;
        RECT  140.1 232.2 141.3 233.4 ;
        RECT  135.9 232.2 137.1 233.4 ;
        RECT  139.8 233.4 141.0 234.0 ;
        RECT  139.2 234.0 141.0 235.2 ;
        RECT  139.8 235.2 141.0 238.8 ;
        RECT  136.2 233.4 137.4 236.7 ;
        RECT  136.2 236.7 138.6 237.9 ;
        RECT  133.5 232.2 134.7 237.9 ;
        RECT  136.2 237.9 137.4 238.8 ;
        RECT  142.5 238.8 143.7 240.9 ;
        RECT  139.5 238.8 140.7 240.0 ;
        RECT  136.5 238.8 137.7 240.0 ;
        RECT  133.5 238.8 134.7 240.9 ;
        RECT  132.3 240.9 143.7 242.1 ;
        RECT  132.3 229.5 143.7 230.7 ;
        RECT  132.3 240.9 143.7 242.1 ;
        RECT  138.6 254.4 141.3 255.6 ;
        RECT  134.4 254.4 137.1 255.6 ;
        RECT  132.3 252.3 143.7 253.5 ;
        RECT  138.0 252.0 139.2 252.3 ;
        RECT  142.5 245.1 143.7 250.8 ;
        RECT  140.1 249.6 141.3 250.8 ;
        RECT  135.9 249.6 137.1 250.8 ;
        RECT  139.8 249.0 141.0 249.6 ;
        RECT  139.2 247.8 141.0 249.0 ;
        RECT  139.8 244.2 141.0 247.8 ;
        RECT  136.2 246.3 137.4 249.6 ;
        RECT  136.2 245.1 138.6 246.3 ;
        RECT  133.5 245.1 134.7 250.8 ;
        RECT  136.2 244.2 137.4 245.1 ;
        RECT  142.5 242.1 143.7 244.2 ;
        RECT  139.5 243.0 140.7 244.2 ;
        RECT  136.5 243.0 137.7 244.2 ;
        RECT  133.5 242.1 134.7 244.2 ;
        RECT  132.3 240.9 143.7 242.1 ;
        RECT  132.3 252.3 143.7 253.5 ;
        RECT  132.3 240.9 143.7 242.1 ;
        RECT  138.6 255.6 141.3 256.8 ;
        RECT  134.4 255.6 137.1 256.8 ;
        RECT  132.3 257.7 143.7 258.9 ;
        RECT  138.0 258.9 139.2 259.2 ;
        RECT  142.5 260.4 143.7 266.1 ;
        RECT  140.1 260.4 141.3 261.6 ;
        RECT  135.9 260.4 137.1 261.6 ;
        RECT  139.8 261.6 141.0 262.2 ;
        RECT  139.2 262.2 141.0 263.4 ;
        RECT  139.8 263.4 141.0 267.0 ;
        RECT  136.2 261.6 137.4 264.9 ;
        RECT  136.2 264.9 138.6 266.1 ;
        RECT  133.5 260.4 134.7 266.1 ;
        RECT  136.2 266.1 137.4 267.0 ;
        RECT  142.5 267.0 143.7 269.1 ;
        RECT  139.5 267.0 140.7 268.2 ;
        RECT  136.5 267.0 137.7 268.2 ;
        RECT  133.5 267.0 134.7 269.1 ;
        RECT  132.3 269.1 143.7 270.3 ;
        RECT  132.3 257.7 143.7 258.9 ;
        RECT  132.3 269.1 143.7 270.3 ;
        RECT  138.6 282.6 141.3 283.8 ;
        RECT  134.4 282.6 137.1 283.8 ;
        RECT  132.3 280.5 143.7 281.7 ;
        RECT  138.0 280.2 139.2 280.5 ;
        RECT  142.5 273.3 143.7 279.0 ;
        RECT  140.1 277.8 141.3 279.0 ;
        RECT  135.9 277.8 137.1 279.0 ;
        RECT  139.8 277.2 141.0 277.8 ;
        RECT  139.2 276.0 141.0 277.2 ;
        RECT  139.8 272.4 141.0 276.0 ;
        RECT  136.2 274.5 137.4 277.8 ;
        RECT  136.2 273.3 138.6 274.5 ;
        RECT  133.5 273.3 134.7 279.0 ;
        RECT  136.2 272.4 137.4 273.3 ;
        RECT  142.5 270.3 143.7 272.4 ;
        RECT  139.5 271.2 140.7 272.4 ;
        RECT  136.5 271.2 137.7 272.4 ;
        RECT  133.5 270.3 134.7 272.4 ;
        RECT  132.3 269.1 143.7 270.3 ;
        RECT  132.3 280.5 143.7 281.7 ;
        RECT  132.3 269.1 143.7 270.3 ;
        RECT  138.6 283.8 141.3 285.0 ;
        RECT  134.4 283.8 137.1 285.0 ;
        RECT  132.3 285.9 143.7 287.1 ;
        RECT  138.0 287.1 139.2 287.4 ;
        RECT  142.5 288.6 143.7 294.3 ;
        RECT  140.1 288.6 141.3 289.8 ;
        RECT  135.9 288.6 137.1 289.8 ;
        RECT  139.8 289.8 141.0 290.4 ;
        RECT  139.2 290.4 141.0 291.6 ;
        RECT  139.8 291.6 141.0 295.2 ;
        RECT  136.2 289.8 137.4 293.1 ;
        RECT  136.2 293.1 138.6 294.3 ;
        RECT  133.5 288.6 134.7 294.3 ;
        RECT  136.2 294.3 137.4 295.2 ;
        RECT  142.5 295.2 143.7 297.3 ;
        RECT  139.5 295.2 140.7 296.4 ;
        RECT  136.5 295.2 137.7 296.4 ;
        RECT  133.5 295.2 134.7 297.3 ;
        RECT  132.3 297.3 143.7 298.5 ;
        RECT  132.3 285.9 143.7 287.1 ;
        RECT  132.3 297.3 143.7 298.5 ;
        RECT  138.6 310.8 141.3 312.0 ;
        RECT  134.4 310.8 137.1 312.0 ;
        RECT  132.3 308.7 143.7 309.9 ;
        RECT  138.0 308.4 139.2 308.7 ;
        RECT  142.5 301.5 143.7 307.2 ;
        RECT  140.1 306.0 141.3 307.2 ;
        RECT  135.9 306.0 137.1 307.2 ;
        RECT  139.8 305.4 141.0 306.0 ;
        RECT  139.2 304.2 141.0 305.4 ;
        RECT  139.8 300.6 141.0 304.2 ;
        RECT  136.2 302.7 137.4 306.0 ;
        RECT  136.2 301.5 138.6 302.7 ;
        RECT  133.5 301.5 134.7 307.2 ;
        RECT  136.2 300.6 137.4 301.5 ;
        RECT  142.5 298.5 143.7 300.6 ;
        RECT  139.5 299.4 140.7 300.6 ;
        RECT  136.5 299.4 137.7 300.6 ;
        RECT  133.5 298.5 134.7 300.6 ;
        RECT  132.3 297.3 143.7 298.5 ;
        RECT  132.3 308.7 143.7 309.9 ;
        RECT  132.3 297.3 143.7 298.5 ;
        RECT  138.6 312.0 141.3 313.2 ;
        RECT  134.4 312.0 137.1 313.2 ;
        RECT  132.3 314.1 143.7 315.3 ;
        RECT  138.0 315.3 139.2 315.6 ;
        RECT  142.5 316.8 143.7 322.5 ;
        RECT  140.1 316.8 141.3 318.0 ;
        RECT  135.9 316.8 137.1 318.0 ;
        RECT  139.8 318.0 141.0 318.6 ;
        RECT  139.2 318.6 141.0 319.8 ;
        RECT  139.8 319.8 141.0 323.4 ;
        RECT  136.2 318.0 137.4 321.3 ;
        RECT  136.2 321.3 138.6 322.5 ;
        RECT  133.5 316.8 134.7 322.5 ;
        RECT  136.2 322.5 137.4 323.4 ;
        RECT  142.5 323.4 143.7 325.5 ;
        RECT  139.5 323.4 140.7 324.6 ;
        RECT  136.5 323.4 137.7 324.6 ;
        RECT  133.5 323.4 134.7 325.5 ;
        RECT  132.3 325.5 143.7 326.7 ;
        RECT  132.3 314.1 143.7 315.3 ;
        RECT  132.3 325.5 143.7 326.7 ;
        RECT  138.6 339.0 141.3 340.2 ;
        RECT  134.4 339.0 137.1 340.2 ;
        RECT  132.3 336.9 143.7 338.1 ;
        RECT  138.0 336.6 139.2 336.9 ;
        RECT  142.5 329.7 143.7 335.4 ;
        RECT  140.1 334.2 141.3 335.4 ;
        RECT  135.9 334.2 137.1 335.4 ;
        RECT  139.8 333.6 141.0 334.2 ;
        RECT  139.2 332.4 141.0 333.6 ;
        RECT  139.8 328.8 141.0 332.4 ;
        RECT  136.2 330.9 137.4 334.2 ;
        RECT  136.2 329.7 138.6 330.9 ;
        RECT  133.5 329.7 134.7 335.4 ;
        RECT  136.2 328.8 137.4 329.7 ;
        RECT  142.5 326.7 143.7 328.8 ;
        RECT  139.5 327.6 140.7 328.8 ;
        RECT  136.5 327.6 137.7 328.8 ;
        RECT  133.5 326.7 134.7 328.8 ;
        RECT  132.3 325.5 143.7 326.7 ;
        RECT  132.3 336.9 143.7 338.1 ;
        RECT  132.3 325.5 143.7 326.7 ;
        RECT  138.6 340.2 141.3 341.4 ;
        RECT  134.4 340.2 137.1 341.4 ;
        RECT  132.3 342.3 143.7 343.5 ;
        RECT  138.0 343.5 139.2 343.8 ;
        RECT  142.5 345.0 143.7 350.7 ;
        RECT  140.1 345.0 141.3 346.2 ;
        RECT  135.9 345.0 137.1 346.2 ;
        RECT  139.8 346.2 141.0 346.8 ;
        RECT  139.2 346.8 141.0 348.0 ;
        RECT  139.8 348.0 141.0 351.6 ;
        RECT  136.2 346.2 137.4 349.5 ;
        RECT  136.2 349.5 138.6 350.7 ;
        RECT  133.5 345.0 134.7 350.7 ;
        RECT  136.2 350.7 137.4 351.6 ;
        RECT  142.5 351.6 143.7 353.7 ;
        RECT  139.5 351.6 140.7 352.8 ;
        RECT  136.5 351.6 137.7 352.8 ;
        RECT  133.5 351.6 134.7 353.7 ;
        RECT  132.3 353.7 143.7 354.9 ;
        RECT  132.3 342.3 143.7 343.5 ;
        RECT  132.3 353.7 143.7 354.9 ;
        RECT  138.6 367.2 141.3 368.4 ;
        RECT  134.4 367.2 137.1 368.4 ;
        RECT  132.3 365.1 143.7 366.3 ;
        RECT  138.0 364.8 139.2 365.1 ;
        RECT  142.5 357.9 143.7 363.6 ;
        RECT  140.1 362.4 141.3 363.6 ;
        RECT  135.9 362.4 137.1 363.6 ;
        RECT  139.8 361.8 141.0 362.4 ;
        RECT  139.2 360.6 141.0 361.8 ;
        RECT  139.8 357.0 141.0 360.6 ;
        RECT  136.2 359.1 137.4 362.4 ;
        RECT  136.2 357.9 138.6 359.1 ;
        RECT  133.5 357.9 134.7 363.6 ;
        RECT  136.2 357.0 137.4 357.9 ;
        RECT  142.5 354.9 143.7 357.0 ;
        RECT  139.5 355.8 140.7 357.0 ;
        RECT  136.5 355.8 137.7 357.0 ;
        RECT  133.5 354.9 134.7 357.0 ;
        RECT  132.3 353.7 143.7 354.9 ;
        RECT  132.3 365.1 143.7 366.3 ;
        RECT  132.3 353.7 143.7 354.9 ;
        RECT  138.6 368.4 141.3 369.6 ;
        RECT  134.4 368.4 137.1 369.6 ;
        RECT  132.3 370.5 143.7 371.7 ;
        RECT  138.0 371.7 139.2 372.0 ;
        RECT  142.5 373.2 143.7 378.9 ;
        RECT  140.1 373.2 141.3 374.4 ;
        RECT  135.9 373.2 137.1 374.4 ;
        RECT  139.8 374.4 141.0 375.0 ;
        RECT  139.2 375.0 141.0 376.2 ;
        RECT  139.8 376.2 141.0 379.8 ;
        RECT  136.2 374.4 137.4 377.7 ;
        RECT  136.2 377.7 138.6 378.9 ;
        RECT  133.5 373.2 134.7 378.9 ;
        RECT  136.2 378.9 137.4 379.8 ;
        RECT  142.5 379.8 143.7 381.9 ;
        RECT  139.5 379.8 140.7 381.0 ;
        RECT  136.5 379.8 137.7 381.0 ;
        RECT  133.5 379.8 134.7 381.9 ;
        RECT  132.3 381.9 143.7 383.1 ;
        RECT  132.3 370.5 143.7 371.7 ;
        RECT  132.3 381.9 143.7 383.1 ;
        RECT  138.6 395.4 141.3 396.6 ;
        RECT  134.4 395.4 137.1 396.6 ;
        RECT  132.3 393.3 143.7 394.5 ;
        RECT  138.0 393.0 139.2 393.3 ;
        RECT  142.5 386.1 143.7 391.8 ;
        RECT  140.1 390.6 141.3 391.8 ;
        RECT  135.9 390.6 137.1 391.8 ;
        RECT  139.8 390.0 141.0 390.6 ;
        RECT  139.2 388.8 141.0 390.0 ;
        RECT  139.8 385.2 141.0 388.8 ;
        RECT  136.2 387.3 137.4 390.6 ;
        RECT  136.2 386.1 138.6 387.3 ;
        RECT  133.5 386.1 134.7 391.8 ;
        RECT  136.2 385.2 137.4 386.1 ;
        RECT  142.5 383.1 143.7 385.2 ;
        RECT  139.5 384.0 140.7 385.2 ;
        RECT  136.5 384.0 137.7 385.2 ;
        RECT  133.5 383.1 134.7 385.2 ;
        RECT  132.3 381.9 143.7 383.1 ;
        RECT  132.3 393.3 143.7 394.5 ;
        RECT  132.3 381.9 143.7 383.1 ;
        RECT  138.6 396.6 141.3 397.8 ;
        RECT  134.4 396.6 137.1 397.8 ;
        RECT  132.3 398.7 143.7 399.9 ;
        RECT  138.0 399.9 139.2 400.2 ;
        RECT  142.5 401.4 143.7 407.1 ;
        RECT  140.1 401.4 141.3 402.6 ;
        RECT  135.9 401.4 137.1 402.6 ;
        RECT  139.8 402.6 141.0 403.2 ;
        RECT  139.2 403.2 141.0 404.4 ;
        RECT  139.8 404.4 141.0 408.0 ;
        RECT  136.2 402.6 137.4 405.9 ;
        RECT  136.2 405.9 138.6 407.1 ;
        RECT  133.5 401.4 134.7 407.1 ;
        RECT  136.2 407.1 137.4 408.0 ;
        RECT  142.5 408.0 143.7 410.1 ;
        RECT  139.5 408.0 140.7 409.2 ;
        RECT  136.5 408.0 137.7 409.2 ;
        RECT  133.5 408.0 134.7 410.1 ;
        RECT  132.3 410.1 143.7 411.3 ;
        RECT  132.3 398.7 143.7 399.9 ;
        RECT  132.3 410.1 143.7 411.3 ;
        RECT  138.6 423.6 141.3 424.8 ;
        RECT  134.4 423.6 137.1 424.8 ;
        RECT  132.3 421.5 143.7 422.7 ;
        RECT  138.0 421.2 139.2 421.5 ;
        RECT  142.5 414.3 143.7 420.0 ;
        RECT  140.1 418.8 141.3 420.0 ;
        RECT  135.9 418.8 137.1 420.0 ;
        RECT  139.8 418.2 141.0 418.8 ;
        RECT  139.2 417.0 141.0 418.2 ;
        RECT  139.8 413.4 141.0 417.0 ;
        RECT  136.2 415.5 137.4 418.8 ;
        RECT  136.2 414.3 138.6 415.5 ;
        RECT  133.5 414.3 134.7 420.0 ;
        RECT  136.2 413.4 137.4 414.3 ;
        RECT  142.5 411.3 143.7 413.4 ;
        RECT  139.5 412.2 140.7 413.4 ;
        RECT  136.5 412.2 137.7 413.4 ;
        RECT  133.5 411.3 134.7 413.4 ;
        RECT  132.3 410.1 143.7 411.3 ;
        RECT  132.3 421.5 143.7 422.7 ;
        RECT  132.3 410.1 143.7 411.3 ;
        RECT  122.7 429.6 143.1 430.5 ;
        RECT  122.7 443.7 143.1 444.6 ;
        RECT  128.1 436.2 129.3 444.6 ;
        RECT  122.7 443.7 132.9 444.6 ;
        RECT  122.7 429.6 132.9 430.5 ;
        RECT  125.7 427.2 126.9 428.4 ;
        RECT  128.1 427.2 129.3 428.4 ;
        RECT  125.7 427.2 126.9 428.4 ;
        RECT  128.1 427.2 129.3 428.4 ;
        RECT  125.7 436.2 126.9 437.4 ;
        RECT  128.1 436.2 129.3 437.4 ;
        RECT  125.7 436.2 126.9 437.4 ;
        RECT  128.1 436.2 129.3 437.4 ;
        RECT  128.1 436.2 129.3 437.4 ;
        RECT  130.5 436.2 131.7 437.4 ;
        RECT  128.1 436.2 129.3 437.4 ;
        RECT  130.5 436.2 131.7 437.4 ;
        RECT  126.6 429.45 127.8 430.65 ;
        RECT  128.1 442.8 129.3 444.0 ;
        RECT  125.7 427.2 126.9 428.4 ;
        RECT  128.1 427.2 129.3 428.4 ;
        RECT  125.7 436.2 126.9 437.4 ;
        RECT  130.5 436.2 131.7 437.4 ;
        RECT  125.7 427.2 126.9 428.4 ;
        RECT  128.1 427.2 129.3 428.4 ;
        RECT  125.7 436.2 126.9 437.4 ;
        RECT  130.5 436.2 131.7 437.4 ;
        RECT  138.3 436.2 139.5 444.6 ;
        RECT  132.9 443.7 143.1 444.6 ;
        RECT  132.9 429.6 143.1 430.5 ;
        RECT  135.9 427.2 137.1 428.4 ;
        RECT  138.3 427.2 139.5 428.4 ;
        RECT  135.9 427.2 137.1 428.4 ;
        RECT  138.3 427.2 139.5 428.4 ;
        RECT  135.9 436.2 137.1 437.4 ;
        RECT  138.3 436.2 139.5 437.4 ;
        RECT  135.9 436.2 137.1 437.4 ;
        RECT  138.3 436.2 139.5 437.4 ;
        RECT  138.3 436.2 139.5 437.4 ;
        RECT  140.7 436.2 141.9 437.4 ;
        RECT  138.3 436.2 139.5 437.4 ;
        RECT  140.7 436.2 141.9 437.4 ;
        RECT  136.8 429.45 138.0 430.65 ;
        RECT  138.3 442.8 139.5 444.0 ;
        RECT  135.9 427.2 137.1 428.4 ;
        RECT  138.3 427.2 139.5 428.4 ;
        RECT  135.9 436.2 137.1 437.4 ;
        RECT  140.7 436.2 141.9 437.4 ;
        RECT  135.9 427.2 137.1 428.4 ;
        RECT  138.3 427.2 139.5 428.4 ;
        RECT  135.9 436.2 137.1 437.4 ;
        RECT  140.7 436.2 141.9 437.4 ;
        RECT  122.7 195.0 143.1 195.9 ;
        RECT  122.7 167.7 143.1 168.6 ;
        RECT  122.7 192.9 143.1 193.8 ;
        RECT  122.1 195.0 133.5 196.2 ;
        RECT  122.1 192.9 133.5 194.1 ;
        RECT  127.5 189.3 128.7 192.0 ;
        RECT  129.9 189.3 131.1 192.9 ;
        RECT  132.3 191.7 133.5 192.9 ;
        RECT  127.5 185.4 128.4 189.3 ;
        RECT  124.8 171.0 126.0 185.4 ;
        RECT  127.2 182.7 128.4 185.4 ;
        RECT  129.6 181.8 130.8 185.4 ;
        RECT  129.6 180.6 131.7 181.8 ;
        RECT  127.2 173.7 128.4 179.1 ;
        RECT  129.6 173.7 130.8 180.6 ;
        RECT  127.2 172.8 128.1 173.7 ;
        RECT  127.2 171.9 129.0 172.8 ;
        RECT  124.8 169.8 126.6 171.0 ;
        RECT  128.1 170.1 129.0 171.9 ;
        RECT  128.1 168.9 129.3 170.1 ;
        RECT  122.1 167.7 133.5 168.9 ;
        RECT  125.4 166.5 126.6 166.8 ;
        RECT  124.5 165.6 126.6 166.5 ;
        RECT  131.4 165.6 132.9 166.8 ;
        RECT  124.5 163.5 125.4 165.6 ;
        RECT  126.6 163.5 127.8 164.7 ;
        RECT  124.5 157.2 125.7 163.5 ;
        RECT  123.6 156.3 125.7 157.2 ;
        RECT  126.9 156.3 128.1 163.5 ;
        RECT  129.3 156.3 130.5 164.7 ;
        RECT  132.0 163.5 132.9 165.6 ;
        RECT  131.7 156.3 132.9 163.5 ;
        RECT  123.6 153.6 124.8 156.3 ;
        RECT  122.1 195.0 133.5 196.2 ;
        RECT  122.1 167.7 133.5 168.9 ;
        RECT  122.1 192.9 133.5 194.1 ;
        RECT  132.3 195.0 143.7 196.2 ;
        RECT  132.3 192.9 143.7 194.1 ;
        RECT  137.7 189.3 138.9 192.0 ;
        RECT  140.1 189.3 141.3 192.9 ;
        RECT  142.5 191.7 143.7 192.9 ;
        RECT  137.7 185.4 138.6 189.3 ;
        RECT  135.0 171.0 136.2 185.4 ;
        RECT  137.4 182.7 138.6 185.4 ;
        RECT  139.8 181.8 141.0 185.4 ;
        RECT  139.8 180.6 141.9 181.8 ;
        RECT  137.4 173.7 138.6 179.1 ;
        RECT  139.8 173.7 141.0 180.6 ;
        RECT  137.4 172.8 138.3 173.7 ;
        RECT  137.4 171.9 139.2 172.8 ;
        RECT  135.0 169.8 136.8 171.0 ;
        RECT  138.3 170.1 139.2 171.9 ;
        RECT  138.3 168.9 139.5 170.1 ;
        RECT  132.3 167.7 143.7 168.9 ;
        RECT  135.6 166.5 136.8 166.8 ;
        RECT  134.7 165.6 136.8 166.5 ;
        RECT  141.6 165.6 143.1 166.8 ;
        RECT  134.7 163.5 135.6 165.6 ;
        RECT  136.8 163.5 138.0 164.7 ;
        RECT  134.7 157.2 135.9 163.5 ;
        RECT  133.8 156.3 135.9 157.2 ;
        RECT  137.1 156.3 138.3 163.5 ;
        RECT  139.5 156.3 140.7 164.7 ;
        RECT  142.2 163.5 143.1 165.6 ;
        RECT  141.9 156.3 143.1 163.5 ;
        RECT  133.8 153.6 135.0 156.3 ;
        RECT  132.3 195.0 143.7 196.2 ;
        RECT  132.3 167.7 143.7 168.9 ;
        RECT  132.3 192.9 143.7 194.1 ;
        RECT  122.7 96.9 143.1 97.8 ;
        RECT  122.7 99.0 143.1 99.9 ;
        RECT  122.7 94.8 143.1 95.7 ;
        RECT  124.2 147.0 125.4 148.2 ;
        RECT  124.2 146.4 125.1 147.0 ;
        RECT  123.9 142.8 125.1 146.4 ;
        RECT  126.3 142.8 127.5 146.4 ;
        RECT  128.7 142.8 129.9 147.6 ;
        RECT  131.1 144.0 132.6 145.2 ;
        RECT  126.6 140.4 127.5 142.8 ;
        RECT  123.9 127.2 125.1 139.8 ;
        RECT  126.6 139.2 130.8 140.4 ;
        RECT  126.0 136.8 130.8 138.0 ;
        RECT  126.3 132.9 127.5 136.8 ;
        RECT  128.7 132.3 129.9 134.1 ;
        RECT  131.7 132.3 132.6 144.0 ;
        RECT  128.7 131.1 132.6 132.3 ;
        RECT  126.3 126.3 127.5 129.3 ;
        RECT  128.7 127.2 129.9 131.1 ;
        RECT  122.7 125.1 133.5 126.3 ;
        RECT  124.2 120.9 125.4 123.9 ;
        RECT  126.6 121.8 127.8 125.1 ;
        RECT  129.0 120.9 130.2 123.9 ;
        RECT  124.2 120.0 130.2 120.9 ;
        RECT  124.2 114.3 125.4 120.0 ;
        RECT  129.0 119.7 130.2 120.0 ;
        RECT  129.0 118.5 130.8 119.7 ;
        RECT  126.6 114.3 127.8 116.4 ;
        RECT  129.0 115.5 130.2 116.4 ;
        RECT  129.0 114.3 132.9 115.5 ;
        RECT  129.6 112.2 132.0 113.4 ;
        RECT  123.6 111.0 124.8 112.2 ;
        RECT  123.9 108.9 124.8 111.0 ;
        RECT  123.6 105.0 124.8 108.9 ;
        RECT  126.0 106.8 127.2 108.9 ;
        RECT  128.4 106.8 129.6 110.1 ;
        RECT  123.6 104.1 127.2 105.0 ;
        RECT  123.6 100.2 124.8 103.2 ;
        RECT  126.0 101.1 127.2 104.1 ;
        RECT  128.4 100.2 129.6 103.2 ;
        RECT  130.8 101.1 132.0 112.2 ;
        RECT  122.7 99.0 133.5 100.2 ;
        RECT  122.7 96.9 133.5 98.1 ;
        RECT  122.7 94.8 133.5 96.0 ;
        RECT  126.3 92.7 128.7 93.9 ;
        RECT  122.7 96.9 133.5 98.1 ;
        RECT  122.7 99.0 133.5 100.2 ;
        RECT  122.7 94.8 133.5 96.0 ;
        RECT  134.4 147.0 135.6 148.2 ;
        RECT  134.4 146.4 135.3 147.0 ;
        RECT  134.1 142.8 135.3 146.4 ;
        RECT  136.5 142.8 137.7 146.4 ;
        RECT  138.9 142.8 140.1 147.6 ;
        RECT  141.3 144.0 142.8 145.2 ;
        RECT  136.8 140.4 137.7 142.8 ;
        RECT  134.1 127.2 135.3 139.8 ;
        RECT  136.8 139.2 141.0 140.4 ;
        RECT  136.2 136.8 141.0 138.0 ;
        RECT  136.5 132.9 137.7 136.8 ;
        RECT  138.9 132.3 140.1 134.1 ;
        RECT  141.9 132.3 142.8 144.0 ;
        RECT  138.9 131.1 142.8 132.3 ;
        RECT  136.5 126.3 137.7 129.3 ;
        RECT  138.9 127.2 140.1 131.1 ;
        RECT  132.9 125.1 143.7 126.3 ;
        RECT  134.4 120.9 135.6 123.9 ;
        RECT  136.8 121.8 138.0 125.1 ;
        RECT  139.2 120.9 140.4 123.9 ;
        RECT  134.4 120.0 140.4 120.9 ;
        RECT  134.4 114.3 135.6 120.0 ;
        RECT  139.2 119.7 140.4 120.0 ;
        RECT  139.2 118.5 141.0 119.7 ;
        RECT  136.8 114.3 138.0 116.4 ;
        RECT  139.2 115.5 140.4 116.4 ;
        RECT  139.2 114.3 143.1 115.5 ;
        RECT  139.8 112.2 142.2 113.4 ;
        RECT  133.8 111.0 135.0 112.2 ;
        RECT  134.1 108.9 135.0 111.0 ;
        RECT  133.8 105.0 135.0 108.9 ;
        RECT  136.2 106.8 137.4 108.9 ;
        RECT  138.6 106.8 139.8 110.1 ;
        RECT  133.8 104.1 137.4 105.0 ;
        RECT  133.8 100.2 135.0 103.2 ;
        RECT  136.2 101.1 137.4 104.1 ;
        RECT  138.6 100.2 139.8 103.2 ;
        RECT  141.0 101.1 142.2 112.2 ;
        RECT  132.9 99.0 143.7 100.2 ;
        RECT  132.9 96.9 143.7 98.1 ;
        RECT  132.9 94.8 143.7 96.0 ;
        RECT  136.5 92.7 138.9 93.9 ;
        RECT  132.9 96.9 143.7 98.1 ;
        RECT  132.9 99.0 143.7 100.2 ;
        RECT  132.9 94.8 143.7 96.0 ;
        RECT  122.7 32.4 143.1 33.3 ;
        RECT  122.7 86.4 143.1 87.3 ;
        RECT  122.1 86.4 133.5 87.3 ;
        RECT  122.1 83.1 123.3 86.4 ;
        RECT  124.5 84.6 131.1 85.5 ;
        RECT  124.5 84.3 127.5 84.6 ;
        RECT  129.9 84.3 131.1 84.6 ;
        RECT  122.1 81.9 126.3 83.1 ;
        RECT  129.9 81.9 133.5 83.1 ;
        RECT  122.1 78.3 123.3 81.9 ;
        RECT  127.5 81.0 128.7 81.9 ;
        RECT  127.5 80.7 129.9 81.0 ;
        RECT  124.5 79.8 131.1 80.7 ;
        RECT  124.5 79.5 126.3 79.8 ;
        RECT  129.9 79.5 131.1 79.8 ;
        RECT  122.1 77.1 126.3 78.3 ;
        RECT  122.1 63.3 123.3 77.1 ;
        RECT  127.8 76.5 129.0 78.9 ;
        RECT  132.6 78.3 133.5 81.9 ;
        RECT  129.9 77.1 133.5 78.3 ;
        RECT  132.3 75.9 133.5 77.1 ;
        RECT  124.5 73.5 125.7 74.7 ;
        RECT  126.6 74.4 129.0 75.6 ;
        RECT  124.5 72.6 131.1 73.5 ;
        RECT  124.5 72.3 126.3 72.6 ;
        RECT  129.9 72.3 131.1 72.6 ;
        RECT  124.5 70.2 131.1 71.1 ;
        RECT  124.5 69.9 126.3 70.2 ;
        RECT  128.7 69.9 131.1 70.2 ;
        RECT  124.5 67.8 131.1 68.7 ;
        RECT  124.5 67.5 126.3 67.8 ;
        RECT  128.7 67.5 131.1 67.8 ;
        RECT  127.5 65.7 128.7 66.6 ;
        RECT  124.5 64.8 131.1 65.7 ;
        RECT  124.5 64.5 127.5 64.8 ;
        RECT  129.9 64.5 131.1 64.8 ;
        RECT  122.1 62.1 126.3 63.3 ;
        RECT  122.1 57.6 123.3 62.1 ;
        RECT  127.2 61.2 128.4 63.6 ;
        RECT  132.6 63.3 133.5 75.9 ;
        RECT  129.9 62.1 133.5 63.3 ;
        RECT  124.5 60.0 125.7 61.2 ;
        RECT  124.5 59.1 131.1 60.0 ;
        RECT  124.5 58.8 126.3 59.1 ;
        RECT  129.9 58.8 131.1 59.1 ;
        RECT  132.6 57.6 133.5 62.1 ;
        RECT  122.1 56.4 126.3 57.6 ;
        RECT  122.1 52.8 123.3 56.4 ;
        RECT  127.8 55.5 129.0 56.7 ;
        RECT  129.9 56.4 133.5 57.6 ;
        RECT  124.5 55.2 129.9 55.5 ;
        RECT  124.5 54.6 131.1 55.2 ;
        RECT  124.5 54.0 126.3 54.6 ;
        RECT  128.7 54.3 131.1 54.6 ;
        RECT  129.9 54.0 131.1 54.3 ;
        RECT  122.1 51.6 126.3 52.8 ;
        RECT  122.1 36.6 123.3 51.6 ;
        RECT  127.8 51.0 129.0 53.4 ;
        RECT  132.6 52.8 133.5 56.4 ;
        RECT  129.9 51.6 133.5 52.8 ;
        RECT  132.3 50.4 133.5 51.6 ;
        RECT  124.5 47.1 125.7 48.3 ;
        RECT  126.6 48.0 129.0 49.2 ;
        RECT  124.5 46.2 131.1 47.1 ;
        RECT  124.5 45.9 126.3 46.2 ;
        RECT  129.9 45.9 131.1 46.2 ;
        RECT  124.5 43.8 131.1 44.7 ;
        RECT  124.5 43.5 126.3 43.8 ;
        RECT  128.7 43.5 131.1 43.8 ;
        RECT  124.5 41.4 131.1 42.3 ;
        RECT  124.5 41.1 126.3 41.4 ;
        RECT  128.7 41.1 131.1 41.4 ;
        RECT  127.5 39.3 128.7 40.2 ;
        RECT  124.5 38.4 131.1 39.3 ;
        RECT  124.5 38.1 127.5 38.4 ;
        RECT  129.9 38.1 131.1 38.4 ;
        RECT  132.6 36.9 133.5 50.4 ;
        RECT  124.5 36.6 126.3 36.9 ;
        RECT  122.1 35.7 126.3 36.6 ;
        RECT  129.9 36.0 133.5 36.9 ;
        RECT  129.9 35.7 131.1 36.0 ;
        RECT  125.1 34.2 126.3 35.7 ;
        RECT  127.2 33.3 128.4 34.2 ;
        RECT  122.1 32.4 133.5 33.3 ;
        RECT  122.1 32.4 133.5 33.3 ;
        RECT  122.1 86.4 133.5 87.3 ;
        RECT  132.3 86.4 143.7 87.3 ;
        RECT  142.5 83.1 143.7 86.4 ;
        RECT  134.7 84.6 141.3 85.5 ;
        RECT  138.3 84.3 141.3 84.6 ;
        RECT  134.7 84.3 135.9 84.6 ;
        RECT  139.5 81.9 143.7 83.1 ;
        RECT  132.3 81.9 135.9 83.1 ;
        RECT  142.5 78.3 143.7 81.9 ;
        RECT  137.1 81.0 138.3 81.9 ;
        RECT  135.9 80.7 138.3 81.0 ;
        RECT  134.7 79.8 141.3 80.7 ;
        RECT  139.5 79.5 141.3 79.8 ;
        RECT  134.7 79.5 135.9 79.8 ;
        RECT  139.5 77.1 143.7 78.3 ;
        RECT  142.5 63.3 143.7 77.1 ;
        RECT  136.8 76.5 138.0 78.9 ;
        RECT  132.3 78.3 133.2 81.9 ;
        RECT  132.3 77.1 135.9 78.3 ;
        RECT  132.3 75.9 133.5 77.1 ;
        RECT  140.1 73.5 141.3 74.7 ;
        RECT  136.8 74.4 139.2 75.6 ;
        RECT  134.7 72.6 141.3 73.5 ;
        RECT  139.5 72.3 141.3 72.6 ;
        RECT  134.7 72.3 135.9 72.6 ;
        RECT  134.7 70.2 141.3 71.1 ;
        RECT  139.5 69.9 141.3 70.2 ;
        RECT  134.7 69.9 137.1 70.2 ;
        RECT  134.7 67.8 141.3 68.7 ;
        RECT  139.5 67.5 141.3 67.8 ;
        RECT  134.7 67.5 137.1 67.8 ;
        RECT  137.1 65.7 138.3 66.6 ;
        RECT  134.7 64.8 141.3 65.7 ;
        RECT  138.3 64.5 141.3 64.8 ;
        RECT  134.7 64.5 135.9 64.8 ;
        RECT  139.5 62.1 143.7 63.3 ;
        RECT  142.5 57.6 143.7 62.1 ;
        RECT  137.4 61.2 138.6 63.6 ;
        RECT  132.3 63.3 133.2 75.9 ;
        RECT  132.3 62.1 135.9 63.3 ;
        RECT  140.1 60.0 141.3 61.2 ;
        RECT  134.7 59.1 141.3 60.0 ;
        RECT  139.5 58.8 141.3 59.1 ;
        RECT  134.7 58.8 135.9 59.1 ;
        RECT  132.3 57.6 133.2 62.1 ;
        RECT  139.5 56.4 143.7 57.6 ;
        RECT  142.5 52.8 143.7 56.4 ;
        RECT  136.8 55.5 138.0 56.7 ;
        RECT  132.3 56.4 135.9 57.6 ;
        RECT  135.9 55.2 141.3 55.5 ;
        RECT  134.7 54.6 141.3 55.2 ;
        RECT  139.5 54.0 141.3 54.6 ;
        RECT  134.7 54.3 137.1 54.6 ;
        RECT  134.7 54.0 135.9 54.3 ;
        RECT  139.5 51.6 143.7 52.8 ;
        RECT  142.5 36.6 143.7 51.6 ;
        RECT  136.8 51.0 138.0 53.4 ;
        RECT  132.3 52.8 133.2 56.4 ;
        RECT  132.3 51.6 135.9 52.8 ;
        RECT  132.3 50.4 133.5 51.6 ;
        RECT  140.1 47.1 141.3 48.3 ;
        RECT  136.8 48.0 139.2 49.2 ;
        RECT  134.7 46.2 141.3 47.1 ;
        RECT  139.5 45.9 141.3 46.2 ;
        RECT  134.7 45.9 135.9 46.2 ;
        RECT  134.7 43.8 141.3 44.7 ;
        RECT  139.5 43.5 141.3 43.8 ;
        RECT  134.7 43.5 137.1 43.8 ;
        RECT  134.7 41.4 141.3 42.3 ;
        RECT  139.5 41.1 141.3 41.4 ;
        RECT  134.7 41.1 137.1 41.4 ;
        RECT  137.1 39.3 138.3 40.2 ;
        RECT  134.7 38.4 141.3 39.3 ;
        RECT  138.3 38.1 141.3 38.4 ;
        RECT  134.7 38.1 135.9 38.4 ;
        RECT  132.3 36.9 133.2 50.4 ;
        RECT  139.5 36.6 141.3 36.9 ;
        RECT  139.5 35.7 143.7 36.6 ;
        RECT  132.3 36.0 135.9 36.9 ;
        RECT  134.7 35.7 135.9 36.0 ;
        RECT  139.5 34.2 140.7 35.7 ;
        RECT  137.4 33.3 138.6 34.2 ;
        RECT  132.3 32.4 143.7 33.3 ;
        RECT  132.3 32.4 143.7 33.3 ;
        RECT  132.3 86.4 143.7 87.3 ;
        RECT  122.7 25.5 143.1 26.4 ;
        RECT  122.7 9.6 143.1 10.5 ;
        RECT  122.7 23.4 143.1 24.3 ;
        RECT  122.7 27.9 143.1 28.8 ;
        RECT  122.7 49.5 133.5 50.7 ;
        RECT  123.6 45.9 125.1 48.3 ;
        RECT  126.3 45.9 127.5 49.5 ;
        RECT  128.7 45.9 129.9 48.3 ;
        RECT  131.1 45.9 132.3 48.3 ;
        RECT  123.6 42.6 124.5 45.9 ;
        RECT  125.4 43.8 126.6 45.0 ;
        RECT  123.6 41.4 128.7 42.6 ;
        RECT  131.4 41.4 132.3 45.9 ;
        RECT  123.6 39.3 124.5 41.4 ;
        RECT  130.2 40.2 132.3 41.4 ;
        RECT  131.4 39.3 132.3 40.2 ;
        RECT  123.6 38.1 125.1 39.3 ;
        RECT  126.3 36.9 127.5 39.3 ;
        RECT  128.7 38.1 129.9 39.3 ;
        RECT  131.1 38.1 132.3 39.3 ;
        RECT  122.7 35.7 133.5 36.9 ;
        RECT  122.7 33.6 133.5 34.8 ;
        RECT  122.7 31.2 133.5 32.4 ;
        RECT  122.7 33.6 133.5 34.8 ;
        RECT  122.7 49.5 133.5 50.7 ;
        RECT  122.7 35.7 133.5 36.9 ;
        RECT  122.7 35.7 133.5 36.9 ;
        RECT  122.7 31.2 133.5 32.4 ;
        RECT  132.9 49.5 143.7 50.7 ;
        RECT  133.8 45.9 135.3 48.3 ;
        RECT  136.5 45.9 137.7 49.5 ;
        RECT  138.9 45.9 140.1 48.3 ;
        RECT  141.3 45.9 142.5 48.3 ;
        RECT  133.8 42.6 134.7 45.9 ;
        RECT  135.6 43.8 136.8 45.0 ;
        RECT  133.8 41.4 138.9 42.6 ;
        RECT  141.6 41.4 142.5 45.9 ;
        RECT  133.8 39.3 134.7 41.4 ;
        RECT  140.4 40.2 142.5 41.4 ;
        RECT  141.6 39.3 142.5 40.2 ;
        RECT  133.8 38.1 135.3 39.3 ;
        RECT  136.5 36.9 137.7 39.3 ;
        RECT  138.9 38.1 140.1 39.3 ;
        RECT  141.3 38.1 142.5 39.3 ;
        RECT  132.9 35.7 143.7 36.9 ;
        RECT  132.9 33.6 143.7 34.8 ;
        RECT  132.9 31.2 143.7 32.4 ;
        RECT  132.9 33.6 143.7 34.8 ;
        RECT  132.9 49.5 143.7 50.7 ;
        RECT  132.9 35.7 143.7 36.9 ;
        RECT  132.9 35.7 143.7 36.9 ;
        RECT  132.9 31.2 143.7 32.4 ;
        RECT  34.95 206.55 35.85 207.45 ;
        RECT  34.95 205.2 35.85 206.1 ;
        RECT  30.9 206.55 35.4 207.45 ;
        RECT  34.95 205.65 35.85 207.0 ;
        RECT  35.4 205.2 39.9 206.1 ;
        RECT  34.95 219.15 35.85 220.05 ;
        RECT  34.95 220.5 35.85 221.4 ;
        RECT  30.9 219.15 35.4 220.05 ;
        RECT  34.95 219.6 35.85 220.95 ;
        RECT  35.4 220.5 39.9 221.4 ;
        RECT  34.95 234.75 35.85 235.65 ;
        RECT  34.95 233.4 35.85 234.3 ;
        RECT  30.9 234.75 35.4 235.65 ;
        RECT  34.95 233.85 35.85 235.2 ;
        RECT  35.4 233.4 39.9 234.3 ;
        RECT  34.95 247.35 35.85 248.25 ;
        RECT  34.95 248.7 35.85 249.6 ;
        RECT  30.9 247.35 35.4 248.25 ;
        RECT  34.95 247.8 35.85 249.15 ;
        RECT  35.4 248.7 39.9 249.6 ;
        RECT  34.95 262.95 35.85 263.85 ;
        RECT  34.95 261.6 35.85 262.5 ;
        RECT  30.9 262.95 35.4 263.85 ;
        RECT  34.95 262.05 35.85 263.4 ;
        RECT  35.4 261.6 39.9 262.5 ;
        RECT  34.95 275.55 35.85 276.45 ;
        RECT  34.95 276.9 35.85 277.8 ;
        RECT  30.9 275.55 35.4 276.45 ;
        RECT  34.95 276.0 35.85 277.35 ;
        RECT  35.4 276.9 39.9 277.8 ;
        RECT  34.95 291.15 35.85 292.05 ;
        RECT  34.95 289.8 35.85 290.7 ;
        RECT  30.9 291.15 35.4 292.05 ;
        RECT  34.95 290.25 35.85 291.6 ;
        RECT  35.4 289.8 39.9 290.7 ;
        RECT  34.95 303.75 35.85 304.65 ;
        RECT  34.95 305.1 35.85 306.0 ;
        RECT  30.9 303.75 35.4 304.65 ;
        RECT  34.95 304.2 35.85 305.55 ;
        RECT  35.4 305.1 39.9 306.0 ;
        RECT  34.95 319.35 35.85 320.25 ;
        RECT  34.95 318.0 35.85 318.9 ;
        RECT  30.9 319.35 35.4 320.25 ;
        RECT  34.95 318.45 35.85 319.8 ;
        RECT  35.4 318.0 39.9 318.9 ;
        RECT  34.95 331.95 35.85 332.85 ;
        RECT  34.95 333.3 35.85 334.2 ;
        RECT  30.9 331.95 35.4 332.85 ;
        RECT  34.95 332.4 35.85 333.75 ;
        RECT  35.4 333.3 39.9 334.2 ;
        RECT  34.95 347.55 35.85 348.45 ;
        RECT  34.95 346.2 35.85 347.1 ;
        RECT  30.9 347.55 35.4 348.45 ;
        RECT  34.95 346.65 35.85 348.0 ;
        RECT  35.4 346.2 39.9 347.1 ;
        RECT  34.95 360.15 35.85 361.05 ;
        RECT  34.95 361.5 35.85 362.4 ;
        RECT  30.9 360.15 35.4 361.05 ;
        RECT  34.95 360.6 35.85 361.95 ;
        RECT  35.4 361.5 39.9 362.4 ;
        RECT  34.95 375.75 35.85 376.65 ;
        RECT  34.95 374.4 35.85 375.3 ;
        RECT  30.9 375.75 35.4 376.65 ;
        RECT  34.95 374.85 35.85 376.2 ;
        RECT  35.4 374.4 39.9 375.3 ;
        RECT  34.95 388.35 35.85 389.25 ;
        RECT  34.95 389.7 35.85 390.6 ;
        RECT  30.9 388.35 35.4 389.25 ;
        RECT  34.95 388.8 35.85 390.15 ;
        RECT  35.4 389.7 39.9 390.6 ;
        RECT  34.95 403.95 35.85 404.85 ;
        RECT  34.95 402.6 35.85 403.5 ;
        RECT  30.9 403.95 35.4 404.85 ;
        RECT  34.95 403.05 35.85 404.4 ;
        RECT  35.4 402.6 39.9 403.5 ;
        RECT  34.95 416.55 35.85 417.45 ;
        RECT  34.95 417.9 35.85 418.8 ;
        RECT  30.9 416.55 35.4 417.45 ;
        RECT  34.95 417.0 35.85 418.35 ;
        RECT  35.4 417.9 39.9 418.8 ;
        RECT  6.75 92.4 23.1 93.3 ;
        RECT  8.85 107.7 23.1 108.6 ;
        RECT  10.95 120.6 23.1 121.5 ;
        RECT  13.05 135.9 23.1 136.8 ;
        RECT  15.15 148.8 23.1 149.7 ;
        RECT  17.25 164.1 23.1 165.0 ;
        RECT  19.35 177.0 23.1 177.9 ;
        RECT  21.45 192.3 23.1 193.2 ;
        RECT  6.75 206.55 25.5 207.45 ;
        RECT  15.15 203.85 28.5 204.75 ;
        RECT  6.75 219.15 25.5 220.05 ;
        RECT  17.25 221.85 28.5 222.75 ;
        RECT  6.75 234.75 25.5 235.65 ;
        RECT  19.35 232.05 28.5 232.95 ;
        RECT  6.75 247.35 25.5 248.25 ;
        RECT  21.45 250.05 28.5 250.95 ;
        RECT  8.85 262.95 25.5 263.85 ;
        RECT  15.15 260.25 28.5 261.15 ;
        RECT  8.85 275.55 25.5 276.45 ;
        RECT  17.25 278.25 28.5 279.15 ;
        RECT  8.85 291.15 25.5 292.05 ;
        RECT  19.35 288.45 28.5 289.35 ;
        RECT  8.85 303.75 25.5 304.65 ;
        RECT  21.45 306.45 28.5 307.35 ;
        RECT  10.95 319.35 25.5 320.25 ;
        RECT  15.15 316.65 28.5 317.55 ;
        RECT  10.95 331.95 25.5 332.85 ;
        RECT  17.25 334.65 28.5 335.55 ;
        RECT  10.95 347.55 25.5 348.45 ;
        RECT  19.35 344.85 28.5 345.75 ;
        RECT  10.95 360.15 25.5 361.05 ;
        RECT  21.45 362.85 28.5 363.75 ;
        RECT  13.05 375.75 25.5 376.65 ;
        RECT  15.15 373.05 28.5 373.95 ;
        RECT  13.05 388.35 25.5 389.25 ;
        RECT  17.25 391.05 28.5 391.95 ;
        RECT  13.05 403.95 25.5 404.85 ;
        RECT  19.35 401.25 28.5 402.15 ;
        RECT  13.05 416.55 25.5 417.45 ;
        RECT  21.45 419.25 28.5 420.15 ;
        RECT  42.45 305.1 43.35 306.0 ;
        RECT  42.45 276.9 43.35 277.8 ;
        RECT  42.45 346.2 43.35 347.1 ;
        RECT  42.45 220.5 43.35 221.4 ;
        RECT  42.45 248.7 43.35 249.6 ;
        RECT  42.45 374.4 43.35 375.3 ;
        RECT  42.45 318.0 43.35 318.9 ;
        RECT  42.45 402.6 43.35 403.5 ;
        RECT  42.45 289.8 43.35 290.7 ;
        RECT  42.45 205.2 43.35 206.1 ;
        RECT  42.45 261.6 43.35 262.5 ;
        RECT  42.45 233.4 43.35 234.3 ;
        RECT  42.45 389.7 43.35 390.6 ;
        RECT  42.45 333.3 43.35 334.2 ;
        RECT  42.45 417.9 43.35 418.8 ;
        RECT  42.45 361.5 43.35 362.4 ;
        RECT  6.3 100.05 77.7 100.95 ;
        RECT  6.3 128.25 77.7 129.15 ;
        RECT  6.3 156.45 77.7 157.35 ;
        RECT  6.3 184.65 77.7 185.55 ;
        RECT  6.3 212.85 77.7 213.75 ;
        RECT  6.3 241.05 77.7 241.95 ;
        RECT  6.3 269.25 77.7 270.15 ;
        RECT  6.3 297.45 77.7 298.35 ;
        RECT  6.3 325.65 77.7 326.55 ;
        RECT  6.3 353.85 77.7 354.75 ;
        RECT  6.3 382.05 77.7 382.95 ;
        RECT  6.3 410.25 77.7 411.15 ;
        RECT  6.3 85.95 77.7 86.85 ;
        RECT  6.3 114.15 77.7 115.05 ;
        RECT  6.3 142.35 77.7 143.25 ;
        RECT  6.3 170.55 77.7 171.45 ;
        RECT  6.3 198.75 77.7 199.65 ;
        RECT  6.3 226.95 77.7 227.85 ;
        RECT  6.3 255.15 77.7 256.05 ;
        RECT  6.3 283.35 77.7 284.25 ;
        RECT  6.3 311.55 77.7 312.45 ;
        RECT  6.3 339.75 77.7 340.65 ;
        RECT  6.3 367.95 77.7 368.85 ;
        RECT  6.3 396.15 77.7 397.05 ;
        RECT  6.3 424.35 77.7 425.25 ;
        RECT  60.75 92.4 61.65 93.3 ;
        RECT  60.75 97.35 61.65 98.25 ;
        RECT  61.2 92.4 65.85 93.3 ;
        RECT  60.75 92.85 61.65 97.8 ;
        RECT  58.65 97.35 61.2 98.25 ;
        RECT  69.3 92.4 77.25 93.3 ;
        RECT  60.75 107.7 61.65 108.6 ;
        RECT  60.75 111.45 61.65 112.35 ;
        RECT  61.2 107.7 65.85 108.6 ;
        RECT  60.75 108.15 61.65 111.9 ;
        RECT  55.65 111.45 61.2 112.35 ;
        RECT  69.3 107.7 74.25 108.6 ;
        RECT  52.65 116.25 77.25 117.15 ;
        RECT  49.65 130.35 74.25 131.25 ;
        RECT  44.7 93.75 58.65 94.65 ;
        RECT  41.7 91.05 55.65 91.95 ;
        RECT  44.7 106.35 52.65 107.25 ;
        RECT  41.7 109.05 55.65 109.95 ;
        RECT  44.7 121.95 58.65 122.85 ;
        RECT  41.7 119.25 49.65 120.15 ;
        RECT  44.7 134.55 52.65 135.45 ;
        RECT  41.7 137.25 49.65 138.15 ;
        RECT  34.35 93.75 35.25 94.65 ;
        RECT  34.35 92.4 35.25 93.3 ;
        RECT  34.8 93.75 39.3 94.65 ;
        RECT  34.35 92.85 35.25 94.2 ;
        RECT  30.3 92.4 34.8 93.3 ;
        RECT  34.35 106.35 35.25 107.25 ;
        RECT  34.35 107.7 35.25 108.6 ;
        RECT  34.8 106.35 39.3 107.25 ;
        RECT  34.35 106.8 35.25 108.15 ;
        RECT  30.3 107.7 34.8 108.6 ;
        RECT  34.35 121.95 35.25 122.85 ;
        RECT  34.35 120.6 35.25 121.5 ;
        RECT  34.8 121.95 39.3 122.85 ;
        RECT  34.35 121.05 35.25 122.4 ;
        RECT  30.3 120.6 34.8 121.5 ;
        RECT  34.35 134.55 35.25 135.45 ;
        RECT  34.35 135.9 35.25 136.8 ;
        RECT  34.8 134.55 39.3 135.45 ;
        RECT  34.35 135.0 35.25 136.35 ;
        RECT  30.3 135.9 34.8 136.8 ;
        RECT  23.1 135.9 26.85 136.8 ;
        RECT  23.1 120.6 26.85 121.5 ;
        RECT  23.1 92.4 26.85 93.3 ;
        RECT  23.1 107.7 26.85 108.6 ;
        RECT  23.1 100.05 77.7 100.95 ;
        RECT  23.1 128.25 77.7 129.15 ;
        RECT  23.1 85.95 77.7 86.85 ;
        RECT  23.1 114.15 77.7 115.05 ;
        RECT  23.1 142.35 77.7 143.25 ;
        RECT  63.9 84.45 65.1 86.4 ;
        RECT  63.9 72.3 65.1 74.25 ;
        RECT  68.7 85.05 69.9 86.85 ;
        RECT  68.7 71.85 69.9 75.45 ;
        RECT  66.3 75.45 67.2 83.85 ;
        RECT  68.1 79.35 69.3 80.55 ;
        RECT  65.85 79.5 66.75 80.4 ;
        RECT  62.1 71.85 71.7 72.75 ;
        RECT  62.1 85.95 71.7 86.85 ;
        RECT  68.7 74.25 69.9 75.45 ;
        RECT  66.3 74.25 67.5 75.45 ;
        RECT  68.7 74.25 69.9 75.45 ;
        RECT  66.3 74.25 67.5 75.45 ;
        RECT  68.7 83.85 69.9 85.05 ;
        RECT  66.3 83.85 67.5 85.05 ;
        RECT  68.7 83.85 69.9 85.05 ;
        RECT  66.3 83.85 67.5 85.05 ;
        RECT  63.9 83.85 65.1 85.05 ;
        RECT  63.9 73.65 65.1 74.85 ;
        RECT  68.1 79.35 69.3 80.55 ;
        RECT  63.9 114.6 65.1 116.55 ;
        RECT  63.9 126.75 65.1 128.7 ;
        RECT  68.7 114.15 69.9 115.95 ;
        RECT  68.7 125.55 69.9 129.15 ;
        RECT  66.3 117.15 67.2 125.55 ;
        RECT  68.1 120.45 69.3 121.65 ;
        RECT  65.85 120.6 66.75 121.5 ;
        RECT  62.1 128.25 71.7 129.15 ;
        RECT  62.1 114.15 71.7 115.05 ;
        RECT  68.7 123.15 69.9 124.35 ;
        RECT  66.3 123.15 67.5 124.35 ;
        RECT  68.7 123.15 69.9 124.35 ;
        RECT  66.3 123.15 67.5 124.35 ;
        RECT  68.7 114.75 69.9 115.95 ;
        RECT  66.3 114.75 67.5 115.95 ;
        RECT  68.7 114.75 69.9 115.95 ;
        RECT  66.3 114.75 67.5 115.95 ;
        RECT  63.9 114.75 65.1 115.95 ;
        RECT  63.9 124.95 65.1 126.15 ;
        RECT  68.1 119.25 69.3 120.45 ;
        RECT  24.9 84.45 26.1 86.4 ;
        RECT  24.9 72.3 26.1 74.25 ;
        RECT  29.7 85.05 30.9 86.85 ;
        RECT  29.7 71.85 30.9 75.45 ;
        RECT  27.3 75.45 28.2 83.85 ;
        RECT  29.1 79.35 30.3 80.55 ;
        RECT  26.85 79.5 27.75 80.4 ;
        RECT  23.1 71.85 32.7 72.75 ;
        RECT  23.1 85.95 32.7 86.85 ;
        RECT  29.7 74.25 30.9 75.45 ;
        RECT  27.3 74.25 28.5 75.45 ;
        RECT  29.7 74.25 30.9 75.45 ;
        RECT  27.3 74.25 28.5 75.45 ;
        RECT  29.7 83.85 30.9 85.05 ;
        RECT  27.3 83.85 28.5 85.05 ;
        RECT  29.7 83.85 30.9 85.05 ;
        RECT  27.3 83.85 28.5 85.05 ;
        RECT  24.9 83.85 26.1 85.05 ;
        RECT  24.9 73.65 26.1 74.85 ;
        RECT  29.1 79.35 30.3 80.55 ;
        RECT  24.9 114.6 26.1 116.55 ;
        RECT  24.9 126.75 26.1 128.7 ;
        RECT  29.7 114.15 30.9 115.95 ;
        RECT  29.7 125.55 30.9 129.15 ;
        RECT  27.3 117.15 28.2 125.55 ;
        RECT  29.1 120.45 30.3 121.65 ;
        RECT  26.85 120.6 27.75 121.5 ;
        RECT  23.1 128.25 32.7 129.15 ;
        RECT  23.1 114.15 32.7 115.05 ;
        RECT  29.7 123.15 30.9 124.35 ;
        RECT  27.3 123.15 28.5 124.35 ;
        RECT  29.7 123.15 30.9 124.35 ;
        RECT  27.3 123.15 28.5 124.35 ;
        RECT  29.7 114.75 30.9 115.95 ;
        RECT  27.3 114.75 28.5 115.95 ;
        RECT  29.7 114.75 30.9 115.95 ;
        RECT  27.3 114.75 28.5 115.95 ;
        RECT  24.9 114.75 26.1 115.95 ;
        RECT  24.9 124.95 26.1 126.15 ;
        RECT  29.1 119.25 30.3 120.45 ;
        RECT  24.9 112.65 26.1 114.6 ;
        RECT  24.9 100.5 26.1 102.45 ;
        RECT  29.7 113.25 30.9 115.05 ;
        RECT  29.7 100.05 30.9 103.65 ;
        RECT  27.3 103.65 28.2 112.05 ;
        RECT  29.1 107.55 30.3 108.75 ;
        RECT  26.85 107.7 27.75 108.6 ;
        RECT  23.1 100.05 32.7 100.95 ;
        RECT  23.1 114.15 32.7 115.05 ;
        RECT  29.7 102.45 30.9 103.65 ;
        RECT  27.3 102.45 28.5 103.65 ;
        RECT  29.7 102.45 30.9 103.65 ;
        RECT  27.3 102.45 28.5 103.65 ;
        RECT  29.7 112.05 30.9 113.25 ;
        RECT  27.3 112.05 28.5 113.25 ;
        RECT  29.7 112.05 30.9 113.25 ;
        RECT  27.3 112.05 28.5 113.25 ;
        RECT  24.9 112.05 26.1 113.25 ;
        RECT  24.9 101.85 26.1 103.05 ;
        RECT  29.1 107.55 30.3 108.75 ;
        RECT  24.9 142.8 26.1 144.75 ;
        RECT  24.9 154.95 26.1 156.9 ;
        RECT  29.7 142.35 30.9 144.15 ;
        RECT  29.7 153.75 30.9 157.35 ;
        RECT  27.3 145.35 28.2 153.75 ;
        RECT  29.1 148.65 30.3 149.85 ;
        RECT  26.85 148.8 27.75 149.7 ;
        RECT  23.1 156.45 32.7 157.35 ;
        RECT  23.1 142.35 32.7 143.25 ;
        RECT  29.7 151.35 30.9 152.55 ;
        RECT  27.3 151.35 28.5 152.55 ;
        RECT  29.7 151.35 30.9 152.55 ;
        RECT  27.3 151.35 28.5 152.55 ;
        RECT  29.7 142.95 30.9 144.15 ;
        RECT  27.3 142.95 28.5 144.15 ;
        RECT  29.7 142.95 30.9 144.15 ;
        RECT  27.3 142.95 28.5 144.15 ;
        RECT  24.9 142.95 26.1 144.15 ;
        RECT  24.9 153.15 26.1 154.35 ;
        RECT  29.1 147.45 30.3 148.65 ;
        RECT  36.9 84.45 38.1 86.4 ;
        RECT  36.9 72.3 38.1 74.25 ;
        RECT  44.1 84.45 45.3 86.85 ;
        RECT  44.1 71.85 45.3 75.45 ;
        RECT  39.3 71.85 40.5 75.45 ;
        RECT  43.5 78.0 44.7 79.2 ;
        RECT  39.3 78.0 40.5 79.2 ;
        RECT  40.5 80.7 41.7 81.9 ;
        RECT  32.7 71.85 47.1 72.75 ;
        RECT  32.7 85.95 47.1 86.85 ;
        RECT  44.1 74.25 45.3 75.45 ;
        RECT  41.7 74.25 42.9 75.45 ;
        RECT  44.1 74.25 45.3 75.45 ;
        RECT  41.7 74.25 42.9 75.45 ;
        RECT  41.7 74.25 42.9 75.45 ;
        RECT  39.3 74.25 40.5 75.45 ;
        RECT  41.7 74.25 42.9 75.45 ;
        RECT  39.3 74.25 40.5 75.45 ;
        RECT  44.1 83.25 45.3 84.45 ;
        RECT  41.7 83.25 42.9 84.45 ;
        RECT  44.1 83.25 45.3 84.45 ;
        RECT  41.7 83.25 42.9 84.45 ;
        RECT  41.7 83.25 42.9 84.45 ;
        RECT  39.3 83.25 40.5 84.45 ;
        RECT  41.7 83.25 42.9 84.45 ;
        RECT  39.3 83.25 40.5 84.45 ;
        RECT  36.9 83.85 38.1 85.05 ;
        RECT  36.9 73.65 38.1 74.85 ;
        RECT  40.5 80.7 41.7 81.9 ;
        RECT  43.5 78.0 44.7 79.2 ;
        RECT  41.7 74.25 42.9 75.45 ;
        RECT  39.3 83.25 40.5 84.45 ;
        RECT  39.3 78.0 40.5 79.2 ;
        RECT  36.9 114.6 38.1 116.55 ;
        RECT  36.9 126.75 38.1 128.7 ;
        RECT  44.1 114.15 45.3 116.55 ;
        RECT  44.1 125.55 45.3 129.15 ;
        RECT  39.3 125.55 40.5 129.15 ;
        RECT  43.5 121.8 44.7 123.0 ;
        RECT  39.3 121.8 40.5 123.0 ;
        RECT  40.5 119.1 41.7 120.3 ;
        RECT  32.7 128.25 47.1 129.15 ;
        RECT  32.7 114.15 47.1 115.05 ;
        RECT  44.1 123.15 45.3 124.35 ;
        RECT  41.7 123.15 42.9 124.35 ;
        RECT  44.1 123.15 45.3 124.35 ;
        RECT  41.7 123.15 42.9 124.35 ;
        RECT  41.7 123.15 42.9 124.35 ;
        RECT  39.3 123.15 40.5 124.35 ;
        RECT  41.7 123.15 42.9 124.35 ;
        RECT  39.3 123.15 40.5 124.35 ;
        RECT  44.1 114.15 45.3 115.35 ;
        RECT  41.7 114.15 42.9 115.35 ;
        RECT  44.1 114.15 45.3 115.35 ;
        RECT  41.7 114.15 42.9 115.35 ;
        RECT  41.7 114.15 42.9 115.35 ;
        RECT  39.3 114.15 40.5 115.35 ;
        RECT  41.7 114.15 42.9 115.35 ;
        RECT  39.3 114.15 40.5 115.35 ;
        RECT  36.9 114.75 38.1 115.95 ;
        RECT  36.9 124.95 38.1 126.15 ;
        RECT  40.5 117.9 41.7 119.1 ;
        RECT  43.5 120.6 44.7 121.8 ;
        RECT  41.7 124.35 42.9 125.55 ;
        RECT  39.3 115.35 40.5 116.55 ;
        RECT  39.3 120.6 40.5 121.8 ;
        RECT  36.9 112.65 38.1 114.6 ;
        RECT  36.9 100.5 38.1 102.45 ;
        RECT  44.1 112.65 45.3 115.05 ;
        RECT  44.1 100.05 45.3 103.65 ;
        RECT  39.3 100.05 40.5 103.65 ;
        RECT  43.5 106.2 44.7 107.4 ;
        RECT  39.3 106.2 40.5 107.4 ;
        RECT  40.5 108.9 41.7 110.1 ;
        RECT  32.7 100.05 47.1 100.95 ;
        RECT  32.7 114.15 47.1 115.05 ;
        RECT  44.1 102.45 45.3 103.65 ;
        RECT  41.7 102.45 42.9 103.65 ;
        RECT  44.1 102.45 45.3 103.65 ;
        RECT  41.7 102.45 42.9 103.65 ;
        RECT  41.7 102.45 42.9 103.65 ;
        RECT  39.3 102.45 40.5 103.65 ;
        RECT  41.7 102.45 42.9 103.65 ;
        RECT  39.3 102.45 40.5 103.65 ;
        RECT  44.1 111.45 45.3 112.65 ;
        RECT  41.7 111.45 42.9 112.65 ;
        RECT  44.1 111.45 45.3 112.65 ;
        RECT  41.7 111.45 42.9 112.65 ;
        RECT  41.7 111.45 42.9 112.65 ;
        RECT  39.3 111.45 40.5 112.65 ;
        RECT  41.7 111.45 42.9 112.65 ;
        RECT  39.3 111.45 40.5 112.65 ;
        RECT  36.9 112.05 38.1 113.25 ;
        RECT  36.9 101.85 38.1 103.05 ;
        RECT  40.5 108.9 41.7 110.1 ;
        RECT  43.5 106.2 44.7 107.4 ;
        RECT  41.7 102.45 42.9 103.65 ;
        RECT  39.3 111.45 40.5 112.65 ;
        RECT  39.3 106.2 40.5 107.4 ;
        RECT  36.9 142.8 38.1 144.75 ;
        RECT  36.9 154.95 38.1 156.9 ;
        RECT  44.1 142.35 45.3 144.75 ;
        RECT  44.1 153.75 45.3 157.35 ;
        RECT  39.3 153.75 40.5 157.35 ;
        RECT  43.5 150.0 44.7 151.2 ;
        RECT  39.3 150.0 40.5 151.2 ;
        RECT  40.5 147.3 41.7 148.5 ;
        RECT  32.7 156.45 47.1 157.35 ;
        RECT  32.7 142.35 47.1 143.25 ;
        RECT  44.1 151.35 45.3 152.55 ;
        RECT  41.7 151.35 42.9 152.55 ;
        RECT  44.1 151.35 45.3 152.55 ;
        RECT  41.7 151.35 42.9 152.55 ;
        RECT  41.7 151.35 42.9 152.55 ;
        RECT  39.3 151.35 40.5 152.55 ;
        RECT  41.7 151.35 42.9 152.55 ;
        RECT  39.3 151.35 40.5 152.55 ;
        RECT  44.1 142.35 45.3 143.55 ;
        RECT  41.7 142.35 42.9 143.55 ;
        RECT  44.1 142.35 45.3 143.55 ;
        RECT  41.7 142.35 42.9 143.55 ;
        RECT  41.7 142.35 42.9 143.55 ;
        RECT  39.3 142.35 40.5 143.55 ;
        RECT  41.7 142.35 42.9 143.55 ;
        RECT  39.3 142.35 40.5 143.55 ;
        RECT  36.9 142.95 38.1 144.15 ;
        RECT  36.9 153.15 38.1 154.35 ;
        RECT  40.5 146.1 41.7 147.3 ;
        RECT  43.5 148.8 44.7 150.0 ;
        RECT  41.7 152.55 42.9 153.75 ;
        RECT  39.3 143.55 40.5 144.75 ;
        RECT  39.3 148.8 40.5 150.0 ;
        RECT  58.05 96.0 59.25 97.2 ;
        RECT  76.65 91.05 77.85 92.25 ;
        RECT  55.05 110.1 56.25 111.3 ;
        RECT  73.65 106.35 74.85 107.55 ;
        RECT  76.65 114.9 77.85 116.1 ;
        RECT  52.05 114.9 53.25 116.1 ;
        RECT  73.65 129.0 74.85 130.2 ;
        RECT  49.05 129.0 50.25 130.2 ;
        RECT  58.05 92.4 59.25 93.6 ;
        RECT  55.05 89.7 56.25 90.9 ;
        RECT  52.05 105.0 53.25 106.2 ;
        RECT  55.05 107.7 56.25 108.9 ;
        RECT  58.05 120.6 59.25 121.8 ;
        RECT  49.05 117.9 50.25 119.1 ;
        RECT  52.05 133.2 53.25 134.4 ;
        RECT  49.05 135.9 50.25 137.1 ;
        RECT  60.75 148.8 61.65 149.7 ;
        RECT  60.75 153.75 61.65 154.65 ;
        RECT  61.2 148.8 65.85 149.7 ;
        RECT  60.75 149.25 61.65 154.2 ;
        RECT  58.65 153.75 61.2 154.65 ;
        RECT  69.3 148.8 77.25 149.7 ;
        RECT  60.75 164.1 61.65 165.0 ;
        RECT  60.75 167.85 61.65 168.75 ;
        RECT  61.2 164.1 65.85 165.0 ;
        RECT  60.75 164.55 61.65 168.3 ;
        RECT  55.65 167.85 61.2 168.75 ;
        RECT  69.3 164.1 74.25 165.0 ;
        RECT  52.65 172.65 77.25 173.55 ;
        RECT  49.65 186.75 74.25 187.65 ;
        RECT  44.7 150.15 58.65 151.05 ;
        RECT  41.7 147.45 55.65 148.35 ;
        RECT  44.7 162.75 52.65 163.65 ;
        RECT  41.7 165.45 55.65 166.35 ;
        RECT  44.7 178.35 58.65 179.25 ;
        RECT  41.7 175.65 49.65 176.55 ;
        RECT  44.7 190.95 52.65 191.85 ;
        RECT  41.7 193.65 49.65 194.55 ;
        RECT  34.35 150.15 35.25 151.05 ;
        RECT  34.35 148.8 35.25 149.7 ;
        RECT  34.8 150.15 39.3 151.05 ;
        RECT  34.35 149.25 35.25 150.6 ;
        RECT  30.3 148.8 34.8 149.7 ;
        RECT  34.35 162.75 35.25 163.65 ;
        RECT  34.35 164.1 35.25 165.0 ;
        RECT  34.8 162.75 39.3 163.65 ;
        RECT  34.35 163.2 35.25 164.55 ;
        RECT  30.3 164.1 34.8 165.0 ;
        RECT  34.35 178.35 35.25 179.25 ;
        RECT  34.35 177.0 35.25 177.9 ;
        RECT  34.8 178.35 39.3 179.25 ;
        RECT  34.35 177.45 35.25 178.8 ;
        RECT  30.3 177.0 34.8 177.9 ;
        RECT  34.35 190.95 35.25 191.85 ;
        RECT  34.35 192.3 35.25 193.2 ;
        RECT  34.8 190.95 39.3 191.85 ;
        RECT  34.35 191.4 35.25 192.75 ;
        RECT  30.3 192.3 34.8 193.2 ;
        RECT  23.1 192.3 26.85 193.2 ;
        RECT  23.1 177.0 26.85 177.9 ;
        RECT  23.1 148.8 26.85 149.7 ;
        RECT  23.1 164.1 26.85 165.0 ;
        RECT  23.1 156.45 77.7 157.35 ;
        RECT  23.1 184.65 77.7 185.55 ;
        RECT  23.1 142.35 77.7 143.25 ;
        RECT  23.1 170.55 77.7 171.45 ;
        RECT  23.1 198.75 77.7 199.65 ;
        RECT  63.9 140.85 65.1 142.8 ;
        RECT  63.9 128.7 65.1 130.65 ;
        RECT  68.7 141.45 69.9 143.25 ;
        RECT  68.7 128.25 69.9 131.85 ;
        RECT  66.3 131.85 67.2 140.25 ;
        RECT  68.1 135.75 69.3 136.95 ;
        RECT  65.85 135.9 66.75 136.8 ;
        RECT  62.1 128.25 71.7 129.15 ;
        RECT  62.1 142.35 71.7 143.25 ;
        RECT  68.7 130.65 69.9 131.85 ;
        RECT  66.3 130.65 67.5 131.85 ;
        RECT  68.7 130.65 69.9 131.85 ;
        RECT  66.3 130.65 67.5 131.85 ;
        RECT  68.7 140.25 69.9 141.45 ;
        RECT  66.3 140.25 67.5 141.45 ;
        RECT  68.7 140.25 69.9 141.45 ;
        RECT  66.3 140.25 67.5 141.45 ;
        RECT  63.9 140.25 65.1 141.45 ;
        RECT  63.9 130.05 65.1 131.25 ;
        RECT  68.1 135.75 69.3 136.95 ;
        RECT  63.9 171.0 65.1 172.95 ;
        RECT  63.9 183.15 65.1 185.1 ;
        RECT  68.7 170.55 69.9 172.35 ;
        RECT  68.7 181.95 69.9 185.55 ;
        RECT  66.3 173.55 67.2 181.95 ;
        RECT  68.1 176.85 69.3 178.05 ;
        RECT  65.85 177.0 66.75 177.9 ;
        RECT  62.1 184.65 71.7 185.55 ;
        RECT  62.1 170.55 71.7 171.45 ;
        RECT  68.7 179.55 69.9 180.75 ;
        RECT  66.3 179.55 67.5 180.75 ;
        RECT  68.7 179.55 69.9 180.75 ;
        RECT  66.3 179.55 67.5 180.75 ;
        RECT  68.7 171.15 69.9 172.35 ;
        RECT  66.3 171.15 67.5 172.35 ;
        RECT  68.7 171.15 69.9 172.35 ;
        RECT  66.3 171.15 67.5 172.35 ;
        RECT  63.9 171.15 65.1 172.35 ;
        RECT  63.9 181.35 65.1 182.55 ;
        RECT  68.1 175.65 69.3 176.85 ;
        RECT  24.9 140.85 26.1 142.8 ;
        RECT  24.9 128.7 26.1 130.65 ;
        RECT  29.7 141.45 30.9 143.25 ;
        RECT  29.7 128.25 30.9 131.85 ;
        RECT  27.3 131.85 28.2 140.25 ;
        RECT  29.1 135.75 30.3 136.95 ;
        RECT  26.85 135.9 27.75 136.8 ;
        RECT  23.1 128.25 32.7 129.15 ;
        RECT  23.1 142.35 32.7 143.25 ;
        RECT  29.7 130.65 30.9 131.85 ;
        RECT  27.3 130.65 28.5 131.85 ;
        RECT  29.7 130.65 30.9 131.85 ;
        RECT  27.3 130.65 28.5 131.85 ;
        RECT  29.7 140.25 30.9 141.45 ;
        RECT  27.3 140.25 28.5 141.45 ;
        RECT  29.7 140.25 30.9 141.45 ;
        RECT  27.3 140.25 28.5 141.45 ;
        RECT  24.9 140.25 26.1 141.45 ;
        RECT  24.9 130.05 26.1 131.25 ;
        RECT  29.1 135.75 30.3 136.95 ;
        RECT  24.9 171.0 26.1 172.95 ;
        RECT  24.9 183.15 26.1 185.1 ;
        RECT  29.7 170.55 30.9 172.35 ;
        RECT  29.7 181.95 30.9 185.55 ;
        RECT  27.3 173.55 28.2 181.95 ;
        RECT  29.1 176.85 30.3 178.05 ;
        RECT  26.85 177.0 27.75 177.9 ;
        RECT  23.1 184.65 32.7 185.55 ;
        RECT  23.1 170.55 32.7 171.45 ;
        RECT  29.7 179.55 30.9 180.75 ;
        RECT  27.3 179.55 28.5 180.75 ;
        RECT  29.7 179.55 30.9 180.75 ;
        RECT  27.3 179.55 28.5 180.75 ;
        RECT  29.7 171.15 30.9 172.35 ;
        RECT  27.3 171.15 28.5 172.35 ;
        RECT  29.7 171.15 30.9 172.35 ;
        RECT  27.3 171.15 28.5 172.35 ;
        RECT  24.9 171.15 26.1 172.35 ;
        RECT  24.9 181.35 26.1 182.55 ;
        RECT  29.1 175.65 30.3 176.85 ;
        RECT  24.9 169.05 26.1 171.0 ;
        RECT  24.9 156.9 26.1 158.85 ;
        RECT  29.7 169.65 30.9 171.45 ;
        RECT  29.7 156.45 30.9 160.05 ;
        RECT  27.3 160.05 28.2 168.45 ;
        RECT  29.1 163.95 30.3 165.15 ;
        RECT  26.85 164.1 27.75 165.0 ;
        RECT  23.1 156.45 32.7 157.35 ;
        RECT  23.1 170.55 32.7 171.45 ;
        RECT  29.7 158.85 30.9 160.05 ;
        RECT  27.3 158.85 28.5 160.05 ;
        RECT  29.7 158.85 30.9 160.05 ;
        RECT  27.3 158.85 28.5 160.05 ;
        RECT  29.7 168.45 30.9 169.65 ;
        RECT  27.3 168.45 28.5 169.65 ;
        RECT  29.7 168.45 30.9 169.65 ;
        RECT  27.3 168.45 28.5 169.65 ;
        RECT  24.9 168.45 26.1 169.65 ;
        RECT  24.9 158.25 26.1 159.45 ;
        RECT  29.1 163.95 30.3 165.15 ;
        RECT  24.9 199.2 26.1 201.15 ;
        RECT  24.9 211.35 26.1 213.3 ;
        RECT  29.7 198.75 30.9 200.55 ;
        RECT  29.7 210.15 30.9 213.75 ;
        RECT  27.3 201.75 28.2 210.15 ;
        RECT  29.1 205.05 30.3 206.25 ;
        RECT  26.85 205.2 27.75 206.1 ;
        RECT  23.1 212.85 32.7 213.75 ;
        RECT  23.1 198.75 32.7 199.65 ;
        RECT  29.7 207.75 30.9 208.95 ;
        RECT  27.3 207.75 28.5 208.95 ;
        RECT  29.7 207.75 30.9 208.95 ;
        RECT  27.3 207.75 28.5 208.95 ;
        RECT  29.7 199.35 30.9 200.55 ;
        RECT  27.3 199.35 28.5 200.55 ;
        RECT  29.7 199.35 30.9 200.55 ;
        RECT  27.3 199.35 28.5 200.55 ;
        RECT  24.9 199.35 26.1 200.55 ;
        RECT  24.9 209.55 26.1 210.75 ;
        RECT  29.1 203.85 30.3 205.05 ;
        RECT  36.9 140.85 38.1 142.8 ;
        RECT  36.9 128.7 38.1 130.65 ;
        RECT  44.1 140.85 45.3 143.25 ;
        RECT  44.1 128.25 45.3 131.85 ;
        RECT  39.3 128.25 40.5 131.85 ;
        RECT  43.5 134.4 44.7 135.6 ;
        RECT  39.3 134.4 40.5 135.6 ;
        RECT  40.5 137.1 41.7 138.3 ;
        RECT  32.7 128.25 47.1 129.15 ;
        RECT  32.7 142.35 47.1 143.25 ;
        RECT  44.1 130.65 45.3 131.85 ;
        RECT  41.7 130.65 42.9 131.85 ;
        RECT  44.1 130.65 45.3 131.85 ;
        RECT  41.7 130.65 42.9 131.85 ;
        RECT  41.7 130.65 42.9 131.85 ;
        RECT  39.3 130.65 40.5 131.85 ;
        RECT  41.7 130.65 42.9 131.85 ;
        RECT  39.3 130.65 40.5 131.85 ;
        RECT  44.1 139.65 45.3 140.85 ;
        RECT  41.7 139.65 42.9 140.85 ;
        RECT  44.1 139.65 45.3 140.85 ;
        RECT  41.7 139.65 42.9 140.85 ;
        RECT  41.7 139.65 42.9 140.85 ;
        RECT  39.3 139.65 40.5 140.85 ;
        RECT  41.7 139.65 42.9 140.85 ;
        RECT  39.3 139.65 40.5 140.85 ;
        RECT  36.9 140.25 38.1 141.45 ;
        RECT  36.9 130.05 38.1 131.25 ;
        RECT  40.5 137.1 41.7 138.3 ;
        RECT  43.5 134.4 44.7 135.6 ;
        RECT  41.7 130.65 42.9 131.85 ;
        RECT  39.3 139.65 40.5 140.85 ;
        RECT  39.3 134.4 40.5 135.6 ;
        RECT  36.9 171.0 38.1 172.95 ;
        RECT  36.9 183.15 38.1 185.1 ;
        RECT  44.1 170.55 45.3 172.95 ;
        RECT  44.1 181.95 45.3 185.55 ;
        RECT  39.3 181.95 40.5 185.55 ;
        RECT  43.5 178.2 44.7 179.4 ;
        RECT  39.3 178.2 40.5 179.4 ;
        RECT  40.5 175.5 41.7 176.7 ;
        RECT  32.7 184.65 47.1 185.55 ;
        RECT  32.7 170.55 47.1 171.45 ;
        RECT  44.1 179.55 45.3 180.75 ;
        RECT  41.7 179.55 42.9 180.75 ;
        RECT  44.1 179.55 45.3 180.75 ;
        RECT  41.7 179.55 42.9 180.75 ;
        RECT  41.7 179.55 42.9 180.75 ;
        RECT  39.3 179.55 40.5 180.75 ;
        RECT  41.7 179.55 42.9 180.75 ;
        RECT  39.3 179.55 40.5 180.75 ;
        RECT  44.1 170.55 45.3 171.75 ;
        RECT  41.7 170.55 42.9 171.75 ;
        RECT  44.1 170.55 45.3 171.75 ;
        RECT  41.7 170.55 42.9 171.75 ;
        RECT  41.7 170.55 42.9 171.75 ;
        RECT  39.3 170.55 40.5 171.75 ;
        RECT  41.7 170.55 42.9 171.75 ;
        RECT  39.3 170.55 40.5 171.75 ;
        RECT  36.9 171.15 38.1 172.35 ;
        RECT  36.9 181.35 38.1 182.55 ;
        RECT  40.5 174.3 41.7 175.5 ;
        RECT  43.5 177.0 44.7 178.2 ;
        RECT  41.7 180.75 42.9 181.95 ;
        RECT  39.3 171.75 40.5 172.95 ;
        RECT  39.3 177.0 40.5 178.2 ;
        RECT  36.9 169.05 38.1 171.0 ;
        RECT  36.9 156.9 38.1 158.85 ;
        RECT  44.1 169.05 45.3 171.45 ;
        RECT  44.1 156.45 45.3 160.05 ;
        RECT  39.3 156.45 40.5 160.05 ;
        RECT  43.5 162.6 44.7 163.8 ;
        RECT  39.3 162.6 40.5 163.8 ;
        RECT  40.5 165.3 41.7 166.5 ;
        RECT  32.7 156.45 47.1 157.35 ;
        RECT  32.7 170.55 47.1 171.45 ;
        RECT  44.1 158.85 45.3 160.05 ;
        RECT  41.7 158.85 42.9 160.05 ;
        RECT  44.1 158.85 45.3 160.05 ;
        RECT  41.7 158.85 42.9 160.05 ;
        RECT  41.7 158.85 42.9 160.05 ;
        RECT  39.3 158.85 40.5 160.05 ;
        RECT  41.7 158.85 42.9 160.05 ;
        RECT  39.3 158.85 40.5 160.05 ;
        RECT  44.1 167.85 45.3 169.05 ;
        RECT  41.7 167.85 42.9 169.05 ;
        RECT  44.1 167.85 45.3 169.05 ;
        RECT  41.7 167.85 42.9 169.05 ;
        RECT  41.7 167.85 42.9 169.05 ;
        RECT  39.3 167.85 40.5 169.05 ;
        RECT  41.7 167.85 42.9 169.05 ;
        RECT  39.3 167.85 40.5 169.05 ;
        RECT  36.9 168.45 38.1 169.65 ;
        RECT  36.9 158.25 38.1 159.45 ;
        RECT  40.5 165.3 41.7 166.5 ;
        RECT  43.5 162.6 44.7 163.8 ;
        RECT  41.7 158.85 42.9 160.05 ;
        RECT  39.3 167.85 40.5 169.05 ;
        RECT  39.3 162.6 40.5 163.8 ;
        RECT  36.9 199.2 38.1 201.15 ;
        RECT  36.9 211.35 38.1 213.3 ;
        RECT  44.1 198.75 45.3 201.15 ;
        RECT  44.1 210.15 45.3 213.75 ;
        RECT  39.3 210.15 40.5 213.75 ;
        RECT  43.5 206.4 44.7 207.6 ;
        RECT  39.3 206.4 40.5 207.6 ;
        RECT  40.5 203.7 41.7 204.9 ;
        RECT  32.7 212.85 47.1 213.75 ;
        RECT  32.7 198.75 47.1 199.65 ;
        RECT  44.1 207.75 45.3 208.95 ;
        RECT  41.7 207.75 42.9 208.95 ;
        RECT  44.1 207.75 45.3 208.95 ;
        RECT  41.7 207.75 42.9 208.95 ;
        RECT  41.7 207.75 42.9 208.95 ;
        RECT  39.3 207.75 40.5 208.95 ;
        RECT  41.7 207.75 42.9 208.95 ;
        RECT  39.3 207.75 40.5 208.95 ;
        RECT  44.1 198.75 45.3 199.95 ;
        RECT  41.7 198.75 42.9 199.95 ;
        RECT  44.1 198.75 45.3 199.95 ;
        RECT  41.7 198.75 42.9 199.95 ;
        RECT  41.7 198.75 42.9 199.95 ;
        RECT  39.3 198.75 40.5 199.95 ;
        RECT  41.7 198.75 42.9 199.95 ;
        RECT  39.3 198.75 40.5 199.95 ;
        RECT  36.9 199.35 38.1 200.55 ;
        RECT  36.9 209.55 38.1 210.75 ;
        RECT  40.5 202.5 41.7 203.7 ;
        RECT  43.5 205.2 44.7 206.4 ;
        RECT  41.7 208.95 42.9 210.15 ;
        RECT  39.3 199.95 40.5 201.15 ;
        RECT  39.3 205.2 40.5 206.4 ;
        RECT  58.05 152.4 59.25 153.6 ;
        RECT  76.65 147.45 77.85 148.65 ;
        RECT  55.05 166.5 56.25 167.7 ;
        RECT  73.65 162.75 74.85 163.95 ;
        RECT  76.65 171.3 77.85 172.5 ;
        RECT  52.05 171.3 53.25 172.5 ;
        RECT  73.65 185.4 74.85 186.6 ;
        RECT  49.05 185.4 50.25 186.6 ;
        RECT  58.05 148.8 59.25 150.0 ;
        RECT  55.05 146.1 56.25 147.3 ;
        RECT  52.05 161.4 53.25 162.6 ;
        RECT  55.05 164.1 56.25 165.3 ;
        RECT  58.05 177.0 59.25 178.2 ;
        RECT  49.05 174.3 50.25 175.5 ;
        RECT  52.05 189.6 53.25 190.8 ;
        RECT  49.05 192.3 50.25 193.5 ;
        RECT  32.1 199.2 33.3 201.15 ;
        RECT  32.1 211.35 33.3 213.3 ;
        RECT  24.9 198.75 26.1 201.15 ;
        RECT  24.9 210.15 26.1 213.75 ;
        RECT  29.7 210.15 30.9 213.75 ;
        RECT  25.5 206.4 26.7 207.6 ;
        RECT  29.7 206.4 30.9 207.6 ;
        RECT  28.5 203.7 29.7 204.9 ;
        RECT  23.1 212.85 37.5 213.75 ;
        RECT  23.1 198.75 37.5 199.65 ;
        RECT  24.9 210.15 26.1 211.35 ;
        RECT  27.3 210.15 28.5 211.35 ;
        RECT  24.9 210.15 26.1 211.35 ;
        RECT  27.3 210.15 28.5 211.35 ;
        RECT  27.3 210.15 28.5 211.35 ;
        RECT  29.7 210.15 30.9 211.35 ;
        RECT  27.3 210.15 28.5 211.35 ;
        RECT  29.7 210.15 30.9 211.35 ;
        RECT  24.9 201.15 26.1 202.35 ;
        RECT  27.3 201.15 28.5 202.35 ;
        RECT  24.9 201.15 26.1 202.35 ;
        RECT  27.3 201.15 28.5 202.35 ;
        RECT  27.3 201.15 28.5 202.35 ;
        RECT  29.7 201.15 30.9 202.35 ;
        RECT  27.3 201.15 28.5 202.35 ;
        RECT  29.7 201.15 30.9 202.35 ;
        RECT  32.1 200.55 33.3 201.75 ;
        RECT  32.1 210.75 33.3 211.95 ;
        RECT  28.5 203.7 29.7 204.9 ;
        RECT  25.5 206.4 26.7 207.6 ;
        RECT  27.3 210.15 28.5 211.35 ;
        RECT  29.7 201.15 30.9 202.35 ;
        RECT  29.7 206.4 30.9 207.6 ;
        RECT  32.1 225.45 33.3 227.4 ;
        RECT  32.1 213.3 33.3 215.25 ;
        RECT  24.9 225.45 26.1 227.85 ;
        RECT  24.9 212.85 26.1 216.45 ;
        RECT  29.7 212.85 30.9 216.45 ;
        RECT  25.5 219.0 26.7 220.2 ;
        RECT  29.7 219.0 30.9 220.2 ;
        RECT  28.5 221.7 29.7 222.9 ;
        RECT  23.1 212.85 37.5 213.75 ;
        RECT  23.1 226.95 37.5 227.85 ;
        RECT  24.9 217.65 26.1 218.85 ;
        RECT  27.3 217.65 28.5 218.85 ;
        RECT  24.9 217.65 26.1 218.85 ;
        RECT  27.3 217.65 28.5 218.85 ;
        RECT  27.3 217.65 28.5 218.85 ;
        RECT  29.7 217.65 30.9 218.85 ;
        RECT  27.3 217.65 28.5 218.85 ;
        RECT  29.7 217.65 30.9 218.85 ;
        RECT  24.9 226.65 26.1 227.85 ;
        RECT  27.3 226.65 28.5 227.85 ;
        RECT  24.9 226.65 26.1 227.85 ;
        RECT  27.3 226.65 28.5 227.85 ;
        RECT  27.3 226.65 28.5 227.85 ;
        RECT  29.7 226.65 30.9 227.85 ;
        RECT  27.3 226.65 28.5 227.85 ;
        RECT  29.7 226.65 30.9 227.85 ;
        RECT  32.1 226.05 33.3 227.25 ;
        RECT  32.1 215.85 33.3 217.05 ;
        RECT  28.5 222.9 29.7 224.1 ;
        RECT  25.5 220.2 26.7 221.4 ;
        RECT  27.3 216.45 28.5 217.65 ;
        RECT  29.7 225.45 30.9 226.65 ;
        RECT  29.7 220.2 30.9 221.4 ;
        RECT  32.1 227.4 33.3 229.35 ;
        RECT  32.1 239.55 33.3 241.5 ;
        RECT  24.9 226.95 26.1 229.35 ;
        RECT  24.9 238.35 26.1 241.95 ;
        RECT  29.7 238.35 30.9 241.95 ;
        RECT  25.5 234.6 26.7 235.8 ;
        RECT  29.7 234.6 30.9 235.8 ;
        RECT  28.5 231.9 29.7 233.1 ;
        RECT  23.1 241.05 37.5 241.95 ;
        RECT  23.1 226.95 37.5 227.85 ;
        RECT  24.9 238.35 26.1 239.55 ;
        RECT  27.3 238.35 28.5 239.55 ;
        RECT  24.9 238.35 26.1 239.55 ;
        RECT  27.3 238.35 28.5 239.55 ;
        RECT  27.3 238.35 28.5 239.55 ;
        RECT  29.7 238.35 30.9 239.55 ;
        RECT  27.3 238.35 28.5 239.55 ;
        RECT  29.7 238.35 30.9 239.55 ;
        RECT  24.9 229.35 26.1 230.55 ;
        RECT  27.3 229.35 28.5 230.55 ;
        RECT  24.9 229.35 26.1 230.55 ;
        RECT  27.3 229.35 28.5 230.55 ;
        RECT  27.3 229.35 28.5 230.55 ;
        RECT  29.7 229.35 30.9 230.55 ;
        RECT  27.3 229.35 28.5 230.55 ;
        RECT  29.7 229.35 30.9 230.55 ;
        RECT  32.1 228.75 33.3 229.95 ;
        RECT  32.1 238.95 33.3 240.15 ;
        RECT  28.5 231.9 29.7 233.1 ;
        RECT  25.5 234.6 26.7 235.8 ;
        RECT  27.3 238.35 28.5 239.55 ;
        RECT  29.7 229.35 30.9 230.55 ;
        RECT  29.7 234.6 30.9 235.8 ;
        RECT  32.1 253.65 33.3 255.6 ;
        RECT  32.1 241.5 33.3 243.45 ;
        RECT  24.9 253.65 26.1 256.05 ;
        RECT  24.9 241.05 26.1 244.65 ;
        RECT  29.7 241.05 30.9 244.65 ;
        RECT  25.5 247.2 26.7 248.4 ;
        RECT  29.7 247.2 30.9 248.4 ;
        RECT  28.5 249.9 29.7 251.1 ;
        RECT  23.1 241.05 37.5 241.95 ;
        RECT  23.1 255.15 37.5 256.05 ;
        RECT  24.9 245.85 26.1 247.05 ;
        RECT  27.3 245.85 28.5 247.05 ;
        RECT  24.9 245.85 26.1 247.05 ;
        RECT  27.3 245.85 28.5 247.05 ;
        RECT  27.3 245.85 28.5 247.05 ;
        RECT  29.7 245.85 30.9 247.05 ;
        RECT  27.3 245.85 28.5 247.05 ;
        RECT  29.7 245.85 30.9 247.05 ;
        RECT  24.9 254.85 26.1 256.05 ;
        RECT  27.3 254.85 28.5 256.05 ;
        RECT  24.9 254.85 26.1 256.05 ;
        RECT  27.3 254.85 28.5 256.05 ;
        RECT  27.3 254.85 28.5 256.05 ;
        RECT  29.7 254.85 30.9 256.05 ;
        RECT  27.3 254.85 28.5 256.05 ;
        RECT  29.7 254.85 30.9 256.05 ;
        RECT  32.1 254.25 33.3 255.45 ;
        RECT  32.1 244.05 33.3 245.25 ;
        RECT  28.5 251.1 29.7 252.3 ;
        RECT  25.5 248.4 26.7 249.6 ;
        RECT  27.3 244.65 28.5 245.85 ;
        RECT  29.7 253.65 30.9 254.85 ;
        RECT  29.7 248.4 30.9 249.6 ;
        RECT  32.1 255.6 33.3 257.55 ;
        RECT  32.1 267.75 33.3 269.7 ;
        RECT  24.9 255.15 26.1 257.55 ;
        RECT  24.9 266.55 26.1 270.15 ;
        RECT  29.7 266.55 30.9 270.15 ;
        RECT  25.5 262.8 26.7 264.0 ;
        RECT  29.7 262.8 30.9 264.0 ;
        RECT  28.5 260.1 29.7 261.3 ;
        RECT  23.1 269.25 37.5 270.15 ;
        RECT  23.1 255.15 37.5 256.05 ;
        RECT  24.9 266.55 26.1 267.75 ;
        RECT  27.3 266.55 28.5 267.75 ;
        RECT  24.9 266.55 26.1 267.75 ;
        RECT  27.3 266.55 28.5 267.75 ;
        RECT  27.3 266.55 28.5 267.75 ;
        RECT  29.7 266.55 30.9 267.75 ;
        RECT  27.3 266.55 28.5 267.75 ;
        RECT  29.7 266.55 30.9 267.75 ;
        RECT  24.9 257.55 26.1 258.75 ;
        RECT  27.3 257.55 28.5 258.75 ;
        RECT  24.9 257.55 26.1 258.75 ;
        RECT  27.3 257.55 28.5 258.75 ;
        RECT  27.3 257.55 28.5 258.75 ;
        RECT  29.7 257.55 30.9 258.75 ;
        RECT  27.3 257.55 28.5 258.75 ;
        RECT  29.7 257.55 30.9 258.75 ;
        RECT  32.1 256.95 33.3 258.15 ;
        RECT  32.1 267.15 33.3 268.35 ;
        RECT  28.5 260.1 29.7 261.3 ;
        RECT  25.5 262.8 26.7 264.0 ;
        RECT  27.3 266.55 28.5 267.75 ;
        RECT  29.7 257.55 30.9 258.75 ;
        RECT  29.7 262.8 30.9 264.0 ;
        RECT  32.1 281.85 33.3 283.8 ;
        RECT  32.1 269.7 33.3 271.65 ;
        RECT  24.9 281.85 26.1 284.25 ;
        RECT  24.9 269.25 26.1 272.85 ;
        RECT  29.7 269.25 30.9 272.85 ;
        RECT  25.5 275.4 26.7 276.6 ;
        RECT  29.7 275.4 30.9 276.6 ;
        RECT  28.5 278.1 29.7 279.3 ;
        RECT  23.1 269.25 37.5 270.15 ;
        RECT  23.1 283.35 37.5 284.25 ;
        RECT  24.9 274.05 26.1 275.25 ;
        RECT  27.3 274.05 28.5 275.25 ;
        RECT  24.9 274.05 26.1 275.25 ;
        RECT  27.3 274.05 28.5 275.25 ;
        RECT  27.3 274.05 28.5 275.25 ;
        RECT  29.7 274.05 30.9 275.25 ;
        RECT  27.3 274.05 28.5 275.25 ;
        RECT  29.7 274.05 30.9 275.25 ;
        RECT  24.9 283.05 26.1 284.25 ;
        RECT  27.3 283.05 28.5 284.25 ;
        RECT  24.9 283.05 26.1 284.25 ;
        RECT  27.3 283.05 28.5 284.25 ;
        RECT  27.3 283.05 28.5 284.25 ;
        RECT  29.7 283.05 30.9 284.25 ;
        RECT  27.3 283.05 28.5 284.25 ;
        RECT  29.7 283.05 30.9 284.25 ;
        RECT  32.1 282.45 33.3 283.65 ;
        RECT  32.1 272.25 33.3 273.45 ;
        RECT  28.5 279.3 29.7 280.5 ;
        RECT  25.5 276.6 26.7 277.8 ;
        RECT  27.3 272.85 28.5 274.05 ;
        RECT  29.7 281.85 30.9 283.05 ;
        RECT  29.7 276.6 30.9 277.8 ;
        RECT  32.1 283.8 33.3 285.75 ;
        RECT  32.1 295.95 33.3 297.9 ;
        RECT  24.9 283.35 26.1 285.75 ;
        RECT  24.9 294.75 26.1 298.35 ;
        RECT  29.7 294.75 30.9 298.35 ;
        RECT  25.5 291.0 26.7 292.2 ;
        RECT  29.7 291.0 30.9 292.2 ;
        RECT  28.5 288.3 29.7 289.5 ;
        RECT  23.1 297.45 37.5 298.35 ;
        RECT  23.1 283.35 37.5 284.25 ;
        RECT  24.9 294.75 26.1 295.95 ;
        RECT  27.3 294.75 28.5 295.95 ;
        RECT  24.9 294.75 26.1 295.95 ;
        RECT  27.3 294.75 28.5 295.95 ;
        RECT  27.3 294.75 28.5 295.95 ;
        RECT  29.7 294.75 30.9 295.95 ;
        RECT  27.3 294.75 28.5 295.95 ;
        RECT  29.7 294.75 30.9 295.95 ;
        RECT  24.9 285.75 26.1 286.95 ;
        RECT  27.3 285.75 28.5 286.95 ;
        RECT  24.9 285.75 26.1 286.95 ;
        RECT  27.3 285.75 28.5 286.95 ;
        RECT  27.3 285.75 28.5 286.95 ;
        RECT  29.7 285.75 30.9 286.95 ;
        RECT  27.3 285.75 28.5 286.95 ;
        RECT  29.7 285.75 30.9 286.95 ;
        RECT  32.1 285.15 33.3 286.35 ;
        RECT  32.1 295.35 33.3 296.55 ;
        RECT  28.5 288.3 29.7 289.5 ;
        RECT  25.5 291.0 26.7 292.2 ;
        RECT  27.3 294.75 28.5 295.95 ;
        RECT  29.7 285.75 30.9 286.95 ;
        RECT  29.7 291.0 30.9 292.2 ;
        RECT  32.1 310.05 33.3 312.0 ;
        RECT  32.1 297.9 33.3 299.85 ;
        RECT  24.9 310.05 26.1 312.45 ;
        RECT  24.9 297.45 26.1 301.05 ;
        RECT  29.7 297.45 30.9 301.05 ;
        RECT  25.5 303.6 26.7 304.8 ;
        RECT  29.7 303.6 30.9 304.8 ;
        RECT  28.5 306.3 29.7 307.5 ;
        RECT  23.1 297.45 37.5 298.35 ;
        RECT  23.1 311.55 37.5 312.45 ;
        RECT  24.9 302.25 26.1 303.45 ;
        RECT  27.3 302.25 28.5 303.45 ;
        RECT  24.9 302.25 26.1 303.45 ;
        RECT  27.3 302.25 28.5 303.45 ;
        RECT  27.3 302.25 28.5 303.45 ;
        RECT  29.7 302.25 30.9 303.45 ;
        RECT  27.3 302.25 28.5 303.45 ;
        RECT  29.7 302.25 30.9 303.45 ;
        RECT  24.9 311.25 26.1 312.45 ;
        RECT  27.3 311.25 28.5 312.45 ;
        RECT  24.9 311.25 26.1 312.45 ;
        RECT  27.3 311.25 28.5 312.45 ;
        RECT  27.3 311.25 28.5 312.45 ;
        RECT  29.7 311.25 30.9 312.45 ;
        RECT  27.3 311.25 28.5 312.45 ;
        RECT  29.7 311.25 30.9 312.45 ;
        RECT  32.1 310.65 33.3 311.85 ;
        RECT  32.1 300.45 33.3 301.65 ;
        RECT  28.5 307.5 29.7 308.7 ;
        RECT  25.5 304.8 26.7 306.0 ;
        RECT  27.3 301.05 28.5 302.25 ;
        RECT  29.7 310.05 30.9 311.25 ;
        RECT  29.7 304.8 30.9 306.0 ;
        RECT  32.1 312.0 33.3 313.95 ;
        RECT  32.1 324.15 33.3 326.1 ;
        RECT  24.9 311.55 26.1 313.95 ;
        RECT  24.9 322.95 26.1 326.55 ;
        RECT  29.7 322.95 30.9 326.55 ;
        RECT  25.5 319.2 26.7 320.4 ;
        RECT  29.7 319.2 30.9 320.4 ;
        RECT  28.5 316.5 29.7 317.7 ;
        RECT  23.1 325.65 37.5 326.55 ;
        RECT  23.1 311.55 37.5 312.45 ;
        RECT  24.9 322.95 26.1 324.15 ;
        RECT  27.3 322.95 28.5 324.15 ;
        RECT  24.9 322.95 26.1 324.15 ;
        RECT  27.3 322.95 28.5 324.15 ;
        RECT  27.3 322.95 28.5 324.15 ;
        RECT  29.7 322.95 30.9 324.15 ;
        RECT  27.3 322.95 28.5 324.15 ;
        RECT  29.7 322.95 30.9 324.15 ;
        RECT  24.9 313.95 26.1 315.15 ;
        RECT  27.3 313.95 28.5 315.15 ;
        RECT  24.9 313.95 26.1 315.15 ;
        RECT  27.3 313.95 28.5 315.15 ;
        RECT  27.3 313.95 28.5 315.15 ;
        RECT  29.7 313.95 30.9 315.15 ;
        RECT  27.3 313.95 28.5 315.15 ;
        RECT  29.7 313.95 30.9 315.15 ;
        RECT  32.1 313.35 33.3 314.55 ;
        RECT  32.1 323.55 33.3 324.75 ;
        RECT  28.5 316.5 29.7 317.7 ;
        RECT  25.5 319.2 26.7 320.4 ;
        RECT  27.3 322.95 28.5 324.15 ;
        RECT  29.7 313.95 30.9 315.15 ;
        RECT  29.7 319.2 30.9 320.4 ;
        RECT  32.1 338.25 33.3 340.2 ;
        RECT  32.1 326.1 33.3 328.05 ;
        RECT  24.9 338.25 26.1 340.65 ;
        RECT  24.9 325.65 26.1 329.25 ;
        RECT  29.7 325.65 30.9 329.25 ;
        RECT  25.5 331.8 26.7 333.0 ;
        RECT  29.7 331.8 30.9 333.0 ;
        RECT  28.5 334.5 29.7 335.7 ;
        RECT  23.1 325.65 37.5 326.55 ;
        RECT  23.1 339.75 37.5 340.65 ;
        RECT  24.9 330.45 26.1 331.65 ;
        RECT  27.3 330.45 28.5 331.65 ;
        RECT  24.9 330.45 26.1 331.65 ;
        RECT  27.3 330.45 28.5 331.65 ;
        RECT  27.3 330.45 28.5 331.65 ;
        RECT  29.7 330.45 30.9 331.65 ;
        RECT  27.3 330.45 28.5 331.65 ;
        RECT  29.7 330.45 30.9 331.65 ;
        RECT  24.9 339.45 26.1 340.65 ;
        RECT  27.3 339.45 28.5 340.65 ;
        RECT  24.9 339.45 26.1 340.65 ;
        RECT  27.3 339.45 28.5 340.65 ;
        RECT  27.3 339.45 28.5 340.65 ;
        RECT  29.7 339.45 30.9 340.65 ;
        RECT  27.3 339.45 28.5 340.65 ;
        RECT  29.7 339.45 30.9 340.65 ;
        RECT  32.1 338.85 33.3 340.05 ;
        RECT  32.1 328.65 33.3 329.85 ;
        RECT  28.5 335.7 29.7 336.9 ;
        RECT  25.5 333.0 26.7 334.2 ;
        RECT  27.3 329.25 28.5 330.45 ;
        RECT  29.7 338.25 30.9 339.45 ;
        RECT  29.7 333.0 30.9 334.2 ;
        RECT  32.1 340.2 33.3 342.15 ;
        RECT  32.1 352.35 33.3 354.3 ;
        RECT  24.9 339.75 26.1 342.15 ;
        RECT  24.9 351.15 26.1 354.75 ;
        RECT  29.7 351.15 30.9 354.75 ;
        RECT  25.5 347.4 26.7 348.6 ;
        RECT  29.7 347.4 30.9 348.6 ;
        RECT  28.5 344.7 29.7 345.9 ;
        RECT  23.1 353.85 37.5 354.75 ;
        RECT  23.1 339.75 37.5 340.65 ;
        RECT  24.9 351.15 26.1 352.35 ;
        RECT  27.3 351.15 28.5 352.35 ;
        RECT  24.9 351.15 26.1 352.35 ;
        RECT  27.3 351.15 28.5 352.35 ;
        RECT  27.3 351.15 28.5 352.35 ;
        RECT  29.7 351.15 30.9 352.35 ;
        RECT  27.3 351.15 28.5 352.35 ;
        RECT  29.7 351.15 30.9 352.35 ;
        RECT  24.9 342.15 26.1 343.35 ;
        RECT  27.3 342.15 28.5 343.35 ;
        RECT  24.9 342.15 26.1 343.35 ;
        RECT  27.3 342.15 28.5 343.35 ;
        RECT  27.3 342.15 28.5 343.35 ;
        RECT  29.7 342.15 30.9 343.35 ;
        RECT  27.3 342.15 28.5 343.35 ;
        RECT  29.7 342.15 30.9 343.35 ;
        RECT  32.1 341.55 33.3 342.75 ;
        RECT  32.1 351.75 33.3 352.95 ;
        RECT  28.5 344.7 29.7 345.9 ;
        RECT  25.5 347.4 26.7 348.6 ;
        RECT  27.3 351.15 28.5 352.35 ;
        RECT  29.7 342.15 30.9 343.35 ;
        RECT  29.7 347.4 30.9 348.6 ;
        RECT  32.1 366.45 33.3 368.4 ;
        RECT  32.1 354.3 33.3 356.25 ;
        RECT  24.9 366.45 26.1 368.85 ;
        RECT  24.9 353.85 26.1 357.45 ;
        RECT  29.7 353.85 30.9 357.45 ;
        RECT  25.5 360.0 26.7 361.2 ;
        RECT  29.7 360.0 30.9 361.2 ;
        RECT  28.5 362.7 29.7 363.9 ;
        RECT  23.1 353.85 37.5 354.75 ;
        RECT  23.1 367.95 37.5 368.85 ;
        RECT  24.9 358.65 26.1 359.85 ;
        RECT  27.3 358.65 28.5 359.85 ;
        RECT  24.9 358.65 26.1 359.85 ;
        RECT  27.3 358.65 28.5 359.85 ;
        RECT  27.3 358.65 28.5 359.85 ;
        RECT  29.7 358.65 30.9 359.85 ;
        RECT  27.3 358.65 28.5 359.85 ;
        RECT  29.7 358.65 30.9 359.85 ;
        RECT  24.9 367.65 26.1 368.85 ;
        RECT  27.3 367.65 28.5 368.85 ;
        RECT  24.9 367.65 26.1 368.85 ;
        RECT  27.3 367.65 28.5 368.85 ;
        RECT  27.3 367.65 28.5 368.85 ;
        RECT  29.7 367.65 30.9 368.85 ;
        RECT  27.3 367.65 28.5 368.85 ;
        RECT  29.7 367.65 30.9 368.85 ;
        RECT  32.1 367.05 33.3 368.25 ;
        RECT  32.1 356.85 33.3 358.05 ;
        RECT  28.5 363.9 29.7 365.1 ;
        RECT  25.5 361.2 26.7 362.4 ;
        RECT  27.3 357.45 28.5 358.65 ;
        RECT  29.7 366.45 30.9 367.65 ;
        RECT  29.7 361.2 30.9 362.4 ;
        RECT  32.1 368.4 33.3 370.35 ;
        RECT  32.1 380.55 33.3 382.5 ;
        RECT  24.9 367.95 26.1 370.35 ;
        RECT  24.9 379.35 26.1 382.95 ;
        RECT  29.7 379.35 30.9 382.95 ;
        RECT  25.5 375.6 26.7 376.8 ;
        RECT  29.7 375.6 30.9 376.8 ;
        RECT  28.5 372.9 29.7 374.1 ;
        RECT  23.1 382.05 37.5 382.95 ;
        RECT  23.1 367.95 37.5 368.85 ;
        RECT  24.9 379.35 26.1 380.55 ;
        RECT  27.3 379.35 28.5 380.55 ;
        RECT  24.9 379.35 26.1 380.55 ;
        RECT  27.3 379.35 28.5 380.55 ;
        RECT  27.3 379.35 28.5 380.55 ;
        RECT  29.7 379.35 30.9 380.55 ;
        RECT  27.3 379.35 28.5 380.55 ;
        RECT  29.7 379.35 30.9 380.55 ;
        RECT  24.9 370.35 26.1 371.55 ;
        RECT  27.3 370.35 28.5 371.55 ;
        RECT  24.9 370.35 26.1 371.55 ;
        RECT  27.3 370.35 28.5 371.55 ;
        RECT  27.3 370.35 28.5 371.55 ;
        RECT  29.7 370.35 30.9 371.55 ;
        RECT  27.3 370.35 28.5 371.55 ;
        RECT  29.7 370.35 30.9 371.55 ;
        RECT  32.1 369.75 33.3 370.95 ;
        RECT  32.1 379.95 33.3 381.15 ;
        RECT  28.5 372.9 29.7 374.1 ;
        RECT  25.5 375.6 26.7 376.8 ;
        RECT  27.3 379.35 28.5 380.55 ;
        RECT  29.7 370.35 30.9 371.55 ;
        RECT  29.7 375.6 30.9 376.8 ;
        RECT  32.1 394.65 33.3 396.6 ;
        RECT  32.1 382.5 33.3 384.45 ;
        RECT  24.9 394.65 26.1 397.05 ;
        RECT  24.9 382.05 26.1 385.65 ;
        RECT  29.7 382.05 30.9 385.65 ;
        RECT  25.5 388.2 26.7 389.4 ;
        RECT  29.7 388.2 30.9 389.4 ;
        RECT  28.5 390.9 29.7 392.1 ;
        RECT  23.1 382.05 37.5 382.95 ;
        RECT  23.1 396.15 37.5 397.05 ;
        RECT  24.9 386.85 26.1 388.05 ;
        RECT  27.3 386.85 28.5 388.05 ;
        RECT  24.9 386.85 26.1 388.05 ;
        RECT  27.3 386.85 28.5 388.05 ;
        RECT  27.3 386.85 28.5 388.05 ;
        RECT  29.7 386.85 30.9 388.05 ;
        RECT  27.3 386.85 28.5 388.05 ;
        RECT  29.7 386.85 30.9 388.05 ;
        RECT  24.9 395.85 26.1 397.05 ;
        RECT  27.3 395.85 28.5 397.05 ;
        RECT  24.9 395.85 26.1 397.05 ;
        RECT  27.3 395.85 28.5 397.05 ;
        RECT  27.3 395.85 28.5 397.05 ;
        RECT  29.7 395.85 30.9 397.05 ;
        RECT  27.3 395.85 28.5 397.05 ;
        RECT  29.7 395.85 30.9 397.05 ;
        RECT  32.1 395.25 33.3 396.45 ;
        RECT  32.1 385.05 33.3 386.25 ;
        RECT  28.5 392.1 29.7 393.3 ;
        RECT  25.5 389.4 26.7 390.6 ;
        RECT  27.3 385.65 28.5 386.85 ;
        RECT  29.7 394.65 30.9 395.85 ;
        RECT  29.7 389.4 30.9 390.6 ;
        RECT  32.1 396.6 33.3 398.55 ;
        RECT  32.1 408.75 33.3 410.7 ;
        RECT  24.9 396.15 26.1 398.55 ;
        RECT  24.9 407.55 26.1 411.15 ;
        RECT  29.7 407.55 30.9 411.15 ;
        RECT  25.5 403.8 26.7 405.0 ;
        RECT  29.7 403.8 30.9 405.0 ;
        RECT  28.5 401.1 29.7 402.3 ;
        RECT  23.1 410.25 37.5 411.15 ;
        RECT  23.1 396.15 37.5 397.05 ;
        RECT  24.9 407.55 26.1 408.75 ;
        RECT  27.3 407.55 28.5 408.75 ;
        RECT  24.9 407.55 26.1 408.75 ;
        RECT  27.3 407.55 28.5 408.75 ;
        RECT  27.3 407.55 28.5 408.75 ;
        RECT  29.7 407.55 30.9 408.75 ;
        RECT  27.3 407.55 28.5 408.75 ;
        RECT  29.7 407.55 30.9 408.75 ;
        RECT  24.9 398.55 26.1 399.75 ;
        RECT  27.3 398.55 28.5 399.75 ;
        RECT  24.9 398.55 26.1 399.75 ;
        RECT  27.3 398.55 28.5 399.75 ;
        RECT  27.3 398.55 28.5 399.75 ;
        RECT  29.7 398.55 30.9 399.75 ;
        RECT  27.3 398.55 28.5 399.75 ;
        RECT  29.7 398.55 30.9 399.75 ;
        RECT  32.1 397.95 33.3 399.15 ;
        RECT  32.1 408.15 33.3 409.35 ;
        RECT  28.5 401.1 29.7 402.3 ;
        RECT  25.5 403.8 26.7 405.0 ;
        RECT  27.3 407.55 28.5 408.75 ;
        RECT  29.7 398.55 30.9 399.75 ;
        RECT  29.7 403.8 30.9 405.0 ;
        RECT  32.1 422.85 33.3 424.8 ;
        RECT  32.1 410.7 33.3 412.65 ;
        RECT  24.9 422.85 26.1 425.25 ;
        RECT  24.9 410.25 26.1 413.85 ;
        RECT  29.7 410.25 30.9 413.85 ;
        RECT  25.5 416.4 26.7 417.6 ;
        RECT  29.7 416.4 30.9 417.6 ;
        RECT  28.5 419.1 29.7 420.3 ;
        RECT  23.1 410.25 37.5 411.15 ;
        RECT  23.1 424.35 37.5 425.25 ;
        RECT  24.9 415.05 26.1 416.25 ;
        RECT  27.3 415.05 28.5 416.25 ;
        RECT  24.9 415.05 26.1 416.25 ;
        RECT  27.3 415.05 28.5 416.25 ;
        RECT  27.3 415.05 28.5 416.25 ;
        RECT  29.7 415.05 30.9 416.25 ;
        RECT  27.3 415.05 28.5 416.25 ;
        RECT  29.7 415.05 30.9 416.25 ;
        RECT  24.9 424.05 26.1 425.25 ;
        RECT  27.3 424.05 28.5 425.25 ;
        RECT  24.9 424.05 26.1 425.25 ;
        RECT  27.3 424.05 28.5 425.25 ;
        RECT  27.3 424.05 28.5 425.25 ;
        RECT  29.7 424.05 30.9 425.25 ;
        RECT  27.3 424.05 28.5 425.25 ;
        RECT  29.7 424.05 30.9 425.25 ;
        RECT  32.1 423.45 33.3 424.65 ;
        RECT  32.1 413.25 33.3 414.45 ;
        RECT  28.5 420.3 29.7 421.5 ;
        RECT  25.5 417.6 26.7 418.8 ;
        RECT  27.3 413.85 28.5 415.05 ;
        RECT  29.7 422.85 30.9 424.05 ;
        RECT  29.7 417.6 30.9 418.8 ;
        RECT  44.1 199.2 45.3 201.15 ;
        RECT  44.1 211.35 45.3 213.3 ;
        RECT  39.3 198.75 40.5 200.55 ;
        RECT  39.3 210.15 40.5 213.75 ;
        RECT  42.0 201.75 42.9 210.15 ;
        RECT  39.9 205.05 41.1 206.25 ;
        RECT  42.45 205.2 43.35 206.1 ;
        RECT  37.5 212.85 47.1 213.75 ;
        RECT  37.5 198.75 47.1 199.65 ;
        RECT  39.3 210.15 40.5 211.35 ;
        RECT  41.7 210.15 42.9 211.35 ;
        RECT  39.3 210.15 40.5 211.35 ;
        RECT  41.7 210.15 42.9 211.35 ;
        RECT  39.3 200.55 40.5 201.75 ;
        RECT  41.7 200.55 42.9 201.75 ;
        RECT  39.3 200.55 40.5 201.75 ;
        RECT  41.7 200.55 42.9 201.75 ;
        RECT  44.1 200.55 45.3 201.75 ;
        RECT  44.1 210.75 45.3 211.95 ;
        RECT  39.9 205.05 41.1 206.25 ;
        RECT  44.1 225.45 45.3 227.4 ;
        RECT  44.1 213.3 45.3 215.25 ;
        RECT  39.3 226.05 40.5 227.85 ;
        RECT  39.3 212.85 40.5 216.45 ;
        RECT  42.0 216.45 42.9 224.85 ;
        RECT  39.9 220.35 41.1 221.55 ;
        RECT  42.45 220.5 43.35 221.4 ;
        RECT  37.5 212.85 47.1 213.75 ;
        RECT  37.5 226.95 47.1 227.85 ;
        RECT  39.3 217.65 40.5 218.85 ;
        RECT  41.7 217.65 42.9 218.85 ;
        RECT  39.3 217.65 40.5 218.85 ;
        RECT  41.7 217.65 42.9 218.85 ;
        RECT  39.3 226.05 40.5 227.25 ;
        RECT  41.7 226.05 42.9 227.25 ;
        RECT  39.3 226.05 40.5 227.25 ;
        RECT  41.7 226.05 42.9 227.25 ;
        RECT  44.1 226.05 45.3 227.25 ;
        RECT  44.1 215.85 45.3 217.05 ;
        RECT  39.9 221.55 41.1 222.75 ;
        RECT  44.1 227.4 45.3 229.35 ;
        RECT  44.1 239.55 45.3 241.5 ;
        RECT  39.3 226.95 40.5 228.75 ;
        RECT  39.3 238.35 40.5 241.95 ;
        RECT  42.0 229.95 42.9 238.35 ;
        RECT  39.9 233.25 41.1 234.45 ;
        RECT  42.45 233.4 43.35 234.3 ;
        RECT  37.5 241.05 47.1 241.95 ;
        RECT  37.5 226.95 47.1 227.85 ;
        RECT  39.3 238.35 40.5 239.55 ;
        RECT  41.7 238.35 42.9 239.55 ;
        RECT  39.3 238.35 40.5 239.55 ;
        RECT  41.7 238.35 42.9 239.55 ;
        RECT  39.3 228.75 40.5 229.95 ;
        RECT  41.7 228.75 42.9 229.95 ;
        RECT  39.3 228.75 40.5 229.95 ;
        RECT  41.7 228.75 42.9 229.95 ;
        RECT  44.1 228.75 45.3 229.95 ;
        RECT  44.1 238.95 45.3 240.15 ;
        RECT  39.9 233.25 41.1 234.45 ;
        RECT  44.1 253.65 45.3 255.6 ;
        RECT  44.1 241.5 45.3 243.45 ;
        RECT  39.3 254.25 40.5 256.05 ;
        RECT  39.3 241.05 40.5 244.65 ;
        RECT  42.0 244.65 42.9 253.05 ;
        RECT  39.9 248.55 41.1 249.75 ;
        RECT  42.45 248.7 43.35 249.6 ;
        RECT  37.5 241.05 47.1 241.95 ;
        RECT  37.5 255.15 47.1 256.05 ;
        RECT  39.3 245.85 40.5 247.05 ;
        RECT  41.7 245.85 42.9 247.05 ;
        RECT  39.3 245.85 40.5 247.05 ;
        RECT  41.7 245.85 42.9 247.05 ;
        RECT  39.3 254.25 40.5 255.45 ;
        RECT  41.7 254.25 42.9 255.45 ;
        RECT  39.3 254.25 40.5 255.45 ;
        RECT  41.7 254.25 42.9 255.45 ;
        RECT  44.1 254.25 45.3 255.45 ;
        RECT  44.1 244.05 45.3 245.25 ;
        RECT  39.9 249.75 41.1 250.95 ;
        RECT  44.1 255.6 45.3 257.55 ;
        RECT  44.1 267.75 45.3 269.7 ;
        RECT  39.3 255.15 40.5 256.95 ;
        RECT  39.3 266.55 40.5 270.15 ;
        RECT  42.0 258.15 42.9 266.55 ;
        RECT  39.9 261.45 41.1 262.65 ;
        RECT  42.45 261.6 43.35 262.5 ;
        RECT  37.5 269.25 47.1 270.15 ;
        RECT  37.5 255.15 47.1 256.05 ;
        RECT  39.3 266.55 40.5 267.75 ;
        RECT  41.7 266.55 42.9 267.75 ;
        RECT  39.3 266.55 40.5 267.75 ;
        RECT  41.7 266.55 42.9 267.75 ;
        RECT  39.3 256.95 40.5 258.15 ;
        RECT  41.7 256.95 42.9 258.15 ;
        RECT  39.3 256.95 40.5 258.15 ;
        RECT  41.7 256.95 42.9 258.15 ;
        RECT  44.1 256.95 45.3 258.15 ;
        RECT  44.1 267.15 45.3 268.35 ;
        RECT  39.9 261.45 41.1 262.65 ;
        RECT  44.1 281.85 45.3 283.8 ;
        RECT  44.1 269.7 45.3 271.65 ;
        RECT  39.3 282.45 40.5 284.25 ;
        RECT  39.3 269.25 40.5 272.85 ;
        RECT  42.0 272.85 42.9 281.25 ;
        RECT  39.9 276.75 41.1 277.95 ;
        RECT  42.45 276.9 43.35 277.8 ;
        RECT  37.5 269.25 47.1 270.15 ;
        RECT  37.5 283.35 47.1 284.25 ;
        RECT  39.3 274.05 40.5 275.25 ;
        RECT  41.7 274.05 42.9 275.25 ;
        RECT  39.3 274.05 40.5 275.25 ;
        RECT  41.7 274.05 42.9 275.25 ;
        RECT  39.3 282.45 40.5 283.65 ;
        RECT  41.7 282.45 42.9 283.65 ;
        RECT  39.3 282.45 40.5 283.65 ;
        RECT  41.7 282.45 42.9 283.65 ;
        RECT  44.1 282.45 45.3 283.65 ;
        RECT  44.1 272.25 45.3 273.45 ;
        RECT  39.9 277.95 41.1 279.15 ;
        RECT  44.1 283.8 45.3 285.75 ;
        RECT  44.1 295.95 45.3 297.9 ;
        RECT  39.3 283.35 40.5 285.15 ;
        RECT  39.3 294.75 40.5 298.35 ;
        RECT  42.0 286.35 42.9 294.75 ;
        RECT  39.9 289.65 41.1 290.85 ;
        RECT  42.45 289.8 43.35 290.7 ;
        RECT  37.5 297.45 47.1 298.35 ;
        RECT  37.5 283.35 47.1 284.25 ;
        RECT  39.3 294.75 40.5 295.95 ;
        RECT  41.7 294.75 42.9 295.95 ;
        RECT  39.3 294.75 40.5 295.95 ;
        RECT  41.7 294.75 42.9 295.95 ;
        RECT  39.3 285.15 40.5 286.35 ;
        RECT  41.7 285.15 42.9 286.35 ;
        RECT  39.3 285.15 40.5 286.35 ;
        RECT  41.7 285.15 42.9 286.35 ;
        RECT  44.1 285.15 45.3 286.35 ;
        RECT  44.1 295.35 45.3 296.55 ;
        RECT  39.9 289.65 41.1 290.85 ;
        RECT  44.1 310.05 45.3 312.0 ;
        RECT  44.1 297.9 45.3 299.85 ;
        RECT  39.3 310.65 40.5 312.45 ;
        RECT  39.3 297.45 40.5 301.05 ;
        RECT  42.0 301.05 42.9 309.45 ;
        RECT  39.9 304.95 41.1 306.15 ;
        RECT  42.45 305.1 43.35 306.0 ;
        RECT  37.5 297.45 47.1 298.35 ;
        RECT  37.5 311.55 47.1 312.45 ;
        RECT  39.3 302.25 40.5 303.45 ;
        RECT  41.7 302.25 42.9 303.45 ;
        RECT  39.3 302.25 40.5 303.45 ;
        RECT  41.7 302.25 42.9 303.45 ;
        RECT  39.3 310.65 40.5 311.85 ;
        RECT  41.7 310.65 42.9 311.85 ;
        RECT  39.3 310.65 40.5 311.85 ;
        RECT  41.7 310.65 42.9 311.85 ;
        RECT  44.1 310.65 45.3 311.85 ;
        RECT  44.1 300.45 45.3 301.65 ;
        RECT  39.9 306.15 41.1 307.35 ;
        RECT  44.1 312.0 45.3 313.95 ;
        RECT  44.1 324.15 45.3 326.1 ;
        RECT  39.3 311.55 40.5 313.35 ;
        RECT  39.3 322.95 40.5 326.55 ;
        RECT  42.0 314.55 42.9 322.95 ;
        RECT  39.9 317.85 41.1 319.05 ;
        RECT  42.45 318.0 43.35 318.9 ;
        RECT  37.5 325.65 47.1 326.55 ;
        RECT  37.5 311.55 47.1 312.45 ;
        RECT  39.3 322.95 40.5 324.15 ;
        RECT  41.7 322.95 42.9 324.15 ;
        RECT  39.3 322.95 40.5 324.15 ;
        RECT  41.7 322.95 42.9 324.15 ;
        RECT  39.3 313.35 40.5 314.55 ;
        RECT  41.7 313.35 42.9 314.55 ;
        RECT  39.3 313.35 40.5 314.55 ;
        RECT  41.7 313.35 42.9 314.55 ;
        RECT  44.1 313.35 45.3 314.55 ;
        RECT  44.1 323.55 45.3 324.75 ;
        RECT  39.9 317.85 41.1 319.05 ;
        RECT  44.1 338.25 45.3 340.2 ;
        RECT  44.1 326.1 45.3 328.05 ;
        RECT  39.3 338.85 40.5 340.65 ;
        RECT  39.3 325.65 40.5 329.25 ;
        RECT  42.0 329.25 42.9 337.65 ;
        RECT  39.9 333.15 41.1 334.35 ;
        RECT  42.45 333.3 43.35 334.2 ;
        RECT  37.5 325.65 47.1 326.55 ;
        RECT  37.5 339.75 47.1 340.65 ;
        RECT  39.3 330.45 40.5 331.65 ;
        RECT  41.7 330.45 42.9 331.65 ;
        RECT  39.3 330.45 40.5 331.65 ;
        RECT  41.7 330.45 42.9 331.65 ;
        RECT  39.3 338.85 40.5 340.05 ;
        RECT  41.7 338.85 42.9 340.05 ;
        RECT  39.3 338.85 40.5 340.05 ;
        RECT  41.7 338.85 42.9 340.05 ;
        RECT  44.1 338.85 45.3 340.05 ;
        RECT  44.1 328.65 45.3 329.85 ;
        RECT  39.9 334.35 41.1 335.55 ;
        RECT  44.1 340.2 45.3 342.15 ;
        RECT  44.1 352.35 45.3 354.3 ;
        RECT  39.3 339.75 40.5 341.55 ;
        RECT  39.3 351.15 40.5 354.75 ;
        RECT  42.0 342.75 42.9 351.15 ;
        RECT  39.9 346.05 41.1 347.25 ;
        RECT  42.45 346.2 43.35 347.1 ;
        RECT  37.5 353.85 47.1 354.75 ;
        RECT  37.5 339.75 47.1 340.65 ;
        RECT  39.3 351.15 40.5 352.35 ;
        RECT  41.7 351.15 42.9 352.35 ;
        RECT  39.3 351.15 40.5 352.35 ;
        RECT  41.7 351.15 42.9 352.35 ;
        RECT  39.3 341.55 40.5 342.75 ;
        RECT  41.7 341.55 42.9 342.75 ;
        RECT  39.3 341.55 40.5 342.75 ;
        RECT  41.7 341.55 42.9 342.75 ;
        RECT  44.1 341.55 45.3 342.75 ;
        RECT  44.1 351.75 45.3 352.95 ;
        RECT  39.9 346.05 41.1 347.25 ;
        RECT  44.1 366.45 45.3 368.4 ;
        RECT  44.1 354.3 45.3 356.25 ;
        RECT  39.3 367.05 40.5 368.85 ;
        RECT  39.3 353.85 40.5 357.45 ;
        RECT  42.0 357.45 42.9 365.85 ;
        RECT  39.9 361.35 41.1 362.55 ;
        RECT  42.45 361.5 43.35 362.4 ;
        RECT  37.5 353.85 47.1 354.75 ;
        RECT  37.5 367.95 47.1 368.85 ;
        RECT  39.3 358.65 40.5 359.85 ;
        RECT  41.7 358.65 42.9 359.85 ;
        RECT  39.3 358.65 40.5 359.85 ;
        RECT  41.7 358.65 42.9 359.85 ;
        RECT  39.3 367.05 40.5 368.25 ;
        RECT  41.7 367.05 42.9 368.25 ;
        RECT  39.3 367.05 40.5 368.25 ;
        RECT  41.7 367.05 42.9 368.25 ;
        RECT  44.1 367.05 45.3 368.25 ;
        RECT  44.1 356.85 45.3 358.05 ;
        RECT  39.9 362.55 41.1 363.75 ;
        RECT  44.1 368.4 45.3 370.35 ;
        RECT  44.1 380.55 45.3 382.5 ;
        RECT  39.3 367.95 40.5 369.75 ;
        RECT  39.3 379.35 40.5 382.95 ;
        RECT  42.0 370.95 42.9 379.35 ;
        RECT  39.9 374.25 41.1 375.45 ;
        RECT  42.45 374.4 43.35 375.3 ;
        RECT  37.5 382.05 47.1 382.95 ;
        RECT  37.5 367.95 47.1 368.85 ;
        RECT  39.3 379.35 40.5 380.55 ;
        RECT  41.7 379.35 42.9 380.55 ;
        RECT  39.3 379.35 40.5 380.55 ;
        RECT  41.7 379.35 42.9 380.55 ;
        RECT  39.3 369.75 40.5 370.95 ;
        RECT  41.7 369.75 42.9 370.95 ;
        RECT  39.3 369.75 40.5 370.95 ;
        RECT  41.7 369.75 42.9 370.95 ;
        RECT  44.1 369.75 45.3 370.95 ;
        RECT  44.1 379.95 45.3 381.15 ;
        RECT  39.9 374.25 41.1 375.45 ;
        RECT  44.1 394.65 45.3 396.6 ;
        RECT  44.1 382.5 45.3 384.45 ;
        RECT  39.3 395.25 40.5 397.05 ;
        RECT  39.3 382.05 40.5 385.65 ;
        RECT  42.0 385.65 42.9 394.05 ;
        RECT  39.9 389.55 41.1 390.75 ;
        RECT  42.45 389.7 43.35 390.6 ;
        RECT  37.5 382.05 47.1 382.95 ;
        RECT  37.5 396.15 47.1 397.05 ;
        RECT  39.3 386.85 40.5 388.05 ;
        RECT  41.7 386.85 42.9 388.05 ;
        RECT  39.3 386.85 40.5 388.05 ;
        RECT  41.7 386.85 42.9 388.05 ;
        RECT  39.3 395.25 40.5 396.45 ;
        RECT  41.7 395.25 42.9 396.45 ;
        RECT  39.3 395.25 40.5 396.45 ;
        RECT  41.7 395.25 42.9 396.45 ;
        RECT  44.1 395.25 45.3 396.45 ;
        RECT  44.1 385.05 45.3 386.25 ;
        RECT  39.9 390.75 41.1 391.95 ;
        RECT  44.1 396.6 45.3 398.55 ;
        RECT  44.1 408.75 45.3 410.7 ;
        RECT  39.3 396.15 40.5 397.95 ;
        RECT  39.3 407.55 40.5 411.15 ;
        RECT  42.0 399.15 42.9 407.55 ;
        RECT  39.9 402.45 41.1 403.65 ;
        RECT  42.45 402.6 43.35 403.5 ;
        RECT  37.5 410.25 47.1 411.15 ;
        RECT  37.5 396.15 47.1 397.05 ;
        RECT  39.3 407.55 40.5 408.75 ;
        RECT  41.7 407.55 42.9 408.75 ;
        RECT  39.3 407.55 40.5 408.75 ;
        RECT  41.7 407.55 42.9 408.75 ;
        RECT  39.3 397.95 40.5 399.15 ;
        RECT  41.7 397.95 42.9 399.15 ;
        RECT  39.3 397.95 40.5 399.15 ;
        RECT  41.7 397.95 42.9 399.15 ;
        RECT  44.1 397.95 45.3 399.15 ;
        RECT  44.1 408.15 45.3 409.35 ;
        RECT  39.9 402.45 41.1 403.65 ;
        RECT  44.1 422.85 45.3 424.8 ;
        RECT  44.1 410.7 45.3 412.65 ;
        RECT  39.3 423.45 40.5 425.25 ;
        RECT  39.3 410.25 40.5 413.85 ;
        RECT  42.0 413.85 42.9 422.25 ;
        RECT  39.9 417.75 41.1 418.95 ;
        RECT  42.45 417.9 43.35 418.8 ;
        RECT  37.5 410.25 47.1 411.15 ;
        RECT  37.5 424.35 47.1 425.25 ;
        RECT  39.3 415.05 40.5 416.25 ;
        RECT  41.7 415.05 42.9 416.25 ;
        RECT  39.3 415.05 40.5 416.25 ;
        RECT  41.7 415.05 42.9 416.25 ;
        RECT  39.3 423.45 40.5 424.65 ;
        RECT  41.7 423.45 42.9 424.65 ;
        RECT  39.3 423.45 40.5 424.65 ;
        RECT  41.7 423.45 42.9 424.65 ;
        RECT  44.1 423.45 45.3 424.65 ;
        RECT  44.1 413.25 45.3 414.45 ;
        RECT  39.9 418.95 41.1 420.15 ;
        RECT  6.15 92.25 7.35 93.45 ;
        RECT  8.25 107.55 9.45 108.75 ;
        RECT  10.35 120.45 11.55 121.65 ;
        RECT  12.45 135.75 13.65 136.95 ;
        RECT  14.55 148.65 15.75 149.85 ;
        RECT  16.65 163.95 17.85 165.15 ;
        RECT  18.75 176.85 19.95 178.05 ;
        RECT  20.85 192.15 22.05 193.35 ;
        RECT  6.15 206.4 7.35 207.6 ;
        RECT  14.55 203.7 15.75 204.9 ;
        RECT  6.15 219.0 7.35 220.2 ;
        RECT  16.65 221.7 17.85 222.9 ;
        RECT  6.15 234.6 7.35 235.8 ;
        RECT  18.75 231.9 19.95 233.1 ;
        RECT  6.15 247.2 7.35 248.4 ;
        RECT  20.85 249.9 22.05 251.1 ;
        RECT  8.25 262.8 9.45 264.0 ;
        RECT  14.55 260.1 15.75 261.3 ;
        RECT  8.25 275.4 9.45 276.6 ;
        RECT  16.65 278.1 17.85 279.3 ;
        RECT  8.25 291.0 9.45 292.2 ;
        RECT  18.75 288.3 19.95 289.5 ;
        RECT  8.25 303.6 9.45 304.8 ;
        RECT  20.85 306.3 22.05 307.5 ;
        RECT  10.35 319.2 11.55 320.4 ;
        RECT  14.55 316.5 15.75 317.7 ;
        RECT  10.35 331.8 11.55 333.0 ;
        RECT  16.65 334.5 17.85 335.7 ;
        RECT  10.35 347.4 11.55 348.6 ;
        RECT  18.75 344.7 19.95 345.9 ;
        RECT  10.35 360.0 11.55 361.2 ;
        RECT  20.85 362.7 22.05 363.9 ;
        RECT  12.45 375.6 13.65 376.8 ;
        RECT  14.55 372.9 15.75 374.1 ;
        RECT  12.45 388.2 13.65 389.4 ;
        RECT  16.65 390.9 17.85 392.1 ;
        RECT  12.45 403.8 13.65 405.0 ;
        RECT  18.75 401.1 19.95 402.3 ;
        RECT  12.45 416.4 13.65 417.6 ;
        RECT  20.85 419.1 22.05 420.3 ;
        RECT  50.25 205.2 55.8 206.1 ;
        RECT  58.35 206.55 59.25 207.45 ;
        RECT  58.35 205.2 59.25 206.1 ;
        RECT  58.35 206.1 59.25 207.0 ;
        RECT  58.8 206.55 65.4 207.45 ;
        RECT  65.4 206.55 66.6 207.45 ;
        RECT  74.85 206.55 75.75 207.45 ;
        RECT  74.85 205.2 75.75 206.1 ;
        RECT  70.8 206.55 75.3 207.45 ;
        RECT  74.85 205.65 75.75 207.0 ;
        RECT  75.3 205.2 79.8 206.1 ;
        RECT  50.25 220.5 55.8 221.4 ;
        RECT  58.35 219.15 59.25 220.05 ;
        RECT  58.35 220.5 59.25 221.4 ;
        RECT  58.35 219.6 59.25 221.4 ;
        RECT  58.8 219.15 65.4 220.05 ;
        RECT  65.4 219.15 66.6 220.05 ;
        RECT  74.85 219.15 75.75 220.05 ;
        RECT  74.85 220.5 75.75 221.4 ;
        RECT  70.8 219.15 75.3 220.05 ;
        RECT  74.85 219.6 75.75 220.95 ;
        RECT  75.3 220.5 79.8 221.4 ;
        RECT  50.25 233.4 55.8 234.3 ;
        RECT  58.35 234.75 59.25 235.65 ;
        RECT  58.35 233.4 59.25 234.3 ;
        RECT  58.35 234.3 59.25 235.2 ;
        RECT  58.8 234.75 65.4 235.65 ;
        RECT  65.4 234.75 66.6 235.65 ;
        RECT  74.85 234.75 75.75 235.65 ;
        RECT  74.85 233.4 75.75 234.3 ;
        RECT  70.8 234.75 75.3 235.65 ;
        RECT  74.85 233.85 75.75 235.2 ;
        RECT  75.3 233.4 79.8 234.3 ;
        RECT  50.25 248.7 55.8 249.6 ;
        RECT  58.35 247.35 59.25 248.25 ;
        RECT  58.35 248.7 59.25 249.6 ;
        RECT  58.35 247.8 59.25 249.6 ;
        RECT  58.8 247.35 65.4 248.25 ;
        RECT  65.4 247.35 66.6 248.25 ;
        RECT  74.85 247.35 75.75 248.25 ;
        RECT  74.85 248.7 75.75 249.6 ;
        RECT  70.8 247.35 75.3 248.25 ;
        RECT  74.85 247.8 75.75 249.15 ;
        RECT  75.3 248.7 79.8 249.6 ;
        RECT  50.25 261.6 55.8 262.5 ;
        RECT  58.35 262.95 59.25 263.85 ;
        RECT  58.35 261.6 59.25 262.5 ;
        RECT  58.35 262.5 59.25 263.4 ;
        RECT  58.8 262.95 65.4 263.85 ;
        RECT  65.4 262.95 66.6 263.85 ;
        RECT  74.85 262.95 75.75 263.85 ;
        RECT  74.85 261.6 75.75 262.5 ;
        RECT  70.8 262.95 75.3 263.85 ;
        RECT  74.85 262.05 75.75 263.4 ;
        RECT  75.3 261.6 79.8 262.5 ;
        RECT  50.25 276.9 55.8 277.8 ;
        RECT  58.35 275.55 59.25 276.45 ;
        RECT  58.35 276.9 59.25 277.8 ;
        RECT  58.35 276.0 59.25 277.8 ;
        RECT  58.8 275.55 65.4 276.45 ;
        RECT  65.4 275.55 66.6 276.45 ;
        RECT  74.85 275.55 75.75 276.45 ;
        RECT  74.85 276.9 75.75 277.8 ;
        RECT  70.8 275.55 75.3 276.45 ;
        RECT  74.85 276.0 75.75 277.35 ;
        RECT  75.3 276.9 79.8 277.8 ;
        RECT  50.25 289.8 55.8 290.7 ;
        RECT  58.35 291.15 59.25 292.05 ;
        RECT  58.35 289.8 59.25 290.7 ;
        RECT  58.35 290.7 59.25 291.6 ;
        RECT  58.8 291.15 65.4 292.05 ;
        RECT  65.4 291.15 66.6 292.05 ;
        RECT  74.85 291.15 75.75 292.05 ;
        RECT  74.85 289.8 75.75 290.7 ;
        RECT  70.8 291.15 75.3 292.05 ;
        RECT  74.85 290.25 75.75 291.6 ;
        RECT  75.3 289.8 79.8 290.7 ;
        RECT  50.25 305.1 55.8 306.0 ;
        RECT  58.35 303.75 59.25 304.65 ;
        RECT  58.35 305.1 59.25 306.0 ;
        RECT  58.35 304.2 59.25 306.0 ;
        RECT  58.8 303.75 65.4 304.65 ;
        RECT  65.4 303.75 66.6 304.65 ;
        RECT  74.85 303.75 75.75 304.65 ;
        RECT  74.85 305.1 75.75 306.0 ;
        RECT  70.8 303.75 75.3 304.65 ;
        RECT  74.85 304.2 75.75 305.55 ;
        RECT  75.3 305.1 79.8 306.0 ;
        RECT  50.25 318.0 55.8 318.9 ;
        RECT  58.35 319.35 59.25 320.25 ;
        RECT  58.35 318.0 59.25 318.9 ;
        RECT  58.35 318.9 59.25 319.8 ;
        RECT  58.8 319.35 65.4 320.25 ;
        RECT  65.4 319.35 66.6 320.25 ;
        RECT  74.85 319.35 75.75 320.25 ;
        RECT  74.85 318.0 75.75 318.9 ;
        RECT  70.8 319.35 75.3 320.25 ;
        RECT  74.85 318.45 75.75 319.8 ;
        RECT  75.3 318.0 79.8 318.9 ;
        RECT  50.25 333.3 55.8 334.2 ;
        RECT  58.35 331.95 59.25 332.85 ;
        RECT  58.35 333.3 59.25 334.2 ;
        RECT  58.35 332.4 59.25 334.2 ;
        RECT  58.8 331.95 65.4 332.85 ;
        RECT  65.4 331.95 66.6 332.85 ;
        RECT  74.85 331.95 75.75 332.85 ;
        RECT  74.85 333.3 75.75 334.2 ;
        RECT  70.8 331.95 75.3 332.85 ;
        RECT  74.85 332.4 75.75 333.75 ;
        RECT  75.3 333.3 79.8 334.2 ;
        RECT  50.25 346.2 55.8 347.1 ;
        RECT  58.35 347.55 59.25 348.45 ;
        RECT  58.35 346.2 59.25 347.1 ;
        RECT  58.35 347.1 59.25 348.0 ;
        RECT  58.8 347.55 65.4 348.45 ;
        RECT  65.4 347.55 66.6 348.45 ;
        RECT  74.85 347.55 75.75 348.45 ;
        RECT  74.85 346.2 75.75 347.1 ;
        RECT  70.8 347.55 75.3 348.45 ;
        RECT  74.85 346.65 75.75 348.0 ;
        RECT  75.3 346.2 79.8 347.1 ;
        RECT  50.25 361.5 55.8 362.4 ;
        RECT  58.35 360.15 59.25 361.05 ;
        RECT  58.35 361.5 59.25 362.4 ;
        RECT  58.35 360.6 59.25 362.4 ;
        RECT  58.8 360.15 65.4 361.05 ;
        RECT  65.4 360.15 66.6 361.05 ;
        RECT  74.85 360.15 75.75 361.05 ;
        RECT  74.85 361.5 75.75 362.4 ;
        RECT  70.8 360.15 75.3 361.05 ;
        RECT  74.85 360.6 75.75 361.95 ;
        RECT  75.3 361.5 79.8 362.4 ;
        RECT  50.25 374.4 55.8 375.3 ;
        RECT  58.35 375.75 59.25 376.65 ;
        RECT  58.35 374.4 59.25 375.3 ;
        RECT  58.35 375.3 59.25 376.2 ;
        RECT  58.8 375.75 65.4 376.65 ;
        RECT  65.4 375.75 66.6 376.65 ;
        RECT  74.85 375.75 75.75 376.65 ;
        RECT  74.85 374.4 75.75 375.3 ;
        RECT  70.8 375.75 75.3 376.65 ;
        RECT  74.85 374.85 75.75 376.2 ;
        RECT  75.3 374.4 79.8 375.3 ;
        RECT  50.25 389.7 55.8 390.6 ;
        RECT  58.35 388.35 59.25 389.25 ;
        RECT  58.35 389.7 59.25 390.6 ;
        RECT  58.35 388.8 59.25 390.6 ;
        RECT  58.8 388.35 65.4 389.25 ;
        RECT  65.4 388.35 66.6 389.25 ;
        RECT  74.85 388.35 75.75 389.25 ;
        RECT  74.85 389.7 75.75 390.6 ;
        RECT  70.8 388.35 75.3 389.25 ;
        RECT  74.85 388.8 75.75 390.15 ;
        RECT  75.3 389.7 79.8 390.6 ;
        RECT  50.25 402.6 55.8 403.5 ;
        RECT  58.35 403.95 59.25 404.85 ;
        RECT  58.35 402.6 59.25 403.5 ;
        RECT  58.35 403.5 59.25 404.4 ;
        RECT  58.8 403.95 65.4 404.85 ;
        RECT  65.4 403.95 66.6 404.85 ;
        RECT  74.85 403.95 75.75 404.85 ;
        RECT  74.85 402.6 75.75 403.5 ;
        RECT  70.8 403.95 75.3 404.85 ;
        RECT  74.85 403.05 75.75 404.4 ;
        RECT  75.3 402.6 79.8 403.5 ;
        RECT  50.25 417.9 55.8 418.8 ;
        RECT  58.35 416.55 59.25 417.45 ;
        RECT  58.35 417.9 59.25 418.8 ;
        RECT  58.35 417.0 59.25 418.8 ;
        RECT  58.8 416.55 65.4 417.45 ;
        RECT  65.4 416.55 66.6 417.45 ;
        RECT  74.85 416.55 75.75 417.45 ;
        RECT  74.85 417.9 75.75 418.8 ;
        RECT  70.8 416.55 75.3 417.45 ;
        RECT  74.85 417.0 75.75 418.35 ;
        RECT  75.3 417.9 79.8 418.8 ;
        RECT  82.35 261.6 83.25 262.5 ;
        RECT  47.1 250.95 52.2 251.85 ;
        RECT  82.35 205.2 83.25 206.1 ;
        RECT  47.1 307.35 52.2 308.25 ;
        RECT  82.35 233.4 83.25 234.3 ;
        RECT  47.1 222.75 52.2 223.65 ;
        RECT  47.1 279.15 52.2 280.05 ;
        RECT  47.1 315.75 52.2 316.65 ;
        RECT  82.35 417.9 83.25 418.8 ;
        RECT  47.1 343.95 52.2 344.85 ;
        RECT  82.35 318.0 83.25 318.9 ;
        RECT  47.1 400.35 52.2 401.25 ;
        RECT  47.1 372.15 52.2 373.05 ;
        RECT  82.35 289.8 83.25 290.7 ;
        RECT  82.35 389.7 83.25 390.6 ;
        RECT  82.35 361.5 83.25 362.4 ;
        RECT  82.35 248.7 83.25 249.6 ;
        RECT  47.1 231.15 52.2 232.05 ;
        RECT  82.35 276.9 83.25 277.8 ;
        RECT  82.35 220.5 83.25 221.4 ;
        RECT  47.1 202.95 52.2 203.85 ;
        RECT  47.1 259.35 52.2 260.25 ;
        RECT  47.1 287.55 52.2 288.45 ;
        RECT  47.1 335.55 52.2 336.45 ;
        RECT  47.1 363.75 52.2 364.65 ;
        RECT  82.35 402.6 83.25 403.5 ;
        RECT  47.1 420.15 52.2 421.05 ;
        RECT  82.35 346.2 83.25 347.1 ;
        RECT  82.35 333.3 83.25 334.2 ;
        RECT  47.1 212.85 53.4 213.75 ;
        RECT  47.1 241.05 53.4 241.95 ;
        RECT  47.1 269.25 53.4 270.15 ;
        RECT  47.1 297.45 53.4 298.35 ;
        RECT  47.1 325.65 53.4 326.55 ;
        RECT  47.1 353.85 53.4 354.75 ;
        RECT  47.1 382.05 53.4 382.95 ;
        RECT  47.1 410.25 53.4 411.15 ;
        RECT  47.1 198.75 53.4 199.65 ;
        RECT  47.1 226.95 53.4 227.85 ;
        RECT  47.1 255.15 53.4 256.05 ;
        RECT  47.1 283.35 53.4 284.25 ;
        RECT  47.1 311.55 53.4 312.45 ;
        RECT  47.1 339.75 53.4 340.65 ;
        RECT  47.1 367.95 53.4 368.85 ;
        RECT  47.1 396.15 53.4 397.05 ;
        RECT  47.1 424.35 53.4 425.25 ;
        RECT  47.1 391.95 52.2 392.85 ;
        RECT  82.35 374.4 83.25 375.3 ;
        RECT  82.35 305.1 83.25 306.0 ;
        RECT  60.0 199.2 61.2 201.15 ;
        RECT  60.0 211.35 61.2 213.3 ;
        RECT  55.2 198.75 56.4 200.55 ;
        RECT  55.2 210.15 56.4 213.75 ;
        RECT  57.9 201.75 58.8 210.15 ;
        RECT  55.8 205.05 57.0 206.25 ;
        RECT  58.35 205.2 59.25 206.1 ;
        RECT  53.4 212.85 63.0 213.75 ;
        RECT  53.4 198.75 63.0 199.65 ;
        RECT  55.2 210.15 56.4 211.35 ;
        RECT  57.6 210.15 58.8 211.35 ;
        RECT  55.2 210.15 56.4 211.35 ;
        RECT  57.6 210.15 58.8 211.35 ;
        RECT  55.2 200.55 56.4 201.75 ;
        RECT  57.6 200.55 58.8 201.75 ;
        RECT  55.2 200.55 56.4 201.75 ;
        RECT  57.6 200.55 58.8 201.75 ;
        RECT  60.0 200.55 61.2 201.75 ;
        RECT  60.0 210.75 61.2 211.95 ;
        RECT  55.8 205.05 57.0 206.25 ;
        RECT  72.0 199.2 73.2 201.15 ;
        RECT  72.0 211.35 73.2 213.3 ;
        RECT  64.8 198.75 66.0 201.15 ;
        RECT  64.8 210.15 66.0 213.75 ;
        RECT  69.6 210.15 70.8 213.75 ;
        RECT  65.4 206.4 66.6 207.6 ;
        RECT  69.6 206.4 70.8 207.6 ;
        RECT  68.4 203.7 69.6 204.9 ;
        RECT  63.0 212.85 77.4 213.75 ;
        RECT  63.0 198.75 77.4 199.65 ;
        RECT  64.8 210.15 66.0 211.35 ;
        RECT  67.2 210.15 68.4 211.35 ;
        RECT  64.8 210.15 66.0 211.35 ;
        RECT  67.2 210.15 68.4 211.35 ;
        RECT  67.2 210.15 68.4 211.35 ;
        RECT  69.6 210.15 70.8 211.35 ;
        RECT  67.2 210.15 68.4 211.35 ;
        RECT  69.6 210.15 70.8 211.35 ;
        RECT  64.8 201.15 66.0 202.35 ;
        RECT  67.2 201.15 68.4 202.35 ;
        RECT  64.8 201.15 66.0 202.35 ;
        RECT  67.2 201.15 68.4 202.35 ;
        RECT  67.2 201.15 68.4 202.35 ;
        RECT  69.6 201.15 70.8 202.35 ;
        RECT  67.2 201.15 68.4 202.35 ;
        RECT  69.6 201.15 70.8 202.35 ;
        RECT  72.0 200.55 73.2 201.75 ;
        RECT  72.0 210.75 73.2 211.95 ;
        RECT  68.4 203.7 69.6 204.9 ;
        RECT  65.4 206.4 66.6 207.6 ;
        RECT  67.2 210.15 68.4 211.35 ;
        RECT  69.6 201.15 70.8 202.35 ;
        RECT  69.6 206.4 70.8 207.6 ;
        RECT  84.0 199.2 85.2 201.15 ;
        RECT  84.0 211.35 85.2 213.3 ;
        RECT  79.2 198.75 80.4 200.55 ;
        RECT  79.2 210.15 80.4 213.75 ;
        RECT  81.9 201.75 82.8 210.15 ;
        RECT  79.8 205.05 81.0 206.25 ;
        RECT  82.35 205.2 83.25 206.1 ;
        RECT  77.4 212.85 87.0 213.75 ;
        RECT  77.4 198.75 87.0 199.65 ;
        RECT  79.2 210.15 80.4 211.35 ;
        RECT  81.6 210.15 82.8 211.35 ;
        RECT  79.2 210.15 80.4 211.35 ;
        RECT  81.6 210.15 82.8 211.35 ;
        RECT  79.2 200.55 80.4 201.75 ;
        RECT  81.6 200.55 82.8 201.75 ;
        RECT  79.2 200.55 80.4 201.75 ;
        RECT  81.6 200.55 82.8 201.75 ;
        RECT  84.0 200.55 85.2 201.75 ;
        RECT  84.0 210.75 85.2 211.95 ;
        RECT  79.8 205.05 81.0 206.25 ;
        RECT  49.65 205.05 50.85 206.25 ;
        RECT  51.6 202.8 52.8 204.0 ;
        RECT  67.2 203.7 68.4 204.9 ;
        RECT  60.0 225.45 61.2 227.4 ;
        RECT  60.0 213.3 61.2 215.25 ;
        RECT  55.2 226.05 56.4 227.85 ;
        RECT  55.2 212.85 56.4 216.45 ;
        RECT  57.9 216.45 58.8 224.85 ;
        RECT  55.8 220.35 57.0 221.55 ;
        RECT  58.35 220.5 59.25 221.4 ;
        RECT  53.4 212.85 63.0 213.75 ;
        RECT  53.4 226.95 63.0 227.85 ;
        RECT  55.2 217.65 56.4 218.85 ;
        RECT  57.6 217.65 58.8 218.85 ;
        RECT  55.2 217.65 56.4 218.85 ;
        RECT  57.6 217.65 58.8 218.85 ;
        RECT  55.2 226.05 56.4 227.25 ;
        RECT  57.6 226.05 58.8 227.25 ;
        RECT  55.2 226.05 56.4 227.25 ;
        RECT  57.6 226.05 58.8 227.25 ;
        RECT  60.0 226.05 61.2 227.25 ;
        RECT  60.0 215.85 61.2 217.05 ;
        RECT  55.8 221.55 57.0 222.75 ;
        RECT  72.0 225.45 73.2 227.4 ;
        RECT  72.0 213.3 73.2 215.25 ;
        RECT  64.8 225.45 66.0 227.85 ;
        RECT  64.8 212.85 66.0 216.45 ;
        RECT  69.6 212.85 70.8 216.45 ;
        RECT  65.4 219.0 66.6 220.2 ;
        RECT  69.6 219.0 70.8 220.2 ;
        RECT  68.4 221.7 69.6 222.9 ;
        RECT  63.0 212.85 77.4 213.75 ;
        RECT  63.0 226.95 77.4 227.85 ;
        RECT  64.8 217.65 66.0 218.85 ;
        RECT  67.2 217.65 68.4 218.85 ;
        RECT  64.8 217.65 66.0 218.85 ;
        RECT  67.2 217.65 68.4 218.85 ;
        RECT  67.2 217.65 68.4 218.85 ;
        RECT  69.6 217.65 70.8 218.85 ;
        RECT  67.2 217.65 68.4 218.85 ;
        RECT  69.6 217.65 70.8 218.85 ;
        RECT  64.8 226.65 66.0 227.85 ;
        RECT  67.2 226.65 68.4 227.85 ;
        RECT  64.8 226.65 66.0 227.85 ;
        RECT  67.2 226.65 68.4 227.85 ;
        RECT  67.2 226.65 68.4 227.85 ;
        RECT  69.6 226.65 70.8 227.85 ;
        RECT  67.2 226.65 68.4 227.85 ;
        RECT  69.6 226.65 70.8 227.85 ;
        RECT  72.0 226.05 73.2 227.25 ;
        RECT  72.0 215.85 73.2 217.05 ;
        RECT  68.4 222.9 69.6 224.1 ;
        RECT  65.4 220.2 66.6 221.4 ;
        RECT  67.2 216.45 68.4 217.65 ;
        RECT  69.6 225.45 70.8 226.65 ;
        RECT  69.6 220.2 70.8 221.4 ;
        RECT  84.0 225.45 85.2 227.4 ;
        RECT  84.0 213.3 85.2 215.25 ;
        RECT  79.2 226.05 80.4 227.85 ;
        RECT  79.2 212.85 80.4 216.45 ;
        RECT  81.9 216.45 82.8 224.85 ;
        RECT  79.8 220.35 81.0 221.55 ;
        RECT  82.35 220.5 83.25 221.4 ;
        RECT  77.4 212.85 87.0 213.75 ;
        RECT  77.4 226.95 87.0 227.85 ;
        RECT  79.2 217.65 80.4 218.85 ;
        RECT  81.6 217.65 82.8 218.85 ;
        RECT  79.2 217.65 80.4 218.85 ;
        RECT  81.6 217.65 82.8 218.85 ;
        RECT  79.2 226.05 80.4 227.25 ;
        RECT  81.6 226.05 82.8 227.25 ;
        RECT  79.2 226.05 80.4 227.25 ;
        RECT  81.6 226.05 82.8 227.25 ;
        RECT  84.0 226.05 85.2 227.25 ;
        RECT  84.0 215.85 85.2 217.05 ;
        RECT  79.8 221.55 81.0 222.75 ;
        RECT  49.65 220.35 50.85 221.55 ;
        RECT  51.6 222.6 52.8 223.8 ;
        RECT  67.2 221.7 68.4 222.9 ;
        RECT  60.0 227.4 61.2 229.35 ;
        RECT  60.0 239.55 61.2 241.5 ;
        RECT  55.2 226.95 56.4 228.75 ;
        RECT  55.2 238.35 56.4 241.95 ;
        RECT  57.9 229.95 58.8 238.35 ;
        RECT  55.8 233.25 57.0 234.45 ;
        RECT  58.35 233.4 59.25 234.3 ;
        RECT  53.4 241.05 63.0 241.95 ;
        RECT  53.4 226.95 63.0 227.85 ;
        RECT  55.2 238.35 56.4 239.55 ;
        RECT  57.6 238.35 58.8 239.55 ;
        RECT  55.2 238.35 56.4 239.55 ;
        RECT  57.6 238.35 58.8 239.55 ;
        RECT  55.2 228.75 56.4 229.95 ;
        RECT  57.6 228.75 58.8 229.95 ;
        RECT  55.2 228.75 56.4 229.95 ;
        RECT  57.6 228.75 58.8 229.95 ;
        RECT  60.0 228.75 61.2 229.95 ;
        RECT  60.0 238.95 61.2 240.15 ;
        RECT  55.8 233.25 57.0 234.45 ;
        RECT  72.0 227.4 73.2 229.35 ;
        RECT  72.0 239.55 73.2 241.5 ;
        RECT  64.8 226.95 66.0 229.35 ;
        RECT  64.8 238.35 66.0 241.95 ;
        RECT  69.6 238.35 70.8 241.95 ;
        RECT  65.4 234.6 66.6 235.8 ;
        RECT  69.6 234.6 70.8 235.8 ;
        RECT  68.4 231.9 69.6 233.1 ;
        RECT  63.0 241.05 77.4 241.95 ;
        RECT  63.0 226.95 77.4 227.85 ;
        RECT  64.8 238.35 66.0 239.55 ;
        RECT  67.2 238.35 68.4 239.55 ;
        RECT  64.8 238.35 66.0 239.55 ;
        RECT  67.2 238.35 68.4 239.55 ;
        RECT  67.2 238.35 68.4 239.55 ;
        RECT  69.6 238.35 70.8 239.55 ;
        RECT  67.2 238.35 68.4 239.55 ;
        RECT  69.6 238.35 70.8 239.55 ;
        RECT  64.8 229.35 66.0 230.55 ;
        RECT  67.2 229.35 68.4 230.55 ;
        RECT  64.8 229.35 66.0 230.55 ;
        RECT  67.2 229.35 68.4 230.55 ;
        RECT  67.2 229.35 68.4 230.55 ;
        RECT  69.6 229.35 70.8 230.55 ;
        RECT  67.2 229.35 68.4 230.55 ;
        RECT  69.6 229.35 70.8 230.55 ;
        RECT  72.0 228.75 73.2 229.95 ;
        RECT  72.0 238.95 73.2 240.15 ;
        RECT  68.4 231.9 69.6 233.1 ;
        RECT  65.4 234.6 66.6 235.8 ;
        RECT  67.2 238.35 68.4 239.55 ;
        RECT  69.6 229.35 70.8 230.55 ;
        RECT  69.6 234.6 70.8 235.8 ;
        RECT  84.0 227.4 85.2 229.35 ;
        RECT  84.0 239.55 85.2 241.5 ;
        RECT  79.2 226.95 80.4 228.75 ;
        RECT  79.2 238.35 80.4 241.95 ;
        RECT  81.9 229.95 82.8 238.35 ;
        RECT  79.8 233.25 81.0 234.45 ;
        RECT  82.35 233.4 83.25 234.3 ;
        RECT  77.4 241.05 87.0 241.95 ;
        RECT  77.4 226.95 87.0 227.85 ;
        RECT  79.2 238.35 80.4 239.55 ;
        RECT  81.6 238.35 82.8 239.55 ;
        RECT  79.2 238.35 80.4 239.55 ;
        RECT  81.6 238.35 82.8 239.55 ;
        RECT  79.2 228.75 80.4 229.95 ;
        RECT  81.6 228.75 82.8 229.95 ;
        RECT  79.2 228.75 80.4 229.95 ;
        RECT  81.6 228.75 82.8 229.95 ;
        RECT  84.0 228.75 85.2 229.95 ;
        RECT  84.0 238.95 85.2 240.15 ;
        RECT  79.8 233.25 81.0 234.45 ;
        RECT  49.65 233.25 50.85 234.45 ;
        RECT  51.6 231.0 52.8 232.2 ;
        RECT  67.2 231.9 68.4 233.1 ;
        RECT  60.0 253.65 61.2 255.6 ;
        RECT  60.0 241.5 61.2 243.45 ;
        RECT  55.2 254.25 56.4 256.05 ;
        RECT  55.2 241.05 56.4 244.65 ;
        RECT  57.9 244.65 58.8 253.05 ;
        RECT  55.8 248.55 57.0 249.75 ;
        RECT  58.35 248.7 59.25 249.6 ;
        RECT  53.4 241.05 63.0 241.95 ;
        RECT  53.4 255.15 63.0 256.05 ;
        RECT  55.2 245.85 56.4 247.05 ;
        RECT  57.6 245.85 58.8 247.05 ;
        RECT  55.2 245.85 56.4 247.05 ;
        RECT  57.6 245.85 58.8 247.05 ;
        RECT  55.2 254.25 56.4 255.45 ;
        RECT  57.6 254.25 58.8 255.45 ;
        RECT  55.2 254.25 56.4 255.45 ;
        RECT  57.6 254.25 58.8 255.45 ;
        RECT  60.0 254.25 61.2 255.45 ;
        RECT  60.0 244.05 61.2 245.25 ;
        RECT  55.8 249.75 57.0 250.95 ;
        RECT  72.0 253.65 73.2 255.6 ;
        RECT  72.0 241.5 73.2 243.45 ;
        RECT  64.8 253.65 66.0 256.05 ;
        RECT  64.8 241.05 66.0 244.65 ;
        RECT  69.6 241.05 70.8 244.65 ;
        RECT  65.4 247.2 66.6 248.4 ;
        RECT  69.6 247.2 70.8 248.4 ;
        RECT  68.4 249.9 69.6 251.1 ;
        RECT  63.0 241.05 77.4 241.95 ;
        RECT  63.0 255.15 77.4 256.05 ;
        RECT  64.8 245.85 66.0 247.05 ;
        RECT  67.2 245.85 68.4 247.05 ;
        RECT  64.8 245.85 66.0 247.05 ;
        RECT  67.2 245.85 68.4 247.05 ;
        RECT  67.2 245.85 68.4 247.05 ;
        RECT  69.6 245.85 70.8 247.05 ;
        RECT  67.2 245.85 68.4 247.05 ;
        RECT  69.6 245.85 70.8 247.05 ;
        RECT  64.8 254.85 66.0 256.05 ;
        RECT  67.2 254.85 68.4 256.05 ;
        RECT  64.8 254.85 66.0 256.05 ;
        RECT  67.2 254.85 68.4 256.05 ;
        RECT  67.2 254.85 68.4 256.05 ;
        RECT  69.6 254.85 70.8 256.05 ;
        RECT  67.2 254.85 68.4 256.05 ;
        RECT  69.6 254.85 70.8 256.05 ;
        RECT  72.0 254.25 73.2 255.45 ;
        RECT  72.0 244.05 73.2 245.25 ;
        RECT  68.4 251.1 69.6 252.3 ;
        RECT  65.4 248.4 66.6 249.6 ;
        RECT  67.2 244.65 68.4 245.85 ;
        RECT  69.6 253.65 70.8 254.85 ;
        RECT  69.6 248.4 70.8 249.6 ;
        RECT  84.0 253.65 85.2 255.6 ;
        RECT  84.0 241.5 85.2 243.45 ;
        RECT  79.2 254.25 80.4 256.05 ;
        RECT  79.2 241.05 80.4 244.65 ;
        RECT  81.9 244.65 82.8 253.05 ;
        RECT  79.8 248.55 81.0 249.75 ;
        RECT  82.35 248.7 83.25 249.6 ;
        RECT  77.4 241.05 87.0 241.95 ;
        RECT  77.4 255.15 87.0 256.05 ;
        RECT  79.2 245.85 80.4 247.05 ;
        RECT  81.6 245.85 82.8 247.05 ;
        RECT  79.2 245.85 80.4 247.05 ;
        RECT  81.6 245.85 82.8 247.05 ;
        RECT  79.2 254.25 80.4 255.45 ;
        RECT  81.6 254.25 82.8 255.45 ;
        RECT  79.2 254.25 80.4 255.45 ;
        RECT  81.6 254.25 82.8 255.45 ;
        RECT  84.0 254.25 85.2 255.45 ;
        RECT  84.0 244.05 85.2 245.25 ;
        RECT  79.8 249.75 81.0 250.95 ;
        RECT  49.65 248.55 50.85 249.75 ;
        RECT  51.6 250.8 52.8 252.0 ;
        RECT  67.2 249.9 68.4 251.1 ;
        RECT  60.0 255.6 61.2 257.55 ;
        RECT  60.0 267.75 61.2 269.7 ;
        RECT  55.2 255.15 56.4 256.95 ;
        RECT  55.2 266.55 56.4 270.15 ;
        RECT  57.9 258.15 58.8 266.55 ;
        RECT  55.8 261.45 57.0 262.65 ;
        RECT  58.35 261.6 59.25 262.5 ;
        RECT  53.4 269.25 63.0 270.15 ;
        RECT  53.4 255.15 63.0 256.05 ;
        RECT  55.2 266.55 56.4 267.75 ;
        RECT  57.6 266.55 58.8 267.75 ;
        RECT  55.2 266.55 56.4 267.75 ;
        RECT  57.6 266.55 58.8 267.75 ;
        RECT  55.2 256.95 56.4 258.15 ;
        RECT  57.6 256.95 58.8 258.15 ;
        RECT  55.2 256.95 56.4 258.15 ;
        RECT  57.6 256.95 58.8 258.15 ;
        RECT  60.0 256.95 61.2 258.15 ;
        RECT  60.0 267.15 61.2 268.35 ;
        RECT  55.8 261.45 57.0 262.65 ;
        RECT  72.0 255.6 73.2 257.55 ;
        RECT  72.0 267.75 73.2 269.7 ;
        RECT  64.8 255.15 66.0 257.55 ;
        RECT  64.8 266.55 66.0 270.15 ;
        RECT  69.6 266.55 70.8 270.15 ;
        RECT  65.4 262.8 66.6 264.0 ;
        RECT  69.6 262.8 70.8 264.0 ;
        RECT  68.4 260.1 69.6 261.3 ;
        RECT  63.0 269.25 77.4 270.15 ;
        RECT  63.0 255.15 77.4 256.05 ;
        RECT  64.8 266.55 66.0 267.75 ;
        RECT  67.2 266.55 68.4 267.75 ;
        RECT  64.8 266.55 66.0 267.75 ;
        RECT  67.2 266.55 68.4 267.75 ;
        RECT  67.2 266.55 68.4 267.75 ;
        RECT  69.6 266.55 70.8 267.75 ;
        RECT  67.2 266.55 68.4 267.75 ;
        RECT  69.6 266.55 70.8 267.75 ;
        RECT  64.8 257.55 66.0 258.75 ;
        RECT  67.2 257.55 68.4 258.75 ;
        RECT  64.8 257.55 66.0 258.75 ;
        RECT  67.2 257.55 68.4 258.75 ;
        RECT  67.2 257.55 68.4 258.75 ;
        RECT  69.6 257.55 70.8 258.75 ;
        RECT  67.2 257.55 68.4 258.75 ;
        RECT  69.6 257.55 70.8 258.75 ;
        RECT  72.0 256.95 73.2 258.15 ;
        RECT  72.0 267.15 73.2 268.35 ;
        RECT  68.4 260.1 69.6 261.3 ;
        RECT  65.4 262.8 66.6 264.0 ;
        RECT  67.2 266.55 68.4 267.75 ;
        RECT  69.6 257.55 70.8 258.75 ;
        RECT  69.6 262.8 70.8 264.0 ;
        RECT  84.0 255.6 85.2 257.55 ;
        RECT  84.0 267.75 85.2 269.7 ;
        RECT  79.2 255.15 80.4 256.95 ;
        RECT  79.2 266.55 80.4 270.15 ;
        RECT  81.9 258.15 82.8 266.55 ;
        RECT  79.8 261.45 81.0 262.65 ;
        RECT  82.35 261.6 83.25 262.5 ;
        RECT  77.4 269.25 87.0 270.15 ;
        RECT  77.4 255.15 87.0 256.05 ;
        RECT  79.2 266.55 80.4 267.75 ;
        RECT  81.6 266.55 82.8 267.75 ;
        RECT  79.2 266.55 80.4 267.75 ;
        RECT  81.6 266.55 82.8 267.75 ;
        RECT  79.2 256.95 80.4 258.15 ;
        RECT  81.6 256.95 82.8 258.15 ;
        RECT  79.2 256.95 80.4 258.15 ;
        RECT  81.6 256.95 82.8 258.15 ;
        RECT  84.0 256.95 85.2 258.15 ;
        RECT  84.0 267.15 85.2 268.35 ;
        RECT  79.8 261.45 81.0 262.65 ;
        RECT  49.65 261.45 50.85 262.65 ;
        RECT  51.6 259.2 52.8 260.4 ;
        RECT  67.2 260.1 68.4 261.3 ;
        RECT  60.0 281.85 61.2 283.8 ;
        RECT  60.0 269.7 61.2 271.65 ;
        RECT  55.2 282.45 56.4 284.25 ;
        RECT  55.2 269.25 56.4 272.85 ;
        RECT  57.9 272.85 58.8 281.25 ;
        RECT  55.8 276.75 57.0 277.95 ;
        RECT  58.35 276.9 59.25 277.8 ;
        RECT  53.4 269.25 63.0 270.15 ;
        RECT  53.4 283.35 63.0 284.25 ;
        RECT  55.2 274.05 56.4 275.25 ;
        RECT  57.6 274.05 58.8 275.25 ;
        RECT  55.2 274.05 56.4 275.25 ;
        RECT  57.6 274.05 58.8 275.25 ;
        RECT  55.2 282.45 56.4 283.65 ;
        RECT  57.6 282.45 58.8 283.65 ;
        RECT  55.2 282.45 56.4 283.65 ;
        RECT  57.6 282.45 58.8 283.65 ;
        RECT  60.0 282.45 61.2 283.65 ;
        RECT  60.0 272.25 61.2 273.45 ;
        RECT  55.8 277.95 57.0 279.15 ;
        RECT  72.0 281.85 73.2 283.8 ;
        RECT  72.0 269.7 73.2 271.65 ;
        RECT  64.8 281.85 66.0 284.25 ;
        RECT  64.8 269.25 66.0 272.85 ;
        RECT  69.6 269.25 70.8 272.85 ;
        RECT  65.4 275.4 66.6 276.6 ;
        RECT  69.6 275.4 70.8 276.6 ;
        RECT  68.4 278.1 69.6 279.3 ;
        RECT  63.0 269.25 77.4 270.15 ;
        RECT  63.0 283.35 77.4 284.25 ;
        RECT  64.8 274.05 66.0 275.25 ;
        RECT  67.2 274.05 68.4 275.25 ;
        RECT  64.8 274.05 66.0 275.25 ;
        RECT  67.2 274.05 68.4 275.25 ;
        RECT  67.2 274.05 68.4 275.25 ;
        RECT  69.6 274.05 70.8 275.25 ;
        RECT  67.2 274.05 68.4 275.25 ;
        RECT  69.6 274.05 70.8 275.25 ;
        RECT  64.8 283.05 66.0 284.25 ;
        RECT  67.2 283.05 68.4 284.25 ;
        RECT  64.8 283.05 66.0 284.25 ;
        RECT  67.2 283.05 68.4 284.25 ;
        RECT  67.2 283.05 68.4 284.25 ;
        RECT  69.6 283.05 70.8 284.25 ;
        RECT  67.2 283.05 68.4 284.25 ;
        RECT  69.6 283.05 70.8 284.25 ;
        RECT  72.0 282.45 73.2 283.65 ;
        RECT  72.0 272.25 73.2 273.45 ;
        RECT  68.4 279.3 69.6 280.5 ;
        RECT  65.4 276.6 66.6 277.8 ;
        RECT  67.2 272.85 68.4 274.05 ;
        RECT  69.6 281.85 70.8 283.05 ;
        RECT  69.6 276.6 70.8 277.8 ;
        RECT  84.0 281.85 85.2 283.8 ;
        RECT  84.0 269.7 85.2 271.65 ;
        RECT  79.2 282.45 80.4 284.25 ;
        RECT  79.2 269.25 80.4 272.85 ;
        RECT  81.9 272.85 82.8 281.25 ;
        RECT  79.8 276.75 81.0 277.95 ;
        RECT  82.35 276.9 83.25 277.8 ;
        RECT  77.4 269.25 87.0 270.15 ;
        RECT  77.4 283.35 87.0 284.25 ;
        RECT  79.2 274.05 80.4 275.25 ;
        RECT  81.6 274.05 82.8 275.25 ;
        RECT  79.2 274.05 80.4 275.25 ;
        RECT  81.6 274.05 82.8 275.25 ;
        RECT  79.2 282.45 80.4 283.65 ;
        RECT  81.6 282.45 82.8 283.65 ;
        RECT  79.2 282.45 80.4 283.65 ;
        RECT  81.6 282.45 82.8 283.65 ;
        RECT  84.0 282.45 85.2 283.65 ;
        RECT  84.0 272.25 85.2 273.45 ;
        RECT  79.8 277.95 81.0 279.15 ;
        RECT  49.65 276.75 50.85 277.95 ;
        RECT  51.6 279.0 52.8 280.2 ;
        RECT  67.2 278.1 68.4 279.3 ;
        RECT  60.0 283.8 61.2 285.75 ;
        RECT  60.0 295.95 61.2 297.9 ;
        RECT  55.2 283.35 56.4 285.15 ;
        RECT  55.2 294.75 56.4 298.35 ;
        RECT  57.9 286.35 58.8 294.75 ;
        RECT  55.8 289.65 57.0 290.85 ;
        RECT  58.35 289.8 59.25 290.7 ;
        RECT  53.4 297.45 63.0 298.35 ;
        RECT  53.4 283.35 63.0 284.25 ;
        RECT  55.2 294.75 56.4 295.95 ;
        RECT  57.6 294.75 58.8 295.95 ;
        RECT  55.2 294.75 56.4 295.95 ;
        RECT  57.6 294.75 58.8 295.95 ;
        RECT  55.2 285.15 56.4 286.35 ;
        RECT  57.6 285.15 58.8 286.35 ;
        RECT  55.2 285.15 56.4 286.35 ;
        RECT  57.6 285.15 58.8 286.35 ;
        RECT  60.0 285.15 61.2 286.35 ;
        RECT  60.0 295.35 61.2 296.55 ;
        RECT  55.8 289.65 57.0 290.85 ;
        RECT  72.0 283.8 73.2 285.75 ;
        RECT  72.0 295.95 73.2 297.9 ;
        RECT  64.8 283.35 66.0 285.75 ;
        RECT  64.8 294.75 66.0 298.35 ;
        RECT  69.6 294.75 70.8 298.35 ;
        RECT  65.4 291.0 66.6 292.2 ;
        RECT  69.6 291.0 70.8 292.2 ;
        RECT  68.4 288.3 69.6 289.5 ;
        RECT  63.0 297.45 77.4 298.35 ;
        RECT  63.0 283.35 77.4 284.25 ;
        RECT  64.8 294.75 66.0 295.95 ;
        RECT  67.2 294.75 68.4 295.95 ;
        RECT  64.8 294.75 66.0 295.95 ;
        RECT  67.2 294.75 68.4 295.95 ;
        RECT  67.2 294.75 68.4 295.95 ;
        RECT  69.6 294.75 70.8 295.95 ;
        RECT  67.2 294.75 68.4 295.95 ;
        RECT  69.6 294.75 70.8 295.95 ;
        RECT  64.8 285.75 66.0 286.95 ;
        RECT  67.2 285.75 68.4 286.95 ;
        RECT  64.8 285.75 66.0 286.95 ;
        RECT  67.2 285.75 68.4 286.95 ;
        RECT  67.2 285.75 68.4 286.95 ;
        RECT  69.6 285.75 70.8 286.95 ;
        RECT  67.2 285.75 68.4 286.95 ;
        RECT  69.6 285.75 70.8 286.95 ;
        RECT  72.0 285.15 73.2 286.35 ;
        RECT  72.0 295.35 73.2 296.55 ;
        RECT  68.4 288.3 69.6 289.5 ;
        RECT  65.4 291.0 66.6 292.2 ;
        RECT  67.2 294.75 68.4 295.95 ;
        RECT  69.6 285.75 70.8 286.95 ;
        RECT  69.6 291.0 70.8 292.2 ;
        RECT  84.0 283.8 85.2 285.75 ;
        RECT  84.0 295.95 85.2 297.9 ;
        RECT  79.2 283.35 80.4 285.15 ;
        RECT  79.2 294.75 80.4 298.35 ;
        RECT  81.9 286.35 82.8 294.75 ;
        RECT  79.8 289.65 81.0 290.85 ;
        RECT  82.35 289.8 83.25 290.7 ;
        RECT  77.4 297.45 87.0 298.35 ;
        RECT  77.4 283.35 87.0 284.25 ;
        RECT  79.2 294.75 80.4 295.95 ;
        RECT  81.6 294.75 82.8 295.95 ;
        RECT  79.2 294.75 80.4 295.95 ;
        RECT  81.6 294.75 82.8 295.95 ;
        RECT  79.2 285.15 80.4 286.35 ;
        RECT  81.6 285.15 82.8 286.35 ;
        RECT  79.2 285.15 80.4 286.35 ;
        RECT  81.6 285.15 82.8 286.35 ;
        RECT  84.0 285.15 85.2 286.35 ;
        RECT  84.0 295.35 85.2 296.55 ;
        RECT  79.8 289.65 81.0 290.85 ;
        RECT  49.65 289.65 50.85 290.85 ;
        RECT  51.6 287.4 52.8 288.6 ;
        RECT  67.2 288.3 68.4 289.5 ;
        RECT  60.0 310.05 61.2 312.0 ;
        RECT  60.0 297.9 61.2 299.85 ;
        RECT  55.2 310.65 56.4 312.45 ;
        RECT  55.2 297.45 56.4 301.05 ;
        RECT  57.9 301.05 58.8 309.45 ;
        RECT  55.8 304.95 57.0 306.15 ;
        RECT  58.35 305.1 59.25 306.0 ;
        RECT  53.4 297.45 63.0 298.35 ;
        RECT  53.4 311.55 63.0 312.45 ;
        RECT  55.2 302.25 56.4 303.45 ;
        RECT  57.6 302.25 58.8 303.45 ;
        RECT  55.2 302.25 56.4 303.45 ;
        RECT  57.6 302.25 58.8 303.45 ;
        RECT  55.2 310.65 56.4 311.85 ;
        RECT  57.6 310.65 58.8 311.85 ;
        RECT  55.2 310.65 56.4 311.85 ;
        RECT  57.6 310.65 58.8 311.85 ;
        RECT  60.0 310.65 61.2 311.85 ;
        RECT  60.0 300.45 61.2 301.65 ;
        RECT  55.8 306.15 57.0 307.35 ;
        RECT  72.0 310.05 73.2 312.0 ;
        RECT  72.0 297.9 73.2 299.85 ;
        RECT  64.8 310.05 66.0 312.45 ;
        RECT  64.8 297.45 66.0 301.05 ;
        RECT  69.6 297.45 70.8 301.05 ;
        RECT  65.4 303.6 66.6 304.8 ;
        RECT  69.6 303.6 70.8 304.8 ;
        RECT  68.4 306.3 69.6 307.5 ;
        RECT  63.0 297.45 77.4 298.35 ;
        RECT  63.0 311.55 77.4 312.45 ;
        RECT  64.8 302.25 66.0 303.45 ;
        RECT  67.2 302.25 68.4 303.45 ;
        RECT  64.8 302.25 66.0 303.45 ;
        RECT  67.2 302.25 68.4 303.45 ;
        RECT  67.2 302.25 68.4 303.45 ;
        RECT  69.6 302.25 70.8 303.45 ;
        RECT  67.2 302.25 68.4 303.45 ;
        RECT  69.6 302.25 70.8 303.45 ;
        RECT  64.8 311.25 66.0 312.45 ;
        RECT  67.2 311.25 68.4 312.45 ;
        RECT  64.8 311.25 66.0 312.45 ;
        RECT  67.2 311.25 68.4 312.45 ;
        RECT  67.2 311.25 68.4 312.45 ;
        RECT  69.6 311.25 70.8 312.45 ;
        RECT  67.2 311.25 68.4 312.45 ;
        RECT  69.6 311.25 70.8 312.45 ;
        RECT  72.0 310.65 73.2 311.85 ;
        RECT  72.0 300.45 73.2 301.65 ;
        RECT  68.4 307.5 69.6 308.7 ;
        RECT  65.4 304.8 66.6 306.0 ;
        RECT  67.2 301.05 68.4 302.25 ;
        RECT  69.6 310.05 70.8 311.25 ;
        RECT  69.6 304.8 70.8 306.0 ;
        RECT  84.0 310.05 85.2 312.0 ;
        RECT  84.0 297.9 85.2 299.85 ;
        RECT  79.2 310.65 80.4 312.45 ;
        RECT  79.2 297.45 80.4 301.05 ;
        RECT  81.9 301.05 82.8 309.45 ;
        RECT  79.8 304.95 81.0 306.15 ;
        RECT  82.35 305.1 83.25 306.0 ;
        RECT  77.4 297.45 87.0 298.35 ;
        RECT  77.4 311.55 87.0 312.45 ;
        RECT  79.2 302.25 80.4 303.45 ;
        RECT  81.6 302.25 82.8 303.45 ;
        RECT  79.2 302.25 80.4 303.45 ;
        RECT  81.6 302.25 82.8 303.45 ;
        RECT  79.2 310.65 80.4 311.85 ;
        RECT  81.6 310.65 82.8 311.85 ;
        RECT  79.2 310.65 80.4 311.85 ;
        RECT  81.6 310.65 82.8 311.85 ;
        RECT  84.0 310.65 85.2 311.85 ;
        RECT  84.0 300.45 85.2 301.65 ;
        RECT  79.8 306.15 81.0 307.35 ;
        RECT  49.65 304.95 50.85 306.15 ;
        RECT  51.6 307.2 52.8 308.4 ;
        RECT  67.2 306.3 68.4 307.5 ;
        RECT  60.0 312.0 61.2 313.95 ;
        RECT  60.0 324.15 61.2 326.1 ;
        RECT  55.2 311.55 56.4 313.35 ;
        RECT  55.2 322.95 56.4 326.55 ;
        RECT  57.9 314.55 58.8 322.95 ;
        RECT  55.8 317.85 57.0 319.05 ;
        RECT  58.35 318.0 59.25 318.9 ;
        RECT  53.4 325.65 63.0 326.55 ;
        RECT  53.4 311.55 63.0 312.45 ;
        RECT  55.2 322.95 56.4 324.15 ;
        RECT  57.6 322.95 58.8 324.15 ;
        RECT  55.2 322.95 56.4 324.15 ;
        RECT  57.6 322.95 58.8 324.15 ;
        RECT  55.2 313.35 56.4 314.55 ;
        RECT  57.6 313.35 58.8 314.55 ;
        RECT  55.2 313.35 56.4 314.55 ;
        RECT  57.6 313.35 58.8 314.55 ;
        RECT  60.0 313.35 61.2 314.55 ;
        RECT  60.0 323.55 61.2 324.75 ;
        RECT  55.8 317.85 57.0 319.05 ;
        RECT  72.0 312.0 73.2 313.95 ;
        RECT  72.0 324.15 73.2 326.1 ;
        RECT  64.8 311.55 66.0 313.95 ;
        RECT  64.8 322.95 66.0 326.55 ;
        RECT  69.6 322.95 70.8 326.55 ;
        RECT  65.4 319.2 66.6 320.4 ;
        RECT  69.6 319.2 70.8 320.4 ;
        RECT  68.4 316.5 69.6 317.7 ;
        RECT  63.0 325.65 77.4 326.55 ;
        RECT  63.0 311.55 77.4 312.45 ;
        RECT  64.8 322.95 66.0 324.15 ;
        RECT  67.2 322.95 68.4 324.15 ;
        RECT  64.8 322.95 66.0 324.15 ;
        RECT  67.2 322.95 68.4 324.15 ;
        RECT  67.2 322.95 68.4 324.15 ;
        RECT  69.6 322.95 70.8 324.15 ;
        RECT  67.2 322.95 68.4 324.15 ;
        RECT  69.6 322.95 70.8 324.15 ;
        RECT  64.8 313.95 66.0 315.15 ;
        RECT  67.2 313.95 68.4 315.15 ;
        RECT  64.8 313.95 66.0 315.15 ;
        RECT  67.2 313.95 68.4 315.15 ;
        RECT  67.2 313.95 68.4 315.15 ;
        RECT  69.6 313.95 70.8 315.15 ;
        RECT  67.2 313.95 68.4 315.15 ;
        RECT  69.6 313.95 70.8 315.15 ;
        RECT  72.0 313.35 73.2 314.55 ;
        RECT  72.0 323.55 73.2 324.75 ;
        RECT  68.4 316.5 69.6 317.7 ;
        RECT  65.4 319.2 66.6 320.4 ;
        RECT  67.2 322.95 68.4 324.15 ;
        RECT  69.6 313.95 70.8 315.15 ;
        RECT  69.6 319.2 70.8 320.4 ;
        RECT  84.0 312.0 85.2 313.95 ;
        RECT  84.0 324.15 85.2 326.1 ;
        RECT  79.2 311.55 80.4 313.35 ;
        RECT  79.2 322.95 80.4 326.55 ;
        RECT  81.9 314.55 82.8 322.95 ;
        RECT  79.8 317.85 81.0 319.05 ;
        RECT  82.35 318.0 83.25 318.9 ;
        RECT  77.4 325.65 87.0 326.55 ;
        RECT  77.4 311.55 87.0 312.45 ;
        RECT  79.2 322.95 80.4 324.15 ;
        RECT  81.6 322.95 82.8 324.15 ;
        RECT  79.2 322.95 80.4 324.15 ;
        RECT  81.6 322.95 82.8 324.15 ;
        RECT  79.2 313.35 80.4 314.55 ;
        RECT  81.6 313.35 82.8 314.55 ;
        RECT  79.2 313.35 80.4 314.55 ;
        RECT  81.6 313.35 82.8 314.55 ;
        RECT  84.0 313.35 85.2 314.55 ;
        RECT  84.0 323.55 85.2 324.75 ;
        RECT  79.8 317.85 81.0 319.05 ;
        RECT  49.65 317.85 50.85 319.05 ;
        RECT  51.6 315.6 52.8 316.8 ;
        RECT  67.2 316.5 68.4 317.7 ;
        RECT  60.0 338.25 61.2 340.2 ;
        RECT  60.0 326.1 61.2 328.05 ;
        RECT  55.2 338.85 56.4 340.65 ;
        RECT  55.2 325.65 56.4 329.25 ;
        RECT  57.9 329.25 58.8 337.65 ;
        RECT  55.8 333.15 57.0 334.35 ;
        RECT  58.35 333.3 59.25 334.2 ;
        RECT  53.4 325.65 63.0 326.55 ;
        RECT  53.4 339.75 63.0 340.65 ;
        RECT  55.2 330.45 56.4 331.65 ;
        RECT  57.6 330.45 58.8 331.65 ;
        RECT  55.2 330.45 56.4 331.65 ;
        RECT  57.6 330.45 58.8 331.65 ;
        RECT  55.2 338.85 56.4 340.05 ;
        RECT  57.6 338.85 58.8 340.05 ;
        RECT  55.2 338.85 56.4 340.05 ;
        RECT  57.6 338.85 58.8 340.05 ;
        RECT  60.0 338.85 61.2 340.05 ;
        RECT  60.0 328.65 61.2 329.85 ;
        RECT  55.8 334.35 57.0 335.55 ;
        RECT  72.0 338.25 73.2 340.2 ;
        RECT  72.0 326.1 73.2 328.05 ;
        RECT  64.8 338.25 66.0 340.65 ;
        RECT  64.8 325.65 66.0 329.25 ;
        RECT  69.6 325.65 70.8 329.25 ;
        RECT  65.4 331.8 66.6 333.0 ;
        RECT  69.6 331.8 70.8 333.0 ;
        RECT  68.4 334.5 69.6 335.7 ;
        RECT  63.0 325.65 77.4 326.55 ;
        RECT  63.0 339.75 77.4 340.65 ;
        RECT  64.8 330.45 66.0 331.65 ;
        RECT  67.2 330.45 68.4 331.65 ;
        RECT  64.8 330.45 66.0 331.65 ;
        RECT  67.2 330.45 68.4 331.65 ;
        RECT  67.2 330.45 68.4 331.65 ;
        RECT  69.6 330.45 70.8 331.65 ;
        RECT  67.2 330.45 68.4 331.65 ;
        RECT  69.6 330.45 70.8 331.65 ;
        RECT  64.8 339.45 66.0 340.65 ;
        RECT  67.2 339.45 68.4 340.65 ;
        RECT  64.8 339.45 66.0 340.65 ;
        RECT  67.2 339.45 68.4 340.65 ;
        RECT  67.2 339.45 68.4 340.65 ;
        RECT  69.6 339.45 70.8 340.65 ;
        RECT  67.2 339.45 68.4 340.65 ;
        RECT  69.6 339.45 70.8 340.65 ;
        RECT  72.0 338.85 73.2 340.05 ;
        RECT  72.0 328.65 73.2 329.85 ;
        RECT  68.4 335.7 69.6 336.9 ;
        RECT  65.4 333.0 66.6 334.2 ;
        RECT  67.2 329.25 68.4 330.45 ;
        RECT  69.6 338.25 70.8 339.45 ;
        RECT  69.6 333.0 70.8 334.2 ;
        RECT  84.0 338.25 85.2 340.2 ;
        RECT  84.0 326.1 85.2 328.05 ;
        RECT  79.2 338.85 80.4 340.65 ;
        RECT  79.2 325.65 80.4 329.25 ;
        RECT  81.9 329.25 82.8 337.65 ;
        RECT  79.8 333.15 81.0 334.35 ;
        RECT  82.35 333.3 83.25 334.2 ;
        RECT  77.4 325.65 87.0 326.55 ;
        RECT  77.4 339.75 87.0 340.65 ;
        RECT  79.2 330.45 80.4 331.65 ;
        RECT  81.6 330.45 82.8 331.65 ;
        RECT  79.2 330.45 80.4 331.65 ;
        RECT  81.6 330.45 82.8 331.65 ;
        RECT  79.2 338.85 80.4 340.05 ;
        RECT  81.6 338.85 82.8 340.05 ;
        RECT  79.2 338.85 80.4 340.05 ;
        RECT  81.6 338.85 82.8 340.05 ;
        RECT  84.0 338.85 85.2 340.05 ;
        RECT  84.0 328.65 85.2 329.85 ;
        RECT  79.8 334.35 81.0 335.55 ;
        RECT  49.65 333.15 50.85 334.35 ;
        RECT  51.6 335.4 52.8 336.6 ;
        RECT  67.2 334.5 68.4 335.7 ;
        RECT  60.0 340.2 61.2 342.15 ;
        RECT  60.0 352.35 61.2 354.3 ;
        RECT  55.2 339.75 56.4 341.55 ;
        RECT  55.2 351.15 56.4 354.75 ;
        RECT  57.9 342.75 58.8 351.15 ;
        RECT  55.8 346.05 57.0 347.25 ;
        RECT  58.35 346.2 59.25 347.1 ;
        RECT  53.4 353.85 63.0 354.75 ;
        RECT  53.4 339.75 63.0 340.65 ;
        RECT  55.2 351.15 56.4 352.35 ;
        RECT  57.6 351.15 58.8 352.35 ;
        RECT  55.2 351.15 56.4 352.35 ;
        RECT  57.6 351.15 58.8 352.35 ;
        RECT  55.2 341.55 56.4 342.75 ;
        RECT  57.6 341.55 58.8 342.75 ;
        RECT  55.2 341.55 56.4 342.75 ;
        RECT  57.6 341.55 58.8 342.75 ;
        RECT  60.0 341.55 61.2 342.75 ;
        RECT  60.0 351.75 61.2 352.95 ;
        RECT  55.8 346.05 57.0 347.25 ;
        RECT  72.0 340.2 73.2 342.15 ;
        RECT  72.0 352.35 73.2 354.3 ;
        RECT  64.8 339.75 66.0 342.15 ;
        RECT  64.8 351.15 66.0 354.75 ;
        RECT  69.6 351.15 70.8 354.75 ;
        RECT  65.4 347.4 66.6 348.6 ;
        RECT  69.6 347.4 70.8 348.6 ;
        RECT  68.4 344.7 69.6 345.9 ;
        RECT  63.0 353.85 77.4 354.75 ;
        RECT  63.0 339.75 77.4 340.65 ;
        RECT  64.8 351.15 66.0 352.35 ;
        RECT  67.2 351.15 68.4 352.35 ;
        RECT  64.8 351.15 66.0 352.35 ;
        RECT  67.2 351.15 68.4 352.35 ;
        RECT  67.2 351.15 68.4 352.35 ;
        RECT  69.6 351.15 70.8 352.35 ;
        RECT  67.2 351.15 68.4 352.35 ;
        RECT  69.6 351.15 70.8 352.35 ;
        RECT  64.8 342.15 66.0 343.35 ;
        RECT  67.2 342.15 68.4 343.35 ;
        RECT  64.8 342.15 66.0 343.35 ;
        RECT  67.2 342.15 68.4 343.35 ;
        RECT  67.2 342.15 68.4 343.35 ;
        RECT  69.6 342.15 70.8 343.35 ;
        RECT  67.2 342.15 68.4 343.35 ;
        RECT  69.6 342.15 70.8 343.35 ;
        RECT  72.0 341.55 73.2 342.75 ;
        RECT  72.0 351.75 73.2 352.95 ;
        RECT  68.4 344.7 69.6 345.9 ;
        RECT  65.4 347.4 66.6 348.6 ;
        RECT  67.2 351.15 68.4 352.35 ;
        RECT  69.6 342.15 70.8 343.35 ;
        RECT  69.6 347.4 70.8 348.6 ;
        RECT  84.0 340.2 85.2 342.15 ;
        RECT  84.0 352.35 85.2 354.3 ;
        RECT  79.2 339.75 80.4 341.55 ;
        RECT  79.2 351.15 80.4 354.75 ;
        RECT  81.9 342.75 82.8 351.15 ;
        RECT  79.8 346.05 81.0 347.25 ;
        RECT  82.35 346.2 83.25 347.1 ;
        RECT  77.4 353.85 87.0 354.75 ;
        RECT  77.4 339.75 87.0 340.65 ;
        RECT  79.2 351.15 80.4 352.35 ;
        RECT  81.6 351.15 82.8 352.35 ;
        RECT  79.2 351.15 80.4 352.35 ;
        RECT  81.6 351.15 82.8 352.35 ;
        RECT  79.2 341.55 80.4 342.75 ;
        RECT  81.6 341.55 82.8 342.75 ;
        RECT  79.2 341.55 80.4 342.75 ;
        RECT  81.6 341.55 82.8 342.75 ;
        RECT  84.0 341.55 85.2 342.75 ;
        RECT  84.0 351.75 85.2 352.95 ;
        RECT  79.8 346.05 81.0 347.25 ;
        RECT  49.65 346.05 50.85 347.25 ;
        RECT  51.6 343.8 52.8 345.0 ;
        RECT  67.2 344.7 68.4 345.9 ;
        RECT  60.0 366.45 61.2 368.4 ;
        RECT  60.0 354.3 61.2 356.25 ;
        RECT  55.2 367.05 56.4 368.85 ;
        RECT  55.2 353.85 56.4 357.45 ;
        RECT  57.9 357.45 58.8 365.85 ;
        RECT  55.8 361.35 57.0 362.55 ;
        RECT  58.35 361.5 59.25 362.4 ;
        RECT  53.4 353.85 63.0 354.75 ;
        RECT  53.4 367.95 63.0 368.85 ;
        RECT  55.2 358.65 56.4 359.85 ;
        RECT  57.6 358.65 58.8 359.85 ;
        RECT  55.2 358.65 56.4 359.85 ;
        RECT  57.6 358.65 58.8 359.85 ;
        RECT  55.2 367.05 56.4 368.25 ;
        RECT  57.6 367.05 58.8 368.25 ;
        RECT  55.2 367.05 56.4 368.25 ;
        RECT  57.6 367.05 58.8 368.25 ;
        RECT  60.0 367.05 61.2 368.25 ;
        RECT  60.0 356.85 61.2 358.05 ;
        RECT  55.8 362.55 57.0 363.75 ;
        RECT  72.0 366.45 73.2 368.4 ;
        RECT  72.0 354.3 73.2 356.25 ;
        RECT  64.8 366.45 66.0 368.85 ;
        RECT  64.8 353.85 66.0 357.45 ;
        RECT  69.6 353.85 70.8 357.45 ;
        RECT  65.4 360.0 66.6 361.2 ;
        RECT  69.6 360.0 70.8 361.2 ;
        RECT  68.4 362.7 69.6 363.9 ;
        RECT  63.0 353.85 77.4 354.75 ;
        RECT  63.0 367.95 77.4 368.85 ;
        RECT  64.8 358.65 66.0 359.85 ;
        RECT  67.2 358.65 68.4 359.85 ;
        RECT  64.8 358.65 66.0 359.85 ;
        RECT  67.2 358.65 68.4 359.85 ;
        RECT  67.2 358.65 68.4 359.85 ;
        RECT  69.6 358.65 70.8 359.85 ;
        RECT  67.2 358.65 68.4 359.85 ;
        RECT  69.6 358.65 70.8 359.85 ;
        RECT  64.8 367.65 66.0 368.85 ;
        RECT  67.2 367.65 68.4 368.85 ;
        RECT  64.8 367.65 66.0 368.85 ;
        RECT  67.2 367.65 68.4 368.85 ;
        RECT  67.2 367.65 68.4 368.85 ;
        RECT  69.6 367.65 70.8 368.85 ;
        RECT  67.2 367.65 68.4 368.85 ;
        RECT  69.6 367.65 70.8 368.85 ;
        RECT  72.0 367.05 73.2 368.25 ;
        RECT  72.0 356.85 73.2 358.05 ;
        RECT  68.4 363.9 69.6 365.1 ;
        RECT  65.4 361.2 66.6 362.4 ;
        RECT  67.2 357.45 68.4 358.65 ;
        RECT  69.6 366.45 70.8 367.65 ;
        RECT  69.6 361.2 70.8 362.4 ;
        RECT  84.0 366.45 85.2 368.4 ;
        RECT  84.0 354.3 85.2 356.25 ;
        RECT  79.2 367.05 80.4 368.85 ;
        RECT  79.2 353.85 80.4 357.45 ;
        RECT  81.9 357.45 82.8 365.85 ;
        RECT  79.8 361.35 81.0 362.55 ;
        RECT  82.35 361.5 83.25 362.4 ;
        RECT  77.4 353.85 87.0 354.75 ;
        RECT  77.4 367.95 87.0 368.85 ;
        RECT  79.2 358.65 80.4 359.85 ;
        RECT  81.6 358.65 82.8 359.85 ;
        RECT  79.2 358.65 80.4 359.85 ;
        RECT  81.6 358.65 82.8 359.85 ;
        RECT  79.2 367.05 80.4 368.25 ;
        RECT  81.6 367.05 82.8 368.25 ;
        RECT  79.2 367.05 80.4 368.25 ;
        RECT  81.6 367.05 82.8 368.25 ;
        RECT  84.0 367.05 85.2 368.25 ;
        RECT  84.0 356.85 85.2 358.05 ;
        RECT  79.8 362.55 81.0 363.75 ;
        RECT  49.65 361.35 50.85 362.55 ;
        RECT  51.6 363.6 52.8 364.8 ;
        RECT  67.2 362.7 68.4 363.9 ;
        RECT  60.0 368.4 61.2 370.35 ;
        RECT  60.0 380.55 61.2 382.5 ;
        RECT  55.2 367.95 56.4 369.75 ;
        RECT  55.2 379.35 56.4 382.95 ;
        RECT  57.9 370.95 58.8 379.35 ;
        RECT  55.8 374.25 57.0 375.45 ;
        RECT  58.35 374.4 59.25 375.3 ;
        RECT  53.4 382.05 63.0 382.95 ;
        RECT  53.4 367.95 63.0 368.85 ;
        RECT  55.2 379.35 56.4 380.55 ;
        RECT  57.6 379.35 58.8 380.55 ;
        RECT  55.2 379.35 56.4 380.55 ;
        RECT  57.6 379.35 58.8 380.55 ;
        RECT  55.2 369.75 56.4 370.95 ;
        RECT  57.6 369.75 58.8 370.95 ;
        RECT  55.2 369.75 56.4 370.95 ;
        RECT  57.6 369.75 58.8 370.95 ;
        RECT  60.0 369.75 61.2 370.95 ;
        RECT  60.0 379.95 61.2 381.15 ;
        RECT  55.8 374.25 57.0 375.45 ;
        RECT  72.0 368.4 73.2 370.35 ;
        RECT  72.0 380.55 73.2 382.5 ;
        RECT  64.8 367.95 66.0 370.35 ;
        RECT  64.8 379.35 66.0 382.95 ;
        RECT  69.6 379.35 70.8 382.95 ;
        RECT  65.4 375.6 66.6 376.8 ;
        RECT  69.6 375.6 70.8 376.8 ;
        RECT  68.4 372.9 69.6 374.1 ;
        RECT  63.0 382.05 77.4 382.95 ;
        RECT  63.0 367.95 77.4 368.85 ;
        RECT  64.8 379.35 66.0 380.55 ;
        RECT  67.2 379.35 68.4 380.55 ;
        RECT  64.8 379.35 66.0 380.55 ;
        RECT  67.2 379.35 68.4 380.55 ;
        RECT  67.2 379.35 68.4 380.55 ;
        RECT  69.6 379.35 70.8 380.55 ;
        RECT  67.2 379.35 68.4 380.55 ;
        RECT  69.6 379.35 70.8 380.55 ;
        RECT  64.8 370.35 66.0 371.55 ;
        RECT  67.2 370.35 68.4 371.55 ;
        RECT  64.8 370.35 66.0 371.55 ;
        RECT  67.2 370.35 68.4 371.55 ;
        RECT  67.2 370.35 68.4 371.55 ;
        RECT  69.6 370.35 70.8 371.55 ;
        RECT  67.2 370.35 68.4 371.55 ;
        RECT  69.6 370.35 70.8 371.55 ;
        RECT  72.0 369.75 73.2 370.95 ;
        RECT  72.0 379.95 73.2 381.15 ;
        RECT  68.4 372.9 69.6 374.1 ;
        RECT  65.4 375.6 66.6 376.8 ;
        RECT  67.2 379.35 68.4 380.55 ;
        RECT  69.6 370.35 70.8 371.55 ;
        RECT  69.6 375.6 70.8 376.8 ;
        RECT  84.0 368.4 85.2 370.35 ;
        RECT  84.0 380.55 85.2 382.5 ;
        RECT  79.2 367.95 80.4 369.75 ;
        RECT  79.2 379.35 80.4 382.95 ;
        RECT  81.9 370.95 82.8 379.35 ;
        RECT  79.8 374.25 81.0 375.45 ;
        RECT  82.35 374.4 83.25 375.3 ;
        RECT  77.4 382.05 87.0 382.95 ;
        RECT  77.4 367.95 87.0 368.85 ;
        RECT  79.2 379.35 80.4 380.55 ;
        RECT  81.6 379.35 82.8 380.55 ;
        RECT  79.2 379.35 80.4 380.55 ;
        RECT  81.6 379.35 82.8 380.55 ;
        RECT  79.2 369.75 80.4 370.95 ;
        RECT  81.6 369.75 82.8 370.95 ;
        RECT  79.2 369.75 80.4 370.95 ;
        RECT  81.6 369.75 82.8 370.95 ;
        RECT  84.0 369.75 85.2 370.95 ;
        RECT  84.0 379.95 85.2 381.15 ;
        RECT  79.8 374.25 81.0 375.45 ;
        RECT  49.65 374.25 50.85 375.45 ;
        RECT  51.6 372.0 52.8 373.2 ;
        RECT  67.2 372.9 68.4 374.1 ;
        RECT  60.0 394.65 61.2 396.6 ;
        RECT  60.0 382.5 61.2 384.45 ;
        RECT  55.2 395.25 56.4 397.05 ;
        RECT  55.2 382.05 56.4 385.65 ;
        RECT  57.9 385.65 58.8 394.05 ;
        RECT  55.8 389.55 57.0 390.75 ;
        RECT  58.35 389.7 59.25 390.6 ;
        RECT  53.4 382.05 63.0 382.95 ;
        RECT  53.4 396.15 63.0 397.05 ;
        RECT  55.2 386.85 56.4 388.05 ;
        RECT  57.6 386.85 58.8 388.05 ;
        RECT  55.2 386.85 56.4 388.05 ;
        RECT  57.6 386.85 58.8 388.05 ;
        RECT  55.2 395.25 56.4 396.45 ;
        RECT  57.6 395.25 58.8 396.45 ;
        RECT  55.2 395.25 56.4 396.45 ;
        RECT  57.6 395.25 58.8 396.45 ;
        RECT  60.0 395.25 61.2 396.45 ;
        RECT  60.0 385.05 61.2 386.25 ;
        RECT  55.8 390.75 57.0 391.95 ;
        RECT  72.0 394.65 73.2 396.6 ;
        RECT  72.0 382.5 73.2 384.45 ;
        RECT  64.8 394.65 66.0 397.05 ;
        RECT  64.8 382.05 66.0 385.65 ;
        RECT  69.6 382.05 70.8 385.65 ;
        RECT  65.4 388.2 66.6 389.4 ;
        RECT  69.6 388.2 70.8 389.4 ;
        RECT  68.4 390.9 69.6 392.1 ;
        RECT  63.0 382.05 77.4 382.95 ;
        RECT  63.0 396.15 77.4 397.05 ;
        RECT  64.8 386.85 66.0 388.05 ;
        RECT  67.2 386.85 68.4 388.05 ;
        RECT  64.8 386.85 66.0 388.05 ;
        RECT  67.2 386.85 68.4 388.05 ;
        RECT  67.2 386.85 68.4 388.05 ;
        RECT  69.6 386.85 70.8 388.05 ;
        RECT  67.2 386.85 68.4 388.05 ;
        RECT  69.6 386.85 70.8 388.05 ;
        RECT  64.8 395.85 66.0 397.05 ;
        RECT  67.2 395.85 68.4 397.05 ;
        RECT  64.8 395.85 66.0 397.05 ;
        RECT  67.2 395.85 68.4 397.05 ;
        RECT  67.2 395.85 68.4 397.05 ;
        RECT  69.6 395.85 70.8 397.05 ;
        RECT  67.2 395.85 68.4 397.05 ;
        RECT  69.6 395.85 70.8 397.05 ;
        RECT  72.0 395.25 73.2 396.45 ;
        RECT  72.0 385.05 73.2 386.25 ;
        RECT  68.4 392.1 69.6 393.3 ;
        RECT  65.4 389.4 66.6 390.6 ;
        RECT  67.2 385.65 68.4 386.85 ;
        RECT  69.6 394.65 70.8 395.85 ;
        RECT  69.6 389.4 70.8 390.6 ;
        RECT  84.0 394.65 85.2 396.6 ;
        RECT  84.0 382.5 85.2 384.45 ;
        RECT  79.2 395.25 80.4 397.05 ;
        RECT  79.2 382.05 80.4 385.65 ;
        RECT  81.9 385.65 82.8 394.05 ;
        RECT  79.8 389.55 81.0 390.75 ;
        RECT  82.35 389.7 83.25 390.6 ;
        RECT  77.4 382.05 87.0 382.95 ;
        RECT  77.4 396.15 87.0 397.05 ;
        RECT  79.2 386.85 80.4 388.05 ;
        RECT  81.6 386.85 82.8 388.05 ;
        RECT  79.2 386.85 80.4 388.05 ;
        RECT  81.6 386.85 82.8 388.05 ;
        RECT  79.2 395.25 80.4 396.45 ;
        RECT  81.6 395.25 82.8 396.45 ;
        RECT  79.2 395.25 80.4 396.45 ;
        RECT  81.6 395.25 82.8 396.45 ;
        RECT  84.0 395.25 85.2 396.45 ;
        RECT  84.0 385.05 85.2 386.25 ;
        RECT  79.8 390.75 81.0 391.95 ;
        RECT  49.65 389.55 50.85 390.75 ;
        RECT  51.6 391.8 52.8 393.0 ;
        RECT  67.2 390.9 68.4 392.1 ;
        RECT  60.0 396.6 61.2 398.55 ;
        RECT  60.0 408.75 61.2 410.7 ;
        RECT  55.2 396.15 56.4 397.95 ;
        RECT  55.2 407.55 56.4 411.15 ;
        RECT  57.9 399.15 58.8 407.55 ;
        RECT  55.8 402.45 57.0 403.65 ;
        RECT  58.35 402.6 59.25 403.5 ;
        RECT  53.4 410.25 63.0 411.15 ;
        RECT  53.4 396.15 63.0 397.05 ;
        RECT  55.2 407.55 56.4 408.75 ;
        RECT  57.6 407.55 58.8 408.75 ;
        RECT  55.2 407.55 56.4 408.75 ;
        RECT  57.6 407.55 58.8 408.75 ;
        RECT  55.2 397.95 56.4 399.15 ;
        RECT  57.6 397.95 58.8 399.15 ;
        RECT  55.2 397.95 56.4 399.15 ;
        RECT  57.6 397.95 58.8 399.15 ;
        RECT  60.0 397.95 61.2 399.15 ;
        RECT  60.0 408.15 61.2 409.35 ;
        RECT  55.8 402.45 57.0 403.65 ;
        RECT  72.0 396.6 73.2 398.55 ;
        RECT  72.0 408.75 73.2 410.7 ;
        RECT  64.8 396.15 66.0 398.55 ;
        RECT  64.8 407.55 66.0 411.15 ;
        RECT  69.6 407.55 70.8 411.15 ;
        RECT  65.4 403.8 66.6 405.0 ;
        RECT  69.6 403.8 70.8 405.0 ;
        RECT  68.4 401.1 69.6 402.3 ;
        RECT  63.0 410.25 77.4 411.15 ;
        RECT  63.0 396.15 77.4 397.05 ;
        RECT  64.8 407.55 66.0 408.75 ;
        RECT  67.2 407.55 68.4 408.75 ;
        RECT  64.8 407.55 66.0 408.75 ;
        RECT  67.2 407.55 68.4 408.75 ;
        RECT  67.2 407.55 68.4 408.75 ;
        RECT  69.6 407.55 70.8 408.75 ;
        RECT  67.2 407.55 68.4 408.75 ;
        RECT  69.6 407.55 70.8 408.75 ;
        RECT  64.8 398.55 66.0 399.75 ;
        RECT  67.2 398.55 68.4 399.75 ;
        RECT  64.8 398.55 66.0 399.75 ;
        RECT  67.2 398.55 68.4 399.75 ;
        RECT  67.2 398.55 68.4 399.75 ;
        RECT  69.6 398.55 70.8 399.75 ;
        RECT  67.2 398.55 68.4 399.75 ;
        RECT  69.6 398.55 70.8 399.75 ;
        RECT  72.0 397.95 73.2 399.15 ;
        RECT  72.0 408.15 73.2 409.35 ;
        RECT  68.4 401.1 69.6 402.3 ;
        RECT  65.4 403.8 66.6 405.0 ;
        RECT  67.2 407.55 68.4 408.75 ;
        RECT  69.6 398.55 70.8 399.75 ;
        RECT  69.6 403.8 70.8 405.0 ;
        RECT  84.0 396.6 85.2 398.55 ;
        RECT  84.0 408.75 85.2 410.7 ;
        RECT  79.2 396.15 80.4 397.95 ;
        RECT  79.2 407.55 80.4 411.15 ;
        RECT  81.9 399.15 82.8 407.55 ;
        RECT  79.8 402.45 81.0 403.65 ;
        RECT  82.35 402.6 83.25 403.5 ;
        RECT  77.4 410.25 87.0 411.15 ;
        RECT  77.4 396.15 87.0 397.05 ;
        RECT  79.2 407.55 80.4 408.75 ;
        RECT  81.6 407.55 82.8 408.75 ;
        RECT  79.2 407.55 80.4 408.75 ;
        RECT  81.6 407.55 82.8 408.75 ;
        RECT  79.2 397.95 80.4 399.15 ;
        RECT  81.6 397.95 82.8 399.15 ;
        RECT  79.2 397.95 80.4 399.15 ;
        RECT  81.6 397.95 82.8 399.15 ;
        RECT  84.0 397.95 85.2 399.15 ;
        RECT  84.0 408.15 85.2 409.35 ;
        RECT  79.8 402.45 81.0 403.65 ;
        RECT  49.65 402.45 50.85 403.65 ;
        RECT  51.6 400.2 52.8 401.4 ;
        RECT  67.2 401.1 68.4 402.3 ;
        RECT  60.0 422.85 61.2 424.8 ;
        RECT  60.0 410.7 61.2 412.65 ;
        RECT  55.2 423.45 56.4 425.25 ;
        RECT  55.2 410.25 56.4 413.85 ;
        RECT  57.9 413.85 58.8 422.25 ;
        RECT  55.8 417.75 57.0 418.95 ;
        RECT  58.35 417.9 59.25 418.8 ;
        RECT  53.4 410.25 63.0 411.15 ;
        RECT  53.4 424.35 63.0 425.25 ;
        RECT  55.2 415.05 56.4 416.25 ;
        RECT  57.6 415.05 58.8 416.25 ;
        RECT  55.2 415.05 56.4 416.25 ;
        RECT  57.6 415.05 58.8 416.25 ;
        RECT  55.2 423.45 56.4 424.65 ;
        RECT  57.6 423.45 58.8 424.65 ;
        RECT  55.2 423.45 56.4 424.65 ;
        RECT  57.6 423.45 58.8 424.65 ;
        RECT  60.0 423.45 61.2 424.65 ;
        RECT  60.0 413.25 61.2 414.45 ;
        RECT  55.8 418.95 57.0 420.15 ;
        RECT  72.0 422.85 73.2 424.8 ;
        RECT  72.0 410.7 73.2 412.65 ;
        RECT  64.8 422.85 66.0 425.25 ;
        RECT  64.8 410.25 66.0 413.85 ;
        RECT  69.6 410.25 70.8 413.85 ;
        RECT  65.4 416.4 66.6 417.6 ;
        RECT  69.6 416.4 70.8 417.6 ;
        RECT  68.4 419.1 69.6 420.3 ;
        RECT  63.0 410.25 77.4 411.15 ;
        RECT  63.0 424.35 77.4 425.25 ;
        RECT  64.8 415.05 66.0 416.25 ;
        RECT  67.2 415.05 68.4 416.25 ;
        RECT  64.8 415.05 66.0 416.25 ;
        RECT  67.2 415.05 68.4 416.25 ;
        RECT  67.2 415.05 68.4 416.25 ;
        RECT  69.6 415.05 70.8 416.25 ;
        RECT  67.2 415.05 68.4 416.25 ;
        RECT  69.6 415.05 70.8 416.25 ;
        RECT  64.8 424.05 66.0 425.25 ;
        RECT  67.2 424.05 68.4 425.25 ;
        RECT  64.8 424.05 66.0 425.25 ;
        RECT  67.2 424.05 68.4 425.25 ;
        RECT  67.2 424.05 68.4 425.25 ;
        RECT  69.6 424.05 70.8 425.25 ;
        RECT  67.2 424.05 68.4 425.25 ;
        RECT  69.6 424.05 70.8 425.25 ;
        RECT  72.0 423.45 73.2 424.65 ;
        RECT  72.0 413.25 73.2 414.45 ;
        RECT  68.4 420.3 69.6 421.5 ;
        RECT  65.4 417.6 66.6 418.8 ;
        RECT  67.2 413.85 68.4 415.05 ;
        RECT  69.6 422.85 70.8 424.05 ;
        RECT  69.6 417.6 70.8 418.8 ;
        RECT  84.0 422.85 85.2 424.8 ;
        RECT  84.0 410.7 85.2 412.65 ;
        RECT  79.2 423.45 80.4 425.25 ;
        RECT  79.2 410.25 80.4 413.85 ;
        RECT  81.9 413.85 82.8 422.25 ;
        RECT  79.8 417.75 81.0 418.95 ;
        RECT  82.35 417.9 83.25 418.8 ;
        RECT  77.4 410.25 87.0 411.15 ;
        RECT  77.4 424.35 87.0 425.25 ;
        RECT  79.2 415.05 80.4 416.25 ;
        RECT  81.6 415.05 82.8 416.25 ;
        RECT  79.2 415.05 80.4 416.25 ;
        RECT  81.6 415.05 82.8 416.25 ;
        RECT  79.2 423.45 80.4 424.65 ;
        RECT  81.6 423.45 82.8 424.65 ;
        RECT  79.2 423.45 80.4 424.65 ;
        RECT  81.6 423.45 82.8 424.65 ;
        RECT  84.0 423.45 85.2 424.65 ;
        RECT  84.0 413.25 85.2 414.45 ;
        RECT  79.8 418.95 81.0 420.15 ;
        RECT  49.65 417.75 50.85 418.95 ;
        RECT  51.6 420.0 52.8 421.2 ;
        RECT  67.2 419.1 68.4 420.3 ;
        RECT  8.7 40.2 9.6 81.0 ;
        RECT  62.7 40.2 63.6 81.0 ;
        RECT  62.7 70.2 63.6 81.6 ;
        RECT  59.4 80.4 62.7 81.6 ;
        RECT  60.9 72.6 61.8 79.2 ;
        RECT  60.6 76.2 60.9 79.2 ;
        RECT  60.6 72.6 60.9 73.8 ;
        RECT  58.2 77.4 59.4 81.6 ;
        RECT  58.2 70.2 59.4 73.8 ;
        RECT  54.6 80.4 58.2 81.6 ;
        RECT  57.3 75.0 58.2 76.2 ;
        RECT  57.0 73.8 57.3 76.2 ;
        RECT  56.1 72.6 57.0 79.2 ;
        RECT  55.8 77.4 56.1 79.2 ;
        RECT  55.8 72.6 56.1 73.8 ;
        RECT  53.4 77.4 54.6 81.6 ;
        RECT  39.6 80.4 53.4 81.6 ;
        RECT  52.8 74.7 55.2 75.9 ;
        RECT  54.6 70.2 58.2 71.1 ;
        RECT  53.4 70.2 54.6 73.8 ;
        RECT  52.2 70.2 53.4 71.4 ;
        RECT  49.8 78.0 51.0 79.2 ;
        RECT  50.7 74.7 51.9 77.1 ;
        RECT  48.9 72.6 49.8 79.2 ;
        RECT  48.6 77.4 48.9 79.2 ;
        RECT  48.6 72.6 48.9 73.8 ;
        RECT  46.5 72.6 47.4 79.2 ;
        RECT  46.2 77.4 46.5 79.2 ;
        RECT  46.2 72.6 46.5 75.0 ;
        RECT  44.1 72.6 45.0 79.2 ;
        RECT  43.8 77.4 44.1 79.2 ;
        RECT  43.8 72.6 44.1 75.0 ;
        RECT  42.0 75.0 42.9 76.2 ;
        RECT  41.1 72.6 42.0 79.2 ;
        RECT  40.8 76.2 41.1 79.2 ;
        RECT  40.8 72.6 41.1 73.8 ;
        RECT  38.4 77.4 39.6 81.6 ;
        RECT  33.9 80.4 38.4 81.6 ;
        RECT  37.5 75.3 39.9 76.5 ;
        RECT  39.6 70.2 52.2 71.1 ;
        RECT  38.4 70.2 39.6 73.8 ;
        RECT  36.3 78.0 37.5 79.2 ;
        RECT  35.4 72.6 36.3 79.2 ;
        RECT  35.1 77.4 35.4 79.2 ;
        RECT  35.1 72.6 35.4 73.8 ;
        RECT  33.9 70.2 38.4 71.1 ;
        RECT  32.7 77.4 33.9 81.6 ;
        RECT  29.1 80.4 32.7 81.6 ;
        RECT  31.8 74.7 33.0 75.9 ;
        RECT  32.7 70.2 33.9 73.8 ;
        RECT  31.5 73.8 31.8 79.2 ;
        RECT  30.9 72.6 31.5 79.2 ;
        RECT  30.3 77.4 30.9 79.2 ;
        RECT  30.6 72.6 30.9 75.0 ;
        RECT  30.3 72.6 30.6 73.8 ;
        RECT  27.9 77.4 29.1 81.6 ;
        RECT  12.9 80.4 27.9 81.6 ;
        RECT  27.3 74.7 29.7 75.9 ;
        RECT  29.1 70.2 32.7 71.1 ;
        RECT  27.9 70.2 29.1 73.8 ;
        RECT  26.7 70.2 27.9 71.4 ;
        RECT  23.4 78.0 24.6 79.2 ;
        RECT  24.3 74.7 25.5 77.1 ;
        RECT  22.5 72.6 23.4 79.2 ;
        RECT  22.2 77.4 22.5 79.2 ;
        RECT  22.2 72.6 22.5 73.8 ;
        RECT  20.1 72.6 21.0 79.2 ;
        RECT  19.8 77.4 20.1 79.2 ;
        RECT  19.8 72.6 20.1 75.0 ;
        RECT  17.7 72.6 18.6 79.2 ;
        RECT  17.4 77.4 17.7 79.2 ;
        RECT  17.4 72.6 17.7 75.0 ;
        RECT  15.6 75.0 16.5 76.2 ;
        RECT  14.7 72.6 15.6 79.2 ;
        RECT  14.4 76.2 14.7 79.2 ;
        RECT  14.4 72.6 14.7 73.8 ;
        RECT  13.2 70.2 26.7 71.1 ;
        RECT  12.9 77.4 13.2 79.2 ;
        RECT  12.0 77.4 12.9 81.6 ;
        RECT  12.3 70.2 13.2 73.8 ;
        RECT  12.0 72.6 12.3 73.8 ;
        RECT  10.5 77.4 12.0 78.6 ;
        RECT  9.6 75.3 10.5 76.5 ;
        RECT  8.7 70.2 9.6 81.6 ;
        RECT  8.7 70.2 9.6 81.6 ;
        RECT  62.7 70.2 63.6 81.6 ;
        RECT  62.7 60.0 63.6 71.4 ;
        RECT  59.4 60.0 62.7 61.2 ;
        RECT  60.9 62.4 61.8 69.0 ;
        RECT  60.6 62.4 60.9 65.4 ;
        RECT  60.6 67.8 60.9 69.0 ;
        RECT  58.2 60.0 59.4 64.2 ;
        RECT  58.2 67.8 59.4 71.4 ;
        RECT  54.6 60.0 58.2 61.2 ;
        RECT  57.3 65.4 58.2 66.6 ;
        RECT  57.0 65.4 57.3 67.8 ;
        RECT  56.1 62.4 57.0 69.0 ;
        RECT  55.8 62.4 56.1 64.2 ;
        RECT  55.8 67.8 56.1 69.0 ;
        RECT  53.4 60.0 54.6 64.2 ;
        RECT  39.6 60.0 53.4 61.2 ;
        RECT  52.8 65.7 55.2 66.9 ;
        RECT  54.6 70.5 58.2 71.4 ;
        RECT  53.4 67.8 54.6 71.4 ;
        RECT  52.2 70.2 53.4 71.4 ;
        RECT  49.8 62.4 51.0 63.6 ;
        RECT  50.7 64.5 51.9 66.9 ;
        RECT  48.9 62.4 49.8 69.0 ;
        RECT  48.6 62.4 48.9 64.2 ;
        RECT  48.6 67.8 48.9 69.0 ;
        RECT  46.5 62.4 47.4 69.0 ;
        RECT  46.2 62.4 46.5 64.2 ;
        RECT  46.2 66.6 46.5 69.0 ;
        RECT  44.1 62.4 45.0 69.0 ;
        RECT  43.8 62.4 44.1 64.2 ;
        RECT  43.8 66.6 44.1 69.0 ;
        RECT  42.0 65.4 42.9 66.6 ;
        RECT  41.1 62.4 42.0 69.0 ;
        RECT  40.8 62.4 41.1 65.4 ;
        RECT  40.8 67.8 41.1 69.0 ;
        RECT  38.4 60.0 39.6 64.2 ;
        RECT  33.9 60.0 38.4 61.2 ;
        RECT  37.5 65.1 39.9 66.3 ;
        RECT  39.6 70.5 52.2 71.4 ;
        RECT  38.4 67.8 39.6 71.4 ;
        RECT  36.3 62.4 37.5 63.6 ;
        RECT  35.4 62.4 36.3 69.0 ;
        RECT  35.1 62.4 35.4 64.2 ;
        RECT  35.1 67.8 35.4 69.0 ;
        RECT  33.9 70.5 38.4 71.4 ;
        RECT  32.7 60.0 33.9 64.2 ;
        RECT  29.1 60.0 32.7 61.2 ;
        RECT  31.8 65.7 33.0 66.9 ;
        RECT  32.7 67.8 33.9 71.4 ;
        RECT  31.5 62.4 31.8 67.8 ;
        RECT  30.9 62.4 31.5 69.0 ;
        RECT  30.3 62.4 30.9 64.2 ;
        RECT  30.6 66.6 30.9 69.0 ;
        RECT  30.3 67.8 30.6 69.0 ;
        RECT  27.9 60.0 29.1 64.2 ;
        RECT  12.9 60.0 27.9 61.2 ;
        RECT  27.3 65.7 29.7 66.9 ;
        RECT  29.1 70.5 32.7 71.4 ;
        RECT  27.9 67.8 29.1 71.4 ;
        RECT  26.7 70.2 27.9 71.4 ;
        RECT  23.4 62.4 24.6 63.6 ;
        RECT  24.3 64.5 25.5 66.9 ;
        RECT  22.5 62.4 23.4 69.0 ;
        RECT  22.2 62.4 22.5 64.2 ;
        RECT  22.2 67.8 22.5 69.0 ;
        RECT  20.1 62.4 21.0 69.0 ;
        RECT  19.8 62.4 20.1 64.2 ;
        RECT  19.8 66.6 20.1 69.0 ;
        RECT  17.7 62.4 18.6 69.0 ;
        RECT  17.4 62.4 17.7 64.2 ;
        RECT  17.4 66.6 17.7 69.0 ;
        RECT  15.6 65.4 16.5 66.6 ;
        RECT  14.7 62.4 15.6 69.0 ;
        RECT  14.4 62.4 14.7 65.4 ;
        RECT  14.4 67.8 14.7 69.0 ;
        RECT  13.2 70.5 26.7 71.4 ;
        RECT  12.9 62.4 13.2 64.2 ;
        RECT  12.0 60.0 12.9 64.2 ;
        RECT  12.3 67.8 13.2 71.4 ;
        RECT  12.0 67.8 12.3 69.0 ;
        RECT  10.5 63.0 12.0 64.2 ;
        RECT  9.6 65.1 10.5 66.3 ;
        RECT  8.7 60.0 9.6 71.4 ;
        RECT  8.7 60.0 9.6 71.4 ;
        RECT  62.7 60.0 63.6 71.4 ;
        RECT  62.7 49.8 63.6 61.2 ;
        RECT  59.4 60.0 62.7 61.2 ;
        RECT  60.9 52.2 61.8 58.8 ;
        RECT  60.6 55.8 60.9 58.8 ;
        RECT  60.6 52.2 60.9 53.4 ;
        RECT  58.2 57.0 59.4 61.2 ;
        RECT  58.2 49.8 59.4 53.4 ;
        RECT  54.6 60.0 58.2 61.2 ;
        RECT  57.3 54.6 58.2 55.8 ;
        RECT  57.0 53.4 57.3 55.8 ;
        RECT  56.1 52.2 57.0 58.8 ;
        RECT  55.8 57.0 56.1 58.8 ;
        RECT  55.8 52.2 56.1 53.4 ;
        RECT  53.4 57.0 54.6 61.2 ;
        RECT  39.6 60.0 53.4 61.2 ;
        RECT  52.8 54.3 55.2 55.5 ;
        RECT  54.6 49.8 58.2 50.7 ;
        RECT  53.4 49.8 54.6 53.4 ;
        RECT  52.2 49.8 53.4 51.0 ;
        RECT  49.8 57.6 51.0 58.8 ;
        RECT  50.7 54.3 51.9 56.7 ;
        RECT  48.9 52.2 49.8 58.8 ;
        RECT  48.6 57.0 48.9 58.8 ;
        RECT  48.6 52.2 48.9 53.4 ;
        RECT  46.5 52.2 47.4 58.8 ;
        RECT  46.2 57.0 46.5 58.8 ;
        RECT  46.2 52.2 46.5 54.6 ;
        RECT  44.1 52.2 45.0 58.8 ;
        RECT  43.8 57.0 44.1 58.8 ;
        RECT  43.8 52.2 44.1 54.6 ;
        RECT  42.0 54.6 42.9 55.8 ;
        RECT  41.1 52.2 42.0 58.8 ;
        RECT  40.8 55.8 41.1 58.8 ;
        RECT  40.8 52.2 41.1 53.4 ;
        RECT  38.4 57.0 39.6 61.2 ;
        RECT  33.9 60.0 38.4 61.2 ;
        RECT  37.5 54.9 39.9 56.1 ;
        RECT  39.6 49.8 52.2 50.7 ;
        RECT  38.4 49.8 39.6 53.4 ;
        RECT  36.3 57.6 37.5 58.8 ;
        RECT  35.4 52.2 36.3 58.8 ;
        RECT  35.1 57.0 35.4 58.8 ;
        RECT  35.1 52.2 35.4 53.4 ;
        RECT  33.9 49.8 38.4 50.7 ;
        RECT  32.7 57.0 33.9 61.2 ;
        RECT  29.1 60.0 32.7 61.2 ;
        RECT  31.8 54.3 33.0 55.5 ;
        RECT  32.7 49.8 33.9 53.4 ;
        RECT  31.5 53.4 31.8 58.8 ;
        RECT  30.9 52.2 31.5 58.8 ;
        RECT  30.3 57.0 30.9 58.8 ;
        RECT  30.6 52.2 30.9 54.6 ;
        RECT  30.3 52.2 30.6 53.4 ;
        RECT  27.9 57.0 29.1 61.2 ;
        RECT  12.9 60.0 27.9 61.2 ;
        RECT  27.3 54.3 29.7 55.5 ;
        RECT  29.1 49.8 32.7 50.7 ;
        RECT  27.9 49.8 29.1 53.4 ;
        RECT  26.7 49.8 27.9 51.0 ;
        RECT  23.4 57.6 24.6 58.8 ;
        RECT  24.3 54.3 25.5 56.7 ;
        RECT  22.5 52.2 23.4 58.8 ;
        RECT  22.2 57.0 22.5 58.8 ;
        RECT  22.2 52.2 22.5 53.4 ;
        RECT  20.1 52.2 21.0 58.8 ;
        RECT  19.8 57.0 20.1 58.8 ;
        RECT  19.8 52.2 20.1 54.6 ;
        RECT  17.7 52.2 18.6 58.8 ;
        RECT  17.4 57.0 17.7 58.8 ;
        RECT  17.4 52.2 17.7 54.6 ;
        RECT  15.6 54.6 16.5 55.8 ;
        RECT  14.7 52.2 15.6 58.8 ;
        RECT  14.4 55.8 14.7 58.8 ;
        RECT  14.4 52.2 14.7 53.4 ;
        RECT  13.2 49.8 26.7 50.7 ;
        RECT  12.9 57.0 13.2 58.8 ;
        RECT  12.0 57.0 12.9 61.2 ;
        RECT  12.3 49.8 13.2 53.4 ;
        RECT  12.0 52.2 12.3 53.4 ;
        RECT  10.5 57.0 12.0 58.2 ;
        RECT  9.6 54.9 10.5 56.1 ;
        RECT  8.7 49.8 9.6 61.2 ;
        RECT  8.7 49.8 9.6 61.2 ;
        RECT  62.7 49.8 63.6 61.2 ;
        RECT  62.7 39.6 63.6 51.0 ;
        RECT  59.4 39.6 62.7 40.8 ;
        RECT  60.9 42.0 61.8 48.6 ;
        RECT  60.6 42.0 60.9 45.0 ;
        RECT  60.6 47.4 60.9 48.6 ;
        RECT  58.2 39.6 59.4 43.8 ;
        RECT  58.2 47.4 59.4 51.0 ;
        RECT  54.6 39.6 58.2 40.8 ;
        RECT  57.3 45.0 58.2 46.2 ;
        RECT  57.0 45.0 57.3 47.4 ;
        RECT  56.1 42.0 57.0 48.6 ;
        RECT  55.8 42.0 56.1 43.8 ;
        RECT  55.8 47.4 56.1 48.6 ;
        RECT  53.4 39.6 54.6 43.8 ;
        RECT  39.6 39.6 53.4 40.8 ;
        RECT  52.8 45.3 55.2 46.5 ;
        RECT  54.6 50.1 58.2 51.0 ;
        RECT  53.4 47.4 54.6 51.0 ;
        RECT  52.2 49.8 53.4 51.0 ;
        RECT  49.8 42.0 51.0 43.2 ;
        RECT  50.7 44.1 51.9 46.5 ;
        RECT  48.9 42.0 49.8 48.6 ;
        RECT  48.6 42.0 48.9 43.8 ;
        RECT  48.6 47.4 48.9 48.6 ;
        RECT  46.5 42.0 47.4 48.6 ;
        RECT  46.2 42.0 46.5 43.8 ;
        RECT  46.2 46.2 46.5 48.6 ;
        RECT  44.1 42.0 45.0 48.6 ;
        RECT  43.8 42.0 44.1 43.8 ;
        RECT  43.8 46.2 44.1 48.6 ;
        RECT  42.0 45.0 42.9 46.2 ;
        RECT  41.1 42.0 42.0 48.6 ;
        RECT  40.8 42.0 41.1 45.0 ;
        RECT  40.8 47.4 41.1 48.6 ;
        RECT  38.4 39.6 39.6 43.8 ;
        RECT  33.9 39.6 38.4 40.8 ;
        RECT  37.5 44.7 39.9 45.9 ;
        RECT  39.6 50.1 52.2 51.0 ;
        RECT  38.4 47.4 39.6 51.0 ;
        RECT  36.3 42.0 37.5 43.2 ;
        RECT  35.4 42.0 36.3 48.6 ;
        RECT  35.1 42.0 35.4 43.8 ;
        RECT  35.1 47.4 35.4 48.6 ;
        RECT  33.9 50.1 38.4 51.0 ;
        RECT  32.7 39.6 33.9 43.8 ;
        RECT  29.1 39.6 32.7 40.8 ;
        RECT  31.8 45.3 33.0 46.5 ;
        RECT  32.7 47.4 33.9 51.0 ;
        RECT  31.5 42.0 31.8 47.4 ;
        RECT  30.9 42.0 31.5 48.6 ;
        RECT  30.3 42.0 30.9 43.8 ;
        RECT  30.6 46.2 30.9 48.6 ;
        RECT  30.3 47.4 30.6 48.6 ;
        RECT  27.9 39.6 29.1 43.8 ;
        RECT  12.9 39.6 27.9 40.8 ;
        RECT  27.3 45.3 29.7 46.5 ;
        RECT  29.1 50.1 32.7 51.0 ;
        RECT  27.9 47.4 29.1 51.0 ;
        RECT  26.7 49.8 27.9 51.0 ;
        RECT  23.4 42.0 24.6 43.2 ;
        RECT  24.3 44.1 25.5 46.5 ;
        RECT  22.5 42.0 23.4 48.6 ;
        RECT  22.2 42.0 22.5 43.8 ;
        RECT  22.2 47.4 22.5 48.6 ;
        RECT  20.1 42.0 21.0 48.6 ;
        RECT  19.8 42.0 20.1 43.8 ;
        RECT  19.8 46.2 20.1 48.6 ;
        RECT  17.7 42.0 18.6 48.6 ;
        RECT  17.4 42.0 17.7 43.8 ;
        RECT  17.4 46.2 17.7 48.6 ;
        RECT  15.6 45.0 16.5 46.2 ;
        RECT  14.7 42.0 15.6 48.6 ;
        RECT  14.4 42.0 14.7 45.0 ;
        RECT  14.4 47.4 14.7 48.6 ;
        RECT  13.2 50.1 26.7 51.0 ;
        RECT  12.9 42.0 13.2 43.8 ;
        RECT  12.0 39.6 12.9 43.8 ;
        RECT  12.3 47.4 13.2 51.0 ;
        RECT  12.0 47.4 12.3 48.6 ;
        RECT  10.5 42.6 12.0 43.8 ;
        RECT  9.6 44.7 10.5 45.9 ;
        RECT  8.7 39.6 9.6 51.0 ;
        RECT  8.7 39.6 9.6 51.0 ;
        RECT  62.7 39.6 63.6 51.0 ;
        RECT  95.25 198.6 96.45 199.8 ;
        RECT  95.25 226.8 96.45 228.0 ;
        RECT  95.25 255.0 96.45 256.2 ;
        RECT  95.25 283.2 96.45 284.4 ;
        RECT  95.25 311.4 96.45 312.6 ;
        RECT  95.25 339.6 96.45 340.8 ;
        RECT  95.25 367.8 96.45 369.0 ;
        RECT  95.25 396.0 96.45 397.2 ;
        RECT  95.25 424.2 96.45 425.4 ;
        RECT  76.5 88.65 77.7 89.85 ;
        RECT  81.6 88.5 82.8 89.7 ;
        RECT  73.5 102.75 74.7 103.95 ;
        RECT  84.3 102.6 85.5 103.8 ;
        RECT  76.5 145.05 77.7 146.25 ;
        RECT  87.0 144.9 88.2 146.1 ;
        RECT  73.5 159.15 74.7 160.35 ;
        RECT  89.7 159.0 90.9 160.2 ;
        RECT  78.6 85.8 79.8 87.0 ;
        RECT  78.6 114.0 79.8 115.2 ;
        RECT  78.6 142.2 79.8 143.4 ;
        RECT  78.6 170.4 79.8 171.6 ;
        RECT  65.7 75.3 66.9 76.5 ;
        RECT  81.6 75.3 82.8 76.5 ;
        RECT  65.7 65.1 66.9 66.3 ;
        RECT  84.3 65.1 85.5 66.3 ;
        RECT  65.7 54.9 66.9 56.1 ;
        RECT  87.0 54.9 88.2 56.1 ;
        RECT  65.7 44.7 66.9 45.9 ;
        RECT  89.7 44.7 90.9 45.9 ;
        RECT  66.3 70.2 67.5 71.4 ;
        RECT  95.25 70.35 96.45 71.55 ;
        RECT  66.3 49.8 67.5 51.0 ;
        RECT  95.25 49.95 96.45 51.15 ;
        RECT  110.4 32.25 111.6 33.45 ;
        RECT  105.0 27.75 106.2 28.95 ;
        RECT  107.7 25.35 108.9 26.55 ;
        RECT  110.4 429.45 111.6 430.65 ;
        RECT  113.1 96.75 114.3 97.95 ;
        RECT  115.8 194.85 117.0 196.05 ;
        RECT  102.3 82.5 103.5 83.7 ;
        RECT  49.65 426.3 50.85 427.5 ;
        RECT  102.3 426.3 103.5 427.5 ;
        RECT  98.55 23.4 99.75 24.6 ;
        RECT  98.55 192.9 99.75 194.1 ;
        RECT  98.55 94.8 99.75 96.0 ;
        RECT  -9.75 207.15 -8.85 208.05 ;
        RECT  -9.45 207.15 -9.3 208.05 ;
        RECT  -9.75 207.6 -8.85 217.2 ;
        RECT  -9.6 223.95 -8.7 224.85 ;
        RECT  -9.3 223.95 -9.15 224.85 ;
        RECT  -9.6 224.4 -8.7 231.6 ;
        RECT  -9.6 243.6 -8.7 250.8 ;
        RECT  -22.5 258.6 -17.55 259.5 ;
        RECT  -9.9 207.15 -9.0 208.05 ;
        RECT  -9.75 223.95 -8.85 224.85 ;
        RECT  -25.2 362.1 -24.3 375.45 ;
        RECT  -9.6 272.85 -8.7 284.85 ;
        RECT  -22.5 204.6 -19.8 205.5 ;
        RECT  -24.6 284.85 -23.7 311.7 ;
        RECT  -27.3 290.25 -26.4 314.7 ;
        RECT  -12.75 303.75 -11.85 312.3 ;
        RECT  -10.8 301.05 -9.9 314.7 ;
        RECT  -8.85 292.95 -7.95 317.1 ;
        RECT  -12.75 326.85 -11.85 327.75 ;
        RECT  -12.75 318.3 -11.85 327.3 ;
        RECT  -12.3 326.85 -9.45 327.75 ;
        RECT  -9.75 329.25 -8.85 330.15 ;
        RECT  -9.45 329.25 -9.3 330.15 ;
        RECT  -9.75 329.7 -8.85 387.3 ;
        RECT  -40.95 303.75 -40.05 321.9 ;
        RECT  -39.0 292.95 -38.1 324.3 ;
        RECT  -37.05 295.65 -36.15 326.7 ;
        RECT  -40.95 336.45 -40.05 337.35 ;
        RECT  -40.95 327.9 -40.05 336.9 ;
        RECT  -40.5 336.45 -37.65 337.35 ;
        RECT  -38.1 339.3 -37.2 346.5 ;
        RECT  -38.1 348.9 -37.2 356.1 ;
        RECT  -25.2 361.65 -24.3 362.55 ;
        RECT  -25.2 361.65 -24.75 362.55 ;
        RECT  -25.2 359.7 -24.3 362.1 ;
        RECT  -25.2 349.5 -24.3 356.7 ;
        RECT  -24.6 316.8 -23.7 323.1 ;
        RECT  -23.85 333.0 -22.95 340.2 ;
        RECT  -38.1 358.5 -37.2 362.7 ;
        RECT  -25.2 342.9 -24.3 347.1 ;
        RECT  -3.45 202.2 -2.55 362.1 ;
        RECT  -3.45 287.55 -2.55 308.7 ;
        RECT  -17.55 202.2 -16.65 362.1 ;
        RECT  -17.55 298.35 -16.65 308.7 ;
        RECT  -31.65 308.7 -30.75 362.1 ;
        RECT  -31.65 287.55 -30.75 308.7 ;
        RECT  -45.75 308.7 -44.85 362.1 ;
        RECT  -45.75 298.35 -44.85 308.7 ;
        RECT  -45.75 361.65 -44.85 362.55 ;
        RECT  -45.75 360.0 -44.85 362.1 ;
        RECT  -49.8 361.65 -45.3 362.55 ;
        RECT  -10.05 204.6 -8.85 205.8 ;
        RECT  -17.55 202.2 -16.65 203.1 ;
        RECT  -3.45 202.2 -2.55 203.1 ;
        RECT  -53.1 204.6 -22.5 205.5 ;
        RECT  -53.1 258.6 -22.5 259.5 ;
        RECT  -53.7 258.6 -42.3 259.5 ;
        RECT  -53.7 255.3 -52.5 258.6 ;
        RECT  -51.3 256.8 -44.7 257.7 ;
        RECT  -51.3 256.5 -48.3 256.8 ;
        RECT  -45.9 256.5 -44.7 256.8 ;
        RECT  -53.7 254.1 -49.5 255.3 ;
        RECT  -45.9 254.1 -42.3 255.3 ;
        RECT  -53.7 250.5 -52.5 254.1 ;
        RECT  -48.3 253.2 -47.1 254.1 ;
        RECT  -48.3 252.9 -45.9 253.2 ;
        RECT  -51.3 252.0 -44.7 252.9 ;
        RECT  -51.3 251.7 -49.5 252.0 ;
        RECT  -45.9 251.7 -44.7 252.0 ;
        RECT  -53.7 249.3 -49.5 250.5 ;
        RECT  -53.7 235.5 -52.5 249.3 ;
        RECT  -48.0 248.7 -46.8 251.1 ;
        RECT  -43.2 250.5 -42.3 254.1 ;
        RECT  -45.9 249.3 -42.3 250.5 ;
        RECT  -43.5 248.1 -42.3 249.3 ;
        RECT  -51.3 245.7 -50.1 246.9 ;
        RECT  -49.2 246.6 -46.8 247.8 ;
        RECT  -51.3 244.8 -44.7 245.7 ;
        RECT  -51.3 244.5 -49.5 244.8 ;
        RECT  -45.9 244.5 -44.7 244.8 ;
        RECT  -51.3 242.4 -44.7 243.3 ;
        RECT  -51.3 242.1 -49.5 242.4 ;
        RECT  -47.1 242.1 -44.7 242.4 ;
        RECT  -51.3 240.0 -44.7 240.9 ;
        RECT  -51.3 239.7 -49.5 240.0 ;
        RECT  -47.1 239.7 -44.7 240.0 ;
        RECT  -48.3 237.9 -47.1 238.8 ;
        RECT  -51.3 237.0 -44.7 237.9 ;
        RECT  -51.3 236.7 -48.3 237.0 ;
        RECT  -45.9 236.7 -44.7 237.0 ;
        RECT  -53.7 234.3 -49.5 235.5 ;
        RECT  -53.7 229.8 -52.5 234.3 ;
        RECT  -48.6 233.4 -47.4 235.8 ;
        RECT  -43.2 235.5 -42.3 248.1 ;
        RECT  -45.9 234.3 -42.3 235.5 ;
        RECT  -51.3 232.2 -50.1 233.4 ;
        RECT  -51.3 231.3 -44.7 232.2 ;
        RECT  -51.3 231.0 -49.5 231.3 ;
        RECT  -45.9 231.0 -44.7 231.3 ;
        RECT  -43.2 229.8 -42.3 234.3 ;
        RECT  -53.7 228.6 -49.5 229.8 ;
        RECT  -53.7 225.0 -52.5 228.6 ;
        RECT  -48.0 227.7 -46.8 228.9 ;
        RECT  -45.9 228.6 -42.3 229.8 ;
        RECT  -51.3 227.4 -45.9 227.7 ;
        RECT  -51.3 226.8 -44.7 227.4 ;
        RECT  -51.3 226.2 -49.5 226.8 ;
        RECT  -47.1 226.5 -44.7 226.8 ;
        RECT  -45.9 226.2 -44.7 226.5 ;
        RECT  -53.7 223.8 -49.5 225.0 ;
        RECT  -53.7 208.8 -52.5 223.8 ;
        RECT  -48.0 223.2 -46.8 225.6 ;
        RECT  -43.2 225.0 -42.3 228.6 ;
        RECT  -45.9 223.8 -42.3 225.0 ;
        RECT  -43.5 222.6 -42.3 223.8 ;
        RECT  -51.3 219.3 -50.1 220.5 ;
        RECT  -49.2 220.2 -46.8 221.4 ;
        RECT  -51.3 218.4 -44.7 219.3 ;
        RECT  -51.3 218.1 -49.5 218.4 ;
        RECT  -45.9 218.1 -44.7 218.4 ;
        RECT  -51.3 216.0 -44.7 216.9 ;
        RECT  -51.3 215.7 -49.5 216.0 ;
        RECT  -47.1 215.7 -44.7 216.0 ;
        RECT  -51.3 213.6 -44.7 214.5 ;
        RECT  -51.3 213.3 -49.5 213.6 ;
        RECT  -47.1 213.3 -44.7 213.6 ;
        RECT  -48.3 211.5 -47.1 212.4 ;
        RECT  -51.3 210.6 -44.7 211.5 ;
        RECT  -51.3 210.3 -48.3 210.6 ;
        RECT  -45.9 210.3 -44.7 210.6 ;
        RECT  -43.2 209.1 -42.3 222.6 ;
        RECT  -51.3 208.8 -49.5 209.1 ;
        RECT  -53.7 207.9 -49.5 208.8 ;
        RECT  -45.9 208.2 -42.3 209.1 ;
        RECT  -45.9 207.9 -44.7 208.2 ;
        RECT  -50.7 206.4 -49.5 207.9 ;
        RECT  -48.6 205.5 -47.4 206.4 ;
        RECT  -53.7 204.6 -42.3 205.5 ;
        RECT  -53.7 204.6 -42.3 205.5 ;
        RECT  -53.7 258.6 -42.3 259.5 ;
        RECT  -43.5 258.6 -32.1 259.5 ;
        RECT  -33.3 255.3 -32.1 258.6 ;
        RECT  -41.1 256.8 -34.5 257.7 ;
        RECT  -37.5 256.5 -34.5 256.8 ;
        RECT  -41.1 256.5 -39.9 256.8 ;
        RECT  -36.3 254.1 -32.1 255.3 ;
        RECT  -43.5 254.1 -39.9 255.3 ;
        RECT  -33.3 250.5 -32.1 254.1 ;
        RECT  -38.7 253.2 -37.5 254.1 ;
        RECT  -39.9 252.9 -37.5 253.2 ;
        RECT  -41.1 252.0 -34.5 252.9 ;
        RECT  -36.3 251.7 -34.5 252.0 ;
        RECT  -41.1 251.7 -39.9 252.0 ;
        RECT  -36.3 249.3 -32.1 250.5 ;
        RECT  -33.3 235.5 -32.1 249.3 ;
        RECT  -39.0 248.7 -37.8 251.1 ;
        RECT  -43.5 250.5 -42.6 254.1 ;
        RECT  -43.5 249.3 -39.9 250.5 ;
        RECT  -43.5 248.1 -42.3 249.3 ;
        RECT  -35.7 245.7 -34.5 246.9 ;
        RECT  -39.0 246.6 -36.6 247.8 ;
        RECT  -41.1 244.8 -34.5 245.7 ;
        RECT  -36.3 244.5 -34.5 244.8 ;
        RECT  -41.1 244.5 -39.9 244.8 ;
        RECT  -41.1 242.4 -34.5 243.3 ;
        RECT  -36.3 242.1 -34.5 242.4 ;
        RECT  -41.1 242.1 -38.7 242.4 ;
        RECT  -41.1 240.0 -34.5 240.9 ;
        RECT  -36.3 239.7 -34.5 240.0 ;
        RECT  -41.1 239.7 -38.7 240.0 ;
        RECT  -38.7 237.9 -37.5 238.8 ;
        RECT  -41.1 237.0 -34.5 237.9 ;
        RECT  -37.5 236.7 -34.5 237.0 ;
        RECT  -41.1 236.7 -39.9 237.0 ;
        RECT  -36.3 234.3 -32.1 235.5 ;
        RECT  -33.3 229.8 -32.1 234.3 ;
        RECT  -38.4 233.4 -37.2 235.8 ;
        RECT  -43.5 235.5 -42.6 248.1 ;
        RECT  -43.5 234.3 -39.9 235.5 ;
        RECT  -35.7 232.2 -34.5 233.4 ;
        RECT  -41.1 231.3 -34.5 232.2 ;
        RECT  -36.3 231.0 -34.5 231.3 ;
        RECT  -41.1 231.0 -39.9 231.3 ;
        RECT  -43.5 229.8 -42.6 234.3 ;
        RECT  -36.3 228.6 -32.1 229.8 ;
        RECT  -33.3 225.0 -32.1 228.6 ;
        RECT  -39.0 227.7 -37.8 228.9 ;
        RECT  -43.5 228.6 -39.9 229.8 ;
        RECT  -39.9 227.4 -34.5 227.7 ;
        RECT  -41.1 226.8 -34.5 227.4 ;
        RECT  -36.3 226.2 -34.5 226.8 ;
        RECT  -41.1 226.5 -38.7 226.8 ;
        RECT  -41.1 226.2 -39.9 226.5 ;
        RECT  -36.3 223.8 -32.1 225.0 ;
        RECT  -33.3 208.8 -32.1 223.8 ;
        RECT  -39.0 223.2 -37.8 225.6 ;
        RECT  -43.5 225.0 -42.6 228.6 ;
        RECT  -43.5 223.8 -39.9 225.0 ;
        RECT  -43.5 222.6 -42.3 223.8 ;
        RECT  -35.7 219.3 -34.5 220.5 ;
        RECT  -39.0 220.2 -36.6 221.4 ;
        RECT  -41.1 218.4 -34.5 219.3 ;
        RECT  -36.3 218.1 -34.5 218.4 ;
        RECT  -41.1 218.1 -39.9 218.4 ;
        RECT  -41.1 216.0 -34.5 216.9 ;
        RECT  -36.3 215.7 -34.5 216.0 ;
        RECT  -41.1 215.7 -38.7 216.0 ;
        RECT  -41.1 213.6 -34.5 214.5 ;
        RECT  -36.3 213.3 -34.5 213.6 ;
        RECT  -41.1 213.3 -38.7 213.6 ;
        RECT  -38.7 211.5 -37.5 212.4 ;
        RECT  -41.1 210.6 -34.5 211.5 ;
        RECT  -37.5 210.3 -34.5 210.6 ;
        RECT  -41.1 210.3 -39.9 210.6 ;
        RECT  -43.5 209.1 -42.6 222.6 ;
        RECT  -36.3 208.8 -34.5 209.1 ;
        RECT  -36.3 207.9 -32.1 208.8 ;
        RECT  -43.5 208.2 -39.9 209.1 ;
        RECT  -41.1 207.9 -39.9 208.2 ;
        RECT  -36.3 206.4 -35.1 207.9 ;
        RECT  -38.4 205.5 -37.2 206.4 ;
        RECT  -43.5 204.6 -32.1 205.5 ;
        RECT  -43.5 204.6 -32.1 205.5 ;
        RECT  -43.5 258.6 -32.1 259.5 ;
        RECT  -33.3 258.6 -21.9 259.5 ;
        RECT  -33.3 255.3 -32.1 258.6 ;
        RECT  -30.9 256.8 -24.3 257.7 ;
        RECT  -30.9 256.5 -27.9 256.8 ;
        RECT  -25.5 256.5 -24.3 256.8 ;
        RECT  -33.3 254.1 -29.1 255.3 ;
        RECT  -25.5 254.1 -21.9 255.3 ;
        RECT  -33.3 250.5 -32.1 254.1 ;
        RECT  -27.9 253.2 -26.7 254.1 ;
        RECT  -27.9 252.9 -25.5 253.2 ;
        RECT  -30.9 252.0 -24.3 252.9 ;
        RECT  -30.9 251.7 -29.1 252.0 ;
        RECT  -25.5 251.7 -24.3 252.0 ;
        RECT  -33.3 249.3 -29.1 250.5 ;
        RECT  -33.3 235.5 -32.1 249.3 ;
        RECT  -27.6 248.7 -26.4 251.1 ;
        RECT  -22.8 250.5 -21.9 254.1 ;
        RECT  -25.5 249.3 -21.9 250.5 ;
        RECT  -23.1 248.1 -21.9 249.3 ;
        RECT  -30.9 245.7 -29.7 246.9 ;
        RECT  -28.8 246.6 -26.4 247.8 ;
        RECT  -30.9 244.8 -24.3 245.7 ;
        RECT  -30.9 244.5 -29.1 244.8 ;
        RECT  -25.5 244.5 -24.3 244.8 ;
        RECT  -30.9 242.4 -24.3 243.3 ;
        RECT  -30.9 242.1 -29.1 242.4 ;
        RECT  -26.7 242.1 -24.3 242.4 ;
        RECT  -30.9 240.0 -24.3 240.9 ;
        RECT  -30.9 239.7 -29.1 240.0 ;
        RECT  -26.7 239.7 -24.3 240.0 ;
        RECT  -27.9 237.9 -26.7 238.8 ;
        RECT  -30.9 237.0 -24.3 237.9 ;
        RECT  -30.9 236.7 -27.9 237.0 ;
        RECT  -25.5 236.7 -24.3 237.0 ;
        RECT  -33.3 234.3 -29.1 235.5 ;
        RECT  -33.3 229.8 -32.1 234.3 ;
        RECT  -28.2 233.4 -27.0 235.8 ;
        RECT  -22.8 235.5 -21.9 248.1 ;
        RECT  -25.5 234.3 -21.9 235.5 ;
        RECT  -30.9 232.2 -29.7 233.4 ;
        RECT  -30.9 231.3 -24.3 232.2 ;
        RECT  -30.9 231.0 -29.1 231.3 ;
        RECT  -25.5 231.0 -24.3 231.3 ;
        RECT  -22.8 229.8 -21.9 234.3 ;
        RECT  -33.3 228.6 -29.1 229.8 ;
        RECT  -33.3 225.0 -32.1 228.6 ;
        RECT  -27.6 227.7 -26.4 228.9 ;
        RECT  -25.5 228.6 -21.9 229.8 ;
        RECT  -30.9 227.4 -25.5 227.7 ;
        RECT  -30.9 226.8 -24.3 227.4 ;
        RECT  -30.9 226.2 -29.1 226.8 ;
        RECT  -26.7 226.5 -24.3 226.8 ;
        RECT  -25.5 226.2 -24.3 226.5 ;
        RECT  -33.3 223.8 -29.1 225.0 ;
        RECT  -33.3 208.8 -32.1 223.8 ;
        RECT  -27.6 223.2 -26.4 225.6 ;
        RECT  -22.8 225.0 -21.9 228.6 ;
        RECT  -25.5 223.8 -21.9 225.0 ;
        RECT  -23.1 222.6 -21.9 223.8 ;
        RECT  -30.9 219.3 -29.7 220.5 ;
        RECT  -28.8 220.2 -26.4 221.4 ;
        RECT  -30.9 218.4 -24.3 219.3 ;
        RECT  -30.9 218.1 -29.1 218.4 ;
        RECT  -25.5 218.1 -24.3 218.4 ;
        RECT  -30.9 216.0 -24.3 216.9 ;
        RECT  -30.9 215.7 -29.1 216.0 ;
        RECT  -26.7 215.7 -24.3 216.0 ;
        RECT  -30.9 213.6 -24.3 214.5 ;
        RECT  -30.9 213.3 -29.1 213.6 ;
        RECT  -26.7 213.3 -24.3 213.6 ;
        RECT  -27.9 211.5 -26.7 212.4 ;
        RECT  -30.9 210.6 -24.3 211.5 ;
        RECT  -30.9 210.3 -27.9 210.6 ;
        RECT  -25.5 210.3 -24.3 210.6 ;
        RECT  -22.8 209.1 -21.9 222.6 ;
        RECT  -30.9 208.8 -29.1 209.1 ;
        RECT  -33.3 207.9 -29.1 208.8 ;
        RECT  -25.5 208.2 -21.9 209.1 ;
        RECT  -25.5 207.9 -24.3 208.2 ;
        RECT  -30.3 206.4 -29.1 207.9 ;
        RECT  -28.2 205.5 -27.0 206.4 ;
        RECT  -33.3 204.6 -21.9 205.5 ;
        RECT  -33.3 204.6 -21.9 205.5 ;
        RECT  -33.3 258.6 -21.9 259.5 ;
        RECT  -4.95 211.2 -3.0 212.4 ;
        RECT  -17.1 211.2 -15.15 212.4 ;
        RECT  -13.95 206.7 -5.55 207.6 ;
        RECT  -10.05 204.6 -8.85 205.8 ;
        RECT  -9.9 207.15 -9.0 208.05 ;
        RECT  -17.55 202.2 -16.65 214.2 ;
        RECT  -3.45 202.2 -2.55 214.2 ;
        RECT  -16.5 204.15 -14.55 205.05 ;
        RECT  -16.5 208.95 -14.55 209.85 ;
        RECT  -16.95 204.0 -16.05 210.0 ;
        RECT  -15.15 206.4 -13.95 207.6 ;
        RECT  -15.15 204.0 -13.95 205.2 ;
        RECT  -15.15 208.8 -13.95 210.0 ;
        RECT  -15.15 206.4 -13.95 207.6 ;
        RECT  -4.95 204.15 -3.0 205.05 ;
        RECT  -4.95 208.95 -3.0 209.85 ;
        RECT  -3.45 204.0 -2.55 210.0 ;
        RECT  -5.55 206.4 -4.35 207.6 ;
        RECT  -5.55 204.0 -4.35 205.2 ;
        RECT  -5.55 208.8 -4.35 210.0 ;
        RECT  -5.55 206.4 -4.35 207.6 ;
        RECT  -5.55 211.2 -4.35 212.4 ;
        RECT  -15.75 211.2 -14.55 212.4 ;
        RECT  -10.05 204.6 -8.85 205.8 ;
        RECT  -4.95 225.6 -3.0 226.8 ;
        RECT  -17.1 225.6 -15.15 226.8 ;
        RECT  -17.55 216.0 -15.75 222.0 ;
        RECT  -11.85 223.5 -7.65 224.4 ;
        RECT  -9.9 216.6 -8.7 217.8 ;
        RECT  -9.75 223.95 -8.85 224.85 ;
        RECT  -17.55 214.2 -16.65 228.6 ;
        RECT  -3.45 214.2 -2.55 228.6 ;
        RECT  -16.2 216.15 -14.25 217.05 ;
        RECT  -16.2 220.95 -14.25 221.85 ;
        RECT  -14.25 218.55 -12.3 219.45 ;
        RECT  -14.25 223.35 -12.3 224.25 ;
        RECT  -16.65 216.0 -15.75 222.0 ;
        RECT  -12.75 218.4 -11.85 224.4 ;
        RECT  -14.85 216.0 -13.65 217.2 ;
        RECT  -14.85 220.8 -13.65 222.0 ;
        RECT  -14.85 218.4 -13.65 219.6 ;
        RECT  -14.85 223.2 -13.65 224.4 ;
        RECT  -5.25 216.15 -3.3 217.05 ;
        RECT  -5.25 220.95 -3.3 221.85 ;
        RECT  -7.2 218.55 -5.25 219.45 ;
        RECT  -7.2 223.35 -5.25 224.25 ;
        RECT  -3.75 216.0 -2.85 222.0 ;
        RECT  -7.65 218.4 -6.75 224.4 ;
        RECT  -5.85 216.0 -4.65 217.2 ;
        RECT  -5.85 220.8 -4.65 222.0 ;
        RECT  -5.85 218.4 -4.65 219.6 ;
        RECT  -5.85 223.2 -4.65 224.4 ;
        RECT  -5.55 225.6 -4.35 226.8 ;
        RECT  -15.75 225.6 -14.55 226.8 ;
        RECT  -9.9 216.6 -8.7 217.8 ;
        RECT  -4.95 244.8 -3.0 246.0 ;
        RECT  -17.1 244.8 -15.15 246.0 ;
        RECT  -17.55 230.4 -15.3 241.2 ;
        RECT  -11.4 242.7 -7.8 243.6 ;
        RECT  -9.75 231.0 -8.55 232.2 ;
        RECT  -9.6 243.15 -8.7 244.05 ;
        RECT  -17.55 228.6 -16.65 247.8 ;
        RECT  -3.45 228.6 -2.55 247.8 ;
        RECT  -15.75 230.55 -13.8 231.45 ;
        RECT  -15.75 235.35 -13.8 236.25 ;
        RECT  -15.75 240.15 -13.8 241.05 ;
        RECT  -13.8 232.95 -11.85 233.85 ;
        RECT  -13.8 237.75 -11.85 238.65 ;
        RECT  -13.8 242.55 -11.85 243.45 ;
        RECT  -16.2 230.4 -15.3 241.2 ;
        RECT  -12.3 232.8 -11.4 243.6 ;
        RECT  -14.4 230.4 -13.2 231.6 ;
        RECT  -14.4 235.2 -13.2 236.4 ;
        RECT  -14.4 240.0 -13.2 241.2 ;
        RECT  -14.4 232.8 -13.2 234.0 ;
        RECT  -14.4 237.6 -13.2 238.8 ;
        RECT  -14.4 242.4 -13.2 243.6 ;
        RECT  -5.4 230.55 -3.45 231.45 ;
        RECT  -5.4 235.35 -3.45 236.25 ;
        RECT  -5.4 240.15 -3.45 241.05 ;
        RECT  -7.35 232.95 -5.4 233.85 ;
        RECT  -7.35 237.75 -5.4 238.65 ;
        RECT  -7.35 242.55 -5.4 243.45 ;
        RECT  -3.9 230.4 -3.0 241.2 ;
        RECT  -7.8 232.8 -6.9 243.6 ;
        RECT  -6.0 230.4 -4.8 231.6 ;
        RECT  -6.0 235.2 -4.8 236.4 ;
        RECT  -6.0 240.0 -4.8 241.2 ;
        RECT  -6.0 232.8 -4.8 234.0 ;
        RECT  -6.0 237.6 -4.8 238.8 ;
        RECT  -6.0 242.4 -4.8 243.6 ;
        RECT  -5.55 244.8 -4.35 246.0 ;
        RECT  -15.75 244.8 -14.55 246.0 ;
        RECT  -9.75 231.0 -8.55 232.2 ;
        RECT  -4.95 276.0 -3.0 277.2 ;
        RECT  -17.1 276.0 -15.15 277.2 ;
        RECT  -17.55 249.6 -15.3 274.8 ;
        RECT  -11.4 271.5 -7.8 272.4 ;
        RECT  -9.75 250.2 -8.55 251.4 ;
        RECT  -9.6 271.95 -8.7 272.85 ;
        RECT  -17.55 247.8 -16.65 279.0 ;
        RECT  -3.45 247.8 -2.55 279.0 ;
        RECT  -15.75 249.75 -13.8 250.65 ;
        RECT  -15.75 254.55 -13.8 255.45 ;
        RECT  -15.75 259.35 -13.8 260.25 ;
        RECT  -15.75 264.15 -13.8 265.05 ;
        RECT  -15.75 268.95 -13.8 269.85 ;
        RECT  -15.75 273.75 -13.8 274.65 ;
        RECT  -13.8 252.15 -11.85 253.05 ;
        RECT  -13.8 256.95 -11.85 257.85 ;
        RECT  -13.8 261.75 -11.85 262.65 ;
        RECT  -13.8 266.55 -11.85 267.45 ;
        RECT  -13.8 271.35 -11.85 272.25 ;
        RECT  -16.2 249.6 -15.3 274.8 ;
        RECT  -12.3 252.0 -11.4 272.4 ;
        RECT  -14.4 249.6 -13.2 250.8 ;
        RECT  -14.4 254.4 -13.2 255.6 ;
        RECT  -14.4 259.2 -13.2 260.4 ;
        RECT  -14.4 264.0 -13.2 265.2 ;
        RECT  -14.4 268.8 -13.2 270.0 ;
        RECT  -14.4 273.6 -13.2 274.8 ;
        RECT  -14.4 252.0 -13.2 253.2 ;
        RECT  -14.4 256.8 -13.2 258.0 ;
        RECT  -14.4 261.6 -13.2 262.8 ;
        RECT  -14.4 266.4 -13.2 267.6 ;
        RECT  -14.4 271.2 -13.2 272.4 ;
        RECT  -5.4 249.75 -3.45 250.65 ;
        RECT  -5.4 254.55 -3.45 255.45 ;
        RECT  -5.4 259.35 -3.45 260.25 ;
        RECT  -5.4 264.15 -3.45 265.05 ;
        RECT  -5.4 268.95 -3.45 269.85 ;
        RECT  -5.4 273.75 -3.45 274.65 ;
        RECT  -7.35 252.15 -5.4 253.05 ;
        RECT  -7.35 256.95 -5.4 257.85 ;
        RECT  -7.35 261.75 -5.4 262.65 ;
        RECT  -7.35 266.55 -5.4 267.45 ;
        RECT  -7.35 271.35 -5.4 272.25 ;
        RECT  -3.9 249.6 -3.0 274.8 ;
        RECT  -7.8 252.0 -6.9 272.4 ;
        RECT  -6.0 249.6 -4.8 250.8 ;
        RECT  -6.0 254.4 -4.8 255.6 ;
        RECT  -6.0 259.2 -4.8 260.4 ;
        RECT  -6.0 264.0 -4.8 265.2 ;
        RECT  -6.0 268.8 -4.8 270.0 ;
        RECT  -6.0 273.6 -4.8 274.8 ;
        RECT  -6.0 252.0 -4.8 253.2 ;
        RECT  -6.0 256.8 -4.8 258.0 ;
        RECT  -6.0 261.6 -4.8 262.8 ;
        RECT  -6.0 266.4 -4.8 267.6 ;
        RECT  -6.0 271.2 -4.8 272.4 ;
        RECT  -5.55 276.0 -4.35 277.2 ;
        RECT  -15.75 276.0 -14.55 277.2 ;
        RECT  -9.75 250.2 -8.55 251.4 ;
        RECT  -4.5 320.1 -3.0 321.3 ;
        RECT  -17.1 320.1 -15.6 321.3 ;
        RECT  -5.1 310.5 -2.55 311.7 ;
        RECT  -17.55 310.5 -14.4 311.7 ;
        RECT  -17.55 315.3 -14.4 316.5 ;
        RECT  -12.9 311.7 -11.7 312.9 ;
        RECT  -9.0 316.5 -7.8 317.7 ;
        RECT  -10.95 314.1 -9.75 315.3 ;
        RECT  -17.55 308.7 -16.65 324.3 ;
        RECT  -3.45 308.7 -2.55 324.3 ;
        RECT  -12.9 317.7 -11.7 318.9 ;
        RECT  -15.6 310.5 -14.4 311.7 ;
        RECT  -15.6 312.9 -14.4 314.1 ;
        RECT  -15.6 310.5 -14.4 311.7 ;
        RECT  -15.6 312.9 -14.4 314.1 ;
        RECT  -15.6 312.9 -14.4 314.1 ;
        RECT  -15.6 315.3 -14.4 316.5 ;
        RECT  -15.6 312.9 -14.4 314.1 ;
        RECT  -15.6 315.3 -14.4 316.5 ;
        RECT  -15.6 315.3 -14.4 316.5 ;
        RECT  -15.6 317.7 -14.4 318.9 ;
        RECT  -15.6 315.3 -14.4 316.5 ;
        RECT  -15.6 317.7 -14.4 318.9 ;
        RECT  -6.3 310.5 -5.1 311.7 ;
        RECT  -6.3 312.9 -5.1 314.1 ;
        RECT  -6.3 310.5 -5.1 311.7 ;
        RECT  -6.3 312.9 -5.1 314.1 ;
        RECT  -6.3 312.9 -5.1 314.1 ;
        RECT  -6.3 315.3 -5.1 316.5 ;
        RECT  -6.3 312.9 -5.1 314.1 ;
        RECT  -6.3 315.3 -5.1 316.5 ;
        RECT  -6.3 315.3 -5.1 316.5 ;
        RECT  -6.3 317.7 -5.1 318.9 ;
        RECT  -6.3 315.3 -5.1 316.5 ;
        RECT  -6.3 317.7 -5.1 318.9 ;
        RECT  -5.1 320.1 -3.9 321.3 ;
        RECT  -16.2 320.1 -15.0 321.3 ;
        RECT  -9.0 316.5 -7.8 317.7 ;
        RECT  -10.95 314.1 -9.75 315.3 ;
        RECT  -12.9 311.7 -11.7 312.9 ;
        RECT  -15.6 312.9 -14.4 314.1 ;
        RECT  -15.6 317.7 -14.4 318.9 ;
        RECT  -6.3 317.7 -5.1 318.9 ;
        RECT  -12.9 317.7 -11.7 318.9 ;
        RECT  -4.95 330.9 -3.0 332.1 ;
        RECT  -17.1 330.9 -15.15 332.1 ;
        RECT  -4.35 326.1 -2.55 327.3 ;
        RECT  -17.55 326.1 -13.95 327.3 ;
        RECT  -13.95 328.8 -5.55 329.7 ;
        RECT  -10.05 326.7 -8.85 327.9 ;
        RECT  -9.9 329.25 -9.0 330.15 ;
        RECT  -17.55 324.3 -16.65 333.9 ;
        RECT  -3.45 324.3 -2.55 333.9 ;
        RECT  -15.15 326.1 -13.95 327.3 ;
        RECT  -15.15 328.5 -13.95 329.7 ;
        RECT  -15.15 326.1 -13.95 327.3 ;
        RECT  -15.15 328.5 -13.95 329.7 ;
        RECT  -5.55 326.1 -4.35 327.3 ;
        RECT  -5.55 328.5 -4.35 329.7 ;
        RECT  -5.55 326.1 -4.35 327.3 ;
        RECT  -5.55 328.5 -4.35 329.7 ;
        RECT  -5.55 330.9 -4.35 332.1 ;
        RECT  -15.75 330.9 -14.55 332.1 ;
        RECT  -10.05 326.7 -8.85 327.9 ;
        RECT  -31.2 317.7 -29.25 318.9 ;
        RECT  -19.05 317.7 -17.1 318.9 ;
        RECT  -31.65 310.5 -29.85 311.7 ;
        RECT  -31.65 315.3 -29.85 316.5 ;
        RECT  -20.85 310.5 -16.65 311.7 ;
        RECT  -24.75 311.1 -23.55 312.3 ;
        RECT  -24.75 316.2 -23.55 317.4 ;
        RECT  -27.45 314.1 -26.25 315.3 ;
        RECT  -17.55 308.7 -16.65 323.1 ;
        RECT  -31.65 308.7 -30.75 323.1 ;
        RECT  -24.45 310.5 -23.25 311.7 ;
        RECT  -24.45 312.9 -23.25 314.1 ;
        RECT  -24.45 310.5 -23.25 311.7 ;
        RECT  -24.45 312.9 -23.25 314.1 ;
        RECT  -24.45 312.9 -23.25 314.1 ;
        RECT  -24.45 315.3 -23.25 316.5 ;
        RECT  -24.45 312.9 -23.25 314.1 ;
        RECT  -24.45 315.3 -23.25 316.5 ;
        RECT  -31.05 310.5 -29.85 311.7 ;
        RECT  -31.05 312.9 -29.85 314.1 ;
        RECT  -31.05 310.5 -29.85 311.7 ;
        RECT  -31.05 312.9 -29.85 314.1 ;
        RECT  -31.05 312.9 -29.85 314.1 ;
        RECT  -31.05 315.3 -29.85 316.5 ;
        RECT  -31.05 312.9 -29.85 314.1 ;
        RECT  -31.05 315.3 -29.85 316.5 ;
        RECT  -31.05 317.7 -29.85 318.9 ;
        RECT  -20.85 317.7 -19.65 318.9 ;
        RECT  -28.65 314.1 -27.45 315.3 ;
        RECT  -25.95 311.1 -24.75 312.3 ;
        RECT  -22.05 315.3 -20.85 316.5 ;
        RECT  -31.05 312.9 -29.85 314.1 ;
        RECT  -25.95 316.2 -24.75 317.4 ;
        RECT  -31.2 334.8 -29.25 336.0 ;
        RECT  -19.05 334.8 -17.1 336.0 ;
        RECT  -31.65 327.6 -29.25 328.8 ;
        RECT  -20.25 327.6 -16.65 328.8 ;
        RECT  -20.25 332.4 -16.65 333.6 ;
        RECT  -24.0 328.2 -22.8 329.4 ;
        RECT  -24.0 332.4 -22.8 333.6 ;
        RECT  -26.7 331.2 -25.5 332.4 ;
        RECT  -17.55 325.8 -16.65 340.2 ;
        RECT  -31.65 325.8 -30.75 340.2 ;
        RECT  -22.65 327.6 -21.45 328.8 ;
        RECT  -22.65 330.0 -21.45 331.2 ;
        RECT  -22.65 327.6 -21.45 328.8 ;
        RECT  -22.65 330.0 -21.45 331.2 ;
        RECT  -22.65 330.0 -21.45 331.2 ;
        RECT  -22.65 332.4 -21.45 333.6 ;
        RECT  -22.65 330.0 -21.45 331.2 ;
        RECT  -22.65 332.4 -21.45 333.6 ;
        RECT  -31.65 327.6 -30.45 328.8 ;
        RECT  -31.65 330.0 -30.45 331.2 ;
        RECT  -31.65 327.6 -30.45 328.8 ;
        RECT  -31.65 330.0 -30.45 331.2 ;
        RECT  -31.65 330.0 -30.45 331.2 ;
        RECT  -31.65 332.4 -30.45 333.6 ;
        RECT  -31.65 330.0 -30.45 331.2 ;
        RECT  -31.65 332.4 -30.45 333.6 ;
        RECT  -31.05 334.8 -29.85 336.0 ;
        RECT  -20.85 334.8 -19.65 336.0 ;
        RECT  -27.9 331.2 -26.7 332.4 ;
        RECT  -25.2 328.2 -24.0 329.4 ;
        RECT  -21.45 330.0 -20.25 331.2 ;
        RECT  -30.45 332.4 -29.25 333.6 ;
        RECT  -25.2 332.4 -24.0 333.6 ;
        RECT  -31.2 344.7 -29.25 345.9 ;
        RECT  -19.05 344.7 -17.1 345.9 ;
        RECT  -31.65 349.5 -29.85 350.7 ;
        RECT  -20.25 349.5 -16.65 350.7 ;
        RECT  -28.65 347.1 -20.25 348.0 ;
        RECT  -25.35 348.9 -24.15 350.1 ;
        RECT  -25.2 346.65 -24.3 347.55 ;
        RECT  -17.55 342.9 -16.65 352.5 ;
        RECT  -31.65 342.9 -30.75 352.5 ;
        RECT  -20.25 349.5 -19.05 350.7 ;
        RECT  -20.25 347.1 -19.05 348.3 ;
        RECT  -20.25 349.5 -19.05 350.7 ;
        RECT  -20.25 347.1 -19.05 348.3 ;
        RECT  -29.85 349.5 -28.65 350.7 ;
        RECT  -29.85 347.1 -28.65 348.3 ;
        RECT  -29.85 349.5 -28.65 350.7 ;
        RECT  -29.85 347.1 -28.65 348.3 ;
        RECT  -29.85 344.7 -28.65 345.9 ;
        RECT  -19.65 344.7 -18.45 345.9 ;
        RECT  -25.35 348.9 -24.15 350.1 ;
        RECT  -31.2 354.3 -29.25 355.5 ;
        RECT  -19.05 354.3 -17.1 355.5 ;
        RECT  -31.65 359.1 -29.85 360.3 ;
        RECT  -20.25 359.1 -16.65 360.3 ;
        RECT  -28.65 356.7 -20.25 357.6 ;
        RECT  -25.35 358.5 -24.15 359.7 ;
        RECT  -25.2 356.25 -24.3 357.15 ;
        RECT  -17.55 352.5 -16.65 362.1 ;
        RECT  -31.65 352.5 -30.75 362.1 ;
        RECT  -20.25 359.1 -19.05 360.3 ;
        RECT  -20.25 356.7 -19.05 357.9 ;
        RECT  -20.25 359.1 -19.05 360.3 ;
        RECT  -20.25 356.7 -19.05 357.9 ;
        RECT  -29.85 359.1 -28.65 360.3 ;
        RECT  -29.85 356.7 -28.65 357.9 ;
        RECT  -29.85 359.1 -28.65 360.3 ;
        RECT  -29.85 356.7 -28.65 357.9 ;
        RECT  -29.85 354.3 -28.65 355.5 ;
        RECT  -19.65 354.3 -18.45 355.5 ;
        RECT  -25.35 358.5 -24.15 359.7 ;
        RECT  -32.7 329.7 -31.2 330.9 ;
        RECT  -45.3 329.7 -43.8 330.9 ;
        RECT  -33.3 320.1 -30.75 321.3 ;
        RECT  -45.75 320.1 -42.6 321.3 ;
        RECT  -45.75 324.9 -42.6 326.1 ;
        RECT  -41.1 321.3 -39.9 322.5 ;
        RECT  -37.2 326.1 -36.0 327.3 ;
        RECT  -39.15 323.7 -37.95 324.9 ;
        RECT  -45.75 318.3 -44.85 333.9 ;
        RECT  -31.65 318.3 -30.75 333.9 ;
        RECT  -41.1 327.3 -39.9 328.5 ;
        RECT  -43.8 320.1 -42.6 321.3 ;
        RECT  -43.8 322.5 -42.6 323.7 ;
        RECT  -43.8 320.1 -42.6 321.3 ;
        RECT  -43.8 322.5 -42.6 323.7 ;
        RECT  -43.8 322.5 -42.6 323.7 ;
        RECT  -43.8 324.9 -42.6 326.1 ;
        RECT  -43.8 322.5 -42.6 323.7 ;
        RECT  -43.8 324.9 -42.6 326.1 ;
        RECT  -43.8 324.9 -42.6 326.1 ;
        RECT  -43.8 327.3 -42.6 328.5 ;
        RECT  -43.8 324.9 -42.6 326.1 ;
        RECT  -43.8 327.3 -42.6 328.5 ;
        RECT  -34.5 320.1 -33.3 321.3 ;
        RECT  -34.5 322.5 -33.3 323.7 ;
        RECT  -34.5 320.1 -33.3 321.3 ;
        RECT  -34.5 322.5 -33.3 323.7 ;
        RECT  -34.5 322.5 -33.3 323.7 ;
        RECT  -34.5 324.9 -33.3 326.1 ;
        RECT  -34.5 322.5 -33.3 323.7 ;
        RECT  -34.5 324.9 -33.3 326.1 ;
        RECT  -34.5 324.9 -33.3 326.1 ;
        RECT  -34.5 327.3 -33.3 328.5 ;
        RECT  -34.5 324.9 -33.3 326.1 ;
        RECT  -34.5 327.3 -33.3 328.5 ;
        RECT  -33.3 329.7 -32.1 330.9 ;
        RECT  -44.4 329.7 -43.2 330.9 ;
        RECT  -37.2 326.1 -36.0 327.3 ;
        RECT  -39.15 323.7 -37.95 324.9 ;
        RECT  -41.1 321.3 -39.9 322.5 ;
        RECT  -43.8 322.5 -42.6 323.7 ;
        RECT  -43.8 327.3 -42.6 328.5 ;
        RECT  -34.5 327.3 -33.3 328.5 ;
        RECT  -41.1 327.3 -39.9 328.5 ;
        RECT  -33.15 340.5 -31.2 341.7 ;
        RECT  -45.3 340.5 -43.35 341.7 ;
        RECT  -32.55 335.7 -30.75 336.9 ;
        RECT  -45.75 335.7 -42.15 336.9 ;
        RECT  -42.15 338.4 -33.75 339.3 ;
        RECT  -38.25 336.3 -37.05 337.5 ;
        RECT  -38.1 338.85 -37.2 339.75 ;
        RECT  -45.75 333.9 -44.85 343.5 ;
        RECT  -31.65 333.9 -30.75 343.5 ;
        RECT  -43.35 335.7 -42.15 336.9 ;
        RECT  -43.35 338.1 -42.15 339.3 ;
        RECT  -43.35 335.7 -42.15 336.9 ;
        RECT  -43.35 338.1 -42.15 339.3 ;
        RECT  -33.75 335.7 -32.55 336.9 ;
        RECT  -33.75 338.1 -32.55 339.3 ;
        RECT  -33.75 335.7 -32.55 336.9 ;
        RECT  -33.75 338.1 -32.55 339.3 ;
        RECT  -33.75 340.5 -32.55 341.7 ;
        RECT  -43.95 340.5 -42.75 341.7 ;
        RECT  -38.25 336.3 -37.05 337.5 ;
        RECT  -33.15 350.1 -31.2 351.3 ;
        RECT  -45.3 350.1 -43.35 351.3 ;
        RECT  -32.55 345.3 -30.75 346.5 ;
        RECT  -45.75 345.3 -42.15 346.5 ;
        RECT  -42.15 348.0 -33.75 348.9 ;
        RECT  -38.25 345.9 -37.05 347.1 ;
        RECT  -38.1 348.45 -37.2 349.35 ;
        RECT  -45.75 343.5 -44.85 353.1 ;
        RECT  -31.65 343.5 -30.75 353.1 ;
        RECT  -43.35 345.3 -42.15 346.5 ;
        RECT  -43.35 347.7 -42.15 348.9 ;
        RECT  -43.35 345.3 -42.15 346.5 ;
        RECT  -43.35 347.7 -42.15 348.9 ;
        RECT  -33.75 345.3 -32.55 346.5 ;
        RECT  -33.75 347.7 -32.55 348.9 ;
        RECT  -33.75 345.3 -32.55 346.5 ;
        RECT  -33.75 347.7 -32.55 348.9 ;
        RECT  -33.75 350.1 -32.55 351.3 ;
        RECT  -43.95 350.1 -42.75 351.3 ;
        RECT  -38.25 345.9 -37.05 347.1 ;
        RECT  -33.15 359.7 -31.2 360.9 ;
        RECT  -45.3 359.7 -43.35 360.9 ;
        RECT  -32.55 354.9 -30.75 356.1 ;
        RECT  -45.75 354.9 -42.15 356.1 ;
        RECT  -42.15 357.6 -33.75 358.5 ;
        RECT  -38.25 355.5 -37.05 356.7 ;
        RECT  -38.1 358.05 -37.2 358.95 ;
        RECT  -45.75 353.1 -44.85 362.7 ;
        RECT  -31.65 353.1 -30.75 362.7 ;
        RECT  -43.35 354.9 -42.15 356.1 ;
        RECT  -43.35 357.3 -42.15 358.5 ;
        RECT  -43.35 354.9 -42.15 356.1 ;
        RECT  -43.35 357.3 -42.15 358.5 ;
        RECT  -33.75 354.9 -32.55 356.1 ;
        RECT  -33.75 357.3 -32.55 358.5 ;
        RECT  -33.75 354.9 -32.55 356.1 ;
        RECT  -33.75 357.3 -32.55 358.5 ;
        RECT  -33.75 359.7 -32.55 360.9 ;
        RECT  -43.95 359.7 -42.75 360.9 ;
        RECT  -38.25 355.5 -37.05 356.7 ;
        RECT  -36.6 398.1 -30.75 399.0 ;
        RECT  -36.6 420.9 -30.75 421.8 ;
        RECT  -46.8 426.45 -31.2 427.35 ;
        RECT  -48.9 409.5 -36.6 410.4 ;
        RECT  -48.9 381.3 -36.6 382.2 ;
        RECT  -25.2 397.5 -24.3 410.1 ;
        RECT  -25.2 392.85 -24.3 393.75 ;
        RECT  -25.2 393.3 -24.3 397.5 ;
        RECT  -36.6 392.85 -24.75 393.75 ;
        RECT  -19.5 398.25 -17.1 399.15 ;
        RECT  -20.55 383.55 -19.65 384.45 ;
        RECT  -25.2 383.55 -24.3 384.45 ;
        RECT  -20.55 384.0 -19.65 395.7 ;
        RECT  -24.75 383.55 -20.1 384.45 ;
        RECT  -25.2 378.9 -24.3 384.0 ;
        RECT  -33.45 383.55 -24.75 384.45 ;
        RECT  -40.2 376.05 -33.45 376.95 ;
        RECT  -25.35 377.7 -24.15 378.9 ;
        RECT  -25.2 410.1 -24.3 413.85 ;
        RECT  -9.75 362.1 -8.85 412.5 ;
        RECT  -49.8 362.1 -48.9 424.65 ;
        RECT  -17.55 362.1 -16.65 410.1 ;
        RECT  -31.65 362.1 -30.75 381.3 ;
        RECT  -3.45 362.1 -2.55 410.1 ;
        RECT  -25.2 362.1 -24.3 375.45 ;
        RECT  -31.2 387.9 -29.25 389.1 ;
        RECT  -19.05 387.9 -17.1 389.1 ;
        RECT  -31.65 383.1 -29.85 384.3 ;
        RECT  -20.25 383.1 -16.65 384.3 ;
        RECT  -28.65 385.8 -20.25 386.7 ;
        RECT  -25.35 383.7 -24.15 384.9 ;
        RECT  -25.2 386.25 -24.3 387.15 ;
        RECT  -17.55 381.3 -16.65 390.9 ;
        RECT  -31.65 381.3 -30.75 390.9 ;
        RECT  -22.65 383.1 -21.45 384.3 ;
        RECT  -22.65 385.5 -21.45 386.7 ;
        RECT  -22.65 383.1 -21.45 384.3 ;
        RECT  -22.65 385.5 -21.45 386.7 ;
        RECT  -31.05 383.1 -29.85 384.3 ;
        RECT  -31.05 385.5 -29.85 386.7 ;
        RECT  -31.05 383.1 -29.85 384.3 ;
        RECT  -31.05 385.5 -29.85 386.7 ;
        RECT  -31.05 387.9 -29.85 389.1 ;
        RECT  -20.85 387.9 -19.65 389.1 ;
        RECT  -26.55 383.7 -25.35 384.9 ;
        RECT  -20.7 394.5 -19.5 395.7 ;
        RECT  -20.7 392.1 -19.5 393.3 ;
        RECT  -20.7 394.5 -19.5 395.7 ;
        RECT  -20.7 392.1 -19.5 393.3 ;
        RECT  -31.65 388.65 -30.75 389.55 ;
        RECT  -3.45 388.65 -2.55 389.55 ;
        RECT  -31.65 389.1 -30.75 390.9 ;
        RECT  -31.2 388.65 -3.0 389.55 ;
        RECT  -3.45 389.1 -2.55 390.9 ;
        RECT  -25.2 406.35 -24.3 410.1 ;
        RECT  -17.55 390.9 -16.65 410.1 ;
        RECT  -31.65 390.9 -30.75 410.1 ;
        RECT  -3.45 390.9 -2.55 410.1 ;
        RECT  -10.05 406.5 -8.85 407.7 ;
        RECT  -4.95 402.3 -3.0 403.5 ;
        RECT  -17.1 402.3 -15.15 403.5 ;
        RECT  -4.35 407.1 -2.55 408.3 ;
        RECT  -17.55 407.1 -13.95 408.3 ;
        RECT  -13.95 404.7 -5.55 405.6 ;
        RECT  -10.05 406.5 -8.85 407.7 ;
        RECT  -9.9 404.25 -9.0 405.15 ;
        RECT  -17.55 400.5 -16.65 410.1 ;
        RECT  -3.45 400.5 -2.55 410.1 ;
        RECT  -12.75 407.1 -11.55 408.3 ;
        RECT  -12.75 404.7 -11.55 405.9 ;
        RECT  -12.75 407.1 -11.55 408.3 ;
        RECT  -12.75 404.7 -11.55 405.9 ;
        RECT  -4.35 407.1 -3.15 408.3 ;
        RECT  -4.35 404.7 -3.15 405.9 ;
        RECT  -4.35 407.1 -3.15 408.3 ;
        RECT  -4.35 404.7 -3.15 405.9 ;
        RECT  -4.35 402.3 -3.15 403.5 ;
        RECT  -14.55 402.3 -13.35 403.5 ;
        RECT  -8.85 406.5 -7.65 407.7 ;
        RECT  -4.95 392.7 -3.0 393.9 ;
        RECT  -17.1 392.7 -15.15 393.9 ;
        RECT  -4.35 397.5 -2.55 398.7 ;
        RECT  -17.55 397.5 -13.95 398.7 ;
        RECT  -13.95 395.1 -5.55 396.0 ;
        RECT  -10.05 396.9 -8.85 398.1 ;
        RECT  -9.9 394.65 -9.0 395.55 ;
        RECT  -17.55 390.9 -16.65 400.5 ;
        RECT  -3.45 390.9 -2.55 400.5 ;
        RECT  -12.75 397.5 -11.55 398.7 ;
        RECT  -12.75 395.1 -11.55 396.3 ;
        RECT  -12.75 397.5 -11.55 398.7 ;
        RECT  -12.75 395.1 -11.55 396.3 ;
        RECT  -4.35 397.5 -3.15 398.7 ;
        RECT  -4.35 395.1 -3.15 396.3 ;
        RECT  -4.35 397.5 -3.15 398.7 ;
        RECT  -4.35 395.1 -3.15 396.3 ;
        RECT  -4.35 392.7 -3.15 393.9 ;
        RECT  -14.55 392.7 -13.35 393.9 ;
        RECT  -8.85 396.9 -7.65 398.1 ;
        RECT  -10.05 396.9 -8.85 398.1 ;
        RECT  -31.2 397.5 -29.25 398.7 ;
        RECT  -19.05 397.5 -17.1 398.7 ;
        RECT  -31.65 392.7 -29.85 393.9 ;
        RECT  -20.25 392.7 -16.65 393.9 ;
        RECT  -28.65 395.4 -20.25 396.3 ;
        RECT  -25.35 393.3 -24.15 394.5 ;
        RECT  -25.2 395.85 -24.3 396.75 ;
        RECT  -17.55 390.9 -16.65 400.5 ;
        RECT  -31.65 390.9 -30.75 400.5 ;
        RECT  -22.65 392.7 -21.45 393.9 ;
        RECT  -22.65 395.1 -21.45 396.3 ;
        RECT  -22.65 392.7 -21.45 393.9 ;
        RECT  -22.65 395.1 -21.45 396.3 ;
        RECT  -31.05 392.7 -29.85 393.9 ;
        RECT  -31.05 395.1 -29.85 396.3 ;
        RECT  -31.05 392.7 -29.85 393.9 ;
        RECT  -31.05 395.1 -29.85 396.3 ;
        RECT  -31.05 397.5 -29.85 398.7 ;
        RECT  -20.85 397.5 -19.65 398.7 ;
        RECT  -26.55 393.3 -25.35 394.5 ;
        RECT  -25.35 393.3 -24.15 394.5 ;
        RECT  -31.2 407.1 -29.25 408.3 ;
        RECT  -19.05 407.1 -17.1 408.3 ;
        RECT  -31.65 402.3 -29.85 403.5 ;
        RECT  -20.25 402.3 -16.65 403.5 ;
        RECT  -28.65 405.0 -20.25 405.9 ;
        RECT  -25.35 402.9 -24.15 404.1 ;
        RECT  -25.2 405.45 -24.3 406.35 ;
        RECT  -17.55 400.5 -16.65 410.1 ;
        RECT  -31.65 400.5 -30.75 410.1 ;
        RECT  -22.65 402.3 -21.45 403.5 ;
        RECT  -22.65 404.7 -21.45 405.9 ;
        RECT  -22.65 402.3 -21.45 403.5 ;
        RECT  -22.65 404.7 -21.45 405.9 ;
        RECT  -31.05 402.3 -29.85 403.5 ;
        RECT  -31.05 404.7 -29.85 405.9 ;
        RECT  -31.05 402.3 -29.85 403.5 ;
        RECT  -31.05 404.7 -29.85 405.9 ;
        RECT  -31.05 407.1 -29.85 408.3 ;
        RECT  -20.85 407.1 -19.65 408.3 ;
        RECT  -26.55 402.9 -25.35 404.1 ;
        RECT  -25.35 402.9 -24.15 404.1 ;
        RECT  -10.05 404.1 -8.85 405.3 ;
        RECT  -10.05 394.5 -8.85 395.7 ;
        RECT  -25.35 395.7 -24.15 396.9 ;
        RECT  -47.4 409.5 -36.6 410.7 ;
        RECT  -38.4 407.4 -37.2 409.5 ;
        RECT  -41.4 407.4 -40.2 408.6 ;
        RECT  -44.4 407.4 -43.2 408.6 ;
        RECT  -47.4 407.4 -46.2 409.5 ;
        RECT  -41.1 406.5 -39.9 407.4 ;
        RECT  -42.3 405.3 -37.2 406.5 ;
        RECT  -38.4 400.2 -37.2 405.3 ;
        RECT  -41.1 402.0 -39.9 405.3 ;
        RECT  -44.7 403.8 -43.5 407.4 ;
        RECT  -44.7 402.6 -42.9 403.8 ;
        RECT  -44.7 402.0 -43.5 402.6 ;
        RECT  -40.8 400.8 -39.6 402.0 ;
        RECT  -45.0 400.8 -43.8 402.0 ;
        RECT  -47.4 400.8 -46.2 406.5 ;
        RECT  -42.9 399.3 -41.7 399.6 ;
        RECT  -47.4 398.1 -36.6 399.3 ;
        RECT  -40.8 396.0 -38.1 397.2 ;
        RECT  -45.0 396.0 -42.3 397.2 ;
        RECT  -47.4 398.1 -36.6 399.3 ;
        RECT  -47.4 409.5 -36.6 410.7 ;
        RECT  -47.4 392.7 -36.0 393.9 ;
        RECT  -47.4 369.9 -36.0 371.1 ;
        RECT  -47.4 381.6 -36.0 382.5 ;
        RECT  -45.0 394.8 -42.3 396.0 ;
        RECT  -40.8 394.8 -38.1 396.0 ;
        RECT  -47.4 392.7 -36.0 393.9 ;
        RECT  -42.9 392.4 -41.7 392.7 ;
        RECT  -47.4 385.5 -46.2 391.2 ;
        RECT  -45.0 390.0 -43.8 391.2 ;
        RECT  -40.8 390.0 -39.6 391.2 ;
        RECT  -44.7 389.4 -43.5 390.0 ;
        RECT  -44.7 388.2 -42.9 389.4 ;
        RECT  -44.7 384.6 -43.5 388.2 ;
        RECT  -41.1 386.7 -39.9 390.0 ;
        RECT  -42.3 385.5 -39.9 386.7 ;
        RECT  -38.4 385.5 -37.2 391.2 ;
        RECT  -41.1 384.6 -39.9 385.5 ;
        RECT  -47.4 382.5 -46.2 384.6 ;
        RECT  -44.4 383.4 -43.2 384.6 ;
        RECT  -41.4 383.4 -40.2 384.6 ;
        RECT  -38.4 382.5 -37.2 384.6 ;
        RECT  -47.4 381.3 -36.0 382.5 ;
        RECT  -47.4 392.7 -36.0 393.9 ;
        RECT  -47.4 381.3 -36.0 382.5 ;
        RECT  -45.0 367.8 -42.3 369.0 ;
        RECT  -40.8 367.8 -38.1 369.0 ;
        RECT  -47.4 369.9 -36.0 371.1 ;
        RECT  -42.9 371.1 -41.7 371.4 ;
        RECT  -47.4 372.6 -46.2 378.3 ;
        RECT  -45.0 372.6 -43.8 373.8 ;
        RECT  -40.8 372.6 -39.6 373.8 ;
        RECT  -44.7 373.8 -43.5 374.4 ;
        RECT  -44.7 374.4 -42.9 375.6 ;
        RECT  -44.7 375.6 -43.5 379.2 ;
        RECT  -41.1 373.8 -39.9 377.1 ;
        RECT  -42.3 377.1 -39.9 378.3 ;
        RECT  -38.4 372.6 -37.2 378.3 ;
        RECT  -41.1 378.3 -39.9 379.2 ;
        RECT  -47.4 379.2 -46.2 381.3 ;
        RECT  -44.4 379.2 -43.2 380.4 ;
        RECT  -41.4 379.2 -40.2 380.4 ;
        RECT  -38.4 379.2 -37.2 381.3 ;
        RECT  -47.4 381.3 -36.0 382.5 ;
        RECT  -47.4 369.9 -36.0 371.1 ;
        RECT  -47.4 381.3 -36.0 382.5 ;
        RECT  -31.95 396.9 -30.75 398.1 ;
        RECT  -31.95 419.7 -30.75 420.9 ;
        RECT  -31.95 408.9 -30.75 410.1 ;
        RECT  -31.95 369.3 -30.75 370.5 ;
        RECT  -31.8 425.1 -30.6 426.3 ;
        RECT  -47.4 425.1 -46.2 426.3 ;
        RECT  -25.35 395.7 -24.15 396.9 ;
        RECT  -34.05 382.2 -32.85 383.4 ;
        RECT  -34.05 374.7 -32.85 375.9 ;
        RECT  -40.8 374.7 -39.6 375.9 ;
        RECT  -9.75 284.25 -8.55 285.45 ;
        RECT  -9.75 243.45 -8.55 244.65 ;
        RECT  -20.4 204.45 -19.2 205.65 ;
        RECT  -24.75 284.25 -23.55 285.45 ;
        RECT  -27.45 289.65 -26.25 290.85 ;
        RECT  -24.0 327.0 -22.8 328.2 ;
        RECT  -26.7 330.0 -25.5 331.2 ;
        RECT  -12.9 303.15 -11.7 304.35 ;
        RECT  -10.95 300.45 -9.75 301.65 ;
        RECT  -9.0 292.35 -7.8 293.55 ;
        RECT  -41.1 303.15 -39.9 304.35 ;
        RECT  -39.15 292.35 -37.95 293.55 ;
        RECT  -37.2 295.05 -36.0 296.25 ;
        RECT  -24.75 322.5 -23.55 323.7 ;
        RECT  -24.0 339.6 -22.8 340.8 ;
        RECT  -38.25 362.1 -37.05 363.3 ;
        RECT  -25.35 342.3 -24.15 343.5 ;
        RECT  -3.6 286.95 -2.4 288.15 ;
        RECT  -17.7 297.75 -16.5 298.95 ;
        RECT  -31.8 286.95 -30.6 288.15 ;
        RECT  -45.9 297.75 -44.7 298.95 ;
        RECT  1.65 297.75 2.85 298.95 ;
        LAYER  via1 ;
        RECT  128.7 199.5 129.3 200.1 ;
        RECT  124.5 199.5 125.1 200.1 ;
        RECT  132.6 208.8 133.2 209.4 ;
        RECT  123.6 208.8 124.2 209.4 ;
        RECT  128.7 226.5 129.3 227.1 ;
        RECT  124.5 226.5 125.1 227.1 ;
        RECT  132.6 217.2 133.2 217.8 ;
        RECT  123.6 217.2 124.2 217.8 ;
        RECT  128.7 227.7 129.3 228.3 ;
        RECT  124.5 227.7 125.1 228.3 ;
        RECT  132.6 237.0 133.2 237.6 ;
        RECT  123.6 237.0 124.2 237.6 ;
        RECT  128.7 254.7 129.3 255.3 ;
        RECT  124.5 254.7 125.1 255.3 ;
        RECT  132.6 245.4 133.2 246.0 ;
        RECT  123.6 245.4 124.2 246.0 ;
        RECT  128.7 255.9 129.3 256.5 ;
        RECT  124.5 255.9 125.1 256.5 ;
        RECT  132.6 265.2 133.2 265.8 ;
        RECT  123.6 265.2 124.2 265.8 ;
        RECT  128.7 282.9 129.3 283.5 ;
        RECT  124.5 282.9 125.1 283.5 ;
        RECT  132.6 273.6 133.2 274.2 ;
        RECT  123.6 273.6 124.2 274.2 ;
        RECT  128.7 284.1 129.3 284.7 ;
        RECT  124.5 284.1 125.1 284.7 ;
        RECT  132.6 293.4 133.2 294.0 ;
        RECT  123.6 293.4 124.2 294.0 ;
        RECT  128.7 311.1 129.3 311.7 ;
        RECT  124.5 311.1 125.1 311.7 ;
        RECT  132.6 301.8 133.2 302.4 ;
        RECT  123.6 301.8 124.2 302.4 ;
        RECT  128.7 312.3 129.3 312.9 ;
        RECT  124.5 312.3 125.1 312.9 ;
        RECT  132.6 321.6 133.2 322.2 ;
        RECT  123.6 321.6 124.2 322.2 ;
        RECT  128.7 339.3 129.3 339.9 ;
        RECT  124.5 339.3 125.1 339.9 ;
        RECT  132.6 330.0 133.2 330.6 ;
        RECT  123.6 330.0 124.2 330.6 ;
        RECT  128.7 340.5 129.3 341.1 ;
        RECT  124.5 340.5 125.1 341.1 ;
        RECT  132.6 349.8 133.2 350.4 ;
        RECT  123.6 349.8 124.2 350.4 ;
        RECT  128.7 367.5 129.3 368.1 ;
        RECT  124.5 367.5 125.1 368.1 ;
        RECT  132.6 358.2 133.2 358.8 ;
        RECT  123.6 358.2 124.2 358.8 ;
        RECT  128.7 368.7 129.3 369.3 ;
        RECT  124.5 368.7 125.1 369.3 ;
        RECT  132.6 378.0 133.2 378.6 ;
        RECT  123.6 378.0 124.2 378.6 ;
        RECT  128.7 395.7 129.3 396.3 ;
        RECT  124.5 395.7 125.1 396.3 ;
        RECT  132.6 386.4 133.2 387.0 ;
        RECT  123.6 386.4 124.2 387.0 ;
        RECT  128.7 396.9 129.3 397.5 ;
        RECT  124.5 396.9 125.1 397.5 ;
        RECT  132.6 406.2 133.2 406.8 ;
        RECT  123.6 406.2 124.2 406.8 ;
        RECT  128.7 423.9 129.3 424.5 ;
        RECT  124.5 423.9 125.1 424.5 ;
        RECT  132.6 414.6 133.2 415.2 ;
        RECT  123.6 414.6 124.2 415.2 ;
        RECT  138.9 199.5 139.5 200.1 ;
        RECT  134.7 199.5 135.3 200.1 ;
        RECT  142.8 208.8 143.4 209.4 ;
        RECT  133.8 208.8 134.4 209.4 ;
        RECT  138.9 226.5 139.5 227.1 ;
        RECT  134.7 226.5 135.3 227.1 ;
        RECT  142.8 217.2 143.4 217.8 ;
        RECT  133.8 217.2 134.4 217.8 ;
        RECT  138.9 227.7 139.5 228.3 ;
        RECT  134.7 227.7 135.3 228.3 ;
        RECT  142.8 237.0 143.4 237.6 ;
        RECT  133.8 237.0 134.4 237.6 ;
        RECT  138.9 254.7 139.5 255.3 ;
        RECT  134.7 254.7 135.3 255.3 ;
        RECT  142.8 245.4 143.4 246.0 ;
        RECT  133.8 245.4 134.4 246.0 ;
        RECT  138.9 255.9 139.5 256.5 ;
        RECT  134.7 255.9 135.3 256.5 ;
        RECT  142.8 265.2 143.4 265.8 ;
        RECT  133.8 265.2 134.4 265.8 ;
        RECT  138.9 282.9 139.5 283.5 ;
        RECT  134.7 282.9 135.3 283.5 ;
        RECT  142.8 273.6 143.4 274.2 ;
        RECT  133.8 273.6 134.4 274.2 ;
        RECT  138.9 284.1 139.5 284.7 ;
        RECT  134.7 284.1 135.3 284.7 ;
        RECT  142.8 293.4 143.4 294.0 ;
        RECT  133.8 293.4 134.4 294.0 ;
        RECT  138.9 311.1 139.5 311.7 ;
        RECT  134.7 311.1 135.3 311.7 ;
        RECT  142.8 301.8 143.4 302.4 ;
        RECT  133.8 301.8 134.4 302.4 ;
        RECT  138.9 312.3 139.5 312.9 ;
        RECT  134.7 312.3 135.3 312.9 ;
        RECT  142.8 321.6 143.4 322.2 ;
        RECT  133.8 321.6 134.4 322.2 ;
        RECT  138.9 339.3 139.5 339.9 ;
        RECT  134.7 339.3 135.3 339.9 ;
        RECT  142.8 330.0 143.4 330.6 ;
        RECT  133.8 330.0 134.4 330.6 ;
        RECT  138.9 340.5 139.5 341.1 ;
        RECT  134.7 340.5 135.3 341.1 ;
        RECT  142.8 349.8 143.4 350.4 ;
        RECT  133.8 349.8 134.4 350.4 ;
        RECT  138.9 367.5 139.5 368.1 ;
        RECT  134.7 367.5 135.3 368.1 ;
        RECT  142.8 358.2 143.4 358.8 ;
        RECT  133.8 358.2 134.4 358.8 ;
        RECT  138.9 368.7 139.5 369.3 ;
        RECT  134.7 368.7 135.3 369.3 ;
        RECT  142.8 378.0 143.4 378.6 ;
        RECT  133.8 378.0 134.4 378.6 ;
        RECT  138.9 395.7 139.5 396.3 ;
        RECT  134.7 395.7 135.3 396.3 ;
        RECT  142.8 386.4 143.4 387.0 ;
        RECT  133.8 386.4 134.4 387.0 ;
        RECT  138.9 396.9 139.5 397.5 ;
        RECT  134.7 396.9 135.3 397.5 ;
        RECT  142.8 406.2 143.4 406.8 ;
        RECT  133.8 406.2 134.4 406.8 ;
        RECT  138.9 423.9 139.5 424.5 ;
        RECT  134.7 423.9 135.3 424.5 ;
        RECT  142.8 414.6 143.4 415.2 ;
        RECT  133.8 414.6 134.4 415.2 ;
        RECT  126.0 427.5 126.6 428.1 ;
        RECT  128.4 427.5 129.0 428.1 ;
        RECT  126.0 436.5 126.6 437.1 ;
        RECT  130.8 436.5 131.4 437.1 ;
        RECT  136.2 427.5 136.8 428.1 ;
        RECT  138.6 427.5 139.2 428.1 ;
        RECT  136.2 436.5 136.8 437.1 ;
        RECT  141.0 436.5 141.6 437.1 ;
        RECT  132.6 193.2 133.2 193.8 ;
        RECT  126.9 163.8 127.5 164.4 ;
        RECT  129.6 163.8 130.2 164.4 ;
        RECT  123.9 153.9 124.5 154.5 ;
        RECT  142.8 193.2 143.4 193.8 ;
        RECT  137.1 163.8 137.7 164.4 ;
        RECT  139.8 163.8 140.4 164.4 ;
        RECT  134.1 153.9 134.7 154.5 ;
        RECT  124.5 147.3 125.1 147.9 ;
        RECT  129.0 146.7 129.6 147.3 ;
        RECT  126.3 137.1 126.9 137.7 ;
        RECT  125.4 125.4 126.0 126.0 ;
        RECT  132.0 114.6 132.6 115.2 ;
        RECT  128.7 109.2 129.3 109.8 ;
        RECT  125.4 99.3 126.0 99.9 ;
        RECT  132.6 95.1 133.2 95.7 ;
        RECT  126.6 93.0 127.2 93.6 ;
        RECT  134.7 147.3 135.3 147.9 ;
        RECT  139.2 146.7 139.8 147.3 ;
        RECT  136.5 137.1 137.1 137.7 ;
        RECT  135.6 125.4 136.2 126.0 ;
        RECT  142.2 114.6 142.8 115.2 ;
        RECT  138.9 109.2 139.5 109.8 ;
        RECT  135.6 99.3 136.2 99.9 ;
        RECT  142.8 95.1 143.4 95.7 ;
        RECT  136.8 93.0 137.4 93.6 ;
        RECT  126.6 84.6 127.2 85.2 ;
        RECT  129.0 80.1 129.6 80.7 ;
        RECT  128.1 76.8 128.7 77.4 ;
        RECT  132.6 76.2 133.2 76.8 ;
        RECT  128.1 74.7 128.7 75.3 ;
        RECT  124.8 73.8 125.4 74.4 ;
        RECT  129.0 70.2 129.6 70.8 ;
        RECT  129.0 67.8 129.6 68.4 ;
        RECT  126.6 64.8 127.2 65.4 ;
        RECT  127.5 61.5 128.1 62.1 ;
        RECT  124.8 60.3 125.4 60.9 ;
        RECT  129.0 54.6 129.6 55.2 ;
        RECT  128.1 51.3 128.7 51.9 ;
        RECT  132.6 50.7 133.2 51.3 ;
        RECT  128.1 48.3 128.7 48.9 ;
        RECT  124.8 47.4 125.4 48.0 ;
        RECT  129.0 43.8 129.6 44.4 ;
        RECT  129.0 41.4 129.6 42.0 ;
        RECT  126.6 38.4 127.2 39.0 ;
        RECT  138.6 84.6 139.2 85.2 ;
        RECT  136.2 80.1 136.8 80.7 ;
        RECT  137.1 76.8 137.7 77.4 ;
        RECT  132.6 76.2 133.2 76.8 ;
        RECT  137.1 74.7 137.7 75.3 ;
        RECT  140.4 73.8 141.0 74.4 ;
        RECT  136.2 70.2 136.8 70.8 ;
        RECT  136.2 67.8 136.8 68.4 ;
        RECT  138.6 64.8 139.2 65.4 ;
        RECT  137.7 61.5 138.3 62.1 ;
        RECT  140.4 60.3 141.0 60.9 ;
        RECT  136.2 54.6 136.8 55.2 ;
        RECT  137.1 51.3 137.7 51.9 ;
        RECT  132.6 50.7 133.2 51.3 ;
        RECT  137.1 48.3 137.7 48.9 ;
        RECT  140.4 47.4 141.0 48.0 ;
        RECT  136.2 43.8 136.8 44.4 ;
        RECT  136.2 41.4 136.8 42.0 ;
        RECT  138.6 38.4 139.2 39.0 ;
        RECT  125.7 44.1 126.3 44.7 ;
        RECT  130.5 40.5 131.1 41.1 ;
        RECT  132.6 36.0 133.2 36.6 ;
        RECT  135.9 44.1 136.5 44.7 ;
        RECT  140.7 40.5 141.3 41.1 ;
        RECT  142.8 36.0 143.4 36.6 ;
        RECT  42.0 74.55 42.6 75.15 ;
        RECT  39.6 83.55 40.2 84.15 ;
        RECT  39.6 78.3 40.2 78.9 ;
        RECT  42.0 124.65 42.6 125.25 ;
        RECT  39.6 115.65 40.2 116.25 ;
        RECT  39.6 120.9 40.2 121.5 ;
        RECT  42.0 102.75 42.6 103.35 ;
        RECT  39.6 111.75 40.2 112.35 ;
        RECT  39.6 106.5 40.2 107.1 ;
        RECT  42.0 152.85 42.6 153.45 ;
        RECT  39.6 143.85 40.2 144.45 ;
        RECT  39.6 149.1 40.2 149.7 ;
        RECT  58.35 96.3 58.95 96.9 ;
        RECT  76.95 91.35 77.55 91.95 ;
        RECT  55.35 110.4 55.95 111.0 ;
        RECT  73.95 106.65 74.55 107.25 ;
        RECT  76.95 115.2 77.55 115.8 ;
        RECT  52.35 115.2 52.95 115.8 ;
        RECT  73.95 129.3 74.55 129.9 ;
        RECT  49.35 129.3 49.95 129.9 ;
        RECT  58.35 92.7 58.95 93.3 ;
        RECT  55.35 90.0 55.95 90.6 ;
        RECT  52.35 105.3 52.95 105.9 ;
        RECT  55.35 108.0 55.95 108.6 ;
        RECT  58.35 120.9 58.95 121.5 ;
        RECT  49.35 118.2 49.95 118.8 ;
        RECT  52.35 133.5 52.95 134.1 ;
        RECT  49.35 136.2 49.95 136.8 ;
        RECT  42.0 130.95 42.6 131.55 ;
        RECT  39.6 139.95 40.2 140.55 ;
        RECT  39.6 134.7 40.2 135.3 ;
        RECT  42.0 181.05 42.6 181.65 ;
        RECT  39.6 172.05 40.2 172.65 ;
        RECT  39.6 177.3 40.2 177.9 ;
        RECT  42.0 159.15 42.6 159.75 ;
        RECT  39.6 168.15 40.2 168.75 ;
        RECT  39.6 162.9 40.2 163.5 ;
        RECT  42.0 209.25 42.6 209.85 ;
        RECT  39.6 200.25 40.2 200.85 ;
        RECT  39.6 205.5 40.2 206.1 ;
        RECT  58.35 152.7 58.95 153.3 ;
        RECT  76.95 147.75 77.55 148.35 ;
        RECT  55.35 166.8 55.95 167.4 ;
        RECT  73.95 163.05 74.55 163.65 ;
        RECT  76.95 171.6 77.55 172.2 ;
        RECT  52.35 171.6 52.95 172.2 ;
        RECT  73.95 185.7 74.55 186.3 ;
        RECT  49.35 185.7 49.95 186.3 ;
        RECT  58.35 149.1 58.95 149.7 ;
        RECT  55.35 146.4 55.95 147.0 ;
        RECT  52.35 161.7 52.95 162.3 ;
        RECT  55.35 164.4 55.95 165.0 ;
        RECT  58.35 177.3 58.95 177.9 ;
        RECT  49.35 174.6 49.95 175.2 ;
        RECT  52.35 189.9 52.95 190.5 ;
        RECT  49.35 192.6 49.95 193.2 ;
        RECT  27.6 210.45 28.2 211.05 ;
        RECT  30.0 201.45 30.6 202.05 ;
        RECT  30.0 206.7 30.6 207.3 ;
        RECT  27.6 216.75 28.2 217.35 ;
        RECT  30.0 225.75 30.6 226.35 ;
        RECT  30.0 220.5 30.6 221.1 ;
        RECT  27.6 238.65 28.2 239.25 ;
        RECT  30.0 229.65 30.6 230.25 ;
        RECT  30.0 234.9 30.6 235.5 ;
        RECT  27.6 244.95 28.2 245.55 ;
        RECT  30.0 253.95 30.6 254.55 ;
        RECT  30.0 248.7 30.6 249.3 ;
        RECT  27.6 266.85 28.2 267.45 ;
        RECT  30.0 257.85 30.6 258.45 ;
        RECT  30.0 263.1 30.6 263.7 ;
        RECT  27.6 273.15 28.2 273.75 ;
        RECT  30.0 282.15 30.6 282.75 ;
        RECT  30.0 276.9 30.6 277.5 ;
        RECT  27.6 295.05 28.2 295.65 ;
        RECT  30.0 286.05 30.6 286.65 ;
        RECT  30.0 291.3 30.6 291.9 ;
        RECT  27.6 301.35 28.2 301.95 ;
        RECT  30.0 310.35 30.6 310.95 ;
        RECT  30.0 305.1 30.6 305.7 ;
        RECT  27.6 323.25 28.2 323.85 ;
        RECT  30.0 314.25 30.6 314.85 ;
        RECT  30.0 319.5 30.6 320.1 ;
        RECT  27.6 329.55 28.2 330.15 ;
        RECT  30.0 338.55 30.6 339.15 ;
        RECT  30.0 333.3 30.6 333.9 ;
        RECT  27.6 351.45 28.2 352.05 ;
        RECT  30.0 342.45 30.6 343.05 ;
        RECT  30.0 347.7 30.6 348.3 ;
        RECT  27.6 357.75 28.2 358.35 ;
        RECT  30.0 366.75 30.6 367.35 ;
        RECT  30.0 361.5 30.6 362.1 ;
        RECT  27.6 379.65 28.2 380.25 ;
        RECT  30.0 370.65 30.6 371.25 ;
        RECT  30.0 375.9 30.6 376.5 ;
        RECT  27.6 385.95 28.2 386.55 ;
        RECT  30.0 394.95 30.6 395.55 ;
        RECT  30.0 389.7 30.6 390.3 ;
        RECT  27.6 407.85 28.2 408.45 ;
        RECT  30.0 398.85 30.6 399.45 ;
        RECT  30.0 404.1 30.6 404.7 ;
        RECT  27.6 414.15 28.2 414.75 ;
        RECT  30.0 423.15 30.6 423.75 ;
        RECT  30.0 417.9 30.6 418.5 ;
        RECT  6.45 92.55 7.05 93.15 ;
        RECT  8.55 107.85 9.15 108.45 ;
        RECT  10.65 120.75 11.25 121.35 ;
        RECT  12.75 136.05 13.35 136.65 ;
        RECT  14.85 148.95 15.45 149.55 ;
        RECT  16.95 164.25 17.55 164.85 ;
        RECT  19.05 177.15 19.65 177.75 ;
        RECT  21.15 192.45 21.75 193.05 ;
        RECT  6.45 206.7 7.05 207.3 ;
        RECT  14.85 204.0 15.45 204.6 ;
        RECT  6.45 219.3 7.05 219.9 ;
        RECT  16.95 222.0 17.55 222.6 ;
        RECT  6.45 234.9 7.05 235.5 ;
        RECT  19.05 232.2 19.65 232.8 ;
        RECT  6.45 247.5 7.05 248.1 ;
        RECT  21.15 250.2 21.75 250.8 ;
        RECT  8.55 263.1 9.15 263.7 ;
        RECT  14.85 260.4 15.45 261.0 ;
        RECT  8.55 275.7 9.15 276.3 ;
        RECT  16.95 278.4 17.55 279.0 ;
        RECT  8.55 291.3 9.15 291.9 ;
        RECT  19.05 288.6 19.65 289.2 ;
        RECT  8.55 303.9 9.15 304.5 ;
        RECT  21.15 306.6 21.75 307.2 ;
        RECT  10.65 319.5 11.25 320.1 ;
        RECT  14.85 316.8 15.45 317.4 ;
        RECT  10.65 332.1 11.25 332.7 ;
        RECT  16.95 334.8 17.55 335.4 ;
        RECT  10.65 347.7 11.25 348.3 ;
        RECT  19.05 345.0 19.65 345.6 ;
        RECT  10.65 360.3 11.25 360.9 ;
        RECT  21.15 363.0 21.75 363.6 ;
        RECT  12.75 375.9 13.35 376.5 ;
        RECT  14.85 373.2 15.45 373.8 ;
        RECT  12.75 388.5 13.35 389.1 ;
        RECT  16.95 391.2 17.55 391.8 ;
        RECT  12.75 404.1 13.35 404.7 ;
        RECT  19.05 401.4 19.65 402.0 ;
        RECT  12.75 416.7 13.35 417.3 ;
        RECT  21.15 419.4 21.75 420.0 ;
        RECT  67.5 210.45 68.1 211.05 ;
        RECT  69.9 201.45 70.5 202.05 ;
        RECT  69.9 206.7 70.5 207.3 ;
        RECT  49.95 205.35 50.55 205.95 ;
        RECT  51.9 203.1 52.5 203.7 ;
        RECT  67.5 204.0 68.1 204.6 ;
        RECT  67.5 216.75 68.1 217.35 ;
        RECT  69.9 225.75 70.5 226.35 ;
        RECT  69.9 220.5 70.5 221.1 ;
        RECT  49.95 220.65 50.55 221.25 ;
        RECT  51.9 222.9 52.5 223.5 ;
        RECT  67.5 222.0 68.1 222.6 ;
        RECT  67.5 238.65 68.1 239.25 ;
        RECT  69.9 229.65 70.5 230.25 ;
        RECT  69.9 234.9 70.5 235.5 ;
        RECT  49.95 233.55 50.55 234.15 ;
        RECT  51.9 231.3 52.5 231.9 ;
        RECT  67.5 232.2 68.1 232.8 ;
        RECT  67.5 244.95 68.1 245.55 ;
        RECT  69.9 253.95 70.5 254.55 ;
        RECT  69.9 248.7 70.5 249.3 ;
        RECT  49.95 248.85 50.55 249.45 ;
        RECT  51.9 251.1 52.5 251.7 ;
        RECT  67.5 250.2 68.1 250.8 ;
        RECT  67.5 266.85 68.1 267.45 ;
        RECT  69.9 257.85 70.5 258.45 ;
        RECT  69.9 263.1 70.5 263.7 ;
        RECT  49.95 261.75 50.55 262.35 ;
        RECT  51.9 259.5 52.5 260.1 ;
        RECT  67.5 260.4 68.1 261.0 ;
        RECT  67.5 273.15 68.1 273.75 ;
        RECT  69.9 282.15 70.5 282.75 ;
        RECT  69.9 276.9 70.5 277.5 ;
        RECT  49.95 277.05 50.55 277.65 ;
        RECT  51.9 279.3 52.5 279.9 ;
        RECT  67.5 278.4 68.1 279.0 ;
        RECT  67.5 295.05 68.1 295.65 ;
        RECT  69.9 286.05 70.5 286.65 ;
        RECT  69.9 291.3 70.5 291.9 ;
        RECT  49.95 289.95 50.55 290.55 ;
        RECT  51.9 287.7 52.5 288.3 ;
        RECT  67.5 288.6 68.1 289.2 ;
        RECT  67.5 301.35 68.1 301.95 ;
        RECT  69.9 310.35 70.5 310.95 ;
        RECT  69.9 305.1 70.5 305.7 ;
        RECT  49.95 305.25 50.55 305.85 ;
        RECT  51.9 307.5 52.5 308.1 ;
        RECT  67.5 306.6 68.1 307.2 ;
        RECT  67.5 323.25 68.1 323.85 ;
        RECT  69.9 314.25 70.5 314.85 ;
        RECT  69.9 319.5 70.5 320.1 ;
        RECT  49.95 318.15 50.55 318.75 ;
        RECT  51.9 315.9 52.5 316.5 ;
        RECT  67.5 316.8 68.1 317.4 ;
        RECT  67.5 329.55 68.1 330.15 ;
        RECT  69.9 338.55 70.5 339.15 ;
        RECT  69.9 333.3 70.5 333.9 ;
        RECT  49.95 333.45 50.55 334.05 ;
        RECT  51.9 335.7 52.5 336.3 ;
        RECT  67.5 334.8 68.1 335.4 ;
        RECT  67.5 351.45 68.1 352.05 ;
        RECT  69.9 342.45 70.5 343.05 ;
        RECT  69.9 347.7 70.5 348.3 ;
        RECT  49.95 346.35 50.55 346.95 ;
        RECT  51.9 344.1 52.5 344.7 ;
        RECT  67.5 345.0 68.1 345.6 ;
        RECT  67.5 357.75 68.1 358.35 ;
        RECT  69.9 366.75 70.5 367.35 ;
        RECT  69.9 361.5 70.5 362.1 ;
        RECT  49.95 361.65 50.55 362.25 ;
        RECT  51.9 363.9 52.5 364.5 ;
        RECT  67.5 363.0 68.1 363.6 ;
        RECT  67.5 379.65 68.1 380.25 ;
        RECT  69.9 370.65 70.5 371.25 ;
        RECT  69.9 375.9 70.5 376.5 ;
        RECT  49.95 374.55 50.55 375.15 ;
        RECT  51.9 372.3 52.5 372.9 ;
        RECT  67.5 373.2 68.1 373.8 ;
        RECT  67.5 385.95 68.1 386.55 ;
        RECT  69.9 394.95 70.5 395.55 ;
        RECT  69.9 389.7 70.5 390.3 ;
        RECT  49.95 389.85 50.55 390.45 ;
        RECT  51.9 392.1 52.5 392.7 ;
        RECT  67.5 391.2 68.1 391.8 ;
        RECT  67.5 407.85 68.1 408.45 ;
        RECT  69.9 398.85 70.5 399.45 ;
        RECT  69.9 404.1 70.5 404.7 ;
        RECT  49.95 402.75 50.55 403.35 ;
        RECT  51.9 400.5 52.5 401.1 ;
        RECT  67.5 401.4 68.1 402.0 ;
        RECT  67.5 414.15 68.1 414.75 ;
        RECT  69.9 423.15 70.5 423.75 ;
        RECT  69.9 417.9 70.5 418.5 ;
        RECT  49.95 418.05 50.55 418.65 ;
        RECT  51.9 420.3 52.5 420.9 ;
        RECT  67.5 419.4 68.1 420.0 ;
        RECT  60.9 76.5 61.5 77.1 ;
        RECT  56.4 74.1 57.0 74.7 ;
        RECT  53.1 75.0 53.7 75.6 ;
        RECT  52.5 70.5 53.1 71.1 ;
        RECT  51.0 75.0 51.6 75.6 ;
        RECT  50.1 78.3 50.7 78.9 ;
        RECT  46.5 74.1 47.1 74.7 ;
        RECT  44.1 74.1 44.7 74.7 ;
        RECT  41.1 76.5 41.7 77.1 ;
        RECT  37.8 75.6 38.4 76.2 ;
        RECT  36.6 78.3 37.2 78.9 ;
        RECT  30.9 74.1 31.5 74.7 ;
        RECT  27.6 75.0 28.2 75.6 ;
        RECT  27.0 70.5 27.6 71.1 ;
        RECT  24.6 75.0 25.2 75.6 ;
        RECT  23.7 78.3 24.3 78.9 ;
        RECT  20.1 74.1 20.7 74.7 ;
        RECT  17.7 74.1 18.3 74.7 ;
        RECT  14.7 76.5 15.3 77.1 ;
        RECT  60.9 64.5 61.5 65.1 ;
        RECT  56.4 66.9 57.0 67.5 ;
        RECT  53.1 66.0 53.7 66.6 ;
        RECT  52.5 70.5 53.1 71.1 ;
        RECT  51.0 66.0 51.6 66.6 ;
        RECT  50.1 62.7 50.7 63.3 ;
        RECT  46.5 66.9 47.1 67.5 ;
        RECT  44.1 66.9 44.7 67.5 ;
        RECT  41.1 64.5 41.7 65.1 ;
        RECT  37.8 65.4 38.4 66.0 ;
        RECT  36.6 62.7 37.2 63.3 ;
        RECT  30.9 66.9 31.5 67.5 ;
        RECT  27.6 66.0 28.2 66.6 ;
        RECT  27.0 70.5 27.6 71.1 ;
        RECT  24.6 66.0 25.2 66.6 ;
        RECT  23.7 62.7 24.3 63.3 ;
        RECT  20.1 66.9 20.7 67.5 ;
        RECT  17.7 66.9 18.3 67.5 ;
        RECT  14.7 64.5 15.3 65.1 ;
        RECT  60.9 56.1 61.5 56.7 ;
        RECT  56.4 53.7 57.0 54.3 ;
        RECT  53.1 54.6 53.7 55.2 ;
        RECT  52.5 50.1 53.1 50.7 ;
        RECT  51.0 54.6 51.6 55.2 ;
        RECT  50.1 57.9 50.7 58.5 ;
        RECT  46.5 53.7 47.1 54.3 ;
        RECT  44.1 53.7 44.7 54.3 ;
        RECT  41.1 56.1 41.7 56.7 ;
        RECT  37.8 55.2 38.4 55.8 ;
        RECT  36.6 57.9 37.2 58.5 ;
        RECT  30.9 53.7 31.5 54.3 ;
        RECT  27.6 54.6 28.2 55.2 ;
        RECT  27.0 50.1 27.6 50.7 ;
        RECT  24.6 54.6 25.2 55.2 ;
        RECT  23.7 57.9 24.3 58.5 ;
        RECT  20.1 53.7 20.7 54.3 ;
        RECT  17.7 53.7 18.3 54.3 ;
        RECT  14.7 56.1 15.3 56.7 ;
        RECT  60.9 44.1 61.5 44.7 ;
        RECT  56.4 46.5 57.0 47.1 ;
        RECT  53.1 45.6 53.7 46.2 ;
        RECT  52.5 50.1 53.1 50.7 ;
        RECT  51.0 45.6 51.6 46.2 ;
        RECT  50.1 42.3 50.7 42.9 ;
        RECT  46.5 46.5 47.1 47.1 ;
        RECT  44.1 46.5 44.7 47.1 ;
        RECT  41.1 44.1 41.7 44.7 ;
        RECT  37.8 45.0 38.4 45.6 ;
        RECT  36.6 42.3 37.2 42.9 ;
        RECT  30.9 46.5 31.5 47.1 ;
        RECT  27.6 45.6 28.2 46.2 ;
        RECT  27.0 50.1 27.6 50.7 ;
        RECT  24.6 45.6 25.2 46.2 ;
        RECT  23.7 42.3 24.3 42.9 ;
        RECT  20.1 46.5 20.7 47.1 ;
        RECT  17.7 46.5 18.3 47.1 ;
        RECT  14.7 44.1 15.3 44.7 ;
        RECT  95.55 198.9 96.15 199.5 ;
        RECT  95.55 227.1 96.15 227.7 ;
        RECT  95.55 255.3 96.15 255.9 ;
        RECT  95.55 283.5 96.15 284.1 ;
        RECT  95.55 311.7 96.15 312.3 ;
        RECT  95.55 339.9 96.15 340.5 ;
        RECT  95.55 368.1 96.15 368.7 ;
        RECT  95.55 396.3 96.15 396.9 ;
        RECT  95.55 424.5 96.15 425.1 ;
        RECT  76.8 88.95 77.4 89.55 ;
        RECT  81.9 88.8 82.5 89.4 ;
        RECT  73.8 103.05 74.4 103.65 ;
        RECT  84.6 102.9 85.2 103.5 ;
        RECT  76.8 145.35 77.4 145.95 ;
        RECT  87.3 145.2 87.9 145.8 ;
        RECT  73.8 159.45 74.4 160.05 ;
        RECT  90.0 159.3 90.6 159.9 ;
        RECT  78.9 86.1 79.5 86.7 ;
        RECT  78.9 114.3 79.5 114.9 ;
        RECT  78.9 142.5 79.5 143.1 ;
        RECT  78.9 170.7 79.5 171.3 ;
        RECT  66.0 75.6 66.6 76.2 ;
        RECT  81.9 75.6 82.5 76.2 ;
        RECT  66.0 65.4 66.6 66.0 ;
        RECT  84.6 65.4 85.2 66.0 ;
        RECT  66.0 55.2 66.6 55.8 ;
        RECT  87.3 55.2 87.9 55.8 ;
        RECT  66.0 45.0 66.6 45.6 ;
        RECT  90.0 45.0 90.6 45.6 ;
        RECT  66.6 70.5 67.2 71.1 ;
        RECT  95.55 70.65 96.15 71.25 ;
        RECT  66.6 50.1 67.2 50.7 ;
        RECT  95.55 50.25 96.15 50.85 ;
        RECT  110.7 32.55 111.3 33.15 ;
        RECT  105.3 28.05 105.9 28.65 ;
        RECT  108.0 25.65 108.6 26.25 ;
        RECT  110.7 429.75 111.3 430.35 ;
        RECT  113.4 97.05 114.0 97.65 ;
        RECT  116.1 195.15 116.7 195.75 ;
        RECT  102.6 82.8 103.2 83.4 ;
        RECT  49.95 426.6 50.55 427.2 ;
        RECT  102.6 426.6 103.2 427.2 ;
        RECT  98.85 23.7 99.45 24.3 ;
        RECT  98.85 193.2 99.45 193.8 ;
        RECT  98.85 95.1 99.45 95.7 ;
        RECT  -49.2 256.8 -48.6 257.4 ;
        RECT  -46.8 252.3 -46.2 252.9 ;
        RECT  -47.7 249.0 -47.1 249.6 ;
        RECT  -43.2 248.4 -42.6 249.0 ;
        RECT  -47.7 246.9 -47.1 247.5 ;
        RECT  -51.0 246.0 -50.4 246.6 ;
        RECT  -46.8 242.4 -46.2 243.0 ;
        RECT  -46.8 240.0 -46.2 240.6 ;
        RECT  -49.2 237.0 -48.6 237.6 ;
        RECT  -48.3 233.7 -47.7 234.3 ;
        RECT  -51.0 232.5 -50.4 233.1 ;
        RECT  -46.8 226.8 -46.2 227.4 ;
        RECT  -47.7 223.5 -47.1 224.1 ;
        RECT  -43.2 222.9 -42.6 223.5 ;
        RECT  -47.7 220.5 -47.1 221.1 ;
        RECT  -51.0 219.6 -50.4 220.2 ;
        RECT  -46.8 216.0 -46.2 216.6 ;
        RECT  -46.8 213.6 -46.2 214.2 ;
        RECT  -49.2 210.6 -48.6 211.2 ;
        RECT  -37.2 256.8 -36.6 257.4 ;
        RECT  -39.6 252.3 -39.0 252.9 ;
        RECT  -38.7 249.0 -38.1 249.6 ;
        RECT  -43.2 248.4 -42.6 249.0 ;
        RECT  -38.7 246.9 -38.1 247.5 ;
        RECT  -35.4 246.0 -34.8 246.6 ;
        RECT  -39.6 242.4 -39.0 243.0 ;
        RECT  -39.6 240.0 -39.0 240.6 ;
        RECT  -37.2 237.0 -36.6 237.6 ;
        RECT  -38.1 233.7 -37.5 234.3 ;
        RECT  -35.4 232.5 -34.8 233.1 ;
        RECT  -39.6 226.8 -39.0 227.4 ;
        RECT  -38.7 223.5 -38.1 224.1 ;
        RECT  -43.2 222.9 -42.6 223.5 ;
        RECT  -38.7 220.5 -38.1 221.1 ;
        RECT  -35.4 219.6 -34.8 220.2 ;
        RECT  -39.6 216.0 -39.0 216.6 ;
        RECT  -39.6 213.6 -39.0 214.2 ;
        RECT  -37.2 210.6 -36.6 211.2 ;
        RECT  -28.8 256.8 -28.2 257.4 ;
        RECT  -26.4 252.3 -25.8 252.9 ;
        RECT  -27.3 249.0 -26.7 249.6 ;
        RECT  -22.8 248.4 -22.2 249.0 ;
        RECT  -27.3 246.9 -26.7 247.5 ;
        RECT  -30.6 246.0 -30.0 246.6 ;
        RECT  -26.4 242.4 -25.8 243.0 ;
        RECT  -26.4 240.0 -25.8 240.6 ;
        RECT  -28.8 237.0 -28.2 237.6 ;
        RECT  -27.9 233.7 -27.3 234.3 ;
        RECT  -30.6 232.5 -30.0 233.1 ;
        RECT  -26.4 226.8 -25.8 227.4 ;
        RECT  -27.3 223.5 -26.7 224.1 ;
        RECT  -22.8 222.9 -22.2 223.5 ;
        RECT  -27.3 220.5 -26.7 221.1 ;
        RECT  -30.6 219.6 -30.0 220.2 ;
        RECT  -26.4 216.0 -25.8 216.6 ;
        RECT  -26.4 213.6 -25.8 214.2 ;
        RECT  -28.8 210.6 -28.2 211.2 ;
        RECT  -15.3 313.2 -14.7 313.8 ;
        RECT  -15.3 318.0 -14.7 318.6 ;
        RECT  -6.0 318.0 -5.4 318.6 ;
        RECT  -12.6 318.0 -12.0 318.6 ;
        RECT  -21.75 315.6 -21.15 316.2 ;
        RECT  -30.75 313.2 -30.15 313.8 ;
        RECT  -25.65 316.5 -25.05 317.1 ;
        RECT  -21.15 330.3 -20.55 330.9 ;
        RECT  -30.15 332.7 -29.55 333.3 ;
        RECT  -24.9 332.7 -24.3 333.3 ;
        RECT  -43.5 322.8 -42.9 323.4 ;
        RECT  -43.5 327.6 -42.9 328.2 ;
        RECT  -34.2 327.6 -33.6 328.2 ;
        RECT  -40.8 327.6 -40.2 328.2 ;
        RECT  -9.75 397.2 -9.15 397.8 ;
        RECT  -25.05 393.6 -24.45 394.2 ;
        RECT  -25.05 403.2 -24.45 403.8 ;
        RECT  -9.75 404.4 -9.15 405.0 ;
        RECT  -9.75 394.8 -9.15 395.4 ;
        RECT  -25.05 396.0 -24.45 396.6 ;
        RECT  -38.1 405.6 -37.5 406.2 ;
        RECT  -47.1 405.6 -46.5 406.2 ;
        RECT  -39.0 396.3 -38.4 396.9 ;
        RECT  -43.2 396.3 -42.6 396.9 ;
        RECT  -43.2 395.1 -42.6 395.7 ;
        RECT  -39.0 395.1 -38.4 395.7 ;
        RECT  -47.1 385.8 -46.5 386.4 ;
        RECT  -38.1 385.8 -37.5 386.4 ;
        RECT  -43.2 368.1 -42.6 368.7 ;
        RECT  -39.0 368.1 -38.4 368.7 ;
        RECT  -47.1 377.4 -46.5 378.0 ;
        RECT  -38.1 377.4 -37.5 378.0 ;
        RECT  -31.65 397.2 -31.05 397.8 ;
        RECT  -31.65 420.0 -31.05 420.6 ;
        RECT  -31.65 409.2 -31.05 409.8 ;
        RECT  -31.65 369.6 -31.05 370.2 ;
        RECT  -31.5 425.4 -30.9 426.0 ;
        RECT  -47.1 425.4 -46.5 426.0 ;
        RECT  -33.75 382.5 -33.15 383.1 ;
        RECT  -33.75 375.0 -33.15 375.6 ;
        RECT  -40.5 375.0 -39.9 375.6 ;
        RECT  -9.45 284.55 -8.85 285.15 ;
        RECT  -9.45 243.75 -8.85 244.35 ;
        RECT  -20.1 204.75 -19.5 205.35 ;
        RECT  -24.45 284.55 -23.85 285.15 ;
        RECT  -27.15 289.95 -26.55 290.55 ;
        RECT  -23.7 327.3 -23.1 327.9 ;
        RECT  -26.4 330.3 -25.8 330.9 ;
        RECT  -12.6 303.45 -12.0 304.05 ;
        RECT  -10.65 300.75 -10.05 301.35 ;
        RECT  -8.7 292.65 -8.1 293.25 ;
        RECT  -40.8 303.45 -40.2 304.05 ;
        RECT  -38.85 292.65 -38.25 293.25 ;
        RECT  -36.9 295.35 -36.3 295.95 ;
        RECT  -24.45 322.8 -23.85 323.4 ;
        RECT  -23.7 339.9 -23.1 340.5 ;
        RECT  -37.95 362.4 -37.35 363.0 ;
        RECT  -25.05 342.6 -24.45 343.2 ;
        RECT  -3.3 287.25 -2.7 287.85 ;
        RECT  -17.4 298.05 -16.8 298.65 ;
        RECT  -31.5 287.25 -30.9 287.85 ;
        RECT  -45.6 298.05 -45.0 298.65 ;
        RECT  1.95 298.05 2.55 298.65 ;
        LAYER  metal2 ;
        RECT  115.95 340.2 116.85 342.9 ;
        RECT  113.25 360.0 114.15 362.7 ;
        RECT  107.85 320.4 108.75 323.1 ;
        RECT  105.15 337.5 106.05 340.2 ;
        RECT  110.55 301.05 111.45 303.75 ;
        RECT  102.45 282.15 103.35 284.85 ;
        RECT  -3.0 297.9 2.25 298.8 ;
        RECT  97.05 284.85 97.95 287.55 ;
        RECT  127.2 0.0 128.1 1.8 ;
        RECT  137.4 0.0 138.3 1.8 ;
        RECT  95.25 0.0 99.75 444.6 ;
        RECT  102.45 0.0 103.35 444.6 ;
        RECT  105.15 0.0 106.05 444.6 ;
        RECT  107.85 0.0 108.75 444.6 ;
        RECT  110.55 0.0 111.45 444.6 ;
        RECT  113.25 0.0 114.15 444.6 ;
        RECT  115.95 0.0 116.85 444.6 ;
        RECT  81.75 34.8 82.65 199.2 ;
        RECT  84.45 34.8 85.35 199.2 ;
        RECT  87.15 34.8 88.05 199.2 ;
        RECT  89.85 34.8 90.75 199.2 ;
        RECT  127.35 5.85 128.25 6.75 ;
        RECT  124.2 5.85 127.8 6.75 ;
        RECT  127.35 6.3 128.25 8.1 ;
        RECT  137.55 5.85 138.45 6.75 ;
        RECT  134.4 5.85 138.0 6.75 ;
        RECT  137.55 6.3 138.45 8.1 ;
        RECT  49.8 424.8 50.7 426.9 ;
        RECT  127.2 0.0 128.1 1.8 ;
        RECT  137.4 0.0 138.3 1.8 ;
        RECT  113.25 0.0 114.15 444.6 ;
        RECT  110.55 0.0 111.45 444.6 ;
        RECT  102.45 0.0 103.35 444.6 ;
        RECT  115.95 0.0 116.85 444.6 ;
        RECT  105.15 0.0 106.05 444.6 ;
        RECT  95.25 0.0 99.75 444.6 ;
        RECT  107.85 0.0 108.75 444.6 ;
        RECT  128.7 199.2 129.9 424.8 ;
        RECT  135.9 199.2 137.1 424.8 ;
        RECT  138.9 199.2 140.1 424.8 ;
        RECT  125.7 199.2 126.9 424.8 ;
        RECT  132.3 199.2 133.5 424.8 ;
        RECT  132.3 199.2 133.5 213.9 ;
        RECT  128.4 199.2 129.9 200.4 ;
        RECT  124.2 199.2 126.9 200.4 ;
        RECT  128.7 199.2 129.9 213.9 ;
        RECT  125.7 199.2 126.9 212.7 ;
        RECT  122.1 203.4 124.5 213.9 ;
        RECT  125.7 199.2 126.9 212.7 ;
        RECT  132.3 199.2 133.5 213.9 ;
        RECT  122.1 203.4 124.5 213.9 ;
        RECT  128.7 199.2 129.9 213.9 ;
        RECT  132.3 212.7 133.5 227.4 ;
        RECT  128.4 226.2 129.9 227.4 ;
        RECT  124.2 226.2 126.9 227.4 ;
        RECT  128.7 212.7 129.9 227.4 ;
        RECT  125.7 213.9 126.9 227.4 ;
        RECT  122.1 212.7 124.5 223.2 ;
        RECT  125.7 213.9 126.9 227.4 ;
        RECT  132.3 212.7 133.5 227.4 ;
        RECT  122.1 212.7 124.5 223.2 ;
        RECT  128.7 212.7 129.9 227.4 ;
        RECT  132.3 227.4 133.5 242.1 ;
        RECT  128.4 227.4 129.9 228.6 ;
        RECT  124.2 227.4 126.9 228.6 ;
        RECT  128.7 227.4 129.9 242.1 ;
        RECT  125.7 227.4 126.9 240.9 ;
        RECT  122.1 231.6 124.5 242.1 ;
        RECT  125.7 227.4 126.9 240.9 ;
        RECT  132.3 227.4 133.5 242.1 ;
        RECT  122.1 231.6 124.5 242.1 ;
        RECT  128.7 227.4 129.9 242.1 ;
        RECT  132.3 240.9 133.5 255.6 ;
        RECT  128.4 254.4 129.9 255.6 ;
        RECT  124.2 254.4 126.9 255.6 ;
        RECT  128.7 240.9 129.9 255.6 ;
        RECT  125.7 242.1 126.9 255.6 ;
        RECT  122.1 240.9 124.5 251.4 ;
        RECT  125.7 242.1 126.9 255.6 ;
        RECT  132.3 240.9 133.5 255.6 ;
        RECT  122.1 240.9 124.5 251.4 ;
        RECT  128.7 240.9 129.9 255.6 ;
        RECT  132.3 255.6 133.5 270.3 ;
        RECT  128.4 255.6 129.9 256.8 ;
        RECT  124.2 255.6 126.9 256.8 ;
        RECT  128.7 255.6 129.9 270.3 ;
        RECT  125.7 255.6 126.9 269.1 ;
        RECT  122.1 259.8 124.5 270.3 ;
        RECT  125.7 255.6 126.9 269.1 ;
        RECT  132.3 255.6 133.5 270.3 ;
        RECT  122.1 259.8 124.5 270.3 ;
        RECT  128.7 255.6 129.9 270.3 ;
        RECT  132.3 269.1 133.5 283.8 ;
        RECT  128.4 282.6 129.9 283.8 ;
        RECT  124.2 282.6 126.9 283.8 ;
        RECT  128.7 269.1 129.9 283.8 ;
        RECT  125.7 270.3 126.9 283.8 ;
        RECT  122.1 269.1 124.5 279.6 ;
        RECT  125.7 270.3 126.9 283.8 ;
        RECT  132.3 269.1 133.5 283.8 ;
        RECT  122.1 269.1 124.5 279.6 ;
        RECT  128.7 269.1 129.9 283.8 ;
        RECT  132.3 283.8 133.5 298.5 ;
        RECT  128.4 283.8 129.9 285.0 ;
        RECT  124.2 283.8 126.9 285.0 ;
        RECT  128.7 283.8 129.9 298.5 ;
        RECT  125.7 283.8 126.9 297.3 ;
        RECT  122.1 288.0 124.5 298.5 ;
        RECT  125.7 283.8 126.9 297.3 ;
        RECT  132.3 283.8 133.5 298.5 ;
        RECT  122.1 288.0 124.5 298.5 ;
        RECT  128.7 283.8 129.9 298.5 ;
        RECT  132.3 297.3 133.5 312.0 ;
        RECT  128.4 310.8 129.9 312.0 ;
        RECT  124.2 310.8 126.9 312.0 ;
        RECT  128.7 297.3 129.9 312.0 ;
        RECT  125.7 298.5 126.9 312.0 ;
        RECT  122.1 297.3 124.5 307.8 ;
        RECT  125.7 298.5 126.9 312.0 ;
        RECT  132.3 297.3 133.5 312.0 ;
        RECT  122.1 297.3 124.5 307.8 ;
        RECT  128.7 297.3 129.9 312.0 ;
        RECT  132.3 312.0 133.5 326.7 ;
        RECT  128.4 312.0 129.9 313.2 ;
        RECT  124.2 312.0 126.9 313.2 ;
        RECT  128.7 312.0 129.9 326.7 ;
        RECT  125.7 312.0 126.9 325.5 ;
        RECT  122.1 316.2 124.5 326.7 ;
        RECT  125.7 312.0 126.9 325.5 ;
        RECT  132.3 312.0 133.5 326.7 ;
        RECT  122.1 316.2 124.5 326.7 ;
        RECT  128.7 312.0 129.9 326.7 ;
        RECT  132.3 325.5 133.5 340.2 ;
        RECT  128.4 339.0 129.9 340.2 ;
        RECT  124.2 339.0 126.9 340.2 ;
        RECT  128.7 325.5 129.9 340.2 ;
        RECT  125.7 326.7 126.9 340.2 ;
        RECT  122.1 325.5 124.5 336.0 ;
        RECT  125.7 326.7 126.9 340.2 ;
        RECT  132.3 325.5 133.5 340.2 ;
        RECT  122.1 325.5 124.5 336.0 ;
        RECT  128.7 325.5 129.9 340.2 ;
        RECT  132.3 340.2 133.5 354.9 ;
        RECT  128.4 340.2 129.9 341.4 ;
        RECT  124.2 340.2 126.9 341.4 ;
        RECT  128.7 340.2 129.9 354.9 ;
        RECT  125.7 340.2 126.9 353.7 ;
        RECT  122.1 344.4 124.5 354.9 ;
        RECT  125.7 340.2 126.9 353.7 ;
        RECT  132.3 340.2 133.5 354.9 ;
        RECT  122.1 344.4 124.5 354.9 ;
        RECT  128.7 340.2 129.9 354.9 ;
        RECT  132.3 353.7 133.5 368.4 ;
        RECT  128.4 367.2 129.9 368.4 ;
        RECT  124.2 367.2 126.9 368.4 ;
        RECT  128.7 353.7 129.9 368.4 ;
        RECT  125.7 354.9 126.9 368.4 ;
        RECT  122.1 353.7 124.5 364.2 ;
        RECT  125.7 354.9 126.9 368.4 ;
        RECT  132.3 353.7 133.5 368.4 ;
        RECT  122.1 353.7 124.5 364.2 ;
        RECT  128.7 353.7 129.9 368.4 ;
        RECT  132.3 368.4 133.5 383.1 ;
        RECT  128.4 368.4 129.9 369.6 ;
        RECT  124.2 368.4 126.9 369.6 ;
        RECT  128.7 368.4 129.9 383.1 ;
        RECT  125.7 368.4 126.9 381.9 ;
        RECT  122.1 372.6 124.5 383.1 ;
        RECT  125.7 368.4 126.9 381.9 ;
        RECT  132.3 368.4 133.5 383.1 ;
        RECT  122.1 372.6 124.5 383.1 ;
        RECT  128.7 368.4 129.9 383.1 ;
        RECT  132.3 381.9 133.5 396.6 ;
        RECT  128.4 395.4 129.9 396.6 ;
        RECT  124.2 395.4 126.9 396.6 ;
        RECT  128.7 381.9 129.9 396.6 ;
        RECT  125.7 383.1 126.9 396.6 ;
        RECT  122.1 381.9 124.5 392.4 ;
        RECT  125.7 383.1 126.9 396.6 ;
        RECT  132.3 381.9 133.5 396.6 ;
        RECT  122.1 381.9 124.5 392.4 ;
        RECT  128.7 381.9 129.9 396.6 ;
        RECT  132.3 396.6 133.5 411.3 ;
        RECT  128.4 396.6 129.9 397.8 ;
        RECT  124.2 396.6 126.9 397.8 ;
        RECT  128.7 396.6 129.9 411.3 ;
        RECT  125.7 396.6 126.9 410.1 ;
        RECT  122.1 400.8 124.5 411.3 ;
        RECT  125.7 396.6 126.9 410.1 ;
        RECT  132.3 396.6 133.5 411.3 ;
        RECT  122.1 400.8 124.5 411.3 ;
        RECT  128.7 396.6 129.9 411.3 ;
        RECT  132.3 410.1 133.5 424.8 ;
        RECT  128.4 423.6 129.9 424.8 ;
        RECT  124.2 423.6 126.9 424.8 ;
        RECT  128.7 410.1 129.9 424.8 ;
        RECT  125.7 411.3 126.9 424.8 ;
        RECT  122.1 410.1 124.5 420.6 ;
        RECT  125.7 411.3 126.9 424.8 ;
        RECT  132.3 410.1 133.5 424.8 ;
        RECT  122.1 410.1 124.5 420.6 ;
        RECT  128.7 410.1 129.9 424.8 ;
        RECT  142.5 199.2 143.7 213.9 ;
        RECT  138.6 199.2 140.1 200.4 ;
        RECT  134.4 199.2 137.1 200.4 ;
        RECT  138.9 199.2 140.1 213.9 ;
        RECT  135.9 199.2 137.1 212.7 ;
        RECT  132.3 203.4 134.7 213.9 ;
        RECT  135.9 199.2 137.1 212.7 ;
        RECT  142.5 199.2 143.7 213.9 ;
        RECT  132.3 203.4 134.7 213.9 ;
        RECT  138.9 199.2 140.1 213.9 ;
        RECT  142.5 212.7 143.7 227.4 ;
        RECT  138.6 226.2 140.1 227.4 ;
        RECT  134.4 226.2 137.1 227.4 ;
        RECT  138.9 212.7 140.1 227.4 ;
        RECT  135.9 213.9 137.1 227.4 ;
        RECT  132.3 212.7 134.7 223.2 ;
        RECT  135.9 213.9 137.1 227.4 ;
        RECT  142.5 212.7 143.7 227.4 ;
        RECT  132.3 212.7 134.7 223.2 ;
        RECT  138.9 212.7 140.1 227.4 ;
        RECT  142.5 227.4 143.7 242.1 ;
        RECT  138.6 227.4 140.1 228.6 ;
        RECT  134.4 227.4 137.1 228.6 ;
        RECT  138.9 227.4 140.1 242.1 ;
        RECT  135.9 227.4 137.1 240.9 ;
        RECT  132.3 231.6 134.7 242.1 ;
        RECT  135.9 227.4 137.1 240.9 ;
        RECT  142.5 227.4 143.7 242.1 ;
        RECT  132.3 231.6 134.7 242.1 ;
        RECT  138.9 227.4 140.1 242.1 ;
        RECT  142.5 240.9 143.7 255.6 ;
        RECT  138.6 254.4 140.1 255.6 ;
        RECT  134.4 254.4 137.1 255.6 ;
        RECT  138.9 240.9 140.1 255.6 ;
        RECT  135.9 242.1 137.1 255.6 ;
        RECT  132.3 240.9 134.7 251.4 ;
        RECT  135.9 242.1 137.1 255.6 ;
        RECT  142.5 240.9 143.7 255.6 ;
        RECT  132.3 240.9 134.7 251.4 ;
        RECT  138.9 240.9 140.1 255.6 ;
        RECT  142.5 255.6 143.7 270.3 ;
        RECT  138.6 255.6 140.1 256.8 ;
        RECT  134.4 255.6 137.1 256.8 ;
        RECT  138.9 255.6 140.1 270.3 ;
        RECT  135.9 255.6 137.1 269.1 ;
        RECT  132.3 259.8 134.7 270.3 ;
        RECT  135.9 255.6 137.1 269.1 ;
        RECT  142.5 255.6 143.7 270.3 ;
        RECT  132.3 259.8 134.7 270.3 ;
        RECT  138.9 255.6 140.1 270.3 ;
        RECT  142.5 269.1 143.7 283.8 ;
        RECT  138.6 282.6 140.1 283.8 ;
        RECT  134.4 282.6 137.1 283.8 ;
        RECT  138.9 269.1 140.1 283.8 ;
        RECT  135.9 270.3 137.1 283.8 ;
        RECT  132.3 269.1 134.7 279.6 ;
        RECT  135.9 270.3 137.1 283.8 ;
        RECT  142.5 269.1 143.7 283.8 ;
        RECT  132.3 269.1 134.7 279.6 ;
        RECT  138.9 269.1 140.1 283.8 ;
        RECT  142.5 283.8 143.7 298.5 ;
        RECT  138.6 283.8 140.1 285.0 ;
        RECT  134.4 283.8 137.1 285.0 ;
        RECT  138.9 283.8 140.1 298.5 ;
        RECT  135.9 283.8 137.1 297.3 ;
        RECT  132.3 288.0 134.7 298.5 ;
        RECT  135.9 283.8 137.1 297.3 ;
        RECT  142.5 283.8 143.7 298.5 ;
        RECT  132.3 288.0 134.7 298.5 ;
        RECT  138.9 283.8 140.1 298.5 ;
        RECT  142.5 297.3 143.7 312.0 ;
        RECT  138.6 310.8 140.1 312.0 ;
        RECT  134.4 310.8 137.1 312.0 ;
        RECT  138.9 297.3 140.1 312.0 ;
        RECT  135.9 298.5 137.1 312.0 ;
        RECT  132.3 297.3 134.7 307.8 ;
        RECT  135.9 298.5 137.1 312.0 ;
        RECT  142.5 297.3 143.7 312.0 ;
        RECT  132.3 297.3 134.7 307.8 ;
        RECT  138.9 297.3 140.1 312.0 ;
        RECT  142.5 312.0 143.7 326.7 ;
        RECT  138.6 312.0 140.1 313.2 ;
        RECT  134.4 312.0 137.1 313.2 ;
        RECT  138.9 312.0 140.1 326.7 ;
        RECT  135.9 312.0 137.1 325.5 ;
        RECT  132.3 316.2 134.7 326.7 ;
        RECT  135.9 312.0 137.1 325.5 ;
        RECT  142.5 312.0 143.7 326.7 ;
        RECT  132.3 316.2 134.7 326.7 ;
        RECT  138.9 312.0 140.1 326.7 ;
        RECT  142.5 325.5 143.7 340.2 ;
        RECT  138.6 339.0 140.1 340.2 ;
        RECT  134.4 339.0 137.1 340.2 ;
        RECT  138.9 325.5 140.1 340.2 ;
        RECT  135.9 326.7 137.1 340.2 ;
        RECT  132.3 325.5 134.7 336.0 ;
        RECT  135.9 326.7 137.1 340.2 ;
        RECT  142.5 325.5 143.7 340.2 ;
        RECT  132.3 325.5 134.7 336.0 ;
        RECT  138.9 325.5 140.1 340.2 ;
        RECT  142.5 340.2 143.7 354.9 ;
        RECT  138.6 340.2 140.1 341.4 ;
        RECT  134.4 340.2 137.1 341.4 ;
        RECT  138.9 340.2 140.1 354.9 ;
        RECT  135.9 340.2 137.1 353.7 ;
        RECT  132.3 344.4 134.7 354.9 ;
        RECT  135.9 340.2 137.1 353.7 ;
        RECT  142.5 340.2 143.7 354.9 ;
        RECT  132.3 344.4 134.7 354.9 ;
        RECT  138.9 340.2 140.1 354.9 ;
        RECT  142.5 353.7 143.7 368.4 ;
        RECT  138.6 367.2 140.1 368.4 ;
        RECT  134.4 367.2 137.1 368.4 ;
        RECT  138.9 353.7 140.1 368.4 ;
        RECT  135.9 354.9 137.1 368.4 ;
        RECT  132.3 353.7 134.7 364.2 ;
        RECT  135.9 354.9 137.1 368.4 ;
        RECT  142.5 353.7 143.7 368.4 ;
        RECT  132.3 353.7 134.7 364.2 ;
        RECT  138.9 353.7 140.1 368.4 ;
        RECT  142.5 368.4 143.7 383.1 ;
        RECT  138.6 368.4 140.1 369.6 ;
        RECT  134.4 368.4 137.1 369.6 ;
        RECT  138.9 368.4 140.1 383.1 ;
        RECT  135.9 368.4 137.1 381.9 ;
        RECT  132.3 372.6 134.7 383.1 ;
        RECT  135.9 368.4 137.1 381.9 ;
        RECT  142.5 368.4 143.7 383.1 ;
        RECT  132.3 372.6 134.7 383.1 ;
        RECT  138.9 368.4 140.1 383.1 ;
        RECT  142.5 381.9 143.7 396.6 ;
        RECT  138.6 395.4 140.1 396.6 ;
        RECT  134.4 395.4 137.1 396.6 ;
        RECT  138.9 381.9 140.1 396.6 ;
        RECT  135.9 383.1 137.1 396.6 ;
        RECT  132.3 381.9 134.7 392.4 ;
        RECT  135.9 383.1 137.1 396.6 ;
        RECT  142.5 381.9 143.7 396.6 ;
        RECT  132.3 381.9 134.7 392.4 ;
        RECT  138.9 381.9 140.1 396.6 ;
        RECT  142.5 396.6 143.7 411.3 ;
        RECT  138.6 396.6 140.1 397.8 ;
        RECT  134.4 396.6 137.1 397.8 ;
        RECT  138.9 396.6 140.1 411.3 ;
        RECT  135.9 396.6 137.1 410.1 ;
        RECT  132.3 400.8 134.7 411.3 ;
        RECT  135.9 396.6 137.1 410.1 ;
        RECT  142.5 396.6 143.7 411.3 ;
        RECT  132.3 400.8 134.7 411.3 ;
        RECT  138.9 396.6 140.1 411.3 ;
        RECT  142.5 410.1 143.7 424.8 ;
        RECT  138.6 423.6 140.1 424.8 ;
        RECT  134.4 423.6 137.1 424.8 ;
        RECT  138.9 410.1 140.1 424.8 ;
        RECT  135.9 411.3 137.1 424.8 ;
        RECT  132.3 410.1 134.7 420.6 ;
        RECT  135.9 411.3 137.1 424.8 ;
        RECT  142.5 410.1 143.7 424.8 ;
        RECT  132.3 410.1 134.7 420.6 ;
        RECT  138.9 410.1 140.1 424.8 ;
        RECT  136.05 424.8 136.95 444.6 ;
        RECT  125.85 424.8 126.75 444.6 ;
        RECT  139.05 424.8 139.95 444.6 ;
        RECT  128.85 424.8 129.75 444.6 ;
        RECT  125.7 427.2 126.9 428.4 ;
        RECT  128.1 427.2 129.75 428.4 ;
        RECT  125.7 436.2 126.9 437.4 ;
        RECT  128.85 436.2 131.7 437.4 ;
        RECT  125.85 424.8 126.75 444.6 ;
        RECT  128.85 424.8 129.75 444.6 ;
        RECT  125.7 427.2 126.9 428.4 ;
        RECT  128.1 427.2 129.3 428.4 ;
        RECT  125.7 436.2 126.9 437.4 ;
        RECT  130.5 436.2 131.7 437.4 ;
        RECT  135.9 427.2 137.1 428.4 ;
        RECT  138.3 427.2 139.95 428.4 ;
        RECT  135.9 436.2 137.1 437.4 ;
        RECT  139.05 436.2 141.9 437.4 ;
        RECT  136.05 424.8 136.95 444.6 ;
        RECT  139.05 424.8 139.95 444.6 ;
        RECT  135.9 427.2 137.1 428.4 ;
        RECT  138.3 427.2 139.5 428.4 ;
        RECT  135.9 436.2 137.1 437.4 ;
        RECT  140.7 436.2 141.9 437.4 ;
        RECT  135.9 150.3 137.1 163.5 ;
        RECT  125.7 150.3 126.9 163.5 ;
        RECT  138.9 150.3 140.1 163.5 ;
        RECT  128.7 150.3 129.9 163.5 ;
        RECT  125.7 164.7 126.9 199.2 ;
        RECT  128.7 164.7 129.9 199.2 ;
        RECT  132.3 191.7 133.5 199.2 ;
        RECT  125.7 163.5 127.8 164.7 ;
        RECT  128.7 163.5 130.5 164.7 ;
        RECT  123.6 150.3 124.8 154.8 ;
        RECT  125.7 150.3 126.9 163.5 ;
        RECT  128.7 150.3 129.9 163.5 ;
        RECT  128.7 150.3 129.9 163.5 ;
        RECT  125.7 150.3 126.9 163.5 ;
        RECT  135.9 164.7 137.1 199.2 ;
        RECT  138.9 164.7 140.1 199.2 ;
        RECT  142.5 191.7 143.7 199.2 ;
        RECT  135.9 163.5 138.0 164.7 ;
        RECT  138.9 163.5 140.7 164.7 ;
        RECT  133.8 150.3 135.0 154.8 ;
        RECT  135.9 150.3 137.1 163.5 ;
        RECT  138.9 150.3 140.1 163.5 ;
        RECT  138.9 150.3 140.1 163.5 ;
        RECT  135.9 150.3 137.1 163.5 ;
        RECT  127.2 90.0 128.4 92.7 ;
        RECT  137.4 90.0 138.6 92.7 ;
        RECT  125.7 148.2 126.9 150.3 ;
        RECT  135.9 148.2 137.1 150.3 ;
        RECT  138.9 142.8 140.1 150.3 ;
        RECT  128.7 142.8 129.9 150.3 ;
        RECT  125.7 148.2 126.9 150.3 ;
        RECT  124.2 147.0 126.9 148.2 ;
        RECT  128.7 142.8 129.9 150.3 ;
        RECT  132.3 138.0 133.5 148.5 ;
        RECT  126.0 136.8 133.5 138.0 ;
        RECT  125.1 99.0 126.3 126.3 ;
        RECT  132.3 115.5 133.5 136.8 ;
        RECT  131.7 114.3 133.5 115.5 ;
        RECT  132.3 111.3 133.5 114.3 ;
        RECT  128.4 110.1 133.5 111.3 ;
        RECT  128.4 108.9 129.6 110.1 ;
        RECT  126.3 92.7 128.7 93.9 ;
        RECT  127.2 90.0 128.4 92.7 ;
        RECT  132.3 90.0 133.5 110.1 ;
        RECT  127.2 90.0 128.4 92.7 ;
        RECT  128.7 142.8 129.9 150.3 ;
        RECT  125.7 148.2 126.9 150.3 ;
        RECT  135.9 148.2 137.1 150.3 ;
        RECT  134.4 147.0 137.1 148.2 ;
        RECT  138.9 142.8 140.1 150.3 ;
        RECT  142.5 138.0 143.7 148.5 ;
        RECT  136.2 136.8 143.7 138.0 ;
        RECT  135.3 99.0 136.5 126.3 ;
        RECT  142.5 115.5 143.7 136.8 ;
        RECT  141.9 114.3 143.7 115.5 ;
        RECT  142.5 111.3 143.7 114.3 ;
        RECT  138.6 110.1 143.7 111.3 ;
        RECT  138.6 108.9 139.8 110.1 ;
        RECT  136.5 92.7 138.9 93.9 ;
        RECT  137.4 90.0 138.6 92.7 ;
        RECT  142.5 90.0 143.7 110.1 ;
        RECT  137.4 90.0 138.6 92.7 ;
        RECT  138.9 142.8 140.1 150.3 ;
        RECT  135.9 148.2 137.1 150.3 ;
        RECT  140.1 85.5 141.3 90.0 ;
        RECT  137.4 30.0 138.6 31.2 ;
        RECT  127.2 30.0 128.4 31.2 ;
        RECT  132.3 30.0 133.5 90.0 ;
        RECT  124.5 85.5 125.7 90.0 ;
        RECT  127.2 88.8 128.4 90.0 ;
        RECT  137.4 88.8 138.6 90.0 ;
        RECT  124.5 85.5 125.7 90.0 ;
        RECT  127.2 88.8 128.4 90.0 ;
        RECT  127.2 87.6 129.9 88.8 ;
        RECT  124.5 84.3 127.5 85.5 ;
        RECT  124.5 74.7 125.4 84.3 ;
        RECT  128.7 79.8 129.9 87.6 ;
        RECT  127.8 76.5 130.8 77.7 ;
        RECT  124.5 73.5 125.7 74.7 ;
        RECT  127.8 74.4 129.0 75.6 ;
        RECT  128.1 72.9 129.0 74.4 ;
        RECT  126.6 72.0 129.0 72.9 ;
        RECT  126.6 65.7 127.5 72.0 ;
        RECT  129.9 71.1 130.8 76.5 ;
        RECT  128.7 69.9 130.8 71.1 ;
        RECT  128.7 67.5 130.8 68.7 ;
        RECT  126.3 64.5 127.5 65.7 ;
        RECT  124.2 60.0 125.7 61.2 ;
        RECT  124.2 48.3 125.1 60.0 ;
        RECT  127.2 57.9 128.4 62.4 ;
        RECT  126.0 57.0 128.4 57.9 ;
        RECT  126.0 50.1 126.9 57.0 ;
        RECT  129.9 55.5 130.8 67.5 ;
        RECT  128.7 54.3 130.8 55.5 ;
        RECT  127.8 51.0 130.8 52.2 ;
        RECT  126.0 49.2 127.5 50.1 ;
        RECT  124.2 47.1 125.7 48.3 ;
        RECT  126.6 48.0 129.0 49.2 ;
        RECT  126.6 39.3 127.5 48.0 ;
        RECT  129.9 44.7 130.8 51.0 ;
        RECT  128.7 43.5 130.8 44.7 ;
        RECT  128.7 41.1 130.8 42.3 ;
        RECT  126.3 38.1 127.5 39.3 ;
        RECT  129.9 32.4 130.8 41.1 ;
        RECT  127.2 31.2 130.8 32.4 ;
        RECT  127.2 30.0 128.4 31.2 ;
        RECT  132.3 30.0 133.5 90.0 ;
        RECT  127.2 30.0 128.4 31.2 ;
        RECT  127.2 88.8 128.4 90.0 ;
        RECT  124.5 85.5 125.7 90.0 ;
        RECT  132.3 30.0 133.5 90.0 ;
        RECT  140.1 85.5 141.3 90.0 ;
        RECT  137.4 88.8 138.6 90.0 ;
        RECT  135.9 87.6 138.6 88.8 ;
        RECT  138.3 84.3 141.3 85.5 ;
        RECT  140.4 74.7 141.3 84.3 ;
        RECT  135.9 79.8 137.1 87.6 ;
        RECT  135.0 76.5 138.0 77.7 ;
        RECT  140.1 73.5 141.3 74.7 ;
        RECT  136.8 74.4 138.0 75.6 ;
        RECT  136.8 72.9 137.7 74.4 ;
        RECT  136.8 72.0 139.2 72.9 ;
        RECT  138.3 65.7 139.2 72.0 ;
        RECT  135.0 71.1 135.9 76.5 ;
        RECT  135.0 69.9 137.1 71.1 ;
        RECT  135.0 67.5 137.1 68.7 ;
        RECT  138.3 64.5 139.5 65.7 ;
        RECT  140.1 60.0 141.6 61.2 ;
        RECT  140.7 48.3 141.6 60.0 ;
        RECT  137.4 57.9 138.6 62.4 ;
        RECT  137.4 57.0 139.8 57.9 ;
        RECT  138.9 50.1 139.8 57.0 ;
        RECT  135.0 55.5 135.9 67.5 ;
        RECT  135.0 54.3 137.1 55.5 ;
        RECT  135.0 51.0 138.0 52.2 ;
        RECT  138.3 49.2 139.8 50.1 ;
        RECT  140.1 47.1 141.6 48.3 ;
        RECT  136.8 48.0 139.2 49.2 ;
        RECT  138.3 39.3 139.2 48.0 ;
        RECT  135.0 44.7 135.9 51.0 ;
        RECT  135.0 43.5 137.1 44.7 ;
        RECT  135.0 41.1 137.1 42.3 ;
        RECT  138.3 38.1 139.5 39.3 ;
        RECT  135.0 32.4 135.9 41.1 ;
        RECT  135.0 31.2 138.6 32.4 ;
        RECT  137.4 30.0 138.6 31.2 ;
        RECT  132.3 30.0 133.5 90.0 ;
        RECT  137.4 30.0 138.6 31.2 ;
        RECT  137.4 88.8 138.6 90.0 ;
        RECT  140.1 85.5 141.3 90.0 ;
        RECT  132.3 30.0 133.5 90.0 ;
        RECT  127.2 8.1 128.4 15.0 ;
        RECT  127.2 28.5 128.4 30.0 ;
        RECT  137.4 28.5 138.6 30.0 ;
        RECT  137.4 8.1 138.6 15.0 ;
        RECT  127.2 45.0 128.4 51.9 ;
        RECT  125.4 43.8 128.4 45.0 ;
        RECT  127.2 40.2 131.4 41.4 ;
        RECT  127.2 32.7 128.4 40.2 ;
        RECT  127.2 31.5 128.7 32.7 ;
        RECT  127.2 30.0 128.4 31.5 ;
        RECT  132.3 30.0 133.5 51.9 ;
        RECT  132.3 30.0 133.5 51.9 ;
        RECT  127.2 45.0 128.4 51.9 ;
        RECT  127.2 30.0 128.4 31.5 ;
        RECT  137.4 45.0 138.6 51.9 ;
        RECT  135.6 43.8 138.6 45.0 ;
        RECT  137.4 40.2 141.6 41.4 ;
        RECT  137.4 32.7 138.6 40.2 ;
        RECT  137.4 31.5 138.9 32.7 ;
        RECT  137.4 30.0 138.6 31.5 ;
        RECT  142.5 30.0 143.7 51.9 ;
        RECT  142.5 30.0 143.7 51.9 ;
        RECT  137.4 45.0 138.6 51.9 ;
        RECT  137.4 30.0 138.6 31.5 ;
        RECT  6.3 86.4 7.2 424.8 ;
        RECT  8.4 86.4 9.3 424.8 ;
        RECT  10.5 86.4 11.4 424.8 ;
        RECT  12.6 86.4 13.5 424.8 ;
        RECT  14.7 86.4 15.6 424.8 ;
        RECT  16.8 86.4 17.7 424.8 ;
        RECT  18.9 86.4 19.8 424.8 ;
        RECT  21.0 86.4 21.9 424.8 ;
        RECT  73.8 142.8 74.7 197.4 ;
        RECT  73.8 86.4 74.7 141.0 ;
        RECT  76.8 86.4 77.7 141.0 ;
        RECT  76.8 142.8 77.7 197.4 ;
        RECT  52.2 86.4 53.1 141.0 ;
        RECT  49.2 86.4 50.1 141.0 ;
        RECT  58.2 86.4 59.1 141.0 ;
        RECT  55.2 86.4 56.1 141.0 ;
        RECT  76.8 86.4 77.7 141.0 ;
        RECT  73.8 86.4 74.7 141.0 ;
        RECT  41.85 78.15 42.75 79.05 ;
        RECT  39.45 78.15 40.35 79.05 ;
        RECT  41.85 75.45 42.75 78.6 ;
        RECT  39.9 78.15 42.3 79.05 ;
        RECT  39.45 78.6 40.35 83.25 ;
        RECT  41.7 74.25 42.9 75.45 ;
        RECT  39.3 83.25 40.5 84.45 ;
        RECT  39.3 78.0 40.5 79.2 ;
        RECT  41.85 121.95 42.75 122.85 ;
        RECT  39.45 121.95 40.35 122.85 ;
        RECT  41.85 122.4 42.75 125.55 ;
        RECT  39.9 121.95 42.3 122.85 ;
        RECT  39.45 117.75 40.35 122.4 ;
        RECT  41.7 124.35 42.9 125.55 ;
        RECT  39.3 115.35 40.5 116.55 ;
        RECT  39.3 120.6 40.5 121.8 ;
        RECT  41.85 106.35 42.75 107.25 ;
        RECT  39.45 106.35 40.35 107.25 ;
        RECT  41.85 103.65 42.75 106.8 ;
        RECT  39.9 106.35 42.3 107.25 ;
        RECT  39.45 106.8 40.35 111.45 ;
        RECT  41.7 102.45 42.9 103.65 ;
        RECT  39.3 111.45 40.5 112.65 ;
        RECT  39.3 106.2 40.5 107.4 ;
        RECT  41.85 150.15 42.75 151.05 ;
        RECT  39.45 150.15 40.35 151.05 ;
        RECT  41.85 150.6 42.75 153.75 ;
        RECT  39.9 150.15 42.3 151.05 ;
        RECT  39.45 145.95 40.35 150.6 ;
        RECT  41.7 152.55 42.9 153.75 ;
        RECT  39.3 143.55 40.5 144.75 ;
        RECT  39.3 148.8 40.5 150.0 ;
        RECT  58.05 96.0 59.25 97.2 ;
        RECT  76.65 91.05 77.85 92.25 ;
        RECT  55.05 110.1 56.25 111.3 ;
        RECT  73.65 106.35 74.85 107.55 ;
        RECT  76.65 114.9 77.85 116.1 ;
        RECT  52.05 114.9 53.25 116.1 ;
        RECT  73.65 129.0 74.85 130.2 ;
        RECT  49.05 129.0 50.25 130.2 ;
        RECT  58.05 92.4 59.25 93.6 ;
        RECT  55.05 89.7 56.25 90.9 ;
        RECT  52.05 105.0 53.25 106.2 ;
        RECT  55.05 107.7 56.25 108.9 ;
        RECT  58.05 120.6 59.25 121.8 ;
        RECT  49.05 117.9 50.25 119.1 ;
        RECT  52.05 133.2 53.25 134.4 ;
        RECT  49.05 135.9 50.25 137.1 ;
        RECT  52.2 142.8 53.1 197.4 ;
        RECT  49.2 142.8 50.1 197.4 ;
        RECT  58.2 142.8 59.1 197.4 ;
        RECT  55.2 142.8 56.1 197.4 ;
        RECT  76.8 142.8 77.7 197.4 ;
        RECT  73.8 142.8 74.7 197.4 ;
        RECT  41.85 134.55 42.75 135.45 ;
        RECT  39.45 134.55 40.35 135.45 ;
        RECT  41.85 131.85 42.75 135.0 ;
        RECT  39.9 134.55 42.3 135.45 ;
        RECT  39.45 135.0 40.35 139.65 ;
        RECT  41.7 130.65 42.9 131.85 ;
        RECT  39.3 139.65 40.5 140.85 ;
        RECT  39.3 134.4 40.5 135.6 ;
        RECT  41.85 178.35 42.75 179.25 ;
        RECT  39.45 178.35 40.35 179.25 ;
        RECT  41.85 178.8 42.75 181.95 ;
        RECT  39.9 178.35 42.3 179.25 ;
        RECT  39.45 174.15 40.35 178.8 ;
        RECT  41.7 180.75 42.9 181.95 ;
        RECT  39.3 171.75 40.5 172.95 ;
        RECT  39.3 177.0 40.5 178.2 ;
        RECT  41.85 162.75 42.75 163.65 ;
        RECT  39.45 162.75 40.35 163.65 ;
        RECT  41.85 160.05 42.75 163.2 ;
        RECT  39.9 162.75 42.3 163.65 ;
        RECT  39.45 163.2 40.35 167.85 ;
        RECT  41.7 158.85 42.9 160.05 ;
        RECT  39.3 167.85 40.5 169.05 ;
        RECT  39.3 162.6 40.5 163.8 ;
        RECT  41.85 206.55 42.75 207.45 ;
        RECT  39.45 206.55 40.35 207.45 ;
        RECT  41.85 207.0 42.75 210.15 ;
        RECT  39.9 206.55 42.3 207.45 ;
        RECT  39.45 202.35 40.35 207.0 ;
        RECT  41.7 208.95 42.9 210.15 ;
        RECT  39.3 199.95 40.5 201.15 ;
        RECT  39.3 205.2 40.5 206.4 ;
        RECT  58.05 152.4 59.25 153.6 ;
        RECT  76.65 147.45 77.85 148.65 ;
        RECT  55.05 166.5 56.25 167.7 ;
        RECT  73.65 162.75 74.85 163.95 ;
        RECT  76.65 171.3 77.85 172.5 ;
        RECT  52.05 171.3 53.25 172.5 ;
        RECT  73.65 185.4 74.85 186.6 ;
        RECT  49.05 185.4 50.25 186.6 ;
        RECT  58.05 148.8 59.25 150.0 ;
        RECT  55.05 146.1 56.25 147.3 ;
        RECT  52.05 161.4 53.25 162.6 ;
        RECT  55.05 164.1 56.25 165.3 ;
        RECT  58.05 177.0 59.25 178.2 ;
        RECT  49.05 174.3 50.25 175.5 ;
        RECT  52.05 189.6 53.25 190.8 ;
        RECT  49.05 192.3 50.25 193.5 ;
        RECT  27.45 206.55 28.35 207.45 ;
        RECT  29.85 206.55 30.75 207.45 ;
        RECT  27.45 207.0 28.35 210.15 ;
        RECT  27.9 206.55 30.3 207.45 ;
        RECT  29.85 202.35 30.75 207.0 ;
        RECT  27.3 210.15 28.5 211.35 ;
        RECT  29.7 201.15 30.9 202.35 ;
        RECT  29.7 206.4 30.9 207.6 ;
        RECT  27.45 219.15 28.35 220.05 ;
        RECT  29.85 219.15 30.75 220.05 ;
        RECT  27.45 216.45 28.35 219.6 ;
        RECT  27.9 219.15 30.3 220.05 ;
        RECT  29.85 219.6 30.75 224.25 ;
        RECT  27.3 216.45 28.5 217.65 ;
        RECT  29.7 225.45 30.9 226.65 ;
        RECT  29.7 220.2 30.9 221.4 ;
        RECT  27.45 234.75 28.35 235.65 ;
        RECT  29.85 234.75 30.75 235.65 ;
        RECT  27.45 235.2 28.35 238.35 ;
        RECT  27.9 234.75 30.3 235.65 ;
        RECT  29.85 230.55 30.75 235.2 ;
        RECT  27.3 238.35 28.5 239.55 ;
        RECT  29.7 229.35 30.9 230.55 ;
        RECT  29.7 234.6 30.9 235.8 ;
        RECT  27.45 247.35 28.35 248.25 ;
        RECT  29.85 247.35 30.75 248.25 ;
        RECT  27.45 244.65 28.35 247.8 ;
        RECT  27.9 247.35 30.3 248.25 ;
        RECT  29.85 247.8 30.75 252.45 ;
        RECT  27.3 244.65 28.5 245.85 ;
        RECT  29.7 253.65 30.9 254.85 ;
        RECT  29.7 248.4 30.9 249.6 ;
        RECT  27.45 262.95 28.35 263.85 ;
        RECT  29.85 262.95 30.75 263.85 ;
        RECT  27.45 263.4 28.35 266.55 ;
        RECT  27.9 262.95 30.3 263.85 ;
        RECT  29.85 258.75 30.75 263.4 ;
        RECT  27.3 266.55 28.5 267.75 ;
        RECT  29.7 257.55 30.9 258.75 ;
        RECT  29.7 262.8 30.9 264.0 ;
        RECT  27.45 275.55 28.35 276.45 ;
        RECT  29.85 275.55 30.75 276.45 ;
        RECT  27.45 272.85 28.35 276.0 ;
        RECT  27.9 275.55 30.3 276.45 ;
        RECT  29.85 276.0 30.75 280.65 ;
        RECT  27.3 272.85 28.5 274.05 ;
        RECT  29.7 281.85 30.9 283.05 ;
        RECT  29.7 276.6 30.9 277.8 ;
        RECT  27.45 291.15 28.35 292.05 ;
        RECT  29.85 291.15 30.75 292.05 ;
        RECT  27.45 291.6 28.35 294.75 ;
        RECT  27.9 291.15 30.3 292.05 ;
        RECT  29.85 286.95 30.75 291.6 ;
        RECT  27.3 294.75 28.5 295.95 ;
        RECT  29.7 285.75 30.9 286.95 ;
        RECT  29.7 291.0 30.9 292.2 ;
        RECT  27.45 303.75 28.35 304.65 ;
        RECT  29.85 303.75 30.75 304.65 ;
        RECT  27.45 301.05 28.35 304.2 ;
        RECT  27.9 303.75 30.3 304.65 ;
        RECT  29.85 304.2 30.75 308.85 ;
        RECT  27.3 301.05 28.5 302.25 ;
        RECT  29.7 310.05 30.9 311.25 ;
        RECT  29.7 304.8 30.9 306.0 ;
        RECT  27.45 319.35 28.35 320.25 ;
        RECT  29.85 319.35 30.75 320.25 ;
        RECT  27.45 319.8 28.35 322.95 ;
        RECT  27.9 319.35 30.3 320.25 ;
        RECT  29.85 315.15 30.75 319.8 ;
        RECT  27.3 322.95 28.5 324.15 ;
        RECT  29.7 313.95 30.9 315.15 ;
        RECT  29.7 319.2 30.9 320.4 ;
        RECT  27.45 331.95 28.35 332.85 ;
        RECT  29.85 331.95 30.75 332.85 ;
        RECT  27.45 329.25 28.35 332.4 ;
        RECT  27.9 331.95 30.3 332.85 ;
        RECT  29.85 332.4 30.75 337.05 ;
        RECT  27.3 329.25 28.5 330.45 ;
        RECT  29.7 338.25 30.9 339.45 ;
        RECT  29.7 333.0 30.9 334.2 ;
        RECT  27.45 347.55 28.35 348.45 ;
        RECT  29.85 347.55 30.75 348.45 ;
        RECT  27.45 348.0 28.35 351.15 ;
        RECT  27.9 347.55 30.3 348.45 ;
        RECT  29.85 343.35 30.75 348.0 ;
        RECT  27.3 351.15 28.5 352.35 ;
        RECT  29.7 342.15 30.9 343.35 ;
        RECT  29.7 347.4 30.9 348.6 ;
        RECT  27.45 360.15 28.35 361.05 ;
        RECT  29.85 360.15 30.75 361.05 ;
        RECT  27.45 357.45 28.35 360.6 ;
        RECT  27.9 360.15 30.3 361.05 ;
        RECT  29.85 360.6 30.75 365.25 ;
        RECT  27.3 357.45 28.5 358.65 ;
        RECT  29.7 366.45 30.9 367.65 ;
        RECT  29.7 361.2 30.9 362.4 ;
        RECT  27.45 375.75 28.35 376.65 ;
        RECT  29.85 375.75 30.75 376.65 ;
        RECT  27.45 376.2 28.35 379.35 ;
        RECT  27.9 375.75 30.3 376.65 ;
        RECT  29.85 371.55 30.75 376.2 ;
        RECT  27.3 379.35 28.5 380.55 ;
        RECT  29.7 370.35 30.9 371.55 ;
        RECT  29.7 375.6 30.9 376.8 ;
        RECT  27.45 388.35 28.35 389.25 ;
        RECT  29.85 388.35 30.75 389.25 ;
        RECT  27.45 385.65 28.35 388.8 ;
        RECT  27.9 388.35 30.3 389.25 ;
        RECT  29.85 388.8 30.75 393.45 ;
        RECT  27.3 385.65 28.5 386.85 ;
        RECT  29.7 394.65 30.9 395.85 ;
        RECT  29.7 389.4 30.9 390.6 ;
        RECT  27.45 403.95 28.35 404.85 ;
        RECT  29.85 403.95 30.75 404.85 ;
        RECT  27.45 404.4 28.35 407.55 ;
        RECT  27.9 403.95 30.3 404.85 ;
        RECT  29.85 399.75 30.75 404.4 ;
        RECT  27.3 407.55 28.5 408.75 ;
        RECT  29.7 398.55 30.9 399.75 ;
        RECT  29.7 403.8 30.9 405.0 ;
        RECT  27.45 416.55 28.35 417.45 ;
        RECT  29.85 416.55 30.75 417.45 ;
        RECT  27.45 413.85 28.35 417.0 ;
        RECT  27.9 416.55 30.3 417.45 ;
        RECT  29.85 417.0 30.75 421.65 ;
        RECT  27.3 413.85 28.5 415.05 ;
        RECT  29.7 422.85 30.9 424.05 ;
        RECT  29.7 417.6 30.9 418.8 ;
        RECT  6.15 92.25 7.35 93.45 ;
        RECT  8.25 107.55 9.45 108.75 ;
        RECT  10.35 120.45 11.55 121.65 ;
        RECT  12.45 135.75 13.65 136.95 ;
        RECT  14.55 148.65 15.75 149.85 ;
        RECT  16.65 163.95 17.85 165.15 ;
        RECT  18.75 176.85 19.95 178.05 ;
        RECT  20.85 192.15 22.05 193.35 ;
        RECT  6.15 206.4 7.35 207.6 ;
        RECT  14.55 203.7 15.75 204.9 ;
        RECT  6.15 219.0 7.35 220.2 ;
        RECT  16.65 221.7 17.85 222.9 ;
        RECT  6.15 234.6 7.35 235.8 ;
        RECT  18.75 231.9 19.95 233.1 ;
        RECT  6.15 247.2 7.35 248.4 ;
        RECT  20.85 249.9 22.05 251.1 ;
        RECT  8.25 262.8 9.45 264.0 ;
        RECT  14.55 260.1 15.75 261.3 ;
        RECT  8.25 275.4 9.45 276.6 ;
        RECT  16.65 278.1 17.85 279.3 ;
        RECT  8.25 291.0 9.45 292.2 ;
        RECT  18.75 288.3 19.95 289.5 ;
        RECT  8.25 303.6 9.45 304.8 ;
        RECT  20.85 306.3 22.05 307.5 ;
        RECT  10.35 319.2 11.55 320.4 ;
        RECT  14.55 316.5 15.75 317.7 ;
        RECT  10.35 331.8 11.55 333.0 ;
        RECT  16.65 334.5 17.85 335.7 ;
        RECT  10.35 347.4 11.55 348.6 ;
        RECT  18.75 344.7 19.95 345.9 ;
        RECT  10.35 360.0 11.55 361.2 ;
        RECT  20.85 362.7 22.05 363.9 ;
        RECT  12.45 375.6 13.65 376.8 ;
        RECT  14.55 372.9 15.75 374.1 ;
        RECT  12.45 388.2 13.65 389.4 ;
        RECT  16.65 390.9 17.85 392.1 ;
        RECT  12.45 403.8 13.65 405.0 ;
        RECT  18.75 401.1 19.95 402.3 ;
        RECT  12.45 416.4 13.65 417.6 ;
        RECT  20.85 419.1 22.05 420.3 ;
        RECT  51.75 203.85 52.65 204.75 ;
        RECT  51.75 203.4 52.65 204.3 ;
        RECT  52.2 203.85 68.4 204.75 ;
        RECT  51.75 221.85 52.65 222.75 ;
        RECT  51.75 222.3 52.65 223.2 ;
        RECT  52.2 221.85 68.4 222.75 ;
        RECT  51.75 232.05 52.65 232.95 ;
        RECT  51.75 231.6 52.65 232.5 ;
        RECT  52.2 232.05 68.4 232.95 ;
        RECT  51.75 250.05 52.65 250.95 ;
        RECT  51.75 250.5 52.65 251.4 ;
        RECT  52.2 250.05 68.4 250.95 ;
        RECT  51.75 260.25 52.65 261.15 ;
        RECT  51.75 259.8 52.65 260.7 ;
        RECT  52.2 260.25 68.4 261.15 ;
        RECT  51.75 278.25 52.65 279.15 ;
        RECT  51.75 278.7 52.65 279.6 ;
        RECT  52.2 278.25 68.4 279.15 ;
        RECT  51.75 288.45 52.65 289.35 ;
        RECT  51.75 288.0 52.65 288.9 ;
        RECT  52.2 288.45 68.4 289.35 ;
        RECT  51.75 306.45 52.65 307.35 ;
        RECT  51.75 306.9 52.65 307.8 ;
        RECT  52.2 306.45 68.4 307.35 ;
        RECT  51.75 316.65 52.65 317.55 ;
        RECT  51.75 316.2 52.65 317.1 ;
        RECT  52.2 316.65 68.4 317.55 ;
        RECT  51.75 334.65 52.65 335.55 ;
        RECT  51.75 335.1 52.65 336.0 ;
        RECT  52.2 334.65 68.4 335.55 ;
        RECT  51.75 344.85 52.65 345.75 ;
        RECT  51.75 344.4 52.65 345.3 ;
        RECT  52.2 344.85 68.4 345.75 ;
        RECT  51.75 362.85 52.65 363.75 ;
        RECT  51.75 363.3 52.65 364.2 ;
        RECT  52.2 362.85 68.4 363.75 ;
        RECT  51.75 373.05 52.65 373.95 ;
        RECT  51.75 372.6 52.65 373.5 ;
        RECT  52.2 373.05 68.4 373.95 ;
        RECT  51.75 391.05 52.65 391.95 ;
        RECT  51.75 391.5 52.65 392.4 ;
        RECT  52.2 391.05 68.4 391.95 ;
        RECT  51.75 401.25 52.65 402.15 ;
        RECT  51.75 400.8 52.65 401.7 ;
        RECT  52.2 401.25 68.4 402.15 ;
        RECT  51.75 419.25 52.65 420.15 ;
        RECT  51.75 419.7 52.65 420.6 ;
        RECT  52.2 419.25 68.4 420.15 ;
        RECT  49.8 199.2 50.7 424.8 ;
        RECT  67.35 206.55 68.25 207.45 ;
        RECT  69.75 206.55 70.65 207.45 ;
        RECT  67.35 207.0 68.25 210.15 ;
        RECT  67.8 206.55 70.2 207.45 ;
        RECT  69.75 202.35 70.65 207.0 ;
        RECT  67.2 210.15 68.4 211.35 ;
        RECT  69.6 201.15 70.8 202.35 ;
        RECT  69.6 206.4 70.8 207.6 ;
        RECT  49.65 205.05 50.85 206.25 ;
        RECT  51.6 202.8 52.8 204.0 ;
        RECT  67.2 203.7 68.4 204.9 ;
        RECT  67.35 219.15 68.25 220.05 ;
        RECT  69.75 219.15 70.65 220.05 ;
        RECT  67.35 216.45 68.25 219.6 ;
        RECT  67.8 219.15 70.2 220.05 ;
        RECT  69.75 219.6 70.65 224.25 ;
        RECT  67.2 216.45 68.4 217.65 ;
        RECT  69.6 225.45 70.8 226.65 ;
        RECT  69.6 220.2 70.8 221.4 ;
        RECT  49.65 220.35 50.85 221.55 ;
        RECT  51.6 222.6 52.8 223.8 ;
        RECT  67.2 221.7 68.4 222.9 ;
        RECT  67.35 234.75 68.25 235.65 ;
        RECT  69.75 234.75 70.65 235.65 ;
        RECT  67.35 235.2 68.25 238.35 ;
        RECT  67.8 234.75 70.2 235.65 ;
        RECT  69.75 230.55 70.65 235.2 ;
        RECT  67.2 238.35 68.4 239.55 ;
        RECT  69.6 229.35 70.8 230.55 ;
        RECT  69.6 234.6 70.8 235.8 ;
        RECT  49.65 233.25 50.85 234.45 ;
        RECT  51.6 231.0 52.8 232.2 ;
        RECT  67.2 231.9 68.4 233.1 ;
        RECT  67.35 247.35 68.25 248.25 ;
        RECT  69.75 247.35 70.65 248.25 ;
        RECT  67.35 244.65 68.25 247.8 ;
        RECT  67.8 247.35 70.2 248.25 ;
        RECT  69.75 247.8 70.65 252.45 ;
        RECT  67.2 244.65 68.4 245.85 ;
        RECT  69.6 253.65 70.8 254.85 ;
        RECT  69.6 248.4 70.8 249.6 ;
        RECT  49.65 248.55 50.85 249.75 ;
        RECT  51.6 250.8 52.8 252.0 ;
        RECT  67.2 249.9 68.4 251.1 ;
        RECT  67.35 262.95 68.25 263.85 ;
        RECT  69.75 262.95 70.65 263.85 ;
        RECT  67.35 263.4 68.25 266.55 ;
        RECT  67.8 262.95 70.2 263.85 ;
        RECT  69.75 258.75 70.65 263.4 ;
        RECT  67.2 266.55 68.4 267.75 ;
        RECT  69.6 257.55 70.8 258.75 ;
        RECT  69.6 262.8 70.8 264.0 ;
        RECT  49.65 261.45 50.85 262.65 ;
        RECT  51.6 259.2 52.8 260.4 ;
        RECT  67.2 260.1 68.4 261.3 ;
        RECT  67.35 275.55 68.25 276.45 ;
        RECT  69.75 275.55 70.65 276.45 ;
        RECT  67.35 272.85 68.25 276.0 ;
        RECT  67.8 275.55 70.2 276.45 ;
        RECT  69.75 276.0 70.65 280.65 ;
        RECT  67.2 272.85 68.4 274.05 ;
        RECT  69.6 281.85 70.8 283.05 ;
        RECT  69.6 276.6 70.8 277.8 ;
        RECT  49.65 276.75 50.85 277.95 ;
        RECT  51.6 279.0 52.8 280.2 ;
        RECT  67.2 278.1 68.4 279.3 ;
        RECT  67.35 291.15 68.25 292.05 ;
        RECT  69.75 291.15 70.65 292.05 ;
        RECT  67.35 291.6 68.25 294.75 ;
        RECT  67.8 291.15 70.2 292.05 ;
        RECT  69.75 286.95 70.65 291.6 ;
        RECT  67.2 294.75 68.4 295.95 ;
        RECT  69.6 285.75 70.8 286.95 ;
        RECT  69.6 291.0 70.8 292.2 ;
        RECT  49.65 289.65 50.85 290.85 ;
        RECT  51.6 287.4 52.8 288.6 ;
        RECT  67.2 288.3 68.4 289.5 ;
        RECT  67.35 303.75 68.25 304.65 ;
        RECT  69.75 303.75 70.65 304.65 ;
        RECT  67.35 301.05 68.25 304.2 ;
        RECT  67.8 303.75 70.2 304.65 ;
        RECT  69.75 304.2 70.65 308.85 ;
        RECT  67.2 301.05 68.4 302.25 ;
        RECT  69.6 310.05 70.8 311.25 ;
        RECT  69.6 304.8 70.8 306.0 ;
        RECT  49.65 304.95 50.85 306.15 ;
        RECT  51.6 307.2 52.8 308.4 ;
        RECT  67.2 306.3 68.4 307.5 ;
        RECT  67.35 319.35 68.25 320.25 ;
        RECT  69.75 319.35 70.65 320.25 ;
        RECT  67.35 319.8 68.25 322.95 ;
        RECT  67.8 319.35 70.2 320.25 ;
        RECT  69.75 315.15 70.65 319.8 ;
        RECT  67.2 322.95 68.4 324.15 ;
        RECT  69.6 313.95 70.8 315.15 ;
        RECT  69.6 319.2 70.8 320.4 ;
        RECT  49.65 317.85 50.85 319.05 ;
        RECT  51.6 315.6 52.8 316.8 ;
        RECT  67.2 316.5 68.4 317.7 ;
        RECT  67.35 331.95 68.25 332.85 ;
        RECT  69.75 331.95 70.65 332.85 ;
        RECT  67.35 329.25 68.25 332.4 ;
        RECT  67.8 331.95 70.2 332.85 ;
        RECT  69.75 332.4 70.65 337.05 ;
        RECT  67.2 329.25 68.4 330.45 ;
        RECT  69.6 338.25 70.8 339.45 ;
        RECT  69.6 333.0 70.8 334.2 ;
        RECT  49.65 333.15 50.85 334.35 ;
        RECT  51.6 335.4 52.8 336.6 ;
        RECT  67.2 334.5 68.4 335.7 ;
        RECT  67.35 347.55 68.25 348.45 ;
        RECT  69.75 347.55 70.65 348.45 ;
        RECT  67.35 348.0 68.25 351.15 ;
        RECT  67.8 347.55 70.2 348.45 ;
        RECT  69.75 343.35 70.65 348.0 ;
        RECT  67.2 351.15 68.4 352.35 ;
        RECT  69.6 342.15 70.8 343.35 ;
        RECT  69.6 347.4 70.8 348.6 ;
        RECT  49.65 346.05 50.85 347.25 ;
        RECT  51.6 343.8 52.8 345.0 ;
        RECT  67.2 344.7 68.4 345.9 ;
        RECT  67.35 360.15 68.25 361.05 ;
        RECT  69.75 360.15 70.65 361.05 ;
        RECT  67.35 357.45 68.25 360.6 ;
        RECT  67.8 360.15 70.2 361.05 ;
        RECT  69.75 360.6 70.65 365.25 ;
        RECT  67.2 357.45 68.4 358.65 ;
        RECT  69.6 366.45 70.8 367.65 ;
        RECT  69.6 361.2 70.8 362.4 ;
        RECT  49.65 361.35 50.85 362.55 ;
        RECT  51.6 363.6 52.8 364.8 ;
        RECT  67.2 362.7 68.4 363.9 ;
        RECT  67.35 375.75 68.25 376.65 ;
        RECT  69.75 375.75 70.65 376.65 ;
        RECT  67.35 376.2 68.25 379.35 ;
        RECT  67.8 375.75 70.2 376.65 ;
        RECT  69.75 371.55 70.65 376.2 ;
        RECT  67.2 379.35 68.4 380.55 ;
        RECT  69.6 370.35 70.8 371.55 ;
        RECT  69.6 375.6 70.8 376.8 ;
        RECT  49.65 374.25 50.85 375.45 ;
        RECT  51.6 372.0 52.8 373.2 ;
        RECT  67.2 372.9 68.4 374.1 ;
        RECT  67.35 388.35 68.25 389.25 ;
        RECT  69.75 388.35 70.65 389.25 ;
        RECT  67.35 385.65 68.25 388.8 ;
        RECT  67.8 388.35 70.2 389.25 ;
        RECT  69.75 388.8 70.65 393.45 ;
        RECT  67.2 385.65 68.4 386.85 ;
        RECT  69.6 394.65 70.8 395.85 ;
        RECT  69.6 389.4 70.8 390.6 ;
        RECT  49.65 389.55 50.85 390.75 ;
        RECT  51.6 391.8 52.8 393.0 ;
        RECT  67.2 390.9 68.4 392.1 ;
        RECT  67.35 403.95 68.25 404.85 ;
        RECT  69.75 403.95 70.65 404.85 ;
        RECT  67.35 404.4 68.25 407.55 ;
        RECT  67.8 403.95 70.2 404.85 ;
        RECT  69.75 399.75 70.65 404.4 ;
        RECT  67.2 407.55 68.4 408.75 ;
        RECT  69.6 398.55 70.8 399.75 ;
        RECT  69.6 403.8 70.8 405.0 ;
        RECT  49.65 402.45 50.85 403.65 ;
        RECT  51.6 400.2 52.8 401.4 ;
        RECT  67.2 401.1 68.4 402.3 ;
        RECT  67.35 416.55 68.25 417.45 ;
        RECT  69.75 416.55 70.65 417.45 ;
        RECT  67.35 413.85 68.25 417.0 ;
        RECT  67.8 416.55 70.2 417.45 ;
        RECT  69.75 417.0 70.65 421.65 ;
        RECT  67.2 413.85 68.4 415.05 ;
        RECT  69.6 422.85 70.8 424.05 ;
        RECT  69.6 417.6 70.8 418.8 ;
        RECT  49.65 417.75 50.85 418.95 ;
        RECT  51.6 420.0 52.8 421.2 ;
        RECT  67.2 419.1 68.4 420.3 ;
        RECT  61.8 62.4 66.3 63.6 ;
        RECT  6.3 44.7 7.5 45.9 ;
        RECT  61.8 57.6 66.3 58.8 ;
        RECT  61.8 42.0 66.3 43.2 ;
        RECT  6.3 65.1 7.5 66.3 ;
        RECT  6.3 75.3 7.5 76.5 ;
        RECT  6.3 54.9 7.5 56.1 ;
        RECT  6.3 70.2 66.3 71.4 ;
        RECT  6.3 49.8 66.3 51.0 ;
        RECT  61.8 78.0 66.3 79.2 ;
        RECT  65.1 75.3 66.3 76.5 ;
        RECT  65.1 65.1 66.3 66.3 ;
        RECT  65.1 44.7 66.3 45.9 ;
        RECT  65.1 54.9 66.3 56.1 ;
        RECT  61.8 78.0 66.3 79.2 ;
        RECT  65.1 75.3 66.3 76.5 ;
        RECT  63.9 73.8 65.1 76.5 ;
        RECT  60.6 76.2 61.8 79.2 ;
        RECT  51.0 78.3 60.6 79.2 ;
        RECT  56.1 73.8 63.9 75.0 ;
        RECT  52.8 72.9 54.0 75.9 ;
        RECT  49.8 78.0 51.0 79.2 ;
        RECT  50.7 74.7 51.9 75.9 ;
        RECT  49.2 74.7 50.7 75.6 ;
        RECT  48.3 74.7 49.2 77.1 ;
        RECT  42.0 76.2 48.3 77.1 ;
        RECT  47.4 72.9 52.8 73.8 ;
        RECT  46.2 72.9 47.4 75.0 ;
        RECT  43.8 72.9 45.0 75.0 ;
        RECT  40.8 76.2 42.0 77.4 ;
        RECT  36.3 78.0 37.5 79.5 ;
        RECT  24.6 78.6 36.3 79.5 ;
        RECT  34.2 75.3 38.7 76.5 ;
        RECT  33.3 75.3 34.2 77.7 ;
        RECT  26.4 76.8 33.3 77.7 ;
        RECT  31.8 72.9 43.8 73.8 ;
        RECT  30.6 72.9 31.8 75.0 ;
        RECT  27.3 72.9 28.5 75.9 ;
        RECT  25.5 76.2 26.4 77.7 ;
        RECT  23.4 78.0 24.6 79.5 ;
        RECT  24.3 74.7 25.5 77.1 ;
        RECT  15.6 76.2 24.3 77.1 ;
        RECT  21.0 72.9 27.3 73.8 ;
        RECT  19.8 72.9 21.0 75.0 ;
        RECT  17.4 72.9 18.6 75.0 ;
        RECT  14.4 76.2 15.6 77.4 ;
        RECT  8.7 72.9 17.4 73.8 ;
        RECT  7.5 72.9 8.7 76.5 ;
        RECT  6.3 75.3 7.5 76.5 ;
        RECT  6.3 70.2 66.3 71.4 ;
        RECT  6.3 75.3 7.5 76.5 ;
        RECT  65.1 75.3 66.3 76.5 ;
        RECT  61.8 78.0 66.3 79.2 ;
        RECT  6.3 70.2 66.3 71.4 ;
        RECT  61.8 62.4 66.3 63.6 ;
        RECT  65.1 65.1 66.3 66.3 ;
        RECT  63.9 65.1 65.1 67.8 ;
        RECT  60.6 62.4 61.8 65.4 ;
        RECT  51.0 62.4 60.6 63.3 ;
        RECT  56.1 66.6 63.9 67.8 ;
        RECT  52.8 65.7 54.0 68.7 ;
        RECT  49.8 62.4 51.0 63.6 ;
        RECT  50.7 65.7 51.9 66.9 ;
        RECT  49.2 66.0 50.7 66.9 ;
        RECT  48.3 64.5 49.2 66.9 ;
        RECT  42.0 64.5 48.3 65.4 ;
        RECT  47.4 67.8 52.8 68.7 ;
        RECT  46.2 66.6 47.4 68.7 ;
        RECT  43.8 66.6 45.0 68.7 ;
        RECT  40.8 64.2 42.0 65.4 ;
        RECT  36.3 62.1 37.5 63.6 ;
        RECT  24.6 62.1 36.3 63.0 ;
        RECT  34.2 65.1 38.7 66.3 ;
        RECT  33.3 63.9 34.2 66.3 ;
        RECT  26.4 63.9 33.3 64.8 ;
        RECT  31.8 67.8 43.8 68.7 ;
        RECT  30.6 66.6 31.8 68.7 ;
        RECT  27.3 65.7 28.5 68.7 ;
        RECT  25.5 63.9 26.4 65.4 ;
        RECT  23.4 62.1 24.6 63.6 ;
        RECT  24.3 64.5 25.5 66.9 ;
        RECT  15.6 64.5 24.3 65.4 ;
        RECT  21.0 67.8 27.3 68.7 ;
        RECT  19.8 66.6 21.0 68.7 ;
        RECT  17.4 66.6 18.6 68.7 ;
        RECT  14.4 64.2 15.6 65.4 ;
        RECT  8.7 67.8 17.4 68.7 ;
        RECT  7.5 65.1 8.7 68.7 ;
        RECT  6.3 65.1 7.5 66.3 ;
        RECT  6.3 70.2 66.3 71.4 ;
        RECT  6.3 65.1 7.5 66.3 ;
        RECT  65.1 65.1 66.3 66.3 ;
        RECT  61.8 62.4 66.3 63.6 ;
        RECT  6.3 70.2 66.3 71.4 ;
        RECT  61.8 57.6 66.3 58.8 ;
        RECT  65.1 54.9 66.3 56.1 ;
        RECT  63.9 53.4 65.1 56.1 ;
        RECT  60.6 55.8 61.8 58.8 ;
        RECT  51.0 57.9 60.6 58.8 ;
        RECT  56.1 53.4 63.9 54.6 ;
        RECT  52.8 52.5 54.0 55.5 ;
        RECT  49.8 57.6 51.0 58.8 ;
        RECT  50.7 54.3 51.9 55.5 ;
        RECT  49.2 54.3 50.7 55.2 ;
        RECT  48.3 54.3 49.2 56.7 ;
        RECT  42.0 55.8 48.3 56.7 ;
        RECT  47.4 52.5 52.8 53.4 ;
        RECT  46.2 52.5 47.4 54.6 ;
        RECT  43.8 52.5 45.0 54.6 ;
        RECT  40.8 55.8 42.0 57.0 ;
        RECT  36.3 57.6 37.5 59.1 ;
        RECT  24.6 58.2 36.3 59.1 ;
        RECT  34.2 54.9 38.7 56.1 ;
        RECT  33.3 54.9 34.2 57.3 ;
        RECT  26.4 56.4 33.3 57.3 ;
        RECT  31.8 52.5 43.8 53.4 ;
        RECT  30.6 52.5 31.8 54.6 ;
        RECT  27.3 52.5 28.5 55.5 ;
        RECT  25.5 55.8 26.4 57.3 ;
        RECT  23.4 57.6 24.6 59.1 ;
        RECT  24.3 54.3 25.5 56.7 ;
        RECT  15.6 55.8 24.3 56.7 ;
        RECT  21.0 52.5 27.3 53.4 ;
        RECT  19.8 52.5 21.0 54.6 ;
        RECT  17.4 52.5 18.6 54.6 ;
        RECT  14.4 55.8 15.6 57.0 ;
        RECT  8.7 52.5 17.4 53.4 ;
        RECT  7.5 52.5 8.7 56.1 ;
        RECT  6.3 54.9 7.5 56.1 ;
        RECT  6.3 49.8 66.3 51.0 ;
        RECT  6.3 54.9 7.5 56.1 ;
        RECT  65.1 54.9 66.3 56.1 ;
        RECT  61.8 57.6 66.3 58.8 ;
        RECT  6.3 49.8 66.3 51.0 ;
        RECT  61.8 42.0 66.3 43.2 ;
        RECT  65.1 44.7 66.3 45.9 ;
        RECT  63.9 44.7 65.1 47.4 ;
        RECT  60.6 42.0 61.8 45.0 ;
        RECT  51.0 42.0 60.6 42.9 ;
        RECT  56.1 46.2 63.9 47.4 ;
        RECT  52.8 45.3 54.0 48.3 ;
        RECT  49.8 42.0 51.0 43.2 ;
        RECT  50.7 45.3 51.9 46.5 ;
        RECT  49.2 45.6 50.7 46.5 ;
        RECT  48.3 44.1 49.2 46.5 ;
        RECT  42.0 44.1 48.3 45.0 ;
        RECT  47.4 47.4 52.8 48.3 ;
        RECT  46.2 46.2 47.4 48.3 ;
        RECT  43.8 46.2 45.0 48.3 ;
        RECT  40.8 43.8 42.0 45.0 ;
        RECT  36.3 41.7 37.5 43.2 ;
        RECT  24.6 41.7 36.3 42.6 ;
        RECT  34.2 44.7 38.7 45.9 ;
        RECT  33.3 43.5 34.2 45.9 ;
        RECT  26.4 43.5 33.3 44.4 ;
        RECT  31.8 47.4 43.8 48.3 ;
        RECT  30.6 46.2 31.8 48.3 ;
        RECT  27.3 45.3 28.5 48.3 ;
        RECT  25.5 43.5 26.4 45.0 ;
        RECT  23.4 41.7 24.6 43.2 ;
        RECT  24.3 44.1 25.5 46.5 ;
        RECT  15.6 44.1 24.3 45.0 ;
        RECT  21.0 47.4 27.3 48.3 ;
        RECT  19.8 46.2 21.0 48.3 ;
        RECT  17.4 46.2 18.6 48.3 ;
        RECT  14.4 43.8 15.6 45.0 ;
        RECT  8.7 47.4 17.4 48.3 ;
        RECT  7.5 44.7 8.7 48.3 ;
        RECT  6.3 44.7 7.5 45.9 ;
        RECT  6.3 49.8 66.3 51.0 ;
        RECT  6.3 44.7 7.5 45.9 ;
        RECT  65.1 44.7 66.3 45.9 ;
        RECT  61.8 42.0 66.3 43.2 ;
        RECT  6.3 49.8 66.3 51.0 ;
        RECT  123.75 5.85 124.95 7.05 ;
        RECT  133.95 5.85 135.15 7.05 ;
        RECT  127.5 0.3 128.7 1.5 ;
        RECT  137.7 0.3 138.9 1.5 ;
        RECT  95.25 198.6 96.45 199.8 ;
        RECT  95.25 226.8 96.45 228.0 ;
        RECT  95.25 255.0 96.45 256.2 ;
        RECT  95.25 283.2 96.45 284.4 ;
        RECT  95.25 311.4 96.45 312.6 ;
        RECT  95.25 339.6 96.45 340.8 ;
        RECT  95.25 367.8 96.45 369.0 ;
        RECT  95.25 396.0 96.45 397.2 ;
        RECT  95.25 424.2 96.45 425.4 ;
        RECT  76.5 88.65 77.7 89.85 ;
        RECT  81.6 88.5 82.8 89.7 ;
        RECT  73.5 102.75 74.7 103.95 ;
        RECT  84.3 102.6 85.5 103.8 ;
        RECT  76.5 145.05 77.7 146.25 ;
        RECT  87.0 144.9 88.2 146.1 ;
        RECT  73.5 159.15 74.7 160.35 ;
        RECT  89.7 159.0 90.9 160.2 ;
        RECT  78.6 85.8 79.8 87.0 ;
        RECT  78.6 85.8 79.8 87.0 ;
        RECT  94.65 85.8 95.85 87.0 ;
        RECT  78.6 114.0 79.8 115.2 ;
        RECT  78.6 114.0 79.8 115.2 ;
        RECT  94.65 114.0 95.85 115.2 ;
        RECT  78.6 142.2 79.8 143.4 ;
        RECT  78.6 142.2 79.8 143.4 ;
        RECT  94.65 142.2 95.85 143.4 ;
        RECT  78.6 170.4 79.8 171.6 ;
        RECT  78.6 170.4 79.8 171.6 ;
        RECT  94.65 170.4 95.85 171.6 ;
        RECT  65.7 75.3 66.9 76.5 ;
        RECT  81.6 75.3 82.8 76.5 ;
        RECT  65.7 65.1 66.9 66.3 ;
        RECT  84.3 65.1 85.5 66.3 ;
        RECT  65.7 54.9 66.9 56.1 ;
        RECT  87.0 54.9 88.2 56.1 ;
        RECT  65.7 44.7 66.9 45.9 ;
        RECT  89.7 44.7 90.9 45.9 ;
        RECT  66.3 70.2 67.5 71.4 ;
        RECT  95.25 70.35 96.45 71.55 ;
        RECT  66.3 49.8 67.5 51.0 ;
        RECT  95.25 49.95 96.45 51.15 ;
        RECT  110.4 32.25 111.6 33.45 ;
        RECT  105.0 27.75 106.2 28.95 ;
        RECT  107.7 25.35 108.9 26.55 ;
        RECT  110.4 429.45 111.6 430.65 ;
        RECT  113.1 96.75 114.3 97.95 ;
        RECT  115.8 194.85 117.0 196.05 ;
        RECT  102.3 82.5 103.5 83.7 ;
        RECT  49.65 426.3 50.85 427.5 ;
        RECT  102.3 426.3 103.5 427.5 ;
        RECT  98.55 23.4 99.75 24.6 ;
        RECT  98.55 192.9 99.75 194.1 ;
        RECT  98.55 94.8 99.75 96.0 ;
        RECT  -53.1 289.8 -3.0 290.7 ;
        RECT  -53.1 292.5 -3.0 293.4 ;
        RECT  -53.1 295.2 -3.0 296.1 ;
        RECT  -53.1 300.6 -3.0 301.5 ;
        RECT  -20.25 205.05 -19.35 284.85 ;
        RECT  -5.7 287.1 -3.0 288.0 ;
        RECT  -17.1 297.9 -14.4 298.8 ;
        RECT  -31.2 287.1 -28.5 288.0 ;
        RECT  -45.3 297.9 -42.6 298.8 ;
        RECT  -53.1 303.3 -3.0 304.2 ;
        RECT  -37.65 362.25 -3.0 363.15 ;
        RECT  -53.1 284.4 -3.0 285.3 ;
        RECT  -23.4 339.75 -3.0 340.65 ;
        RECT  -53.1 297.9 -3.0 298.8 ;
        RECT  -53.1 287.1 -3.0 288.0 ;
        RECT  -24.75 342.45 -3.0 343.35 ;
        RECT  -24.15 322.65 -3.0 323.55 ;
        RECT  -35.7 257.7 -34.5 262.2 ;
        RECT  -30.9 257.7 -29.7 262.2 ;
        RECT  -38.4 202.2 -37.2 203.4 ;
        RECT  -48.6 202.2 -47.4 203.4 ;
        RECT  -28.2 202.2 -27.0 203.4 ;
        RECT  -43.5 202.2 -42.3 262.2 ;
        RECT  -23.1 202.2 -21.9 262.2 ;
        RECT  -51.3 257.7 -50.1 262.2 ;
        RECT  -48.6 261.0 -47.4 262.2 ;
        RECT  -38.4 261.0 -37.2 262.2 ;
        RECT  -28.2 261.0 -27.0 262.2 ;
        RECT  -51.3 257.7 -50.1 262.2 ;
        RECT  -48.6 261.0 -47.4 262.2 ;
        RECT  -48.6 259.8 -45.9 261.0 ;
        RECT  -51.3 256.5 -48.3 257.7 ;
        RECT  -51.3 246.9 -50.4 256.5 ;
        RECT  -47.1 252.0 -45.9 259.8 ;
        RECT  -48.0 248.7 -45.0 249.9 ;
        RECT  -51.3 245.7 -50.1 246.9 ;
        RECT  -48.0 246.6 -46.8 247.8 ;
        RECT  -47.7 245.1 -46.8 246.6 ;
        RECT  -49.2 244.2 -46.8 245.1 ;
        RECT  -49.2 237.9 -48.3 244.2 ;
        RECT  -45.9 243.3 -45.0 248.7 ;
        RECT  -47.1 242.1 -45.0 243.3 ;
        RECT  -47.1 239.7 -45.0 240.9 ;
        RECT  -49.5 236.7 -48.3 237.9 ;
        RECT  -51.6 232.2 -50.1 233.4 ;
        RECT  -51.6 220.5 -50.7 232.2 ;
        RECT  -48.6 230.1 -47.4 234.6 ;
        RECT  -49.8 229.2 -47.4 230.1 ;
        RECT  -49.8 222.3 -48.9 229.2 ;
        RECT  -45.9 227.7 -45.0 239.7 ;
        RECT  -47.1 226.5 -45.0 227.7 ;
        RECT  -48.0 223.2 -45.0 224.4 ;
        RECT  -49.8 221.4 -48.3 222.3 ;
        RECT  -51.6 219.3 -50.1 220.5 ;
        RECT  -49.2 220.2 -46.8 221.4 ;
        RECT  -49.2 211.5 -48.3 220.2 ;
        RECT  -45.9 216.9 -45.0 223.2 ;
        RECT  -47.1 215.7 -45.0 216.9 ;
        RECT  -47.1 213.3 -45.0 214.5 ;
        RECT  -49.5 210.3 -48.3 211.5 ;
        RECT  -45.9 204.6 -45.0 213.3 ;
        RECT  -48.6 203.4 -45.0 204.6 ;
        RECT  -48.6 202.2 -47.4 203.4 ;
        RECT  -43.5 202.2 -42.3 262.2 ;
        RECT  -48.6 202.2 -47.4 203.4 ;
        RECT  -48.6 261.0 -47.4 262.2 ;
        RECT  -51.3 257.7 -50.1 262.2 ;
        RECT  -43.5 202.2 -42.3 262.2 ;
        RECT  -35.7 257.7 -34.5 262.2 ;
        RECT  -38.4 261.0 -37.2 262.2 ;
        RECT  -39.9 259.8 -37.2 261.0 ;
        RECT  -37.5 256.5 -34.5 257.7 ;
        RECT  -35.4 246.9 -34.5 256.5 ;
        RECT  -39.9 252.0 -38.7 259.8 ;
        RECT  -40.8 248.7 -37.8 249.9 ;
        RECT  -35.7 245.7 -34.5 246.9 ;
        RECT  -39.0 246.6 -37.8 247.8 ;
        RECT  -39.0 245.1 -38.1 246.6 ;
        RECT  -39.0 244.2 -36.6 245.1 ;
        RECT  -37.5 237.9 -36.6 244.2 ;
        RECT  -40.8 243.3 -39.9 248.7 ;
        RECT  -40.8 242.1 -38.7 243.3 ;
        RECT  -40.8 239.7 -38.7 240.9 ;
        RECT  -37.5 236.7 -36.3 237.9 ;
        RECT  -35.7 232.2 -34.2 233.4 ;
        RECT  -35.1 220.5 -34.2 232.2 ;
        RECT  -38.4 230.1 -37.2 234.6 ;
        RECT  -38.4 229.2 -36.0 230.1 ;
        RECT  -36.9 222.3 -36.0 229.2 ;
        RECT  -40.8 227.7 -39.9 239.7 ;
        RECT  -40.8 226.5 -38.7 227.7 ;
        RECT  -40.8 223.2 -37.8 224.4 ;
        RECT  -37.5 221.4 -36.0 222.3 ;
        RECT  -35.7 219.3 -34.2 220.5 ;
        RECT  -39.0 220.2 -36.6 221.4 ;
        RECT  -37.5 211.5 -36.6 220.2 ;
        RECT  -40.8 216.9 -39.9 223.2 ;
        RECT  -40.8 215.7 -38.7 216.9 ;
        RECT  -40.8 213.3 -38.7 214.5 ;
        RECT  -37.5 210.3 -36.3 211.5 ;
        RECT  -40.8 204.6 -39.9 213.3 ;
        RECT  -40.8 203.4 -37.2 204.6 ;
        RECT  -38.4 202.2 -37.2 203.4 ;
        RECT  -43.5 202.2 -42.3 262.2 ;
        RECT  -38.4 202.2 -37.2 203.4 ;
        RECT  -38.4 261.0 -37.2 262.2 ;
        RECT  -35.7 257.7 -34.5 262.2 ;
        RECT  -43.5 202.2 -42.3 262.2 ;
        RECT  -30.9 257.7 -29.7 262.2 ;
        RECT  -28.2 261.0 -27.0 262.2 ;
        RECT  -28.2 259.8 -25.5 261.0 ;
        RECT  -30.9 256.5 -27.9 257.7 ;
        RECT  -30.9 246.9 -30.0 256.5 ;
        RECT  -26.7 252.0 -25.5 259.8 ;
        RECT  -27.6 248.7 -24.6 249.9 ;
        RECT  -30.9 245.7 -29.7 246.9 ;
        RECT  -27.6 246.6 -26.4 247.8 ;
        RECT  -27.3 245.1 -26.4 246.6 ;
        RECT  -28.8 244.2 -26.4 245.1 ;
        RECT  -28.8 237.9 -27.9 244.2 ;
        RECT  -25.5 243.3 -24.6 248.7 ;
        RECT  -26.7 242.1 -24.6 243.3 ;
        RECT  -26.7 239.7 -24.6 240.9 ;
        RECT  -29.1 236.7 -27.9 237.9 ;
        RECT  -31.2 232.2 -29.7 233.4 ;
        RECT  -31.2 220.5 -30.3 232.2 ;
        RECT  -28.2 230.1 -27.0 234.6 ;
        RECT  -29.4 229.2 -27.0 230.1 ;
        RECT  -29.4 222.3 -28.5 229.2 ;
        RECT  -25.5 227.7 -24.6 239.7 ;
        RECT  -26.7 226.5 -24.6 227.7 ;
        RECT  -27.6 223.2 -24.6 224.4 ;
        RECT  -29.4 221.4 -27.9 222.3 ;
        RECT  -31.2 219.3 -29.7 220.5 ;
        RECT  -28.8 220.2 -26.4 221.4 ;
        RECT  -28.8 211.5 -27.9 220.2 ;
        RECT  -25.5 216.9 -24.6 223.2 ;
        RECT  -26.7 215.7 -24.6 216.9 ;
        RECT  -26.7 213.3 -24.6 214.5 ;
        RECT  -29.1 210.3 -27.9 211.5 ;
        RECT  -25.5 204.6 -24.6 213.3 ;
        RECT  -28.2 203.4 -24.6 204.6 ;
        RECT  -28.2 202.2 -27.0 203.4 ;
        RECT  -23.1 202.2 -21.9 262.2 ;
        RECT  -28.2 202.2 -27.0 203.4 ;
        RECT  -28.2 261.0 -27.0 262.2 ;
        RECT  -30.9 257.7 -29.7 262.2 ;
        RECT  -23.1 202.2 -21.9 262.2 ;
        RECT  -14.4 317.85 -6.3 318.75 ;
        RECT  -12.75 313.05 -11.85 313.95 ;
        RECT  -12.75 317.85 -11.85 318.75 ;
        RECT  -14.4 313.05 -12.3 313.95 ;
        RECT  -12.75 313.5 -11.85 318.3 ;
        RECT  -12.3 317.85 -6.3 318.75 ;
        RECT  -15.6 312.9 -14.4 314.1 ;
        RECT  -15.6 317.7 -14.4 318.9 ;
        RECT  -6.3 317.7 -5.1 318.9 ;
        RECT  -12.9 317.7 -11.7 318.9 ;
        RECT  -24.6 315.45 -23.7 316.35 ;
        RECT  -24.15 315.45 -20.85 316.35 ;
        RECT  -24.6 315.9 -23.7 316.8 ;
        RECT  -29.7 315.45 -28.8 316.35 ;
        RECT  -29.7 314.1 -28.8 315.9 ;
        RECT  -29.25 315.45 -24.15 316.35 ;
        RECT  -22.05 315.3 -20.85 316.5 ;
        RECT  -31.05 312.9 -29.85 314.1 ;
        RECT  -25.95 316.2 -24.75 317.4 ;
        RECT  -23.85 330.15 -22.95 331.05 ;
        RECT  -23.85 332.55 -22.95 333.45 ;
        RECT  -23.4 330.15 -20.25 331.05 ;
        RECT  -23.85 330.6 -22.95 333.0 ;
        RECT  -28.05 332.55 -23.4 333.45 ;
        RECT  -21.45 330.0 -20.25 331.2 ;
        RECT  -30.45 332.4 -29.25 333.6 ;
        RECT  -25.2 332.4 -24.0 333.6 ;
        RECT  -42.6 327.45 -34.5 328.35 ;
        RECT  -40.95 322.65 -40.05 323.55 ;
        RECT  -40.95 327.45 -40.05 328.35 ;
        RECT  -42.6 322.65 -40.5 323.55 ;
        RECT  -40.95 323.1 -40.05 327.9 ;
        RECT  -40.5 327.45 -34.5 328.35 ;
        RECT  -43.8 322.5 -42.6 323.7 ;
        RECT  -43.8 327.3 -42.6 328.5 ;
        RECT  -34.5 327.3 -33.3 328.5 ;
        RECT  -41.1 327.3 -39.9 328.5 ;
        RECT  -51.3 261.6 -50.1 262.8 ;
        RECT  -51.3 300.45 -50.1 301.65 ;
        RECT  -48.6 261.6 -47.4 262.8 ;
        RECT  -48.6 289.65 -47.4 290.85 ;
        RECT  -35.7 261.6 -34.5 262.8 ;
        RECT  -35.7 292.35 -34.5 293.55 ;
        RECT  -30.9 261.6 -29.7 262.8 ;
        RECT  -30.9 295.05 -29.7 296.25 ;
        RECT  -43.5 261.6 -42.3 262.8 ;
        RECT  -43.5 286.95 -42.3 288.15 ;
        RECT  -23.1 261.6 -21.9 262.8 ;
        RECT  -23.1 286.95 -21.9 288.15 ;
        RECT  -31.65 371.7 -30.75 426.9 ;
        RECT  -31.65 381.3 -30.75 384.0 ;
        RECT  -31.65 384.0 -30.75 426.9 ;
        RECT  -47.25 424.2 -46.35 426.9 ;
        RECT  -33.9 376.5 -33.0 384.0 ;
        RECT  -40.65 376.5 -39.75 381.3 ;
        RECT  -9.9 397.5 -9.0 404.7 ;
        RECT  -17.55 394.65 -16.65 395.55 ;
        RECT  -17.55 393.45 -16.65 394.35 ;
        RECT  -17.1 394.65 -9.45 395.55 ;
        RECT  -17.55 393.9 -16.65 395.1 ;
        RECT  -24.75 393.45 -17.1 394.35 ;
        RECT  -25.2 396.3 -24.3 403.5 ;
        RECT  -10.05 396.9 -8.85 398.1 ;
        RECT  -25.35 393.3 -24.15 394.5 ;
        RECT  -25.35 402.9 -24.15 404.1 ;
        RECT  -10.05 404.1 -8.85 405.3 ;
        RECT  -10.05 394.5 -8.85 395.7 ;
        RECT  -25.35 395.7 -24.15 396.9 ;
        RECT  -38.4 400.2 -36.6 410.7 ;
        RECT  -40.8 397.2 -39.6 410.7 ;
        RECT  -43.8 397.2 -42.6 410.7 ;
        RECT  -40.8 396.0 -38.1 397.2 ;
        RECT  -43.8 396.0 -42.3 397.2 ;
        RECT  -47.4 396.0 -46.2 410.7 ;
        RECT  -40.8 397.2 -39.6 410.7 ;
        RECT  -38.4 400.2 -36.6 410.7 ;
        RECT  -47.4 396.0 -46.2 410.7 ;
        RECT  -43.8 397.2 -42.6 410.7 ;
        RECT  -40.8 367.8 -39.6 396.0 ;
        RECT  -47.4 367.8 -46.2 396.0 ;
        RECT  -43.8 367.8 -42.6 396.0 ;
        RECT  -47.4 381.3 -46.2 396.0 ;
        RECT  -43.8 394.8 -42.3 396.0 ;
        RECT  -40.8 394.8 -38.1 396.0 ;
        RECT  -43.8 381.3 -42.6 396.0 ;
        RECT  -40.8 382.5 -39.6 396.0 ;
        RECT  -38.4 381.3 -36.0 391.8 ;
        RECT  -40.8 382.5 -39.6 396.0 ;
        RECT  -47.4 381.3 -46.2 396.0 ;
        RECT  -38.4 381.3 -36.0 391.8 ;
        RECT  -43.8 381.3 -42.6 396.0 ;
        RECT  -47.4 367.8 -46.2 382.5 ;
        RECT  -43.8 367.8 -42.3 369.0 ;
        RECT  -40.8 367.8 -38.1 369.0 ;
        RECT  -43.8 367.8 -42.6 382.5 ;
        RECT  -40.8 367.8 -39.6 381.3 ;
        RECT  -38.4 372.0 -36.0 382.5 ;
        RECT  -40.8 367.8 -39.6 381.3 ;
        RECT  -47.4 367.8 -46.2 382.5 ;
        RECT  -38.4 372.0 -36.0 382.5 ;
        RECT  -43.8 367.8 -42.6 382.5 ;
        RECT  -31.95 396.9 -30.75 398.1 ;
        RECT  -31.95 419.7 -30.75 420.9 ;
        RECT  -31.95 408.9 -30.75 410.1 ;
        RECT  -31.95 369.3 -30.75 370.5 ;
        RECT  -31.8 425.1 -30.6 426.3 ;
        RECT  -47.4 425.1 -46.2 426.3 ;
        RECT  -34.05 382.2 -32.85 383.4 ;
        RECT  -34.05 374.7 -32.85 375.9 ;
        RECT  -40.8 374.7 -39.6 375.9 ;
        RECT  -9.75 284.25 -8.55 285.45 ;
        RECT  -9.75 243.45 -8.55 244.65 ;
        RECT  -9.75 303.15 -8.55 304.35 ;
        RECT  -9.75 243.45 -8.55 244.65 ;
        RECT  -20.4 204.45 -19.2 205.65 ;
        RECT  -24.75 284.25 -23.55 285.45 ;
        RECT  -27.45 289.65 -26.25 290.85 ;
        RECT  -24.0 327.0 -22.8 328.2 ;
        RECT  -24.0 327.0 -22.8 328.2 ;
        RECT  -24.0 303.15 -22.8 304.35 ;
        RECT  -26.7 330.0 -25.5 331.2 ;
        RECT  -26.7 330.0 -25.5 331.2 ;
        RECT  -26.7 300.45 -25.5 301.65 ;
        RECT  -12.9 303.15 -11.7 304.35 ;
        RECT  -10.95 300.45 -9.75 301.65 ;
        RECT  -9.0 292.35 -7.8 293.55 ;
        RECT  -41.1 303.15 -39.9 304.35 ;
        RECT  -39.15 292.35 -37.95 293.55 ;
        RECT  -37.2 295.05 -36.0 296.25 ;
        RECT  -24.75 322.5 -23.55 323.7 ;
        RECT  -24.0 339.6 -22.8 340.8 ;
        RECT  -38.25 362.1 -37.05 363.3 ;
        RECT  -25.35 342.3 -24.15 343.5 ;
        RECT  -3.6 286.95 -2.4 288.15 ;
        RECT  -17.7 297.75 -16.5 298.95 ;
        RECT  -31.8 286.95 -30.6 288.15 ;
        RECT  -45.9 297.75 -44.7 298.95 ;
        RECT  115.8 342.3 117.0 343.5 ;
        RECT  -4.5 342.45 -3.3 343.65 ;
        RECT  113.1 362.1 114.3 363.3 ;
        RECT  -4.5 362.25 -3.3 363.45 ;
        RECT  107.7 322.5 108.9 323.7 ;
        RECT  -4.5 322.65 -3.3 323.85 ;
        RECT  105.0 339.6 106.2 340.8 ;
        RECT  -4.5 339.75 -3.3 340.95 ;
        RECT  110.4 303.15 111.6 304.35 ;
        RECT  -4.5 303.3 -3.3 304.5 ;
        RECT  102.3 284.25 103.5 285.45 ;
        RECT  -4.5 284.4 -3.3 285.6 ;
        RECT  1.65 297.75 2.85 298.95 ;
        RECT  96.9 286.95 98.1 288.15 ;
        RECT  -4.5 287.1 -3.3 288.3 ;
        LAYER  via2 ;
        RECT  123.9 151.8 124.5 152.4 ;
        RECT  134.1 151.8 134.7 152.4 ;
        RECT  127.5 31.5 128.1 32.1 ;
        RECT  137.7 31.5 138.3 32.1 ;
        RECT  127.5 31.8 128.1 32.4 ;
        RECT  137.7 31.8 138.3 32.4 ;
        RECT  7.8 75.6 8.4 76.2 ;
        RECT  7.8 65.4 8.4 66.0 ;
        RECT  7.8 55.2 8.4 55.8 ;
        RECT  7.8 45.0 8.4 45.6 ;
        RECT  124.05 6.15 124.65 6.75 ;
        RECT  134.25 6.15 134.85 6.75 ;
        RECT  127.8 0.6 128.4 1.2 ;
        RECT  138.0 0.6 138.6 1.2 ;
        RECT  78.9 86.1 79.5 86.7 ;
        RECT  94.95 86.1 95.55 86.7 ;
        RECT  78.9 114.3 79.5 114.9 ;
        RECT  94.95 114.3 95.55 114.9 ;
        RECT  78.9 142.5 79.5 143.1 ;
        RECT  94.95 142.5 95.55 143.1 ;
        RECT  78.9 170.7 79.5 171.3 ;
        RECT  94.95 170.7 95.55 171.3 ;
        RECT  -48.3 203.7 -47.7 204.3 ;
        RECT  -38.1 203.7 -37.5 204.3 ;
        RECT  -27.9 203.7 -27.3 204.3 ;
        RECT  -51.0 261.9 -50.4 262.5 ;
        RECT  -51.0 300.75 -50.4 301.35 ;
        RECT  -48.3 261.9 -47.7 262.5 ;
        RECT  -48.3 289.95 -47.7 290.55 ;
        RECT  -35.4 261.9 -34.8 262.5 ;
        RECT  -35.4 292.65 -34.8 293.25 ;
        RECT  -30.6 261.9 -30.0 262.5 ;
        RECT  -30.6 295.35 -30.0 295.95 ;
        RECT  -43.2 261.9 -42.6 262.5 ;
        RECT  -43.2 287.25 -42.6 287.85 ;
        RECT  -22.8 261.9 -22.2 262.5 ;
        RECT  -22.8 287.25 -22.2 287.85 ;
        RECT  -9.45 243.75 -8.85 244.35 ;
        RECT  -9.45 303.45 -8.85 304.05 ;
        RECT  -23.7 327.3 -23.1 327.9 ;
        RECT  -23.7 303.45 -23.1 304.05 ;
        RECT  -26.4 330.3 -25.8 330.9 ;
        RECT  -26.4 300.75 -25.8 301.35 ;
        RECT  116.1 342.6 116.7 343.2 ;
        RECT  -4.2 342.75 -3.6 343.35 ;
        RECT  113.4 362.4 114.0 363.0 ;
        RECT  -4.2 362.55 -3.6 363.15 ;
        RECT  108.0 322.8 108.6 323.4 ;
        RECT  -4.2 322.95 -3.6 323.55 ;
        RECT  105.3 339.9 105.9 340.5 ;
        RECT  -4.2 340.05 -3.6 340.65 ;
        RECT  110.7 303.45 111.3 304.05 ;
        RECT  -4.2 303.6 -3.6 304.2 ;
        RECT  102.6 284.55 103.2 285.15 ;
        RECT  -4.2 284.7 -3.6 285.3 ;
        RECT  97.2 287.25 97.8 287.85 ;
        RECT  -4.2 287.4 -3.6 288.0 ;
        LAYER  metal3 ;
        RECT  -3.0 342.15 116.4 343.65 ;
        RECT  -3.0 361.95 113.7 363.45 ;
        RECT  -3.0 322.35 108.3 323.85 ;
        RECT  -3.0 339.45 105.6 340.95 ;
        RECT  -3.0 303.0 111.0 304.5 ;
        RECT  -3.0 284.1 102.9 285.6 ;
        RECT  -3.0 286.8 97.5 288.3 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  0.0 44.4 7.2 45.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  0.0 64.8 7.2 66.3 ;
        RECT  0.0 75.0 7.2 76.5 ;
        RECT  0.0 54.6 7.2 56.1 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  123.45 6.3 124.95 151.2 ;
        RECT  133.65 6.3 135.15 151.2 ;
        RECT  127.2 0.0 128.7 30.0 ;
        RECT  137.4 0.0 138.9 30.0 ;
        RECT  79.2 85.65 95.25 87.15 ;
        RECT  79.2 113.85 95.25 115.35 ;
        RECT  79.2 142.05 95.25 143.55 ;
        RECT  79.2 170.25 95.25 171.75 ;
        RECT  0.0 44.4 7.2 45.9 ;
        RECT  0.0 64.8 7.2 66.3 ;
        RECT  0.0 75.0 7.2 76.5 ;
        RECT  0.0 54.6 7.2 56.1 ;
        RECT  123.3 151.2 125.1 153.0 ;
        RECT  133.5 151.2 135.3 153.0 ;
        RECT  123.3 151.2 125.1 153.0 ;
        RECT  123.3 151.2 125.1 153.0 ;
        RECT  133.5 151.2 135.3 153.0 ;
        RECT  133.5 151.2 135.3 153.0 ;
        RECT  137.1 30.9 138.9 32.7 ;
        RECT  126.9 30.9 128.7 32.7 ;
        RECT  126.9 30.9 128.7 32.7 ;
        RECT  126.9 30.9 128.7 32.7 ;
        RECT  137.1 30.9 138.9 32.7 ;
        RECT  137.1 30.9 138.9 32.7 ;
        RECT  126.9 31.2 128.7 33.0 ;
        RECT  137.1 31.2 138.9 33.0 ;
        RECT  7.2 44.4 9.0 46.2 ;
        RECT  7.2 64.8 9.0 66.6 ;
        RECT  7.2 75.0 9.0 76.8 ;
        RECT  7.2 54.6 9.0 56.4 ;
        RECT  7.2 75.0 9.0 76.8 ;
        RECT  7.2 75.0 9.0 76.8 ;
        RECT  7.2 64.8 9.0 66.6 ;
        RECT  7.2 64.8 9.0 66.6 ;
        RECT  7.2 54.6 9.0 56.4 ;
        RECT  7.2 54.6 9.0 56.4 ;
        RECT  7.2 44.4 9.0 46.2 ;
        RECT  7.2 44.4 9.0 46.2 ;
        RECT  123.45 5.55 125.25 7.35 ;
        RECT  133.65 5.55 135.45 7.35 ;
        RECT  127.2 0.0 129.0 1.8 ;
        RECT  137.4 0.0 139.2 1.8 ;
        RECT  78.3 85.5 80.1 87.3 ;
        RECT  94.35 85.5 96.15 87.3 ;
        RECT  78.3 113.7 80.1 115.5 ;
        RECT  94.35 113.7 96.15 115.5 ;
        RECT  78.3 141.9 80.1 143.7 ;
        RECT  94.35 141.9 96.15 143.7 ;
        RECT  78.3 170.1 80.1 171.9 ;
        RECT  94.35 170.1 96.15 171.9 ;
        RECT  -51.45 262.2 -49.95 301.05 ;
        RECT  -48.75 262.2 -47.25 290.25 ;
        RECT  -35.85 262.2 -34.35 292.95 ;
        RECT  -31.05 262.2 -29.55 295.65 ;
        RECT  -43.65 262.2 -42.15 287.55 ;
        RECT  -23.25 262.2 -21.75 287.55 ;
        RECT  -9.9 244.05 -8.4 303.75 ;
        RECT  -24.15 303.75 -22.65 327.6 ;
        RECT  -26.85 301.05 -25.35 330.6 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -48.9 203.1 -47.1 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -38.7 203.1 -36.9 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -28.5 203.1 -26.7 204.9 ;
        RECT  -51.6 261.3 -49.8 263.1 ;
        RECT  -51.6 300.15 -49.8 301.95 ;
        RECT  -48.9 261.3 -47.1 263.1 ;
        RECT  -48.9 289.35 -47.1 291.15 ;
        RECT  -36.0 261.3 -34.2 263.1 ;
        RECT  -36.0 292.05 -34.2 293.85 ;
        RECT  -31.2 261.3 -29.4 263.1 ;
        RECT  -31.2 294.75 -29.4 296.55 ;
        RECT  -43.8 261.3 -42.0 263.1 ;
        RECT  -43.8 286.65 -42.0 288.45 ;
        RECT  -23.4 261.3 -21.6 263.1 ;
        RECT  -23.4 286.65 -21.6 288.45 ;
        RECT  -10.05 243.15 -8.25 244.95 ;
        RECT  -10.05 302.85 -8.25 304.65 ;
        RECT  -24.3 326.7 -22.5 328.5 ;
        RECT  -24.3 302.85 -22.5 304.65 ;
        RECT  -27.0 329.7 -25.2 331.5 ;
        RECT  -27.0 300.15 -25.2 301.95 ;
        RECT  115.5 342.0 117.3 343.8 ;
        RECT  -4.8 342.15 -3.0 343.95 ;
        RECT  112.8 361.8 114.6 363.6 ;
        RECT  -4.8 361.95 -3.0 363.75 ;
        RECT  107.4 322.2 109.2 324.0 ;
        RECT  -4.8 322.35 -3.0 324.15 ;
        RECT  104.7 339.3 106.5 341.1 ;
        RECT  -4.8 339.45 -3.0 341.25 ;
        RECT  110.1 302.85 111.9 304.65 ;
        RECT  -4.8 303.0 -3.0 304.8 ;
        RECT  102.0 283.95 103.8 285.75 ;
        RECT  -4.8 284.1 -3.0 285.9 ;
        RECT  96.6 286.65 98.4 288.45 ;
        RECT  -4.8 286.8 -3.0 288.6 ;
    END
END    sram_2_16_1_scn3me_subm
END    LIBRARY
