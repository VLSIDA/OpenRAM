magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1260 -1286 1410 1358
<< scnmos >>
rect 60 0 90 72
<< ndiff >>
rect 0 0 60 72
rect 90 0 150 72
<< poly >>
rect 60 72 90 98
rect 60 -26 90 0
<< locali >>
rect 8 3 42 69
rect 108 3 142 69
use contact_17  contact_17_0
timestamp 1595931502
transform 1 0 100 0 1 3
box 0 0 50 66
use contact_17  contact_17_1
timestamp 1595931502
transform 1 0 0 0 1 3
box 0 0 50 66
<< labels >>
rlabel poly s 75 36 75 36 4 G
rlabel corelocali s 25 36 25 36 4 S
rlabel corelocali s 125 36 125 36 4 D
<< properties >>
string FIXED_BBOX -25 -26 175 98
<< end >>
