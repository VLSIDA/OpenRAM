magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1296 -1277 3416 2731
<< nwell >>
rect -36 679 2156 1471
<< locali >>
rect 0 1397 2120 1431
rect 64 636 98 702
rect 547 690 707 724
rect 196 652 449 686
rect 547 669 581 690
rect 915 674 1187 708
rect 1613 674 1647 708
rect 0 -17 2120 17
use pinv_4  pinv_4_0
timestamp 1595931502
transform 1 0 0 0 1 0
box -36 -17 404 1471
use pinv_12  pinv_12_0
timestamp 1595931502
transform 1 0 1106 0 1 0
box -36 -17 1050 1471
use pinv_11  pinv_11_0
timestamp 1595931502
transform 1 0 626 0 1 0
box -36 -17 516 1471
use pinv_7  pinv_7_0
timestamp 1595931502
transform 1 0 368 0 1 0
box -36 -17 294 1471
<< labels >>
rlabel corelocali s 1060 0 1060 0 4 gnd
rlabel corelocali s 1630 691 1630 691 4 Z
rlabel corelocali s 1060 1414 1060 1414 4 vdd
rlabel corelocali s 81 669 81 669 4 A
<< properties >>
string FIXED_BBOX 0 0 2120 1414
<< end >>
